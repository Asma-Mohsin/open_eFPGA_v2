magic
tech sky130A
magscale 1 2
timestamp 1733616289
<< viali >>
rect 1593 43401 1627 43435
rect 2329 43401 2363 43435
rect 6101 43401 6135 43435
rect 7205 43401 7239 43435
rect 8217 43401 8251 43435
rect 8677 43401 8711 43435
rect 9137 43401 9171 43435
rect 9689 43401 9723 43435
rect 10057 43401 10091 43435
rect 14289 43401 14323 43435
rect 18337 43401 18371 43435
rect 20361 43401 20395 43435
rect 20729 43401 20763 43435
rect 22385 43401 22419 43435
rect 23765 43401 23799 43435
rect 2697 43333 2731 43367
rect 3065 43333 3099 43367
rect 3617 43333 3651 43367
rect 12449 43333 12483 43367
rect 13185 43333 13219 43367
rect 13553 43333 13587 43367
rect 15853 43333 15887 43367
rect 16773 43333 16807 43367
rect 16957 43333 16991 43367
rect 17141 43333 17175 43367
rect 21649 43333 21683 43367
rect 1409 43265 1443 43299
rect 2053 43265 2087 43299
rect 3249 43265 3283 43299
rect 4075 43265 4109 43299
rect 5273 43265 5307 43299
rect 5825 43265 5859 43299
rect 6377 43265 6411 43299
rect 6929 43265 6963 43299
rect 7481 43265 7515 43299
rect 8493 43265 8527 43299
rect 8953 43265 8987 43299
rect 9413 43265 9447 43299
rect 9965 43265 9999 43299
rect 10425 43265 10459 43299
rect 10977 43265 11011 43299
rect 11529 43265 11563 43299
rect 12081 43265 12115 43299
rect 12817 43265 12851 43299
rect 14105 43265 14139 43299
rect 14473 43265 14507 43299
rect 14841 43265 14875 43299
rect 16129 43265 16163 43299
rect 17417 43265 17451 43299
rect 17969 43265 18003 43299
rect 18245 43265 18279 43299
rect 18521 43265 18555 43299
rect 18797 43265 18831 43299
rect 19073 43265 19107 43299
rect 19441 43265 19475 43299
rect 19717 43265 19751 43299
rect 19993 43265 20027 43299
rect 20177 43265 20211 43299
rect 20637 43265 20671 43299
rect 21281 43265 21315 43299
rect 21833 43265 21867 43299
rect 22293 43265 22327 43299
rect 22845 43265 22879 43299
rect 23489 43265 23523 43299
rect 23673 43265 23707 43299
rect 3801 43197 3835 43231
rect 5549 43197 5583 43231
rect 10609 43197 10643 43231
rect 15117 43197 15151 43231
rect 4813 43129 4847 43163
rect 6561 43129 6595 43163
rect 7757 43129 7791 43163
rect 11161 43129 11195 43163
rect 13001 43129 13035 43163
rect 13369 43129 13403 43163
rect 18889 43129 18923 43163
rect 22017 43129 22051 43163
rect 23305 43129 23339 43163
rect 11713 43061 11747 43095
rect 12265 43061 12299 43095
rect 12541 43061 12575 43095
rect 13645 43061 13679 43095
rect 14657 43061 14691 43095
rect 15945 43061 15979 43095
rect 16313 43061 16347 43095
rect 17233 43061 17267 43095
rect 17601 43061 17635 43095
rect 17785 43061 17819 43095
rect 18061 43061 18095 43095
rect 18613 43061 18647 43095
rect 19257 43061 19291 43095
rect 19533 43061 19567 43095
rect 19809 43061 19843 43095
rect 22937 43061 22971 43095
rect 2973 42857 3007 42891
rect 7941 42857 7975 42891
rect 8493 42857 8527 42891
rect 9505 42857 9539 42891
rect 20269 42857 20303 42891
rect 20545 42857 20579 42891
rect 22017 42857 22051 42891
rect 23489 42857 23523 42891
rect 3801 42789 3835 42823
rect 10793 42789 10827 42823
rect 14473 42789 14507 42823
rect 19993 42789 20027 42823
rect 1869 42721 1903 42755
rect 7389 42721 7423 42755
rect 22569 42721 22603 42755
rect 3985 42653 4019 42687
rect 4077 42653 4111 42687
rect 4351 42653 4385 42687
rect 5457 42653 5491 42687
rect 5731 42653 5765 42687
rect 7849 42653 7883 42687
rect 8953 42653 8987 42687
rect 9873 42653 9907 42687
rect 10241 42653 10275 42687
rect 10609 42653 10643 42687
rect 11713 42653 11747 42687
rect 11805 42653 11839 42687
rect 12633 42653 12667 42687
rect 13737 42653 13771 42687
rect 14289 42653 14323 42687
rect 15117 42653 15151 42687
rect 16313 42653 16347 42687
rect 17049 42653 17083 42687
rect 17417 42653 17451 42687
rect 17785 42653 17819 42687
rect 18153 42653 18187 42687
rect 18337 42653 18371 42687
rect 18889 42653 18923 42687
rect 19349 42653 19383 42687
rect 20177 42653 20211 42687
rect 20453 42653 20487 42687
rect 20729 42653 20763 42687
rect 21005 42653 21039 42687
rect 22845 42653 22879 42687
rect 23949 42653 23983 42687
rect 1593 42585 1627 42619
rect 2329 42585 2363 42619
rect 2697 42585 2731 42619
rect 3249 42585 3283 42619
rect 7113 42585 7147 42619
rect 8401 42585 8435 42619
rect 9413 42585 9447 42619
rect 16497 42585 16531 42619
rect 16681 42585 16715 42619
rect 17969 42585 18003 42619
rect 18521 42585 18555 42619
rect 19533 42585 19567 42619
rect 19717 42585 19751 42619
rect 21189 42585 21223 42619
rect 21557 42585 21591 42619
rect 21741 42585 21775 42619
rect 22293 42585 22327 42619
rect 23397 42585 23431 42619
rect 3525 42517 3559 42551
rect 5089 42517 5123 42551
rect 6469 42517 6503 42551
rect 9137 42517 9171 42551
rect 10057 42517 10091 42551
rect 10425 42517 10459 42551
rect 11529 42517 11563 42551
rect 11989 42517 12023 42551
rect 12817 42517 12851 42551
rect 13921 42517 13955 42551
rect 15301 42517 15335 42551
rect 16773 42517 16807 42551
rect 17141 42517 17175 42551
rect 17509 42517 17543 42551
rect 18613 42517 18647 42551
rect 18981 42517 19015 42551
rect 19809 42517 19843 42551
rect 20821 42517 20855 42551
rect 22937 42517 22971 42551
rect 24133 42517 24167 42551
rect 2329 42313 2363 42347
rect 5917 42313 5951 42347
rect 6653 42313 6687 42347
rect 9137 42313 9171 42347
rect 9965 42313 9999 42347
rect 10241 42313 10275 42347
rect 21557 42313 21591 42347
rect 22293 42313 22327 42347
rect 22845 42313 22879 42347
rect 23949 42313 23983 42347
rect 2697 42245 2731 42279
rect 3801 42245 3835 42279
rect 18429 42245 18463 42279
rect 20453 42245 20487 42279
rect 23489 42245 23523 42279
rect 1409 42177 1443 42211
rect 2053 42177 2087 42211
rect 2973 42177 3007 42211
rect 3065 42177 3099 42211
rect 3433 42177 3467 42211
rect 4443 42177 4477 42211
rect 5825 42177 5859 42211
rect 6469 42177 6503 42211
rect 7111 42177 7145 42211
rect 8309 42177 8343 42211
rect 9045 42177 9079 42211
rect 9321 42177 9355 42211
rect 9689 42177 9723 42211
rect 10149 42177 10183 42211
rect 10425 42177 10459 42211
rect 18705 42177 18739 42211
rect 20729 42177 20763 42211
rect 21005 42177 21039 42211
rect 21281 42177 21315 42211
rect 21373 42177 21407 42211
rect 22017 42177 22051 42211
rect 22569 42177 22603 42211
rect 23121 42177 23155 42211
rect 23673 42177 23707 42211
rect 1593 42109 1627 42143
rect 4169 42109 4203 42143
rect 6837 42109 6871 42143
rect 8861 42041 8895 42075
rect 20545 42041 20579 42075
rect 3985 41973 4019 42007
rect 5181 41973 5215 42007
rect 7849 41973 7883 42007
rect 8401 41973 8435 42007
rect 18521 41973 18555 42007
rect 20821 41973 20855 42007
rect 21097 41973 21131 42007
rect 3341 41769 3375 41803
rect 4077 41769 4111 41803
rect 7297 41769 7331 41803
rect 8953 41769 8987 41803
rect 9229 41769 9263 41803
rect 19901 41769 19935 41803
rect 20637 41769 20671 41803
rect 21189 41769 21223 41803
rect 21741 41769 21775 41803
rect 23949 41769 23983 41803
rect 20361 41701 20395 41735
rect 21465 41701 21499 41735
rect 22477 41701 22511 41735
rect 23581 41701 23615 41735
rect 2329 41633 2363 41667
rect 7481 41633 7515 41667
rect 1409 41565 1443 41599
rect 1777 41565 1811 41599
rect 2603 41565 2637 41599
rect 3893 41565 3927 41599
rect 4537 41565 4571 41599
rect 5445 41565 5479 41599
rect 7113 41565 7147 41599
rect 7755 41565 7789 41599
rect 9137 41565 9171 41599
rect 9413 41565 9447 41599
rect 19809 41565 19843 41599
rect 20085 41565 20119 41599
rect 20545 41565 20579 41599
rect 20821 41565 20855 41599
rect 21097 41565 21131 41599
rect 21373 41565 21407 41599
rect 21649 41565 21683 41599
rect 21925 41565 21959 41599
rect 23121 41565 23155 41599
rect 2053 41497 2087 41531
rect 5089 41497 5123 41531
rect 5365 41497 5399 41531
rect 5825 41497 5859 41531
rect 6653 41497 6687 41531
rect 19349 41497 19383 41531
rect 22201 41497 22235 41531
rect 22753 41497 22787 41531
rect 23305 41497 23339 41531
rect 23857 41497 23891 41531
rect 1593 41429 1627 41463
rect 6193 41429 6227 41463
rect 6377 41429 6411 41463
rect 6745 41429 6779 41463
rect 8493 41429 8527 41463
rect 19441 41429 19475 41463
rect 19625 41429 19659 41463
rect 20913 41429 20947 41463
rect 2789 41225 2823 41259
rect 4537 41225 4571 41259
rect 5825 41225 5859 41259
rect 6009 41225 6043 41259
rect 8677 41225 8711 41259
rect 20361 41225 20395 41259
rect 20913 41225 20947 41259
rect 21189 41225 21223 41259
rect 21465 41225 21499 41259
rect 22293 41225 22327 41259
rect 23397 41225 23431 41259
rect 23949 41225 23983 41259
rect 4905 41157 4939 41191
rect 5273 41157 5307 41191
rect 5641 41157 5675 41191
rect 7573 41157 7607 41191
rect 7941 41157 7975 41191
rect 1409 41089 1443 41123
rect 2513 41089 2547 41123
rect 3247 41089 3281 41123
rect 4813 41089 4847 41123
rect 6193 41089 6227 41123
rect 6469 41089 6503 41123
rect 7297 41089 7331 41123
rect 7849 41089 7883 41123
rect 8309 41089 8343 41123
rect 19257 41089 19291 41123
rect 20545 41089 20579 41123
rect 20821 41089 20855 41123
rect 21097 41089 21131 41123
rect 21373 41089 21407 41123
rect 21649 41089 21683 41123
rect 22201 41089 22235 41123
rect 22477 41089 22511 41123
rect 22661 41089 22695 41123
rect 23121 41089 23155 41123
rect 23673 41089 23707 41123
rect 2145 41021 2179 41055
rect 2973 41021 3007 41055
rect 3985 40953 4019 40987
rect 20637 40953 20671 40987
rect 22017 40953 22051 40987
rect 6561 40885 6595 40919
rect 8861 40885 8895 40919
rect 19073 40885 19107 40919
rect 22845 40885 22879 40919
rect 3433 40681 3467 40715
rect 3985 40681 4019 40715
rect 4537 40681 4571 40715
rect 5641 40681 5675 40715
rect 6009 40681 6043 40715
rect 7205 40681 7239 40715
rect 18429 40681 18463 40715
rect 21557 40681 21591 40715
rect 21649 40681 21683 40715
rect 21925 40681 21959 40715
rect 22201 40681 22235 40715
rect 23121 40681 23155 40715
rect 24133 40681 24167 40715
rect 6929 40613 6963 40647
rect 21097 40613 21131 40647
rect 23581 40613 23615 40647
rect 2145 40545 2179 40579
rect 2421 40545 2455 40579
rect 2559 40545 2593 40579
rect 3341 40545 3375 40579
rect 1501 40477 1535 40511
rect 1685 40477 1719 40511
rect 2697 40477 2731 40511
rect 3617 40477 3651 40511
rect 6193 40477 6227 40511
rect 7113 40477 7147 40511
rect 7389 40477 7423 40511
rect 18613 40477 18647 40511
rect 21281 40477 21315 40511
rect 21373 40477 21407 40511
rect 21833 40477 21867 40511
rect 22109 40477 22143 40511
rect 22385 40477 22419 40511
rect 22845 40477 22879 40511
rect 23305 40477 23339 40511
rect 23397 40477 23431 40511
rect 3893 40409 3927 40443
rect 4445 40409 4479 40443
rect 4997 40409 5031 40443
rect 5549 40409 5583 40443
rect 23857 40409 23891 40443
rect 5089 40341 5123 40375
rect 6561 40341 6595 40375
rect 22661 40341 22695 40375
rect 2605 40137 2639 40171
rect 21465 40137 21499 40171
rect 22017 40137 22051 40171
rect 22293 40137 22327 40171
rect 22937 40137 22971 40171
rect 23213 40137 23247 40171
rect 2973 40069 3007 40103
rect 5917 40069 5951 40103
rect 23857 40069 23891 40103
rect 1867 40001 1901 40035
rect 4227 40001 4261 40035
rect 6651 40001 6685 40035
rect 21649 40001 21683 40035
rect 22201 40001 22235 40035
rect 22477 40001 22511 40035
rect 22753 40001 22787 40035
rect 23121 40001 23155 40035
rect 23397 40001 23431 40035
rect 23673 40001 23707 40035
rect 1593 39933 1627 39967
rect 3801 39933 3835 39967
rect 3985 39933 4019 39967
rect 6377 39933 6411 39967
rect 5641 39865 5675 39899
rect 23489 39865 23523 39899
rect 4997 39797 5031 39831
rect 7389 39797 7423 39831
rect 24133 39797 24167 39831
rect 1685 39593 1719 39627
rect 4353 39593 4387 39627
rect 9137 39593 9171 39627
rect 22845 39593 22879 39627
rect 23673 39593 23707 39627
rect 2053 39525 2087 39559
rect 9045 39525 9079 39559
rect 9689 39525 9723 39559
rect 19349 39525 19383 39559
rect 22385 39525 22419 39559
rect 23397 39525 23431 39559
rect 3985 39457 4019 39491
rect 9229 39457 9263 39491
rect 9413 39457 9447 39491
rect 9873 39457 9907 39491
rect 2329 39389 2363 39423
rect 2603 39389 2637 39423
rect 3801 39389 3835 39423
rect 4537 39389 4571 39423
rect 5549 39389 5583 39423
rect 6837 39389 6871 39423
rect 7111 39389 7145 39423
rect 8953 39389 8987 39423
rect 9321 39389 9355 39423
rect 9505 39389 9539 39423
rect 9597 39389 9631 39423
rect 10147 39389 10181 39423
rect 19533 39389 19567 39423
rect 22569 39389 22603 39423
rect 23029 39389 23063 39423
rect 23305 39389 23339 39423
rect 23581 39389 23615 39423
rect 23857 39389 23891 39423
rect 23949 39389 23983 39423
rect 1869 39321 1903 39355
rect 5089 39321 5123 39355
rect 5181 39321 5215 39355
rect 3341 39253 3375 39287
rect 4813 39253 4847 39287
rect 5917 39253 5951 39287
rect 6101 39253 6135 39287
rect 7849 39253 7883 39287
rect 10885 39253 10919 39287
rect 23121 39253 23155 39287
rect 24133 39253 24167 39287
rect 5917 39049 5951 39083
rect 8769 39049 8803 39083
rect 9781 39049 9815 39083
rect 20361 39049 20395 39083
rect 21833 39049 21867 39083
rect 22937 39049 22971 39083
rect 10057 38981 10091 39015
rect 10149 38981 10183 39015
rect 10885 38981 10919 39015
rect 23857 38981 23891 39015
rect 1667 38943 1701 38977
rect 2789 38913 2823 38947
rect 3801 38913 3835 38947
rect 4077 38913 4111 38947
rect 4353 38913 4387 38947
rect 4905 38913 4939 38947
rect 5179 38923 5213 38957
rect 6929 38913 6963 38947
rect 7665 38913 7699 38947
rect 7782 38913 7816 38947
rect 7941 38913 7975 38947
rect 8953 38913 8987 38947
rect 9321 38913 9355 38947
rect 10517 38913 10551 38947
rect 11529 38913 11563 38947
rect 20545 38913 20579 38947
rect 22017 38913 22051 38947
rect 23121 38913 23155 38947
rect 23397 38913 23431 38947
rect 1409 38845 1443 38879
rect 3617 38845 3651 38879
rect 4629 38845 4663 38879
rect 6745 38845 6779 38879
rect 7389 38845 7423 38879
rect 2421 38777 2455 38811
rect 23213 38777 23247 38811
rect 8585 38709 8619 38743
rect 11069 38709 11103 38743
rect 11713 38709 11747 38743
rect 24133 38709 24167 38743
rect 8309 38505 8343 38539
rect 10241 38505 10275 38539
rect 18613 38505 18647 38539
rect 19717 38505 19751 38539
rect 22661 38505 22695 38539
rect 4813 38437 4847 38471
rect 7113 38437 7147 38471
rect 2237 38369 2271 38403
rect 3801 38369 3835 38403
rect 7389 38369 7423 38403
rect 7665 38369 7699 38403
rect 9229 38369 9263 38403
rect 2421 38301 2455 38335
rect 2973 38301 3007 38335
rect 4075 38301 4109 38335
rect 5181 38301 5215 38335
rect 6469 38301 6503 38335
rect 6653 38301 6687 38335
rect 7506 38301 7540 38335
rect 9137 38301 9171 38335
rect 9503 38301 9537 38335
rect 18797 38301 18831 38335
rect 19901 38301 19935 38335
rect 22845 38301 22879 38335
rect 23949 38301 23983 38335
rect 1409 38233 1443 38267
rect 2697 38233 2731 38267
rect 3249 38233 3283 38267
rect 5457 38233 5491 38267
rect 8953 38165 8987 38199
rect 24133 38165 24167 38199
rect 9413 37961 9447 37995
rect 21925 37961 21959 37995
rect 23397 37961 23431 37995
rect 23673 37961 23707 37995
rect 1775 37825 1809 37859
rect 3247 37825 3281 37859
rect 4353 37825 4387 37859
rect 4627 37825 4661 37859
rect 8643 37825 8677 37859
rect 11803 37825 11837 37859
rect 22109 37825 22143 37859
rect 23581 37825 23615 37859
rect 23857 37825 23891 37859
rect 23949 37825 23983 37859
rect 1501 37757 1535 37791
rect 2973 37757 3007 37791
rect 8401 37757 8435 37791
rect 11529 37757 11563 37791
rect 2513 37621 2547 37655
rect 3985 37621 4019 37655
rect 5365 37621 5399 37655
rect 12541 37621 12575 37655
rect 24133 37621 24167 37655
rect 3249 37417 3283 37451
rect 23397 37417 23431 37451
rect 23673 37417 23707 37451
rect 6285 37349 6319 37383
rect 11989 37349 12023 37383
rect 21741 37349 21775 37383
rect 2053 37281 2087 37315
rect 2329 37281 2363 37315
rect 2446 37281 2480 37315
rect 2605 37281 2639 37315
rect 1409 37213 1443 37247
rect 1593 37213 1627 37247
rect 3801 37213 3835 37247
rect 5273 37213 5307 37247
rect 6929 37213 6963 37247
rect 7203 37213 7237 37247
rect 11069 37213 11103 37247
rect 21005 37213 21039 37247
rect 21925 37213 21959 37247
rect 23581 37213 23615 37247
rect 23857 37213 23891 37247
rect 23949 37213 23983 37247
rect 4077 37145 4111 37179
rect 4997 37145 5031 37179
rect 5365 37145 5399 37179
rect 5733 37145 5767 37179
rect 6101 37145 6135 37179
rect 10701 37145 10735 37179
rect 10977 37145 11011 37179
rect 11437 37145 11471 37179
rect 11805 37145 11839 37179
rect 7941 37077 7975 37111
rect 20821 37077 20855 37111
rect 24133 37077 24167 37111
rect 2421 36873 2455 36907
rect 5917 36873 5951 36907
rect 10977 36873 11011 36907
rect 20177 36873 20211 36907
rect 4169 36805 4203 36839
rect 7481 36805 7515 36839
rect 7757 36805 7791 36839
rect 7849 36805 7883 36839
rect 8585 36805 8619 36839
rect 1683 36737 1717 36771
rect 2789 36737 2823 36771
rect 3341 36737 3375 36771
rect 3893 36737 3927 36771
rect 5179 36737 5213 36771
rect 8217 36737 8251 36771
rect 9965 36737 9999 36771
rect 10239 36737 10273 36771
rect 20361 36737 20395 36771
rect 21189 36737 21223 36771
rect 23673 36737 23707 36771
rect 23949 36737 23983 36771
rect 1409 36669 1443 36703
rect 2973 36669 3007 36703
rect 3525 36669 3559 36703
rect 4629 36669 4663 36703
rect 4905 36669 4939 36703
rect 21005 36601 21039 36635
rect 23489 36601 23523 36635
rect 8769 36533 8803 36567
rect 24133 36533 24167 36567
rect 21281 36329 21315 36363
rect 3341 36261 3375 36295
rect 23397 36261 23431 36295
rect 1685 36193 1719 36227
rect 2329 36193 2363 36227
rect 7481 36193 7515 36227
rect 9045 36193 9079 36227
rect 10425 36193 10459 36227
rect 1409 36125 1443 36159
rect 2587 36095 2621 36129
rect 4353 36125 4387 36159
rect 5457 36125 5491 36159
rect 7723 36125 7757 36159
rect 9287 36125 9321 36159
rect 10699 36125 10733 36159
rect 14565 36125 14599 36159
rect 14749 36125 14783 36159
rect 20637 36125 20671 36159
rect 21465 36125 21499 36159
rect 23305 36125 23339 36159
rect 23581 36125 23615 36159
rect 4261 36057 4295 36091
rect 4721 36057 4755 36091
rect 5733 36057 5767 36091
rect 23857 36057 23891 36091
rect 24225 36057 24259 36091
rect 3985 35989 4019 36023
rect 5089 35989 5123 36023
rect 5273 35989 5307 36023
rect 8493 35989 8527 36023
rect 10057 35989 10091 36023
rect 11437 35989 11471 36023
rect 14749 35989 14783 36023
rect 20453 35989 20487 36023
rect 23121 35989 23155 36023
rect 3065 35785 3099 35819
rect 8401 35785 8435 35819
rect 14473 35785 14507 35819
rect 15117 35785 15151 35819
rect 21833 35785 21867 35819
rect 22661 35785 22695 35819
rect 23673 35785 23707 35819
rect 3341 35717 3375 35751
rect 3433 35717 3467 35751
rect 3801 35717 3835 35751
rect 8953 35717 8987 35751
rect 9321 35717 9355 35751
rect 10057 35717 10091 35751
rect 1683 35649 1717 35683
rect 4193 35649 4227 35683
rect 5179 35649 5213 35683
rect 7631 35649 7665 35683
rect 9229 35649 9263 35683
rect 9689 35649 9723 35683
rect 11529 35649 11563 35683
rect 13461 35649 13495 35683
rect 13719 35679 13753 35713
rect 14841 35649 14875 35683
rect 15209 35649 15243 35683
rect 20545 35649 20579 35683
rect 22017 35649 22051 35683
rect 22569 35649 22603 35683
rect 22845 35649 22879 35683
rect 23581 35649 23615 35683
rect 23857 35649 23891 35683
rect 23949 35649 23983 35683
rect 1409 35581 1443 35615
rect 4905 35581 4939 35615
rect 7389 35581 7423 35615
rect 11345 35581 11379 35615
rect 11713 35581 11747 35615
rect 12173 35581 12207 35615
rect 12449 35581 12483 35615
rect 12566 35581 12600 35615
rect 12725 35581 12759 35615
rect 15117 35581 15151 35615
rect 10241 35513 10275 35547
rect 14933 35513 14967 35547
rect 15301 35513 15335 35547
rect 2421 35445 2455 35479
rect 4353 35445 4387 35479
rect 5917 35445 5951 35479
rect 13369 35445 13403 35479
rect 20361 35445 20395 35479
rect 22385 35445 22419 35479
rect 23305 35445 23339 35479
rect 23397 35445 23431 35479
rect 24133 35445 24167 35479
rect 12173 35241 12207 35275
rect 14749 35241 14783 35275
rect 15025 35241 15059 35275
rect 22845 35241 22879 35275
rect 23673 35241 23707 35275
rect 2329 35173 2363 35207
rect 19349 35173 19383 35207
rect 2605 35105 2639 35139
rect 2722 35105 2756 35139
rect 11161 35105 11195 35139
rect 1685 35037 1719 35071
rect 1869 35037 1903 35071
rect 2881 35037 2915 35071
rect 3525 35037 3559 35071
rect 3801 35037 3835 35071
rect 4353 35037 4387 35071
rect 5641 35037 5675 35071
rect 6009 35037 6043 35071
rect 6745 35037 6779 35071
rect 7019 35037 7053 35071
rect 11435 35037 11469 35071
rect 14933 35037 14967 35071
rect 15209 35037 15243 35071
rect 19533 35037 19567 35071
rect 19993 35037 20027 35071
rect 20545 35037 20579 35071
rect 23029 35037 23063 35071
rect 23857 35037 23891 35071
rect 23949 35037 23983 35071
rect 4077 34969 4111 35003
rect 4629 34969 4663 35003
rect 5549 34969 5583 35003
rect 5273 34901 5307 34935
rect 6377 34901 6411 34935
rect 6561 34901 6595 34935
rect 7757 34901 7791 34935
rect 20085 34901 20119 34935
rect 20361 34901 20395 34935
rect 23305 34901 23339 34935
rect 24133 34901 24167 34935
rect 2789 34697 2823 34731
rect 5733 34697 5767 34731
rect 9873 34697 9907 34731
rect 20269 34697 20303 34731
rect 21833 34697 21867 34731
rect 22661 34697 22695 34731
rect 23397 34697 23431 34731
rect 19156 34629 19190 34663
rect 20913 34629 20947 34663
rect 21097 34629 21131 34663
rect 23857 34629 23891 34663
rect 2035 34591 2069 34625
rect 3415 34591 3449 34625
rect 4721 34561 4755 34595
rect 4995 34561 5029 34595
rect 6895 34561 6929 34595
rect 9597 34561 9631 34595
rect 18889 34561 18923 34595
rect 20545 34561 20579 34595
rect 20729 34561 20763 34595
rect 21005 34561 21039 34595
rect 21189 34561 21223 34595
rect 22017 34561 22051 34595
rect 22845 34561 22879 34595
rect 23581 34561 23615 34595
rect 1777 34493 1811 34527
rect 3157 34493 3191 34527
rect 6653 34493 6687 34527
rect 9873 34493 9907 34527
rect 24133 34493 24167 34527
rect 20545 34425 20579 34459
rect 4169 34357 4203 34391
rect 7665 34357 7699 34391
rect 9689 34357 9723 34391
rect 5365 34153 5399 34187
rect 8677 34153 8711 34187
rect 10333 34153 10367 34187
rect 10793 34153 10827 34187
rect 20453 34153 20487 34187
rect 21465 34153 21499 34187
rect 9045 34085 9079 34119
rect 23673 34085 23707 34119
rect 3341 34017 3375 34051
rect 11253 34017 11287 34051
rect 19441 34017 19475 34051
rect 1409 33949 1443 33983
rect 1961 33949 1995 33983
rect 2513 33949 2547 33983
rect 3065 33949 3099 33983
rect 6837 33949 6871 33983
rect 6929 33949 6963 33983
rect 8585 33949 8619 33983
rect 9229 33949 9263 33983
rect 9321 33949 9355 33983
rect 9595 33949 9629 33983
rect 10701 33949 10735 33983
rect 10885 33949 10919 33983
rect 11527 33949 11561 33983
rect 14841 33949 14875 33983
rect 15115 33949 15149 33983
rect 19715 33949 19749 33983
rect 21649 33949 21683 33983
rect 23857 33949 23891 33983
rect 23949 33949 23983 33983
rect 1685 33881 1719 33915
rect 2237 33881 2271 33915
rect 2789 33881 2823 33915
rect 4353 33881 4387 33915
rect 4445 33881 4479 33915
rect 4813 33881 4847 33915
rect 7297 33881 7331 33915
rect 4077 33813 4111 33847
rect 5181 33813 5215 33847
rect 6561 33813 6595 33847
rect 7665 33813 7699 33847
rect 7849 33813 7883 33847
rect 12265 33813 12299 33847
rect 15853 33813 15887 33847
rect 24133 33813 24167 33847
rect 4169 33609 4203 33643
rect 5273 33609 5307 33643
rect 9689 33609 9723 33643
rect 11713 33609 11747 33643
rect 16497 33609 16531 33643
rect 21649 33609 21683 33643
rect 23213 33609 23247 33643
rect 11989 33541 12023 33575
rect 12081 33541 12115 33575
rect 12817 33541 12851 33575
rect 20514 33541 20548 33575
rect 1683 33473 1717 33507
rect 2789 33473 2823 33507
rect 3985 33473 4019 33507
rect 4261 33473 4295 33507
rect 4503 33483 4537 33517
rect 7907 33473 7941 33507
rect 9873 33473 9907 33507
rect 10331 33473 10365 33507
rect 12449 33473 12483 33507
rect 13551 33473 13585 33507
rect 15577 33473 15611 33507
rect 20269 33473 20303 33507
rect 22017 33473 22051 33507
rect 22109 33473 22143 33507
rect 22569 33473 22603 33507
rect 23121 33473 23155 33507
rect 23397 33473 23431 33507
rect 23765 33473 23799 33507
rect 23949 33473 23983 33507
rect 1409 33405 1443 33439
rect 3065 33405 3099 33439
rect 7665 33405 7699 33439
rect 10057 33405 10091 33439
rect 13277 33405 13311 33439
rect 14657 33405 14691 33439
rect 14841 33405 14875 33439
rect 15301 33405 15335 33439
rect 15694 33405 15728 33439
rect 15853 33405 15887 33439
rect 11069 33337 11103 33371
rect 21833 33337 21867 33371
rect 22937 33337 22971 33371
rect 23581 33337 23615 33371
rect 2421 33269 2455 33303
rect 8677 33269 8711 33303
rect 13001 33269 13035 33303
rect 14289 33269 14323 33303
rect 22201 33269 22235 33303
rect 22385 33269 22419 33303
rect 24133 33269 24167 33303
rect 3157 33065 3191 33099
rect 13553 33065 13587 33099
rect 15945 33065 15979 33099
rect 17049 33065 17083 33099
rect 22569 33065 22603 33099
rect 22661 33065 22695 33099
rect 14749 32997 14783 33031
rect 22109 32997 22143 33031
rect 23673 32997 23707 33031
rect 7113 32929 7147 32963
rect 12541 32929 12575 32963
rect 15025 32929 15059 32963
rect 15142 32929 15176 32963
rect 16037 32929 16071 32963
rect 21097 32929 21131 32963
rect 22753 32929 22787 32963
rect 22937 32929 22971 32963
rect 1593 32861 1627 32895
rect 1851 32831 1885 32865
rect 2973 32861 3007 32895
rect 4629 32861 4663 32895
rect 7355 32861 7389 32895
rect 12081 32861 12115 32895
rect 12799 32861 12833 32895
rect 14105 32861 14139 32895
rect 14289 32861 14323 32895
rect 15301 32861 15335 32895
rect 16311 32861 16345 32895
rect 21371 32861 21405 32895
rect 22477 32861 22511 32895
rect 22845 32861 22879 32895
rect 23029 32861 23063 32895
rect 23305 32861 23339 32895
rect 23857 32861 23891 32895
rect 23949 32861 23983 32895
rect 3801 32793 3835 32827
rect 2605 32725 2639 32759
rect 8125 32725 8159 32759
rect 12173 32725 12207 32759
rect 23121 32725 23155 32759
rect 24133 32725 24167 32759
rect 9413 32521 9447 32555
rect 15025 32521 15059 32555
rect 22569 32521 22603 32555
rect 23213 32521 23247 32555
rect 3617 32453 3651 32487
rect 1593 32385 1627 32419
rect 2329 32385 2363 32419
rect 2605 32385 2639 32419
rect 3341 32385 3375 32419
rect 3893 32385 3927 32419
rect 5147 32385 5181 32419
rect 7573 32385 7607 32419
rect 8769 32385 8803 32419
rect 13369 32385 13403 32419
rect 14381 32385 14415 32419
rect 18889 32385 18923 32419
rect 19145 32385 19179 32419
rect 22753 32385 22787 32419
rect 23397 32385 23431 32419
rect 23673 32385 23707 32419
rect 23949 32385 23983 32419
rect 1409 32317 1443 32351
rect 2053 32317 2087 32351
rect 2467 32317 2501 32351
rect 4905 32317 4939 32351
rect 7757 32317 7791 32351
rect 8217 32317 8251 32351
rect 8493 32317 8527 32351
rect 8631 32317 8665 32351
rect 13185 32317 13219 32351
rect 13829 32317 13863 32351
rect 14105 32317 14139 32351
rect 14222 32317 14256 32351
rect 23857 32249 23891 32283
rect 3249 32181 3283 32215
rect 4077 32181 4111 32215
rect 5917 32181 5951 32215
rect 20269 32181 20303 32215
rect 24133 32181 24167 32215
rect 6745 31977 6779 32011
rect 8769 31977 8803 32011
rect 23213 31977 23247 32011
rect 2237 31909 2271 31943
rect 4813 31909 4847 31943
rect 7573 31909 7607 31943
rect 10425 31909 10459 31943
rect 17693 31909 17727 31943
rect 18797 31909 18831 31943
rect 19349 31909 19383 31943
rect 20361 31909 20395 31943
rect 21097 31909 21131 31943
rect 22753 31909 22787 31943
rect 23489 31909 23523 31943
rect 3801 31841 3835 31875
rect 8125 31841 8159 31875
rect 12357 31841 12391 31875
rect 16313 31841 16347 31875
rect 19993 31841 20027 31875
rect 20913 31841 20947 31875
rect 1409 31773 1443 31807
rect 1685 31773 1719 31807
rect 2053 31773 2087 31807
rect 2329 31773 2363 31807
rect 2603 31773 2637 31807
rect 4043 31773 4077 31807
rect 5733 31773 5767 31807
rect 5825 31773 5859 31807
rect 6929 31773 6963 31807
rect 7113 31773 7147 31807
rect 7849 31773 7883 31807
rect 7987 31773 8021 31807
rect 9413 31773 9447 31807
rect 9873 31773 9907 31807
rect 12599 31773 12633 31807
rect 14933 31773 14967 31807
rect 15207 31773 15241 31807
rect 16587 31773 16621 31807
rect 17877 31773 17911 31807
rect 18337 31773 18371 31807
rect 18429 31773 18463 31807
rect 18981 31773 19015 31807
rect 19533 31773 19567 31807
rect 19901 31773 19935 31807
rect 20177 31773 20211 31807
rect 20361 31773 20395 31807
rect 20729 31773 20763 31807
rect 20821 31773 20855 31807
rect 21005 31773 21039 31807
rect 21281 31773 21315 31807
rect 22937 31773 22971 31807
rect 23397 31773 23431 31807
rect 23673 31773 23707 31807
rect 23857 31773 23891 31807
rect 24225 31773 24259 31807
rect 5457 31705 5491 31739
rect 6193 31705 6227 31739
rect 6561 31705 6595 31739
rect 9505 31705 9539 31739
rect 3341 31637 3375 31671
rect 9137 31637 9171 31671
rect 10241 31637 10275 31671
rect 13369 31637 13403 31671
rect 15945 31637 15979 31671
rect 17325 31637 17359 31671
rect 3157 31433 3191 31467
rect 4537 31433 4571 31467
rect 4721 31433 4755 31467
rect 8493 31433 8527 31467
rect 10425 31433 10459 31467
rect 18613 31433 18647 31467
rect 19901 31433 19935 31467
rect 23397 31433 23431 31467
rect 1409 31365 1443 31399
rect 2697 31365 2731 31399
rect 3433 31365 3467 31399
rect 2421 31297 2455 31331
rect 2973 31297 3007 31331
rect 3709 31297 3743 31331
rect 3801 31297 3835 31331
rect 4169 31297 4203 31331
rect 5179 31297 5213 31331
rect 7481 31297 7515 31331
rect 7755 31297 7789 31331
rect 9655 31297 9689 31331
rect 11713 31297 11747 31331
rect 13091 31297 13125 31331
rect 14197 31297 14231 31331
rect 14455 31327 14489 31361
rect 17233 31297 17267 31331
rect 17500 31297 17534 31331
rect 19163 31297 19197 31331
rect 20269 31297 20303 31331
rect 20525 31297 20559 31331
rect 23581 31297 23615 31331
rect 23857 31297 23891 31331
rect 23949 31297 23983 31331
rect 2145 31229 2179 31263
rect 4905 31229 4939 31263
rect 9413 31229 9447 31263
rect 12817 31229 12851 31263
rect 18889 31229 18923 31263
rect 11897 31161 11931 31195
rect 5917 31093 5951 31127
rect 9045 31093 9079 31127
rect 13829 31093 13863 31127
rect 15209 31093 15243 31127
rect 21649 31093 21683 31127
rect 23673 31093 23707 31127
rect 24133 31093 24167 31127
rect 7389 30889 7423 30923
rect 17049 30889 17083 30923
rect 19349 30889 19383 30923
rect 19441 30889 19475 30923
rect 23305 30889 23339 30923
rect 15853 30821 15887 30855
rect 18797 30821 18831 30855
rect 23029 30821 23063 30855
rect 1409 30753 1443 30787
rect 3065 30753 3099 30787
rect 6377 30753 6411 30787
rect 10701 30753 10735 30787
rect 16246 30753 16280 30787
rect 16405 30753 16439 30787
rect 19533 30753 19567 30787
rect 19717 30753 19751 30787
rect 21373 30753 21407 30787
rect 1683 30685 1717 30719
rect 2789 30685 2823 30719
rect 4997 30685 5031 30719
rect 6619 30685 6653 30719
rect 10943 30685 10977 30719
rect 12725 30685 12759 30719
rect 15209 30685 15243 30719
rect 15393 30685 15427 30719
rect 16129 30685 16163 30719
rect 17785 30685 17819 30719
rect 18059 30685 18093 30719
rect 19257 30685 19291 30719
rect 19625 30685 19659 30719
rect 19809 30685 19843 30719
rect 21281 30685 21315 30719
rect 21631 30655 21665 30689
rect 22753 30685 22787 30719
rect 22937 30685 22971 30719
rect 23213 30685 23247 30719
rect 23489 30685 23523 30719
rect 23857 30685 23891 30719
rect 4905 30617 4939 30651
rect 5365 30617 5399 30651
rect 5733 30617 5767 30651
rect 12357 30617 12391 30651
rect 12633 30617 12667 30651
rect 13093 30617 13127 30651
rect 24225 30617 24259 30651
rect 2421 30549 2455 30583
rect 4169 30549 4203 30583
rect 4629 30549 4663 30583
rect 5917 30549 5951 30583
rect 11713 30549 11747 30583
rect 13461 30549 13495 30583
rect 13645 30549 13679 30583
rect 21097 30549 21131 30583
rect 22385 30549 22419 30583
rect 22845 30549 22879 30583
rect 4997 30345 5031 30379
rect 14105 30345 14139 30379
rect 15209 30345 15243 30379
rect 22753 30345 22787 30379
rect 3525 30277 3559 30311
rect 13369 30277 13403 30311
rect 14473 30277 14507 30311
rect 1685 30209 1719 30243
rect 2605 30209 2639 30243
rect 2722 30209 2756 30243
rect 3709 30209 3743 30243
rect 4259 30219 4293 30253
rect 5365 30209 5399 30243
rect 5917 30209 5951 30243
rect 7663 30209 7697 30243
rect 10057 30209 10091 30243
rect 10331 30209 10365 30243
rect 11897 30209 11931 30243
rect 12155 30239 12189 30273
rect 14381 30209 14415 30243
rect 14841 30209 14875 30243
rect 21833 30209 21867 30243
rect 22201 30209 22235 30243
rect 22937 30209 22971 30243
rect 23213 30209 23247 30243
rect 23489 30209 23523 30243
rect 23857 30209 23891 30243
rect 23949 30209 23983 30243
rect 1869 30141 1903 30175
rect 2329 30141 2363 30175
rect 2881 30141 2915 30175
rect 3985 30141 4019 30175
rect 5641 30141 5675 30175
rect 7389 30141 7423 30175
rect 22488 30152 22522 30186
rect 6101 30073 6135 30107
rect 12909 30073 12943 30107
rect 23305 30073 23339 30107
rect 3801 30005 3835 30039
rect 8401 30005 8435 30039
rect 11069 30005 11103 30039
rect 13461 30005 13495 30039
rect 15393 30005 15427 30039
rect 21925 30005 21959 30039
rect 22293 30005 22327 30039
rect 22385 30005 22419 30039
rect 23029 30005 23063 30039
rect 23673 30005 23707 30039
rect 24133 30005 24167 30039
rect 2881 29801 2915 29835
rect 23213 29801 23247 29835
rect 5917 29733 5951 29767
rect 16773 29733 16807 29767
rect 19533 29733 19567 29767
rect 1869 29665 1903 29699
rect 3801 29665 3835 29699
rect 1501 29597 1535 29631
rect 2143 29597 2177 29631
rect 3249 29597 3283 29631
rect 4077 29597 4111 29631
rect 4905 29597 4939 29631
rect 5163 29567 5197 29601
rect 7205 29597 7239 29631
rect 8953 29597 8987 29631
rect 9227 29597 9261 29631
rect 10793 29597 10827 29631
rect 10885 29597 10919 29631
rect 15761 29597 15795 29631
rect 16035 29597 16069 29631
rect 17141 29597 17175 29631
rect 17415 29597 17449 29631
rect 19717 29597 19751 29631
rect 20637 29597 20671 29631
rect 23397 29597 23431 29631
rect 23857 29597 23891 29631
rect 23949 29597 23983 29631
rect 6469 29529 6503 29563
rect 6745 29529 6779 29563
rect 6837 29529 6871 29563
rect 7573 29529 7607 29563
rect 10517 29529 10551 29563
rect 11253 29529 11287 29563
rect 1593 29461 1627 29495
rect 3433 29461 3467 29495
rect 7757 29461 7791 29495
rect 9965 29461 9999 29495
rect 11621 29461 11655 29495
rect 11805 29461 11839 29495
rect 18153 29461 18187 29495
rect 20453 29461 20487 29495
rect 23673 29461 23707 29495
rect 24133 29461 24167 29495
rect 7389 29257 7423 29291
rect 10149 29257 10183 29291
rect 20361 29257 20395 29291
rect 20913 29257 20947 29291
rect 23489 29257 23523 29291
rect 14749 29189 14783 29223
rect 19248 29189 19282 29223
rect 23857 29189 23891 29223
rect 2421 29121 2455 29155
rect 3433 29121 3467 29155
rect 3707 29121 3741 29155
rect 6619 29121 6653 29155
rect 8677 29121 8711 29155
rect 8953 29121 8987 29155
rect 9597 29121 9631 29155
rect 10057 29121 10091 29155
rect 10333 29121 10367 29155
rect 10425 29121 10459 29155
rect 10609 29121 10643 29155
rect 10701 29121 10735 29155
rect 12909 29121 12943 29155
rect 16497 29121 16531 29155
rect 16865 29121 16899 29155
rect 17718 29121 17752 29155
rect 17877 29121 17911 29155
rect 18981 29121 19015 29155
rect 20453 29121 20487 29155
rect 20821 29119 20855 29153
rect 21097 29121 21131 29155
rect 21281 29121 21315 29155
rect 23397 29121 23431 29155
rect 23673 29121 23707 29155
rect 1409 29053 1443 29087
rect 1685 29053 1719 29087
rect 6377 29053 6411 29087
rect 7757 29053 7791 29087
rect 7941 29053 7975 29087
rect 8401 29053 8435 29087
rect 8794 29053 8828 29087
rect 13093 29053 13127 29087
rect 13829 29053 13863 29087
rect 13946 29053 13980 29087
rect 14105 29053 14139 29087
rect 16681 29053 16715 29087
rect 17325 29053 17359 29087
rect 17601 29053 17635 29087
rect 20545 29053 20579 29087
rect 20729 29053 20763 29087
rect 21189 29053 21223 29087
rect 2605 28985 2639 29019
rect 9873 28985 9907 29019
rect 13553 28985 13587 29019
rect 18521 28985 18555 29019
rect 23213 28985 23247 29019
rect 24133 28985 24167 29019
rect 4445 28917 4479 28951
rect 10517 28917 10551 28951
rect 10793 28917 10827 28951
rect 20637 28917 20671 28951
rect 10609 28713 10643 28747
rect 13461 28713 13495 28747
rect 14289 28713 14323 28747
rect 20637 28713 20671 28747
rect 3341 28645 3375 28679
rect 12081 28645 12115 28679
rect 18705 28645 18739 28679
rect 23121 28645 23155 28679
rect 23489 28645 23523 28679
rect 2329 28577 2363 28611
rect 9597 28577 9631 28611
rect 2603 28509 2637 28543
rect 4353 28509 4387 28543
rect 5457 28509 5491 28543
rect 5731 28509 5765 28543
rect 9839 28509 9873 28543
rect 11069 28509 11103 28543
rect 11343 28509 11377 28543
rect 12449 28509 12483 28543
rect 12723 28509 12757 28543
rect 14657 28509 14691 28543
rect 14899 28509 14933 28543
rect 17325 28509 17359 28543
rect 18981 28509 19015 28543
rect 19625 28509 19659 28543
rect 19899 28509 19933 28543
rect 22109 28509 22143 28543
rect 22845 28509 22879 28543
rect 23673 28509 23707 28543
rect 23949 28509 23983 28543
rect 1501 28441 1535 28475
rect 1685 28441 1719 28475
rect 4261 28441 4295 28475
rect 4721 28441 4755 28475
rect 17592 28441 17626 28475
rect 3985 28373 4019 28407
rect 5089 28373 5123 28407
rect 5273 28373 5307 28407
rect 6469 28373 6503 28407
rect 15669 28373 15703 28407
rect 18797 28373 18831 28407
rect 22201 28373 22235 28407
rect 22661 28373 22695 28407
rect 24133 28373 24167 28407
rect 3249 28169 3283 28203
rect 3893 28169 3927 28203
rect 6101 28169 6135 28203
rect 9689 28169 9723 28203
rect 14197 28169 14231 28203
rect 17693 28169 17727 28203
rect 21465 28169 21499 28203
rect 4813 28101 4847 28135
rect 5181 28101 5215 28135
rect 5917 28101 5951 28135
rect 10977 28101 11011 28135
rect 11713 28101 11747 28135
rect 12817 28101 12851 28135
rect 16497 28101 16531 28135
rect 2329 28033 2363 28067
rect 2446 28033 2480 28067
rect 3433 28033 3467 28067
rect 3709 28033 3743 28067
rect 5089 28033 5123 28067
rect 5549 28033 5583 28067
rect 8769 28033 8803 28067
rect 9045 28033 9079 28067
rect 10609 28033 10643 28067
rect 11989 28033 12023 28067
rect 12081 28033 12115 28067
rect 12449 28033 12483 28067
rect 13185 28033 13219 28067
rect 13443 28063 13477 28097
rect 14657 28033 14691 28067
rect 15715 28033 15749 28067
rect 17877 28033 17911 28067
rect 18245 28033 18279 28067
rect 18521 28033 18555 28067
rect 18889 28033 18923 28067
rect 19073 28033 19107 28067
rect 21649 28033 21683 28067
rect 22291 28033 22325 28067
rect 23397 28033 23431 28067
rect 23489 28033 23523 28067
rect 23949 28033 23983 28067
rect 1409 27965 1443 27999
rect 1593 27965 1627 27999
rect 2605 27965 2639 27999
rect 7849 27965 7883 27999
rect 8033 27965 8067 27999
rect 8493 27965 8527 27999
rect 8886 27965 8920 27999
rect 10701 27965 10735 27999
rect 14841 27965 14875 27999
rect 15301 27965 15335 27999
rect 15577 27965 15611 27999
rect 15853 27965 15887 27999
rect 18797 27965 18831 27999
rect 18981 27965 19015 27999
rect 22017 27965 22051 27999
rect 23673 27965 23707 27999
rect 2053 27897 2087 27931
rect 13001 27897 13035 27931
rect 3525 27829 3559 27863
rect 10885 27829 10919 27863
rect 18337 27829 18371 27863
rect 18613 27829 18647 27863
rect 18705 27829 18739 27863
rect 23029 27829 23063 27863
rect 23581 27829 23615 27863
rect 24133 27829 24167 27863
rect 2605 27625 2639 27659
rect 16497 27625 16531 27659
rect 18613 27625 18647 27659
rect 3433 27557 3467 27591
rect 6101 27557 6135 27591
rect 11805 27557 11839 27591
rect 22201 27557 22235 27591
rect 22385 27557 22419 27591
rect 22753 27557 22787 27591
rect 22937 27557 22971 27591
rect 5089 27489 5123 27523
rect 7021 27489 7055 27523
rect 10793 27489 10827 27523
rect 17601 27489 17635 27523
rect 1593 27421 1627 27455
rect 1867 27421 1901 27455
rect 2973 27421 3007 27455
rect 3249 27421 3283 27455
rect 3801 27421 3835 27455
rect 5331 27421 5365 27455
rect 7295 27421 7329 27455
rect 11067 27421 11101 27455
rect 14105 27421 14139 27455
rect 14379 27411 14413 27445
rect 15485 27421 15519 27455
rect 15727 27421 15761 27455
rect 17843 27421 17877 27455
rect 20821 27421 20855 27455
rect 21088 27421 21122 27455
rect 22569 27421 22603 27455
rect 22661 27421 22695 27455
rect 22845 27421 22879 27455
rect 23121 27421 23155 27455
rect 23397 27421 23431 27455
rect 23857 27421 23891 27455
rect 23949 27421 23983 27455
rect 3157 27285 3191 27319
rect 3985 27285 4019 27319
rect 8033 27285 8067 27319
rect 15117 27285 15151 27319
rect 23213 27285 23247 27319
rect 23673 27285 23707 27319
rect 24133 27285 24167 27319
rect 2421 27081 2455 27115
rect 3249 27081 3283 27115
rect 3525 27081 3559 27115
rect 7021 27081 7055 27115
rect 7297 27013 7331 27047
rect 7389 27013 7423 27047
rect 8125 27013 8159 27047
rect 1683 26945 1717 26979
rect 2789 26945 2823 26979
rect 3065 26945 3099 26979
rect 3341 26945 3375 26979
rect 3617 26945 3651 26979
rect 3891 26945 3925 26979
rect 7757 26945 7791 26979
rect 9011 26945 9045 26979
rect 12539 26945 12573 26979
rect 19255 26945 19289 26979
rect 20361 26945 20395 26979
rect 20545 26945 20579 26979
rect 20913 26945 20947 26979
rect 23305 26945 23339 26979
rect 23857 26945 23891 26979
rect 23949 26945 23983 26979
rect 1409 26877 1443 26911
rect 8769 26877 8803 26911
rect 12265 26877 12299 26911
rect 18981 26877 19015 26911
rect 23121 26809 23155 26843
rect 23673 26809 23707 26843
rect 2973 26741 3007 26775
rect 4629 26741 4663 26775
rect 8309 26741 8343 26775
rect 9781 26741 9815 26775
rect 13277 26741 13311 26775
rect 19993 26741 20027 26775
rect 20453 26741 20487 26775
rect 20729 26741 20763 26775
rect 24133 26741 24167 26775
rect 1869 26537 1903 26571
rect 7113 26537 7147 26571
rect 10425 26537 10459 26571
rect 1593 26469 1627 26503
rect 3157 26469 3191 26503
rect 4445 26469 4479 26503
rect 8493 26469 8527 26503
rect 10701 26469 10735 26503
rect 11069 26469 11103 26503
rect 21649 26469 21683 26503
rect 21741 26469 21775 26503
rect 2145 26401 2179 26435
rect 3801 26401 3835 26435
rect 4721 26401 4755 26435
rect 4859 26401 4893 26435
rect 6101 26401 6135 26435
rect 7481 26401 7515 26435
rect 10885 26401 10919 26435
rect 11345 26401 11379 26435
rect 14565 26401 14599 26435
rect 16221 26401 16255 26435
rect 16681 26401 16715 26435
rect 19533 26401 19567 26435
rect 19901 26401 19935 26435
rect 20085 26401 20119 26435
rect 20269 26401 20303 26435
rect 1409 26333 1443 26367
rect 1685 26333 1719 26367
rect 2419 26333 2453 26367
rect 3985 26333 4019 26367
rect 4997 26333 5031 26367
rect 6343 26333 6377 26367
rect 7723 26333 7757 26367
rect 9873 26333 9907 26367
rect 10609 26333 10643 26367
rect 10977 26333 11011 26367
rect 11253 26333 11287 26367
rect 11437 26333 11471 26367
rect 11897 26333 11931 26367
rect 12171 26333 12205 26367
rect 14823 26303 14857 26337
rect 16037 26333 16071 26367
rect 16975 26333 17009 26367
rect 17074 26333 17108 26367
rect 17233 26333 17267 26367
rect 17877 26333 17911 26367
rect 18981 26333 19015 26367
rect 19441 26333 19475 26367
rect 19809 26333 19843 26367
rect 20536 26333 20570 26367
rect 21925 26333 21959 26367
rect 23857 26333 23891 26367
rect 5641 26265 5675 26299
rect 9137 26265 9171 26299
rect 9413 26265 9447 26299
rect 9505 26265 9539 26299
rect 10241 26265 10275 26299
rect 20085 26265 20119 26299
rect 24225 26265 24259 26299
rect 10885 26197 10919 26231
rect 12909 26197 12943 26231
rect 15577 26197 15611 26231
rect 18797 26197 18831 26231
rect 2973 25993 3007 26027
rect 4169 25993 4203 26027
rect 10701 25993 10735 26027
rect 11069 25993 11103 26027
rect 17693 25993 17727 26027
rect 19717 25993 19751 26027
rect 19901 25993 19935 26027
rect 18582 25925 18616 25959
rect 1683 25857 1717 25891
rect 2789 25857 2823 25891
rect 3399 25857 3433 25891
rect 5163 25887 5197 25921
rect 9963 25857 9997 25891
rect 11253 25857 11287 25891
rect 11529 25857 11563 25891
rect 11803 25857 11837 25891
rect 13921 25857 13955 25891
rect 14195 25857 14229 25891
rect 16923 25857 16957 25891
rect 18337 25857 18371 25891
rect 20085 25857 20119 25891
rect 20603 25857 20637 25891
rect 21833 25857 21867 25891
rect 22201 25857 22235 25891
rect 22385 25857 22419 25891
rect 22845 25857 22879 25891
rect 23305 25857 23339 25891
rect 23489 25857 23523 25891
rect 23581 25857 23615 25891
rect 23949 25857 23983 25891
rect 1409 25789 1443 25823
rect 3157 25789 3191 25823
rect 4905 25789 4939 25823
rect 9689 25789 9723 25823
rect 16681 25789 16715 25823
rect 20361 25789 20395 25823
rect 22109 25789 22143 25823
rect 22293 25789 22327 25823
rect 21373 25721 21407 25755
rect 22017 25721 22051 25755
rect 2421 25653 2455 25687
rect 5917 25653 5951 25687
rect 12541 25653 12575 25687
rect 14933 25653 14967 25687
rect 21925 25653 21959 25687
rect 22661 25653 22695 25687
rect 23397 25653 23431 25687
rect 23765 25653 23799 25687
rect 24133 25653 24167 25687
rect 10793 25449 10827 25483
rect 13369 25449 13403 25483
rect 17049 25449 17083 25483
rect 21373 25449 21407 25483
rect 12173 25381 12207 25415
rect 14749 25381 14783 25415
rect 23765 25381 23799 25415
rect 24133 25381 24167 25415
rect 11529 25313 11563 25347
rect 12449 25313 12483 25347
rect 12566 25313 12600 25347
rect 12725 25313 12759 25347
rect 14289 25313 14323 25347
rect 15301 25313 15335 25347
rect 16037 25313 16071 25347
rect 23949 25313 23983 25347
rect 3065 25245 3099 25279
rect 5641 25245 5675 25279
rect 5915 25245 5949 25279
rect 10977 25245 11011 25279
rect 11713 25245 11747 25279
rect 14105 25245 14139 25279
rect 15025 25245 15059 25279
rect 15142 25245 15176 25279
rect 16279 25245 16313 25279
rect 21281 25245 21315 25279
rect 22109 25245 22143 25279
rect 23673 25245 23707 25279
rect 24041 25245 24075 25279
rect 1593 25177 1627 25211
rect 1869 25177 1903 25211
rect 1961 25177 1995 25211
rect 2329 25177 2363 25211
rect 2697 25177 2731 25211
rect 22354 25177 22388 25211
rect 2881 25109 2915 25143
rect 3249 25109 3283 25143
rect 6653 25109 6687 25143
rect 15945 25109 15979 25143
rect 23489 25109 23523 25143
rect 23949 25109 23983 25143
rect 2697 24905 2731 24939
rect 7665 24905 7699 24939
rect 23673 24905 23707 24939
rect 24041 24905 24075 24939
rect 6561 24837 6595 24871
rect 7297 24837 7331 24871
rect 1409 24769 1443 24803
rect 1927 24769 1961 24803
rect 4075 24769 4109 24803
rect 6837 24769 6871 24803
rect 6929 24769 6963 24803
rect 8033 24769 8067 24803
rect 8307 24769 8341 24803
rect 9871 24769 9905 24803
rect 12539 24769 12573 24803
rect 13645 24769 13679 24803
rect 14682 24769 14716 24803
rect 14841 24769 14875 24803
rect 17141 24769 17175 24803
rect 17408 24769 17442 24803
rect 18613 24769 18647 24803
rect 19073 24769 19107 24803
rect 19165 24769 19199 24803
rect 19349 24769 19383 24803
rect 19625 24769 19659 24803
rect 20085 24769 20119 24803
rect 22935 24769 22969 24803
rect 24225 24769 24259 24803
rect 1685 24701 1719 24735
rect 3801 24701 3835 24735
rect 9597 24701 9631 24735
rect 12265 24701 12299 24735
rect 13829 24701 13863 24735
rect 14565 24701 14599 24735
rect 22661 24701 22695 24735
rect 1593 24633 1627 24667
rect 7849 24633 7883 24667
rect 13277 24633 13311 24667
rect 14289 24633 14323 24667
rect 18521 24633 18555 24667
rect 19441 24633 19475 24667
rect 4813 24565 4847 24599
rect 9045 24565 9079 24599
rect 10609 24565 10643 24599
rect 15485 24565 15519 24599
rect 18705 24565 18739 24599
rect 18889 24565 18923 24599
rect 19257 24565 19291 24599
rect 20177 24565 20211 24599
rect 6101 24361 6135 24395
rect 10977 24361 11011 24395
rect 17325 24361 17359 24395
rect 18613 24361 18647 24395
rect 20821 24361 20855 24395
rect 23765 24361 23799 24395
rect 2789 24293 2823 24327
rect 4905 24293 4939 24327
rect 21373 24293 21407 24327
rect 1409 24225 1443 24259
rect 1685 24225 1719 24259
rect 4261 24225 4295 24259
rect 5319 24225 5353 24259
rect 9321 24225 9355 24259
rect 9781 24225 9815 24259
rect 10057 24225 10091 24259
rect 10195 24225 10229 24259
rect 11805 24225 11839 24259
rect 12449 24225 12483 24259
rect 12842 24225 12876 24259
rect 13001 24225 13035 24259
rect 17601 24225 17635 24259
rect 21005 24225 21039 24259
rect 21189 24225 21223 24259
rect 2329 24157 2363 24191
rect 2605 24157 2639 24191
rect 4445 24157 4479 24191
rect 5181 24157 5215 24191
rect 5457 24157 5491 24191
rect 7573 24157 7607 24191
rect 9137 24157 9171 24191
rect 10333 24157 10367 24191
rect 11989 24157 12023 24191
rect 12725 24157 12759 24191
rect 13645 24157 13679 24191
rect 17509 24157 17543 24191
rect 17859 24127 17893 24161
rect 19257 24157 19291 24191
rect 19524 24157 19558 24191
rect 20729 24157 20763 24191
rect 21097 24157 21131 24191
rect 21281 24157 21315 24191
rect 21557 24157 21591 24191
rect 22753 24157 22787 24191
rect 23489 24157 23523 24191
rect 23949 24157 23983 24191
rect 7481 24089 7515 24123
rect 7941 24089 7975 24123
rect 2513 24021 2547 24055
rect 7205 24021 7239 24055
rect 8309 24021 8343 24055
rect 8493 24021 8527 24055
rect 20637 24021 20671 24055
rect 21005 24021 21039 24055
rect 22569 24021 22603 24055
rect 24133 24021 24167 24055
rect 1593 23817 1627 23851
rect 1869 23817 1903 23851
rect 10977 23817 11011 23851
rect 12633 23817 12667 23851
rect 20453 23817 20487 23851
rect 2605 23749 2639 23783
rect 3709 23749 3743 23783
rect 22262 23749 22296 23783
rect 23857 23749 23891 23783
rect 1409 23681 1443 23715
rect 1685 23681 1719 23715
rect 1961 23681 1995 23715
rect 2881 23681 2915 23715
rect 2973 23681 3007 23715
rect 3341 23681 3375 23715
rect 4687 23681 4721 23715
rect 6619 23681 6653 23715
rect 7757 23681 7791 23715
rect 8015 23681 8049 23715
rect 9137 23681 9171 23715
rect 11621 23681 11655 23715
rect 11895 23681 11929 23715
rect 15483 23681 15517 23715
rect 16681 23681 16715 23715
rect 16865 23681 16899 23715
rect 17718 23681 17752 23715
rect 18613 23681 18647 23715
rect 18705 23681 18739 23715
rect 19683 23681 19717 23715
rect 21373 23681 21407 23715
rect 22017 23681 22051 23715
rect 23673 23681 23707 23715
rect 4445 23613 4479 23647
rect 6377 23613 6411 23647
rect 9321 23613 9355 23647
rect 10057 23613 10091 23647
rect 10195 23613 10229 23647
rect 10333 23613 10367 23647
rect 15209 23613 15243 23647
rect 17601 23613 17635 23647
rect 17877 23613 17911 23647
rect 18889 23613 18923 23647
rect 19441 23613 19475 23647
rect 2145 23545 2179 23579
rect 7389 23545 7423 23579
rect 8769 23545 8803 23579
rect 9761 23545 9795 23579
rect 16221 23545 16255 23579
rect 17325 23545 17359 23579
rect 23397 23545 23431 23579
rect 3893 23477 3927 23511
rect 5457 23477 5491 23511
rect 18521 23477 18555 23511
rect 18797 23477 18831 23511
rect 21465 23477 21499 23511
rect 23489 23477 23523 23511
rect 24133 23477 24167 23511
rect 1961 23273 1995 23307
rect 3341 23273 3375 23307
rect 17141 23273 17175 23307
rect 20729 23273 20763 23307
rect 2329 23137 2363 23171
rect 16129 23137 16163 23171
rect 21005 23137 21039 23171
rect 22569 23137 22603 23171
rect 24225 23137 24259 23171
rect 2603 23069 2637 23103
rect 14473 23069 14507 23103
rect 14747 23069 14781 23103
rect 16403 23069 16437 23103
rect 20913 23069 20947 23103
rect 21279 23069 21313 23103
rect 22811 23069 22845 23103
rect 23949 23069 23983 23103
rect 24041 23069 24075 23103
rect 1501 23001 1535 23035
rect 1685 23001 1719 23035
rect 1869 23001 1903 23035
rect 15485 22933 15519 22967
rect 22017 22933 22051 22967
rect 23581 22933 23615 22967
rect 24225 22933 24259 22967
rect 2973 22729 3007 22763
rect 5917 22729 5951 22763
rect 23121 22729 23155 22763
rect 2881 22661 2915 22695
rect 1683 22593 1717 22627
rect 3341 22593 3375 22627
rect 3583 22593 3617 22627
rect 5163 22593 5197 22627
rect 6561 22593 6595 22627
rect 6745 22593 6779 22627
rect 7598 22593 7632 22627
rect 8401 22593 8435 22627
rect 8861 22593 8895 22627
rect 10055 22593 10089 22627
rect 12449 22593 12483 22627
rect 12707 22623 12741 22657
rect 14866 22593 14900 22627
rect 15669 22593 15703 22627
rect 16865 22593 16899 22627
rect 18153 22593 18187 22627
rect 18420 22593 18454 22627
rect 19809 22593 19843 22627
rect 20276 22593 20310 22627
rect 20525 22593 20559 22627
rect 21833 22593 21867 22627
rect 21925 22593 21959 22627
rect 22385 22593 22419 22627
rect 22477 22593 22511 22627
rect 22661 22593 22695 22627
rect 22937 22593 22971 22627
rect 23121 22593 23155 22627
rect 23213 22593 23247 22627
rect 23305 22593 23339 22627
rect 23581 22593 23615 22627
rect 23949 22593 23983 22627
rect 1409 22525 1443 22559
rect 4905 22525 4939 22559
rect 7481 22525 7515 22559
rect 7757 22525 7791 22559
rect 9781 22525 9815 22559
rect 13829 22525 13863 22559
rect 14013 22525 14047 22559
rect 14749 22525 14783 22559
rect 15025 22525 15059 22559
rect 22109 22525 22143 22559
rect 22569 22525 22603 22559
rect 7205 22457 7239 22491
rect 13461 22457 13495 22491
rect 14473 22457 14507 22491
rect 19533 22457 19567 22491
rect 21649 22457 21683 22491
rect 22201 22457 22235 22491
rect 2421 22389 2455 22423
rect 4353 22389 4387 22423
rect 8677 22389 8711 22423
rect 10793 22389 10827 22423
rect 16681 22389 16715 22423
rect 19625 22389 19659 22423
rect 22017 22389 22051 22423
rect 23765 22389 23799 22423
rect 24133 22389 24167 22423
rect 11529 22185 11563 22219
rect 13277 22117 13311 22151
rect 14749 22117 14783 22151
rect 2145 22049 2179 22083
rect 2421 22049 2455 22083
rect 2559 22049 2593 22083
rect 2697 22049 2731 22083
rect 7481 22049 7515 22083
rect 14105 22049 14139 22083
rect 14289 22049 14323 22083
rect 15142 22049 15176 22083
rect 15301 22049 15335 22083
rect 15945 22049 15979 22083
rect 19257 22049 19291 22083
rect 1501 21981 1535 22015
rect 1685 21981 1719 22015
rect 3985 21981 4019 22015
rect 4243 21951 4277 21985
rect 5457 21981 5491 22015
rect 5731 21981 5765 22015
rect 6837 21981 6871 22015
rect 7021 21981 7055 22015
rect 7757 21981 7791 22015
rect 7895 21981 7929 22015
rect 8033 21981 8067 22015
rect 8677 21981 8711 22015
rect 9229 21981 9263 22015
rect 9413 21981 9447 22015
rect 9597 21981 9631 22015
rect 10977 21981 11011 22015
rect 12265 21981 12299 22015
rect 15025 21981 15059 22015
rect 17233 21981 17267 22015
rect 17509 21981 17543 22015
rect 17601 21981 17635 22015
rect 17969 21981 18003 22015
rect 18153 21981 18187 22015
rect 18337 21981 18371 22015
rect 18797 21981 18831 22015
rect 18889 21981 18923 22015
rect 19515 21951 19549 21985
rect 20637 21981 20671 22015
rect 20821 21981 20855 22015
rect 21189 21981 21223 22015
rect 23949 21981 23983 22015
rect 10517 21913 10551 21947
rect 10609 21913 10643 21947
rect 11345 21913 11379 21947
rect 12357 21913 12391 21947
rect 12725 21913 12759 21947
rect 3341 21845 3375 21879
rect 4997 21845 5031 21879
rect 6469 21845 6503 21879
rect 9045 21845 9079 21879
rect 9597 21845 9631 21879
rect 10241 21845 10275 21879
rect 11989 21845 12023 21879
rect 13093 21845 13127 21879
rect 17785 21845 17819 21879
rect 18337 21845 18371 21879
rect 18613 21845 18647 21879
rect 18981 21845 19015 21879
rect 20269 21845 20303 21879
rect 20729 21845 20763 21879
rect 21373 21845 21407 21879
rect 24133 21845 24167 21879
rect 2421 21641 2455 21675
rect 8033 21641 8067 21675
rect 11069 21641 11103 21675
rect 13093 21641 13127 21675
rect 19073 21641 19107 21675
rect 22753 21641 22787 21675
rect 5641 21573 5675 21607
rect 1683 21505 1717 21539
rect 2789 21505 2823 21539
rect 3065 21505 3099 21539
rect 4997 21505 5031 21539
rect 7295 21505 7329 21539
rect 8951 21505 8985 21539
rect 10331 21505 10365 21539
rect 12081 21505 12115 21539
rect 12355 21505 12389 21539
rect 15209 21505 15243 21539
rect 15483 21505 15517 21539
rect 16681 21505 16715 21539
rect 16923 21505 16957 21539
rect 18335 21505 18369 21539
rect 19625 21505 19659 21539
rect 19717 21505 19751 21539
rect 22937 21505 22971 21539
rect 23397 21505 23431 21539
rect 23857 21505 23891 21539
rect 23949 21505 23983 21539
rect 1409 21437 1443 21471
rect 3801 21437 3835 21471
rect 3985 21437 4019 21471
rect 4721 21437 4755 21471
rect 4859 21437 4893 21471
rect 7021 21437 7055 21471
rect 8677 21437 8711 21471
rect 10057 21437 10091 21471
rect 18061 21437 18095 21471
rect 19901 21437 19935 21471
rect 4445 21369 4479 21403
rect 23673 21369 23707 21403
rect 2973 21301 3007 21335
rect 3249 21301 3283 21335
rect 9689 21301 9723 21335
rect 16221 21301 16255 21335
rect 17693 21301 17727 21335
rect 19809 21301 19843 21335
rect 23489 21301 23523 21335
rect 24133 21301 24167 21335
rect 3525 21097 3559 21131
rect 8033 21097 8067 21131
rect 12449 21097 12483 21131
rect 18153 21097 18187 21131
rect 23581 21097 23615 21131
rect 5733 21029 5767 21063
rect 6929 21029 6963 21063
rect 16773 21029 16807 21063
rect 5273 20961 5307 20995
rect 6009 20961 6043 20995
rect 6285 20961 6319 20995
rect 9229 20961 9263 20995
rect 11437 20961 11471 20995
rect 16313 20961 16347 20995
rect 17049 20961 17083 20995
rect 17325 20961 17359 20995
rect 18337 20961 18371 20995
rect 1501 20893 1535 20927
rect 1777 20893 1811 20927
rect 2973 20893 3007 20927
rect 5089 20893 5123 20927
rect 6147 20893 6181 20927
rect 7021 20893 7055 20927
rect 7295 20893 7329 20927
rect 9137 20893 9171 20927
rect 9413 20893 9447 20927
rect 9597 20893 9631 20927
rect 9965 20893 9999 20927
rect 11679 20893 11713 20927
rect 16129 20893 16163 20927
rect 17187 20893 17221 20927
rect 18061 20893 18095 20927
rect 20085 20893 20119 20927
rect 22201 20893 22235 20927
rect 23857 20893 23891 20927
rect 2513 20825 2547 20859
rect 2605 20825 2639 20859
rect 3341 20825 3375 20859
rect 9873 20825 9907 20859
rect 20330 20825 20364 20859
rect 22446 20825 22480 20859
rect 24225 20825 24259 20859
rect 1593 20757 1627 20791
rect 1961 20757 1995 20791
rect 2237 20757 2271 20791
rect 17969 20757 18003 20791
rect 18337 20757 18371 20791
rect 21465 20757 21499 20791
rect 1593 20553 1627 20587
rect 1961 20553 1995 20587
rect 2329 20553 2363 20587
rect 3709 20553 3743 20587
rect 20637 20553 20671 20587
rect 21833 20553 21867 20587
rect 13001 20485 13035 20519
rect 14105 20485 14139 20519
rect 1501 20417 1535 20451
rect 1869 20417 1903 20451
rect 2237 20417 2271 20451
rect 2697 20417 2731 20451
rect 2955 20447 2989 20481
rect 4353 20417 4387 20451
rect 7847 20417 7881 20451
rect 12357 20417 12391 20451
rect 13277 20417 13311 20451
rect 13369 20417 13403 20451
rect 13737 20417 13771 20451
rect 14473 20417 14507 20451
rect 14715 20427 14749 20461
rect 19717 20417 19751 20451
rect 20361 20417 20395 20451
rect 20821 20417 20855 20451
rect 21189 20417 21223 20451
rect 22017 20417 22051 20451
rect 22109 20417 22143 20451
rect 22293 20417 22327 20451
rect 23087 20417 23121 20451
rect 4077 20349 4111 20383
rect 7573 20349 7607 20383
rect 22845 20349 22879 20383
rect 8585 20213 8619 20247
rect 11897 20213 11931 20247
rect 12541 20213 12575 20247
rect 14289 20213 14323 20247
rect 15485 20213 15519 20247
rect 16037 20213 16071 20247
rect 19809 20213 19843 20247
rect 20177 20213 20211 20247
rect 21281 20213 21315 20247
rect 22201 20213 22235 20247
rect 23857 20213 23891 20247
rect 2973 20009 3007 20043
rect 3525 20009 3559 20043
rect 8677 20009 8711 20043
rect 13645 20009 13679 20043
rect 18889 20009 18923 20043
rect 20637 20009 20671 20043
rect 23765 20009 23799 20043
rect 24041 20009 24075 20043
rect 1685 19941 1719 19975
rect 10333 19941 10367 19975
rect 15301 19941 15335 19975
rect 21741 19941 21775 19975
rect 23213 19941 23247 19975
rect 1961 19873 1995 19907
rect 12633 19873 12667 19907
rect 14657 19873 14691 19907
rect 14841 19873 14875 19907
rect 15577 19873 15611 19907
rect 19257 19873 19291 19907
rect 20729 19873 20763 19907
rect 22385 19873 22419 19907
rect 24225 19873 24259 19907
rect 1501 19805 1535 19839
rect 2203 19805 2237 19839
rect 3341 19805 3375 19839
rect 5825 19805 5859 19839
rect 6083 19775 6117 19809
rect 7665 19805 7699 19839
rect 7757 19805 7791 19839
rect 9321 19805 9355 19839
rect 9579 19805 9613 19839
rect 11161 19805 11195 19839
rect 11621 19805 11655 19839
rect 12875 19805 12909 19839
rect 15694 19805 15728 19839
rect 15853 19805 15887 19839
rect 19073 19805 19107 19839
rect 19513 19805 19547 19839
rect 20971 19805 21005 19839
rect 22109 19805 22143 19839
rect 22201 19805 22235 19839
rect 23121 19805 23155 19839
rect 23305 19805 23339 19839
rect 23489 19805 23523 19839
rect 23949 19805 23983 19839
rect 7389 19737 7423 19771
rect 8125 19737 8159 19771
rect 8493 19737 8527 19771
rect 11253 19737 11287 19771
rect 11989 19737 12023 19771
rect 22385 19737 22419 19771
rect 6837 19669 6871 19703
rect 10885 19669 10919 19703
rect 12173 19669 12207 19703
rect 16497 19669 16531 19703
rect 24225 19669 24259 19703
rect 7941 19465 7975 19499
rect 13461 19465 13495 19499
rect 15945 19465 15979 19499
rect 23213 19465 23247 19499
rect 23673 19397 23707 19431
rect 1683 19329 1717 19363
rect 2789 19329 2823 19363
rect 3523 19329 3557 19363
rect 4905 19329 4939 19363
rect 5179 19329 5213 19363
rect 6929 19329 6963 19363
rect 7171 19329 7205 19363
rect 8677 19329 8711 19363
rect 8951 19329 8985 19363
rect 12449 19329 12483 19363
rect 12707 19359 12741 19393
rect 14933 19329 14967 19363
rect 15207 19329 15241 19363
rect 16681 19329 16715 19363
rect 17601 19329 17635 19363
rect 18855 19329 18889 19363
rect 20235 19329 20269 19363
rect 21833 19329 21867 19363
rect 22100 19329 22134 19363
rect 23489 19329 23523 19363
rect 1409 19261 1443 19295
rect 3249 19261 3283 19295
rect 10241 19261 10275 19295
rect 16865 19261 16899 19295
rect 17718 19261 17752 19295
rect 17877 19261 17911 19295
rect 18613 19261 18647 19295
rect 19993 19261 20027 19295
rect 2973 19193 3007 19227
rect 17325 19193 17359 19227
rect 2421 19125 2455 19159
rect 4261 19125 4295 19159
rect 5917 19125 5951 19159
rect 9689 19125 9723 19159
rect 18521 19125 18555 19159
rect 19625 19125 19659 19159
rect 21005 19125 21039 19159
rect 23305 19125 23339 19159
rect 23949 19125 23983 19159
rect 1593 18921 1627 18955
rect 11897 18921 11931 18955
rect 18429 18921 18463 18955
rect 20269 18921 20303 18955
rect 2329 18853 2363 18887
rect 6009 18853 6043 18887
rect 18153 18853 18187 18887
rect 18797 18853 18831 18887
rect 19349 18853 19383 18887
rect 2722 18785 2756 18819
rect 3801 18785 3835 18819
rect 5365 18785 5399 18819
rect 6402 18785 6436 18819
rect 6561 18785 6595 18819
rect 18981 18785 19015 18819
rect 19625 18785 19659 18819
rect 20453 18785 20487 18819
rect 20637 18785 20671 18819
rect 22477 18785 22511 18819
rect 24133 18785 24167 18819
rect 1409 18717 1443 18751
rect 1685 18717 1719 18751
rect 1869 18717 1903 18751
rect 2605 18717 2639 18751
rect 2881 18717 2915 18751
rect 4075 18717 4109 18751
rect 5549 18717 5583 18751
rect 6285 18717 6319 18751
rect 9413 18717 9447 18751
rect 9505 18717 9539 18751
rect 9919 18717 9953 18751
rect 10885 18717 10919 18751
rect 11159 18717 11193 18751
rect 18337 18717 18371 18751
rect 18613 18717 18647 18751
rect 18705 18717 18739 18751
rect 19257 18717 19291 18751
rect 19533 18717 19567 18751
rect 19717 18717 19751 18751
rect 20177 18717 20211 18751
rect 20545 18717 20579 18751
rect 20729 18717 20763 18751
rect 22385 18717 22419 18751
rect 22719 18717 22753 18751
rect 23857 18717 23891 18751
rect 23949 18717 23983 18751
rect 10241 18649 10275 18683
rect 3525 18581 3559 18615
rect 4813 18581 4847 18615
rect 7205 18581 7239 18615
rect 9137 18581 9171 18615
rect 10425 18581 10459 18615
rect 18981 18581 19015 18615
rect 20453 18581 20487 18615
rect 22201 18581 22235 18615
rect 23489 18581 23523 18615
rect 24133 18581 24167 18615
rect 2697 18377 2731 18411
rect 10425 18377 10459 18411
rect 18521 18377 18555 18411
rect 22753 18377 22787 18411
rect 23029 18377 23063 18411
rect 24133 18377 24167 18411
rect 1409 18241 1443 18275
rect 1959 18241 1993 18275
rect 3157 18241 3191 18275
rect 3617 18241 3651 18275
rect 3801 18241 3835 18275
rect 4813 18241 4847 18275
rect 9687 18241 9721 18275
rect 11989 18241 12023 18275
rect 12263 18251 12297 18285
rect 13553 18241 13587 18275
rect 14406 18241 14440 18275
rect 14565 18241 14599 18275
rect 16681 18241 16715 18275
rect 16865 18241 16899 18275
rect 17877 18241 17911 18275
rect 20913 18241 20947 18275
rect 22661 18241 22695 18275
rect 22845 18241 22879 18275
rect 22937 18241 22971 18275
rect 23305 18241 23339 18275
rect 23857 18241 23891 18275
rect 1685 18173 1719 18207
rect 4261 18173 4295 18207
rect 4537 18173 4571 18207
rect 4675 18173 4709 18207
rect 9413 18173 9447 18207
rect 13369 18173 13403 18207
rect 14289 18173 14323 18207
rect 17325 18173 17359 18207
rect 17601 18173 17635 18207
rect 17718 18173 17752 18207
rect 13001 18105 13035 18139
rect 14013 18105 14047 18139
rect 1593 18037 1627 18071
rect 3249 18037 3283 18071
rect 5457 18037 5491 18071
rect 11897 18037 11931 18071
rect 15209 18037 15243 18071
rect 20729 18037 20763 18071
rect 23581 18037 23615 18071
rect 15117 17833 15151 17867
rect 17693 17833 17727 17867
rect 24133 17833 24167 17867
rect 2973 17765 3007 17799
rect 10885 17765 10919 17799
rect 23765 17765 23799 17799
rect 11897 17697 11931 17731
rect 12173 17697 12207 17731
rect 16681 17697 16715 17731
rect 1409 17629 1443 17663
rect 1683 17629 1717 17663
rect 2789 17629 2823 17663
rect 3249 17629 3283 17663
rect 4629 17629 4663 17663
rect 4813 17629 4847 17663
rect 7205 17629 7239 17663
rect 7479 17629 7513 17663
rect 9873 17629 9907 17663
rect 10115 17629 10149 17663
rect 11253 17629 11287 17663
rect 11437 17629 11471 17663
rect 12290 17629 12324 17663
rect 12449 17629 12483 17663
rect 14105 17629 14139 17663
rect 14379 17629 14413 17663
rect 15761 17629 15795 17663
rect 16955 17629 16989 17663
rect 19533 17629 19567 17663
rect 20453 17629 20487 17663
rect 22017 17629 22051 17663
rect 23581 17629 23615 17663
rect 23949 17629 23983 17663
rect 4077 17561 4111 17595
rect 13093 17561 13127 17595
rect 20698 17561 20732 17595
rect 22284 17561 22318 17595
rect 2421 17493 2455 17527
rect 3341 17493 3375 17527
rect 4169 17493 4203 17527
rect 8217 17493 8251 17527
rect 19349 17493 19383 17527
rect 21833 17493 21867 17527
rect 23397 17493 23431 17527
rect 7941 17289 7975 17323
rect 12541 17289 12575 17323
rect 17693 17289 17727 17323
rect 22569 17289 22603 17323
rect 9045 17221 9079 17255
rect 19156 17221 19190 17255
rect 24041 17221 24075 17255
rect 1501 17153 1535 17187
rect 1961 17153 1995 17187
rect 2235 17153 2269 17187
rect 3615 17153 3649 17187
rect 5163 17183 5197 17217
rect 6377 17153 6411 17187
rect 6635 17183 6669 17217
rect 8217 17153 8251 17187
rect 8309 17153 8343 17187
rect 8677 17153 8711 17187
rect 9747 17153 9781 17187
rect 11771 17153 11805 17187
rect 14841 17153 14875 17187
rect 15577 17153 15611 17187
rect 16923 17153 16957 17187
rect 20603 17153 20637 17187
rect 22017 17153 22051 17187
rect 22293 17153 22327 17187
rect 22753 17153 22787 17187
rect 23029 17153 23063 17187
rect 23305 17153 23339 17187
rect 23765 17153 23799 17187
rect 3341 17085 3375 17119
rect 4905 17085 4939 17119
rect 9505 17085 9539 17119
rect 11529 17085 11563 17119
rect 14657 17085 14691 17119
rect 15694 17085 15728 17119
rect 15853 17085 15887 17119
rect 16681 17085 16715 17119
rect 18889 17085 18923 17119
rect 20361 17085 20395 17119
rect 24041 17085 24075 17119
rect 15301 17017 15335 17051
rect 23857 17017 23891 17051
rect 1593 16949 1627 16983
rect 2973 16949 3007 16983
rect 4353 16949 4387 16983
rect 5917 16949 5951 16983
rect 7389 16949 7423 16983
rect 9229 16949 9263 16983
rect 10517 16949 10551 16983
rect 16497 16949 16531 16983
rect 20269 16949 20303 16983
rect 21373 16949 21407 16983
rect 21833 16949 21867 16983
rect 22385 16949 22419 16983
rect 22845 16949 22879 16983
rect 23581 16949 23615 16983
rect 15393 16745 15427 16779
rect 18705 16745 18739 16779
rect 21833 16745 21867 16779
rect 22201 16745 22235 16779
rect 23673 16745 23707 16779
rect 24133 16745 24167 16779
rect 2237 16677 2271 16711
rect 4905 16677 4939 16711
rect 6837 16677 6871 16711
rect 11161 16677 11195 16711
rect 18613 16677 18647 16711
rect 18981 16677 19015 16711
rect 19625 16677 19659 16711
rect 1593 16609 1627 16643
rect 2513 16609 2547 16643
rect 2630 16609 2664 16643
rect 3433 16609 3467 16643
rect 5181 16609 5215 16643
rect 5319 16609 5353 16643
rect 5457 16609 5491 16643
rect 6193 16609 6227 16643
rect 6377 16609 6411 16643
rect 7230 16609 7264 16643
rect 10149 16609 10183 16643
rect 11897 16609 11931 16643
rect 16957 16609 16991 16643
rect 18797 16609 18831 16643
rect 20085 16609 20119 16643
rect 20453 16609 20487 16643
rect 20637 16609 20671 16643
rect 21097 16609 21131 16643
rect 22017 16609 22051 16643
rect 22477 16609 22511 16643
rect 1777 16541 1811 16575
rect 2789 16541 2823 16575
rect 3801 16541 3835 16575
rect 4261 16541 4295 16575
rect 4445 16541 4479 16575
rect 7113 16541 7147 16575
rect 7387 16541 7421 16575
rect 10391 16541 10425 16575
rect 12171 16541 12205 16575
rect 13645 16541 13679 16575
rect 14381 16541 14415 16575
rect 14655 16541 14689 16575
rect 17213 16541 17247 16575
rect 18521 16541 18555 16575
rect 18889 16541 18923 16575
rect 19441 16541 19475 16575
rect 19533 16541 19567 16575
rect 19717 16541 19751 16575
rect 19993 16541 20027 16575
rect 20361 16541 20395 16575
rect 20913 16541 20947 16575
rect 21005 16541 21039 16575
rect 21189 16541 21223 16575
rect 21741 16541 21775 16575
rect 22109 16541 22143 16575
rect 22385 16541 22419 16575
rect 22569 16541 22603 16575
rect 22661 16541 22695 16575
rect 22919 16511 22953 16545
rect 24041 16541 24075 16575
rect 24225 16541 24259 16575
rect 20637 16473 20671 16507
rect 3985 16405 4019 16439
rect 6101 16405 6135 16439
rect 8033 16405 8067 16439
rect 12909 16405 12943 16439
rect 18337 16405 18371 16439
rect 19257 16405 19291 16439
rect 20729 16405 20763 16439
rect 22017 16405 22051 16439
rect 2697 16201 2731 16235
rect 7665 16201 7699 16235
rect 9045 16201 9079 16235
rect 12081 16201 12115 16235
rect 16129 16201 16163 16235
rect 17417 16201 17451 16235
rect 18797 16201 18831 16235
rect 22845 16201 22879 16235
rect 24133 16201 24167 16235
rect 1943 16095 1977 16129
rect 3433 16065 3467 16099
rect 4169 16065 4203 16099
rect 4445 16065 4479 16099
rect 6653 16065 6687 16099
rect 6927 16065 6961 16099
rect 8033 16065 8067 16099
rect 8307 16065 8341 16099
rect 9505 16065 9539 16099
rect 12633 16065 12667 16099
rect 13369 16065 13403 16099
rect 13645 16065 13679 16099
rect 15391 16065 15425 16099
rect 17601 16065 17635 16099
rect 18027 16065 18061 16099
rect 22075 16065 22109 16099
rect 23581 16065 23615 16099
rect 23949 16065 23983 16099
rect 1685 15997 1719 16031
rect 3249 15997 3283 16031
rect 3893 15997 3927 16031
rect 4307 15997 4341 16031
rect 9689 15997 9723 16031
rect 10149 15997 10183 16031
rect 10425 15997 10459 16031
rect 10563 15997 10597 16031
rect 10701 15997 10735 16031
rect 12449 15997 12483 16031
rect 13093 15997 13127 16031
rect 13507 15997 13541 16031
rect 15117 15997 15151 16031
rect 17785 15997 17819 16031
rect 21833 15997 21867 16031
rect 5089 15861 5123 15895
rect 11345 15861 11379 15895
rect 14289 15861 14323 15895
rect 23765 15861 23799 15895
rect 2145 15657 2179 15691
rect 3249 15657 3283 15691
rect 3985 15657 4019 15691
rect 5549 15657 5583 15691
rect 13645 15657 13679 15691
rect 12633 15521 12667 15555
rect 1685 15453 1719 15487
rect 2053 15453 2087 15487
rect 3157 15453 3191 15487
rect 4537 15453 4571 15487
rect 4811 15453 4845 15487
rect 9689 15453 9723 15487
rect 12907 15453 12941 15487
rect 14565 15453 14599 15487
rect 14839 15453 14873 15487
rect 17693 15453 17727 15487
rect 19809 15453 19843 15487
rect 23857 15453 23891 15487
rect 2605 15385 2639 15419
rect 3893 15385 3927 15419
rect 24225 15385 24259 15419
rect 2697 15317 2731 15351
rect 15577 15317 15611 15351
rect 17509 15317 17543 15351
rect 19625 15317 19659 15351
rect 3157 15113 3191 15147
rect 3709 15113 3743 15147
rect 10333 15113 10367 15147
rect 20913 15113 20947 15147
rect 1651 14977 1685 15011
rect 3065 14977 3099 15011
rect 3617 14977 3651 15011
rect 4887 15007 4921 15041
rect 7387 14977 7421 15011
rect 8493 14977 8527 15011
rect 9413 14977 9447 15011
rect 14289 14977 14323 15011
rect 15485 14977 15519 15011
rect 17213 14977 17247 15011
rect 18705 14977 18739 15011
rect 18889 14977 18923 15011
rect 19432 14977 19466 15011
rect 20637 14977 20671 15011
rect 21189 14977 21223 15011
rect 22293 14977 22327 15011
rect 22560 14977 22594 15011
rect 23949 14977 23983 15011
rect 1409 14909 1443 14943
rect 4629 14909 4663 14943
rect 7113 14909 7147 14943
rect 8677 14909 8711 14943
rect 9530 14909 9564 14943
rect 9689 14909 9723 14943
rect 14473 14909 14507 14943
rect 15209 14909 15243 14943
rect 15347 14909 15381 14943
rect 16957 14909 16991 14943
rect 19165 14909 19199 14943
rect 20913 14909 20947 14943
rect 8125 14841 8159 14875
rect 9137 14841 9171 14875
rect 14933 14841 14967 14875
rect 20545 14841 20579 14875
rect 20729 14841 20763 14875
rect 2421 14773 2455 14807
rect 5641 14773 5675 14807
rect 16129 14773 16163 14807
rect 18337 14773 18371 14807
rect 18797 14773 18831 14807
rect 21005 14773 21039 14807
rect 23673 14773 23707 14807
rect 24133 14773 24167 14807
rect 1593 14569 1627 14603
rect 3065 14569 3099 14603
rect 3985 14569 4019 14603
rect 9965 14569 9999 14603
rect 15117 14569 15151 14603
rect 18705 14569 18739 14603
rect 20637 14569 20671 14603
rect 21097 14569 21131 14603
rect 21373 14569 21407 14603
rect 22569 14501 22603 14535
rect 22845 14501 22879 14535
rect 4537 14433 4571 14467
rect 4997 14433 5031 14467
rect 5273 14433 5307 14467
rect 5549 14433 5583 14467
rect 7389 14433 7423 14467
rect 8953 14433 8987 14467
rect 12081 14433 12115 14467
rect 19533 14433 19567 14467
rect 24041 14433 24075 14467
rect 2605 14365 2639 14399
rect 2973 14365 3007 14399
rect 4353 14365 4387 14399
rect 5411 14365 5445 14399
rect 7663 14365 7697 14399
rect 9195 14365 9229 14399
rect 11897 14365 11931 14399
rect 12323 14365 12357 14399
rect 14105 14365 14139 14399
rect 14347 14365 14381 14399
rect 17693 14365 17727 14399
rect 17967 14355 18001 14389
rect 19257 14365 19291 14399
rect 19349 14365 19383 14399
rect 19625 14365 19659 14399
rect 19899 14365 19933 14399
rect 21005 14365 21039 14399
rect 21281 14365 21315 14399
rect 21465 14365 21499 14399
rect 22293 14365 22327 14399
rect 22477 14365 22511 14399
rect 22753 14365 22787 14399
rect 23029 14365 23063 14399
rect 23765 14365 23799 14399
rect 23857 14365 23891 14399
rect 1501 14297 1535 14331
rect 3893 14297 3927 14331
rect 19533 14297 19567 14331
rect 22385 14297 22419 14331
rect 23305 14297 23339 14331
rect 24041 14297 24075 14331
rect 6193 14229 6227 14263
rect 8401 14229 8435 14263
rect 13093 14229 13127 14263
rect 23581 14229 23615 14263
rect 8953 14025 8987 14059
rect 13645 14025 13679 14059
rect 18153 14025 18187 14059
rect 18613 14025 18647 14059
rect 22385 14025 22419 14059
rect 22753 14025 22787 14059
rect 23949 14025 23983 14059
rect 14749 13957 14783 13991
rect 2421 13889 2455 13923
rect 2559 13889 2593 13923
rect 3691 13919 3725 13953
rect 4905 13889 4939 13923
rect 5179 13889 5213 13923
rect 7297 13889 7331 13923
rect 8309 13889 8343 13923
rect 10315 13919 10349 13953
rect 11529 13889 11563 13923
rect 12449 13889 12483 13923
rect 12725 13889 12759 13923
rect 13369 13889 13403 13923
rect 13921 13889 13955 13923
rect 14013 13889 14047 13923
rect 14381 13889 14415 13923
rect 15451 13889 15485 13923
rect 16923 13889 16957 13923
rect 18061 13889 18095 13923
rect 18797 13889 18831 13923
rect 21557 13889 21591 13923
rect 22109 13889 22143 13923
rect 22293 13889 22327 13923
rect 22569 13889 22603 13923
rect 22685 13879 22719 13913
rect 22937 13889 22971 13923
rect 23195 13919 23229 13953
rect 1501 13821 1535 13855
rect 1685 13821 1719 13855
rect 2145 13821 2179 13855
rect 2697 13821 2731 13855
rect 3433 13821 3467 13855
rect 7113 13821 7147 13855
rect 8033 13821 8067 13855
rect 8171 13821 8205 13855
rect 10057 13821 10091 13855
rect 11713 13821 11747 13855
rect 12173 13821 12207 13855
rect 12587 13821 12621 13855
rect 15209 13821 15243 13855
rect 16681 13821 16715 13855
rect 7757 13753 7791 13787
rect 11069 13753 11103 13787
rect 3341 13685 3375 13719
rect 4445 13685 4479 13719
rect 5917 13685 5951 13719
rect 14933 13685 14967 13719
rect 16221 13685 16255 13719
rect 17693 13685 17727 13719
rect 21373 13685 21407 13719
rect 22201 13685 22235 13719
rect 2513 13481 2547 13515
rect 5089 13481 5123 13515
rect 7665 13481 7699 13515
rect 11989 13481 12023 13515
rect 13645 13481 13679 13515
rect 22201 13481 22235 13515
rect 24133 13481 24167 13515
rect 6469 13413 6503 13447
rect 16129 13413 16163 13447
rect 4077 13345 4111 13379
rect 6862 13345 6896 13379
rect 8953 13345 8987 13379
rect 12633 13345 12667 13379
rect 15669 13345 15703 13379
rect 16405 13345 16439 13379
rect 16522 13345 16556 13379
rect 16681 13345 16715 13379
rect 1501 13277 1535 13311
rect 1775 13277 1809 13311
rect 4335 13247 4369 13281
rect 5825 13277 5859 13311
rect 6009 13277 6043 13311
rect 6745 13277 6779 13311
rect 7021 13277 7055 13311
rect 9227 13277 9261 13311
rect 10517 13277 10551 13311
rect 10977 13277 11011 13311
rect 11251 13277 11285 13311
rect 12907 13277 12941 13311
rect 15485 13277 15519 13311
rect 20821 13277 20855 13311
rect 22293 13277 22327 13311
rect 22535 13267 22569 13301
rect 23949 13277 23983 13311
rect 21088 13209 21122 13243
rect 9965 13141 9999 13175
rect 17325 13141 17359 13175
rect 23305 13141 23339 13175
rect 2329 12937 2363 12971
rect 4813 12937 4847 12971
rect 7849 12937 7883 12971
rect 22753 12937 22787 12971
rect 23397 12937 23431 12971
rect 1685 12869 1719 12903
rect 2237 12869 2271 12903
rect 4721 12869 4755 12903
rect 9505 12869 9539 12903
rect 9781 12869 9815 12903
rect 10609 12869 10643 12903
rect 19901 12869 19935 12903
rect 23673 12869 23707 12903
rect 2697 12801 2731 12835
rect 2881 12801 2915 12835
rect 3734 12801 3768 12835
rect 6837 12801 6871 12835
rect 7111 12801 7145 12835
rect 9873 12801 9907 12835
rect 10241 12801 10275 12835
rect 11771 12801 11805 12835
rect 14807 12801 14841 12835
rect 17323 12801 17357 12835
rect 19625 12801 19659 12835
rect 19993 12801 20027 12835
rect 20361 12801 20395 12835
rect 20603 12801 20637 12835
rect 22017 12801 22051 12835
rect 22477 12801 22511 12835
rect 22937 12801 22971 12835
rect 23213 12801 23247 12835
rect 3617 12733 3651 12767
rect 3893 12733 3927 12767
rect 11529 12733 11563 12767
rect 14565 12733 14599 12767
rect 17049 12733 17083 12767
rect 19809 12733 19843 12767
rect 22753 12733 22787 12767
rect 3341 12665 3375 12699
rect 1777 12597 1811 12631
rect 4537 12597 4571 12631
rect 10793 12597 10827 12631
rect 12541 12597 12575 12631
rect 15577 12597 15611 12631
rect 18061 12597 18095 12631
rect 21373 12597 21407 12631
rect 22109 12597 22143 12631
rect 22569 12597 22603 12631
rect 23029 12597 23063 12631
rect 23949 12597 23983 12631
rect 1593 12393 1627 12427
rect 3341 12393 3375 12427
rect 4721 12393 4755 12427
rect 10609 12393 10643 12427
rect 13921 12393 13955 12427
rect 18981 12393 19015 12427
rect 20269 12393 20303 12427
rect 20729 12393 20763 12427
rect 17969 12325 18003 12359
rect 23397 12325 23431 12359
rect 9597 12257 9631 12291
rect 12081 12257 12115 12291
rect 12265 12257 12299 12291
rect 12725 12257 12759 12291
rect 13001 12257 13035 12291
rect 19257 12257 19291 12291
rect 22201 12257 22235 12291
rect 1501 12189 1535 12223
rect 2329 12189 2363 12223
rect 2603 12189 2637 12223
rect 5457 12189 5491 12223
rect 5715 12159 5749 12193
rect 9871 12189 9905 12223
rect 13118 12189 13152 12223
rect 13277 12189 13311 12223
rect 14749 12189 14783 12223
rect 17969 12189 18003 12223
rect 18153 12189 18187 12223
rect 18429 12189 18463 12223
rect 18613 12189 18647 12223
rect 18889 12189 18923 12223
rect 19531 12189 19565 12223
rect 20637 12189 20671 12223
rect 20821 12189 20855 12223
rect 21465 12189 21499 12223
rect 21833 12189 21867 12223
rect 22109 12189 22143 12223
rect 23213 12189 23247 12223
rect 23673 12189 23707 12223
rect 4077 12121 4111 12155
rect 4629 12121 4663 12155
rect 14657 12121 14691 12155
rect 15117 12121 15151 12155
rect 18337 12121 18371 12155
rect 18521 12121 18555 12155
rect 24041 12121 24075 12155
rect 4169 12053 4203 12087
rect 6469 12053 6503 12087
rect 14381 12053 14415 12087
rect 15485 12053 15519 12087
rect 15669 12053 15703 12087
rect 7389 11849 7423 11883
rect 9689 11849 9723 11883
rect 13461 11849 13495 11883
rect 14933 11849 14967 11883
rect 20637 11849 20671 11883
rect 22017 11849 22051 11883
rect 1685 11713 1719 11747
rect 2421 11713 2455 11747
rect 2538 11713 2572 11747
rect 4813 11713 4847 11747
rect 6377 11713 6411 11747
rect 6635 11743 6669 11777
rect 7849 11713 7883 11747
rect 9045 11713 9079 11747
rect 12723 11713 12757 11747
rect 14179 11743 14213 11777
rect 17325 11713 17359 11747
rect 17417 11713 17451 11747
rect 17673 11713 17707 11747
rect 19073 11713 19107 11747
rect 19165 11713 19199 11747
rect 19432 11713 19466 11747
rect 20821 11713 20855 11747
rect 21833 11713 21867 11747
rect 22017 11711 22051 11745
rect 22385 11713 22419 11747
rect 23087 11713 23121 11747
rect 1501 11645 1535 11679
rect 2697 11645 2731 11679
rect 3617 11645 3651 11679
rect 3801 11645 3835 11679
rect 4537 11645 4571 11679
rect 4675 11645 4709 11679
rect 8033 11645 8067 11679
rect 8769 11645 8803 11679
rect 8907 11645 8941 11679
rect 12449 11645 12483 11679
rect 13921 11645 13955 11679
rect 22845 11645 22879 11679
rect 2145 11577 2179 11611
rect 4261 11577 4295 11611
rect 8493 11577 8527 11611
rect 18797 11577 18831 11611
rect 18889 11577 18923 11611
rect 20545 11577 20579 11611
rect 22201 11577 22235 11611
rect 3341 11509 3375 11543
rect 5457 11509 5491 11543
rect 17141 11509 17175 11543
rect 23857 11509 23891 11543
rect 2697 11305 2731 11339
rect 3341 11305 3375 11339
rect 4537 11305 4571 11339
rect 6929 11305 6963 11339
rect 8493 11305 8527 11339
rect 9965 11305 9999 11339
rect 12265 11305 12299 11339
rect 18061 11305 18095 11339
rect 19533 11305 19567 11339
rect 22569 11305 22603 11339
rect 5733 11169 5767 11203
rect 6009 11169 6043 11203
rect 6126 11169 6160 11203
rect 6285 11169 6319 11203
rect 7481 11169 7515 11203
rect 8953 11169 8987 11203
rect 10609 11169 10643 11203
rect 11069 11169 11103 11203
rect 11483 11169 11517 11203
rect 15853 11169 15887 11203
rect 16313 11169 16347 11203
rect 16706 11169 16740 11203
rect 19809 11169 19843 11203
rect 22753 11169 22787 11203
rect 1685 11101 1719 11135
rect 1959 11101 1993 11135
rect 3893 11101 3927 11135
rect 4445 11101 4479 11135
rect 5089 11101 5123 11135
rect 5273 11101 5307 11135
rect 7755 11101 7789 11135
rect 9195 11101 9229 11135
rect 10425 11101 10459 11135
rect 11345 11101 11379 11135
rect 11621 11101 11655 11135
rect 15669 11101 15703 11135
rect 16589 11101 16623 11135
rect 16865 11101 16899 11135
rect 17969 11101 18003 11135
rect 19717 11101 19751 11135
rect 20051 11101 20085 11135
rect 21189 11101 21223 11135
rect 23027 11101 23061 11135
rect 3249 11033 3283 11067
rect 17509 11033 17543 11067
rect 21456 11033 21490 11067
rect 3985 10965 4019 10999
rect 20821 10965 20855 10999
rect 23765 10965 23799 10999
rect 1593 10761 1627 10795
rect 2973 10761 3007 10795
rect 4353 10761 4387 10795
rect 5733 10761 5767 10795
rect 11069 10761 11103 10795
rect 12541 10761 12575 10795
rect 16221 10761 16255 10795
rect 17693 10761 17727 10795
rect 21925 10761 21959 10795
rect 1501 10625 1535 10659
rect 1961 10625 1995 10659
rect 2235 10625 2269 10659
rect 3341 10625 3375 10659
rect 3599 10655 3633 10689
rect 4721 10625 4755 10659
rect 4995 10625 5029 10659
rect 10057 10625 10091 10659
rect 10331 10625 10365 10659
rect 11771 10625 11805 10659
rect 13461 10625 13495 10659
rect 13735 10625 13769 10659
rect 15451 10625 15485 10659
rect 16681 10625 16715 10659
rect 16955 10625 16989 10659
rect 21833 10625 21867 10659
rect 22293 10625 22327 10659
rect 22661 10625 22695 10659
rect 22935 10625 22969 10659
rect 24225 10625 24259 10659
rect 11529 10557 11563 10591
rect 15209 10557 15243 10591
rect 22109 10489 22143 10523
rect 14473 10421 14507 10455
rect 23673 10421 23707 10455
rect 24041 10421 24075 10455
rect 2421 10217 2455 10251
rect 2973 10217 3007 10251
rect 5089 10217 5123 10251
rect 5641 10217 5675 10251
rect 8769 10217 8803 10251
rect 22569 10217 22603 10251
rect 24133 10217 24167 10251
rect 7573 10149 7607 10183
rect 13461 10149 13495 10183
rect 18705 10149 18739 10183
rect 20913 10149 20947 10183
rect 22293 10149 22327 10183
rect 4169 10081 4203 10115
rect 6929 10081 6963 10115
rect 7113 10081 7147 10115
rect 7849 10081 7883 10115
rect 8125 10081 8159 10115
rect 14289 10081 14323 10115
rect 14749 10081 14783 10115
rect 20821 10081 20855 10115
rect 1409 10013 1443 10047
rect 1683 10013 1717 10047
rect 4445 10013 4479 10047
rect 5549 10013 5583 10047
rect 7987 10013 8021 10047
rect 8953 10013 8987 10047
rect 9211 9983 9245 10017
rect 12909 10013 12943 10047
rect 14105 10013 14139 10047
rect 15025 10013 15059 10047
rect 15163 10013 15197 10047
rect 15301 10013 15335 10047
rect 18061 10013 18095 10047
rect 18245 10013 18279 10047
rect 18705 10013 18739 10047
rect 19809 10013 19843 10047
rect 19993 10013 20027 10047
rect 20913 10013 20947 10047
rect 22477 10013 22511 10047
rect 22753 10013 22787 10047
rect 22845 10013 22879 10047
rect 23857 10013 23891 10047
rect 2881 9945 2915 9979
rect 3893 9945 3927 9979
rect 4997 9945 5031 9979
rect 12173 9945 12207 9979
rect 12449 9945 12483 9979
rect 12541 9945 12575 9979
rect 21281 9945 21315 9979
rect 23305 9945 23339 9979
rect 23673 9945 23707 9979
rect 4537 9877 4571 9911
rect 9965 9877 9999 9911
rect 13281 9877 13315 9911
rect 15945 9877 15979 9911
rect 19993 9877 20027 9911
rect 23029 9877 23063 9911
rect 1777 9673 1811 9707
rect 8309 9673 8343 9707
rect 10793 9673 10827 9707
rect 13369 9673 13403 9707
rect 15117 9673 15151 9707
rect 21281 9673 21315 9707
rect 21557 9673 21591 9707
rect 9505 9605 9539 9639
rect 9873 9605 9907 9639
rect 10609 9605 10643 9639
rect 1685 9537 1719 9571
rect 2605 9537 2639 9571
rect 3617 9537 3651 9571
rect 4445 9537 4479 9571
rect 5179 9537 5213 9571
rect 7297 9537 7331 9571
rect 7571 9537 7605 9571
rect 9781 9537 9815 9571
rect 10241 9537 10275 9571
rect 12631 9537 12665 9571
rect 14105 9537 14139 9571
rect 14379 9537 14413 9571
rect 17323 9537 17357 9571
rect 18871 9567 18905 9601
rect 20361 9537 20395 9571
rect 20821 9537 20855 9571
rect 21189 9537 21223 9571
rect 21465 9537 21499 9571
rect 21649 9537 21683 9571
rect 22017 9537 22051 9571
rect 23087 9537 23121 9571
rect 2421 9469 2455 9503
rect 3341 9469 3375 9503
rect 3479 9469 3513 9503
rect 4905 9469 4939 9503
rect 12357 9469 12391 9503
rect 17049 9469 17083 9503
rect 18613 9469 18647 9503
rect 20085 9469 20119 9503
rect 22845 9469 22879 9503
rect 3065 9401 3099 9435
rect 4721 9401 4755 9435
rect 19625 9401 19659 9435
rect 20821 9401 20855 9435
rect 21833 9401 21867 9435
rect 4261 9333 4295 9367
rect 5917 9333 5951 9367
rect 18061 9333 18095 9367
rect 23857 9333 23891 9367
rect 2881 9129 2915 9163
rect 8493 9129 8527 9163
rect 10609 9129 10643 9163
rect 12449 9129 12483 9163
rect 22109 9129 22143 9163
rect 24133 9129 24167 9163
rect 6193 9061 6227 9095
rect 17509 9061 17543 9095
rect 7389 8993 7423 9027
rect 11437 8993 11471 9027
rect 15853 8993 15887 9027
rect 16313 8993 16347 9027
rect 16589 8993 16623 9027
rect 16727 8993 16761 9027
rect 23121 8993 23155 9027
rect 1869 8925 1903 8959
rect 2143 8925 2177 8959
rect 4169 8925 4203 8959
rect 4443 8925 4477 8959
rect 5549 8925 5583 8959
rect 5733 8925 5767 8959
rect 6469 8925 6503 8959
rect 6586 8925 6620 8959
rect 6745 8925 6779 8959
rect 7481 8925 7515 8959
rect 7755 8925 7789 8959
rect 9597 8925 9631 8959
rect 9871 8925 9905 8959
rect 11711 8925 11745 8959
rect 15669 8925 15703 8959
rect 16865 8925 16899 8959
rect 17601 8925 17635 8959
rect 19257 8925 19291 8959
rect 20729 8925 20763 8959
rect 22293 8925 22327 8959
rect 22569 8925 22603 8959
rect 23029 8925 23063 8959
rect 23581 8925 23615 8959
rect 23857 8925 23891 8959
rect 23949 8925 23983 8959
rect 17868 8857 17902 8891
rect 19524 8857 19558 8891
rect 20996 8857 21030 8891
rect 5181 8789 5215 8823
rect 18981 8789 19015 8823
rect 20637 8789 20671 8823
rect 23397 8789 23431 8823
rect 23673 8789 23707 8823
rect 5733 8585 5767 8619
rect 7389 8585 7423 8619
rect 17693 8585 17727 8619
rect 18153 8585 18187 8619
rect 18429 8585 18463 8619
rect 19625 8585 19659 8619
rect 20177 8585 20211 8619
rect 20821 8585 20855 8619
rect 23765 8585 23799 8619
rect 24041 8585 24075 8619
rect 22560 8517 22594 8551
rect 1685 8449 1719 8483
rect 2421 8449 2455 8483
rect 2697 8449 2731 8483
rect 3893 8449 3927 8483
rect 4077 8449 4111 8483
rect 5089 8449 5123 8483
rect 6635 8479 6669 8513
rect 8307 8449 8341 8483
rect 15483 8449 15517 8483
rect 16955 8449 16989 8483
rect 18061 8449 18095 8483
rect 18337 8449 18371 8483
rect 18521 8449 18555 8483
rect 18797 8449 18831 8483
rect 19073 8449 19107 8483
rect 19533 8449 19567 8483
rect 19993 8449 20027 8483
rect 20361 8449 20395 8483
rect 21005 8449 21039 8483
rect 22017 8447 22051 8481
rect 23949 8449 23983 8483
rect 24225 8449 24259 8483
rect 1501 8381 1535 8415
rect 2559 8381 2593 8415
rect 4813 8381 4847 8415
rect 4951 8381 4985 8415
rect 6377 8381 6411 8415
rect 8033 8381 8067 8415
rect 15209 8381 15243 8415
rect 16681 8381 16715 8415
rect 22109 8381 22143 8415
rect 22293 8381 22327 8415
rect 2145 8313 2179 8347
rect 4537 8313 4571 8347
rect 18613 8313 18647 8347
rect 18889 8313 18923 8347
rect 19809 8313 19843 8347
rect 23673 8313 23707 8347
rect 3341 8245 3375 8279
rect 3617 8245 3651 8279
rect 9045 8245 9079 8279
rect 16221 8245 16255 8279
rect 1961 8041 1995 8075
rect 3341 8041 3375 8075
rect 4813 8041 4847 8075
rect 5917 8041 5951 8075
rect 13829 8041 13863 8075
rect 22845 8041 22879 8075
rect 23213 8041 23247 8075
rect 24225 8041 24259 8075
rect 22477 7973 22511 8007
rect 23581 7973 23615 8007
rect 2329 7905 2363 7939
rect 3801 7905 3835 7939
rect 10977 7905 11011 7939
rect 2603 7837 2637 7871
rect 4075 7837 4109 7871
rect 5825 7837 5859 7871
rect 7297 7837 7331 7871
rect 7571 7837 7605 7871
rect 9137 7837 9171 7871
rect 9411 7837 9445 7871
rect 11219 7837 11253 7871
rect 12909 7837 12943 7871
rect 14841 7837 14875 7871
rect 15115 7837 15149 7871
rect 21465 7837 21499 7871
rect 21707 7837 21741 7871
rect 23029 7837 23063 7871
rect 23121 7837 23155 7871
rect 23305 7837 23339 7871
rect 23397 7837 23431 7871
rect 23857 7837 23891 7871
rect 24041 7837 24075 7871
rect 1869 7769 1903 7803
rect 5273 7769 5307 7803
rect 12817 7769 12851 7803
rect 13277 7769 13311 7803
rect 13645 7769 13679 7803
rect 5365 7701 5399 7735
rect 8309 7701 8343 7735
rect 10149 7701 10183 7735
rect 11989 7701 12023 7735
rect 12541 7701 12575 7735
rect 15853 7701 15887 7735
rect 23673 7701 23707 7735
rect 2513 7497 2547 7531
rect 5825 7497 5859 7531
rect 16313 7497 16347 7531
rect 23949 7497 23983 7531
rect 24225 7497 24259 7531
rect 4629 7429 4663 7463
rect 9873 7429 9907 7463
rect 10977 7429 11011 7463
rect 11713 7429 11747 7463
rect 12081 7429 12115 7463
rect 12449 7429 12483 7463
rect 12817 7429 12851 7463
rect 1501 7361 1535 7395
rect 1775 7361 1809 7395
rect 3415 7371 3449 7405
rect 5181 7361 5215 7395
rect 5733 7361 5767 7395
rect 7757 7361 7791 7395
rect 8677 7361 8711 7395
rect 8953 7361 8987 7395
rect 10149 7361 10183 7395
rect 10241 7361 10275 7395
rect 10609 7361 10643 7395
rect 11989 7361 12023 7395
rect 14657 7361 14691 7395
rect 15669 7361 15703 7395
rect 17417 7361 17451 7395
rect 17969 7361 18003 7395
rect 19809 7361 19843 7395
rect 20083 7361 20117 7395
rect 23305 7365 23339 7399
rect 23673 7361 23707 7395
rect 23765 7361 23799 7395
rect 24041 7361 24075 7395
rect 3157 7293 3191 7327
rect 7941 7293 7975 7327
rect 8401 7293 8435 7327
rect 8815 7293 8849 7327
rect 14473 7293 14507 7327
rect 15393 7293 15427 7327
rect 15531 7293 15565 7327
rect 17233 7293 17267 7327
rect 11161 7225 11195 7259
rect 15117 7225 15151 7259
rect 17877 7225 17911 7259
rect 23489 7225 23523 7259
rect 4169 7157 4203 7191
rect 4721 7157 4755 7191
rect 5273 7157 5307 7191
rect 9597 7157 9631 7191
rect 13001 7157 13035 7191
rect 20821 7157 20855 7191
rect 23121 7157 23155 7191
rect 1593 6953 1627 6987
rect 7481 6953 7515 6987
rect 10885 6953 10919 6987
rect 12265 6953 12299 6987
rect 13645 6953 13679 6987
rect 15209 6953 15243 6987
rect 16497 6953 16531 6987
rect 18429 6885 18463 6919
rect 21465 6885 21499 6919
rect 23765 6885 23799 6919
rect 5641 6817 5675 6851
rect 5825 6817 5859 6851
rect 6285 6817 6319 6851
rect 6678 6817 6712 6851
rect 6837 6817 6871 6851
rect 11253 6817 11287 6851
rect 14197 6817 14231 6851
rect 20821 6817 20855 6851
rect 21925 6817 21959 6851
rect 2329 6749 2363 6783
rect 2571 6749 2605 6783
rect 4261 6749 4295 6783
rect 4535 6749 4569 6783
rect 6561 6749 6595 6783
rect 9873 6749 9907 6783
rect 10147 6749 10181 6783
rect 11511 6719 11545 6753
rect 12633 6749 12667 6783
rect 12907 6749 12941 6783
rect 14455 6719 14489 6753
rect 16405 6749 16439 6783
rect 16865 6749 16899 6783
rect 16957 6749 16991 6783
rect 18613 6749 18647 6783
rect 19257 6749 19291 6783
rect 20545 6749 20579 6783
rect 21005 6749 21039 6783
rect 21557 6749 21591 6783
rect 21833 6749 21867 6783
rect 22017 6749 22051 6783
rect 22293 6749 22327 6783
rect 22569 6749 22603 6783
rect 23121 6749 23155 6783
rect 23489 6749 23523 6783
rect 23857 6749 23891 6783
rect 1501 6681 1535 6715
rect 17224 6681 17258 6715
rect 3341 6613 3375 6647
rect 5273 6613 5307 6647
rect 16681 6613 16715 6647
rect 18337 6613 18371 6647
rect 19349 6613 19383 6647
rect 20361 6613 20395 6647
rect 22109 6613 22143 6647
rect 22753 6613 22787 6647
rect 2421 6409 2455 6443
rect 5917 6409 5951 6443
rect 14197 6409 14231 6443
rect 17693 6409 17727 6443
rect 18153 6409 18187 6443
rect 18337 6409 18371 6443
rect 20361 6409 20395 6443
rect 21005 6409 21039 6443
rect 21833 6409 21867 6443
rect 23121 6409 23155 6443
rect 23581 6409 23615 6443
rect 23857 6409 23891 6443
rect 24225 6409 24259 6443
rect 18880 6341 18914 6375
rect 1683 6273 1717 6307
rect 2973 6273 3007 6307
rect 3826 6273 3860 6307
rect 5179 6273 5213 6307
rect 6911 6303 6945 6337
rect 8307 6273 8341 6307
rect 13459 6273 13493 6307
rect 16923 6273 16957 6307
rect 18061 6273 18095 6307
rect 18245 6273 18279 6307
rect 18521 6273 18555 6307
rect 20085 6273 20119 6307
rect 20269 6273 20303 6307
rect 20545 6273 20579 6307
rect 20913 6273 20947 6307
rect 21189 6273 21223 6307
rect 21373 6273 21407 6307
rect 21465 6273 21499 6307
rect 22017 6273 22051 6307
rect 22109 6273 22143 6307
rect 22383 6273 22417 6307
rect 23489 6273 23523 6307
rect 23765 6273 23799 6307
rect 23949 6273 23983 6307
rect 24041 6273 24075 6307
rect 1409 6205 1443 6239
rect 2789 6205 2823 6239
rect 3433 6205 3467 6239
rect 3709 6205 3743 6239
rect 3985 6205 4019 6239
rect 4905 6205 4939 6239
rect 6653 6205 6687 6239
rect 8033 6205 8067 6239
rect 13185 6205 13219 6239
rect 16681 6205 16715 6239
rect 18613 6205 18647 6239
rect 19993 6137 20027 6171
rect 21281 6137 21315 6171
rect 4629 6069 4663 6103
rect 7665 6069 7699 6103
rect 9045 6069 9079 6103
rect 20177 6069 20211 6103
rect 21649 6069 21683 6103
rect 3341 5865 3375 5899
rect 7389 5865 7423 5899
rect 22201 5865 22235 5899
rect 24225 5865 24259 5899
rect 20085 5797 20119 5831
rect 22477 5797 22511 5831
rect 22569 5797 22603 5831
rect 1685 5729 1719 5763
rect 2145 5729 2179 5763
rect 2421 5729 2455 5763
rect 2559 5729 2593 5763
rect 4629 5729 4663 5763
rect 5089 5729 5123 5763
rect 5482 5729 5516 5763
rect 5641 5729 5675 5763
rect 14657 5729 14691 5763
rect 15117 5729 15151 5763
rect 15393 5729 15427 5763
rect 15510 5729 15544 5763
rect 15669 5729 15703 5763
rect 17785 5729 17819 5763
rect 20821 5729 20855 5763
rect 22845 5729 22879 5763
rect 1501 5661 1535 5695
rect 2697 5661 2731 5695
rect 3433 5661 3467 5695
rect 4077 5661 4111 5695
rect 4445 5661 4479 5695
rect 5365 5661 5399 5695
rect 6377 5661 6411 5695
rect 6651 5661 6685 5695
rect 9965 5661 9999 5695
rect 10239 5661 10273 5695
rect 14473 5661 14507 5695
rect 18027 5661 18061 5695
rect 19441 5661 19475 5695
rect 19625 5661 19659 5695
rect 20177 5661 20211 5695
rect 20545 5661 20579 5695
rect 20729 5661 20763 5695
rect 22293 5661 22327 5695
rect 22753 5661 22787 5695
rect 21088 5593 21122 5627
rect 23112 5593 23146 5627
rect 3617 5525 3651 5559
rect 6285 5525 6319 5559
rect 10977 5525 11011 5559
rect 16313 5525 16347 5559
rect 18797 5525 18831 5559
rect 20729 5525 20763 5559
rect 2421 5321 2455 5355
rect 3249 5321 3283 5355
rect 3801 5321 3835 5355
rect 5181 5321 5215 5355
rect 9781 5321 9815 5355
rect 15761 5321 15795 5355
rect 20453 5321 20487 5355
rect 21097 5321 21131 5355
rect 21649 5321 21683 5355
rect 3157 5253 3191 5287
rect 10517 5253 10551 5287
rect 10885 5253 10919 5287
rect 23857 5253 23891 5287
rect 1409 5185 1443 5219
rect 1667 5215 1701 5249
rect 2789 5185 2823 5219
rect 3709 5185 3743 5219
rect 4169 5185 4203 5219
rect 4443 5185 4477 5219
rect 7665 5185 7699 5219
rect 8585 5185 8619 5219
rect 8861 5185 8895 5219
rect 9505 5185 9539 5219
rect 10057 5185 10091 5219
rect 10149 5185 10183 5219
rect 12817 5185 12851 5219
rect 14013 5185 14047 5219
rect 14749 5185 14783 5219
rect 15023 5185 15057 5219
rect 19349 5185 19383 5219
rect 19436 5185 19470 5219
rect 19683 5195 19717 5229
rect 20913 5185 20947 5219
rect 21373 5185 21407 5219
rect 21465 5185 21499 5219
rect 21649 5185 21683 5219
rect 21833 5185 21867 5219
rect 22201 5185 22235 5219
rect 22661 5185 22695 5219
rect 23029 5185 23063 5219
rect 7849 5117 7883 5151
rect 8309 5117 8343 5151
rect 8723 5117 8757 5151
rect 13001 5117 13035 5151
rect 13737 5117 13771 5151
rect 13875 5117 13909 5151
rect 13461 5049 13495 5083
rect 22661 5049 22695 5083
rect 2973 4981 3007 5015
rect 11069 4981 11103 5015
rect 14657 4981 14691 5015
rect 19165 4981 19199 5015
rect 21189 4981 21223 5015
rect 3249 4777 3283 4811
rect 4537 4777 4571 4811
rect 5089 4777 5123 4811
rect 5549 4777 5583 4811
rect 10149 4777 10183 4811
rect 12633 4777 12667 4811
rect 15761 4777 15795 4811
rect 19349 4777 19383 4811
rect 20269 4777 20303 4811
rect 24133 4777 24167 4811
rect 2421 4709 2455 4743
rect 4077 4709 4111 4743
rect 8309 4709 8343 4743
rect 19625 4709 19659 4743
rect 1409 4641 1443 4675
rect 5917 4641 5951 4675
rect 14749 4641 14783 4675
rect 22201 4641 22235 4675
rect 23213 4641 23247 4675
rect 1683 4573 1717 4607
rect 2789 4573 2823 4607
rect 3893 4573 3927 4607
rect 4905 4573 4939 4607
rect 5273 4573 5307 4607
rect 5733 4573 5767 4607
rect 6191 4573 6225 4607
rect 7297 4573 7331 4607
rect 7571 4573 7605 4607
rect 9137 4573 9171 4607
rect 9411 4573 9445 4607
rect 11621 4573 11655 4607
rect 11713 4573 11747 4607
rect 15023 4573 15057 4607
rect 17233 4573 17267 4607
rect 17507 4573 17541 4607
rect 18797 4573 18831 4607
rect 18889 4573 18923 4607
rect 19533 4573 19567 4607
rect 19809 4573 19843 4607
rect 20085 4573 20119 4607
rect 20177 4573 20211 4607
rect 20453 4573 20487 4607
rect 21925 4573 21959 4607
rect 22845 4573 22879 4607
rect 3157 4505 3191 4539
rect 4445 4505 4479 4539
rect 12081 4505 12115 4539
rect 20720 4505 20754 4539
rect 24041 4505 24075 4539
rect 2973 4437 3007 4471
rect 5457 4437 5491 4471
rect 6929 4437 6963 4471
rect 11345 4437 11379 4471
rect 12449 4437 12483 4471
rect 18245 4437 18279 4471
rect 18613 4437 18647 4471
rect 18981 4437 19015 4471
rect 19901 4437 19935 4471
rect 21833 4437 21867 4471
rect 8953 4233 8987 4267
rect 12541 4233 12575 4267
rect 14105 4233 14139 4267
rect 1869 4165 1903 4199
rect 2421 4165 2455 4199
rect 10149 4165 10183 4199
rect 10517 4165 10551 4199
rect 20177 4165 20211 4199
rect 21465 4165 21499 4199
rect 21649 4165 21683 4199
rect 24041 4165 24075 4199
rect 1409 4097 1443 4131
rect 2697 4097 2731 4131
rect 3617 4097 3651 4131
rect 4629 4097 4663 4131
rect 4903 4097 4937 4131
rect 6193 4097 6227 4131
rect 7297 4097 7331 4131
rect 8309 4097 8343 4131
rect 11771 4097 11805 4131
rect 13367 4097 13401 4131
rect 17693 4097 17727 4131
rect 17877 4097 17911 4131
rect 18245 4097 18279 4131
rect 18521 4097 18555 4131
rect 18795 4097 18829 4131
rect 20821 4097 20855 4131
rect 22017 4097 22051 4131
rect 22383 4097 22417 4131
rect 23581 4097 23615 4131
rect 23765 4097 23799 4131
rect 24225 4097 24259 4131
rect 2605 4029 2639 4063
rect 2881 4029 2915 4063
rect 3734 4029 3768 4063
rect 3893 4029 3927 4063
rect 7113 4029 7147 4063
rect 7757 4029 7791 4063
rect 8033 4029 8067 4063
rect 8171 4029 8205 4063
rect 11529 4029 11563 4063
rect 13093 4029 13127 4063
rect 22109 4029 22143 4063
rect 2145 3961 2179 3995
rect 3341 3961 3375 3995
rect 17877 3961 17911 3995
rect 1593 3893 1627 3927
rect 4537 3893 4571 3927
rect 5641 3893 5675 3927
rect 6009 3893 6043 3927
rect 10609 3893 10643 3927
rect 19533 3893 19567 3927
rect 20269 3893 20303 3927
rect 20913 3893 20947 3927
rect 21833 3893 21867 3927
rect 23121 3893 23155 3927
rect 1593 3689 1627 3723
rect 2789 3689 2823 3723
rect 7573 3689 7607 3723
rect 11897 3689 11931 3723
rect 13553 3689 13587 3723
rect 17785 3689 17819 3723
rect 19717 3689 19751 3723
rect 3433 3621 3467 3655
rect 4445 3621 4479 3655
rect 17509 3621 17543 3655
rect 21741 3621 21775 3655
rect 22293 3621 22327 3655
rect 23857 3621 23891 3655
rect 1777 3553 1811 3587
rect 3801 3553 3835 3587
rect 5733 3553 5767 3587
rect 5917 3553 5951 3587
rect 6377 3553 6411 3587
rect 6653 3553 6687 3587
rect 6791 3553 6825 3587
rect 12541 3553 12575 3587
rect 17233 3553 17267 3587
rect 20729 3553 20763 3587
rect 23121 3553 23155 3587
rect 1409 3485 1443 3519
rect 2051 3485 2085 3519
rect 3985 3485 4019 3519
rect 4721 3485 4755 3519
rect 4838 3485 4872 3519
rect 4997 3485 5031 3519
rect 6929 3485 6963 3519
rect 7849 3485 7883 3519
rect 8125 3485 8159 3519
rect 8769 3485 8803 3519
rect 9413 3485 9447 3519
rect 10885 3485 10919 3519
rect 11159 3485 11193 3519
rect 12783 3485 12817 3519
rect 17141 3485 17175 3519
rect 17417 3485 17451 3519
rect 17601 3485 17635 3519
rect 17693 3485 17727 3519
rect 18613 3485 18647 3519
rect 19257 3485 19291 3519
rect 19441 3485 19475 3519
rect 19809 3485 19843 3519
rect 19993 3485 20027 3519
rect 20637 3485 20671 3519
rect 21003 3485 21037 3519
rect 22109 3485 22143 3519
rect 22293 3485 22327 3519
rect 22661 3485 22695 3519
rect 23305 3485 23339 3519
rect 23765 3485 23799 3519
rect 3249 3417 3283 3451
rect 9505 3417 9539 3451
rect 9873 3417 9907 3451
rect 10241 3417 10275 3451
rect 18061 3417 18095 3451
rect 5641 3349 5675 3383
rect 7665 3349 7699 3383
rect 7941 3349 7975 3383
rect 8585 3349 8619 3383
rect 9137 3349 9171 3383
rect 10425 3349 10459 3383
rect 18153 3349 18187 3383
rect 18705 3349 18739 3383
rect 20085 3349 20119 3383
rect 20453 3349 20487 3383
rect 1777 3145 1811 3179
rect 4629 3145 4663 3179
rect 5917 3145 5951 3179
rect 6561 3145 6595 3179
rect 8585 3145 8619 3179
rect 9965 3145 9999 3179
rect 16957 3145 16991 3179
rect 17325 3145 17359 3179
rect 21465 3145 21499 3179
rect 1685 3077 1719 3111
rect 10885 3077 10919 3111
rect 16497 3077 16531 3111
rect 19073 3077 19107 3111
rect 19625 3077 19659 3111
rect 22998 3077 23032 3111
rect 2237 3009 2271 3043
rect 2605 3009 2639 3043
rect 3985 3009 4019 3043
rect 5163 3039 5197 3073
rect 6469 3009 6503 3043
rect 6929 3009 6963 3043
rect 7205 3009 7239 3043
rect 7481 3009 7515 3043
rect 7847 3009 7881 3043
rect 9227 3009 9261 3043
rect 11621 3009 11655 3043
rect 11895 3019 11929 3053
rect 16773 3009 16807 3043
rect 16957 3009 16991 3043
rect 17233 3009 17267 3043
rect 17509 3009 17543 3043
rect 17693 3009 17727 3043
rect 18337 3009 18371 3043
rect 18521 3009 18555 3043
rect 20269 3009 20303 3043
rect 20361 3009 20395 3043
rect 21649 3009 21683 3043
rect 22109 3009 22143 3043
rect 22753 3009 22787 3043
rect 2789 2941 2823 2975
rect 2973 2941 3007 2975
rect 3709 2941 3743 2975
rect 3847 2941 3881 2975
rect 4905 2941 4939 2975
rect 7573 2941 7607 2975
rect 8953 2941 8987 2975
rect 20913 2941 20947 2975
rect 21833 2941 21867 2975
rect 3433 2873 3467 2907
rect 18705 2873 18739 2907
rect 20085 2873 20119 2907
rect 6745 2805 6779 2839
rect 7021 2805 7055 2839
rect 7297 2805 7331 2839
rect 10977 2805 11011 2839
rect 12633 2805 12667 2839
rect 17049 2805 17083 2839
rect 17785 2805 17819 2839
rect 18153 2805 18187 2839
rect 19165 2805 19199 2839
rect 19717 2805 19751 2839
rect 24133 2805 24167 2839
rect 1777 2601 1811 2635
rect 5365 2601 5399 2635
rect 6929 2601 6963 2635
rect 13461 2601 13495 2635
rect 15853 2601 15887 2635
rect 23857 2601 23891 2635
rect 3341 2533 3375 2567
rect 5825 2533 5859 2567
rect 8953 2533 8987 2567
rect 18705 2533 18739 2567
rect 21925 2533 21959 2567
rect 24041 2533 24075 2567
rect 2329 2465 2363 2499
rect 3801 2465 3835 2499
rect 5917 2465 5951 2499
rect 7573 2465 7607 2499
rect 19901 2465 19935 2499
rect 23305 2465 23339 2499
rect 1685 2397 1719 2431
rect 2603 2397 2637 2431
rect 4059 2367 4093 2401
rect 5641 2397 5675 2431
rect 6191 2397 6225 2431
rect 8401 2397 8435 2431
rect 8677 2397 8711 2431
rect 9137 2397 9171 2431
rect 9413 2397 9447 2431
rect 9689 2397 9723 2431
rect 10701 2397 10735 2431
rect 13829 2397 13863 2431
rect 16037 2397 16071 2431
rect 16313 2397 16347 2431
rect 16589 2397 16623 2431
rect 16865 2397 16899 2431
rect 17141 2397 17175 2431
rect 17325 2397 17359 2431
rect 18797 2397 18831 2431
rect 19441 2397 19475 2431
rect 19717 2397 19751 2431
rect 22569 2397 22603 2431
rect 24225 2397 24259 2431
rect 5273 2329 5307 2363
rect 7389 2329 7423 2363
rect 7757 2329 7791 2363
rect 10241 2329 10275 2363
rect 10333 2329 10367 2363
rect 12173 2329 12207 2363
rect 12445 2329 12479 2363
rect 12541 2329 12575 2363
rect 12909 2329 12943 2363
rect 13277 2329 13311 2363
rect 15761 2329 15795 2363
rect 17570 2329 17604 2363
rect 20637 2329 20671 2363
rect 23765 2329 23799 2363
rect 4813 2261 4847 2295
rect 7849 2261 7883 2295
rect 8217 2261 8251 2295
rect 8493 2261 8527 2295
rect 9229 2261 9263 2295
rect 9505 2261 9539 2295
rect 9965 2261 9999 2295
rect 11069 2261 11103 2295
rect 11253 2261 11287 2295
rect 11713 2261 11747 2295
rect 13645 2261 13679 2295
rect 16129 2261 16163 2295
rect 16405 2261 16439 2295
rect 16681 2261 16715 2295
rect 16957 2261 16991 2295
rect 18981 2261 19015 2295
rect 19257 2261 19291 2295
rect 3893 2057 3927 2091
rect 5273 2057 5307 2091
rect 6101 2057 6135 2091
rect 6929 2057 6963 2091
rect 7665 2057 7699 2091
rect 8033 2057 8067 2091
rect 8769 2057 8803 2091
rect 11069 2057 11103 2091
rect 13369 2057 13403 2091
rect 14473 2057 14507 2091
rect 19073 2057 19107 2091
rect 20637 2057 20671 2091
rect 23213 2057 23247 2091
rect 24041 2057 24075 2091
rect 1501 1989 1535 2023
rect 1869 1989 1903 2023
rect 6469 1989 6503 2023
rect 6837 1989 6871 2023
rect 7573 1989 7607 2023
rect 7941 1989 7975 2023
rect 11897 1989 11931 2023
rect 15485 1989 15519 2023
rect 16773 1989 16807 2023
rect 17325 1989 17359 2023
rect 17877 1989 17911 2023
rect 18429 1989 18463 2023
rect 22078 1989 22112 2023
rect 2237 1921 2271 1955
rect 2881 1921 2915 1955
rect 3155 1921 3189 1955
rect 4261 1921 4295 1955
rect 4535 1921 4569 1955
rect 5825 1921 5859 1955
rect 6009 1921 6043 1955
rect 7205 1921 7239 1955
rect 7389 1921 7423 1955
rect 8217 1921 8251 1955
rect 8677 1921 8711 1955
rect 9597 1921 9631 1955
rect 10299 1931 10333 1965
rect 11713 1921 11747 1955
rect 12615 1951 12649 1985
rect 13921 1921 13955 1955
rect 14841 1921 14875 1955
rect 16037 1921 16071 1955
rect 18797 1921 18831 1955
rect 18889 1921 18923 1955
rect 19257 1921 19291 1955
rect 19524 1921 19558 1955
rect 21833 1921 21867 1955
rect 23765 1921 23799 1955
rect 24225 1921 24259 1955
rect 9229 1853 9263 1887
rect 10057 1853 10091 1887
rect 12357 1853 12391 1887
rect 18153 1853 18187 1887
rect 20821 1853 20855 1887
rect 21097 1853 21131 1887
rect 2513 1785 2547 1819
rect 5641 1785 5675 1819
rect 8401 1785 8435 1819
rect 6561 1717 6595 1751
rect 9873 1717 9907 1751
rect 11529 1717 11563 1751
rect 11989 1717 12023 1751
rect 13737 1717 13771 1751
rect 15025 1717 15059 1751
rect 15577 1717 15611 1751
rect 16129 1717 16163 1751
rect 16865 1717 16899 1751
rect 17417 1717 17451 1751
rect 8677 1513 8711 1547
rect 9321 1513 9355 1547
rect 10609 1513 10643 1547
rect 11253 1513 11287 1547
rect 15393 1513 15427 1547
rect 15945 1513 15979 1547
rect 16313 1513 16347 1547
rect 23121 1513 23155 1547
rect 23857 1513 23891 1547
rect 6193 1445 6227 1479
rect 14749 1445 14783 1479
rect 17509 1445 17543 1479
rect 9597 1377 9631 1411
rect 12541 1377 12575 1411
rect 19901 1377 19935 1411
rect 1501 1309 1535 1343
rect 2237 1309 2271 1343
rect 2605 1309 2639 1343
rect 3341 1309 3375 1343
rect 3801 1309 3835 1343
rect 4169 1309 4203 1343
rect 4445 1309 4479 1343
rect 5825 1309 5859 1343
rect 6009 1309 6043 1343
rect 6377 1309 6411 1343
rect 6653 1309 6687 1343
rect 7297 1309 7331 1343
rect 7573 1309 7607 1343
rect 7941 1309 7975 1343
rect 9045 1309 9079 1343
rect 9839 1309 9873 1343
rect 11069 1309 11103 1343
rect 11713 1309 11747 1343
rect 11805 1309 11839 1343
rect 12265 1309 12299 1343
rect 12725 1309 12759 1343
rect 13093 1309 13127 1343
rect 13461 1309 13495 1343
rect 14105 1309 14139 1343
rect 14565 1309 14599 1343
rect 15301 1309 15335 1343
rect 16497 1309 16531 1343
rect 16773 1309 16807 1343
rect 17785 1309 17819 1343
rect 18245 1309 18279 1343
rect 19257 1309 19291 1343
rect 19349 1309 19383 1343
rect 19717 1309 19751 1343
rect 20821 1309 20855 1343
rect 24225 1309 24259 1343
rect 1961 1241 1995 1275
rect 3065 1241 3099 1275
rect 5273 1241 5307 1275
rect 5457 1241 5491 1275
rect 5641 1241 5675 1275
rect 8401 1241 8435 1275
rect 15853 1241 15887 1275
rect 17325 1241 17359 1275
rect 18889 1241 18923 1275
rect 21465 1241 21499 1275
rect 21833 1241 21867 1275
rect 23765 1241 23799 1275
rect 1685 1173 1719 1207
rect 2053 1173 2087 1207
rect 2421 1173 2455 1207
rect 2789 1173 2823 1207
rect 3157 1173 3191 1207
rect 3525 1173 3559 1207
rect 3985 1173 4019 1207
rect 7481 1173 7515 1207
rect 7757 1173 7791 1207
rect 8125 1173 8159 1207
rect 11529 1173 11563 1207
rect 11989 1173 12023 1207
rect 12909 1173 12943 1207
rect 13277 1173 13311 1207
rect 13645 1173 13679 1207
rect 14289 1173 14323 1207
rect 16865 1173 16899 1207
rect 17969 1173 18003 1207
rect 24041 1173 24075 1207
<< metal1 >>
rect 658 44276 664 44328
rect 716 44316 722 44328
rect 7742 44316 7748 44328
rect 716 44288 7748 44316
rect 716 44276 722 44288
rect 7742 44276 7748 44288
rect 7800 44276 7806 44328
rect 6178 44208 6184 44260
rect 6236 44248 6242 44260
rect 6546 44248 6552 44260
rect 6236 44220 6552 44248
rect 6236 44208 6242 44220
rect 6546 44208 6552 44220
rect 6604 44208 6610 44260
rect 3050 44140 3056 44192
rect 3108 44180 3114 44192
rect 4522 44180 4528 44192
rect 3108 44152 4528 44180
rect 3108 44140 3114 44152
rect 4522 44140 4528 44152
rect 4580 44140 4586 44192
rect 5442 44140 5448 44192
rect 5500 44180 5506 44192
rect 5500 44152 12434 44180
rect 5500 44140 5506 44152
rect 3510 44072 3516 44124
rect 3568 44112 3574 44124
rect 10686 44112 10692 44124
rect 3568 44084 10692 44112
rect 3568 44072 3574 44084
rect 10686 44072 10692 44084
rect 10744 44072 10750 44124
rect 5810 44044 5816 44056
rect 1412 44016 5816 44044
rect 1412 43852 1440 44016
rect 5810 44004 5816 44016
rect 5868 44004 5874 44056
rect 6270 43976 6276 43988
rect 2746 43948 6276 43976
rect 2746 43852 2774 43948
rect 6270 43936 6276 43948
rect 6328 43936 6334 43988
rect 1394 43800 1400 43852
rect 1452 43800 1458 43852
rect 2682 43800 2688 43852
rect 2740 43812 2774 43852
rect 2740 43800 2746 43812
rect 3234 43800 3240 43852
rect 3292 43840 3298 43852
rect 5994 43840 6000 43852
rect 3292 43812 6000 43840
rect 3292 43800 3298 43812
rect 5994 43800 6000 43812
rect 6052 43800 6058 43852
rect 106 43732 112 43784
rect 164 43772 170 43784
rect 164 43744 9904 43772
rect 164 43732 170 43744
rect 9876 43716 9904 43744
rect 1578 43664 1584 43716
rect 1636 43704 1642 43716
rect 6178 43704 6184 43716
rect 1636 43676 6184 43704
rect 1636 43664 1642 43676
rect 6178 43664 6184 43676
rect 6236 43664 6242 43716
rect 9858 43664 9864 43716
rect 9916 43664 9922 43716
rect 2314 43596 2320 43648
rect 2372 43636 2378 43648
rect 5534 43636 5540 43648
rect 2372 43608 5540 43636
rect 2372 43596 2378 43608
rect 5534 43596 5540 43608
rect 5592 43596 5598 43648
rect 5718 43596 5724 43648
rect 5776 43636 5782 43648
rect 11054 43636 11060 43648
rect 5776 43608 11060 43636
rect 5776 43596 5782 43608
rect 11054 43596 11060 43608
rect 11112 43596 11118 43648
rect 12406 43636 12434 44152
rect 18046 44072 18052 44124
rect 18104 44112 18110 44124
rect 19150 44112 19156 44124
rect 18104 44084 19156 44112
rect 18104 44072 18110 44084
rect 19150 44072 19156 44084
rect 19208 44072 19214 44124
rect 17954 44004 17960 44056
rect 18012 44044 18018 44056
rect 19058 44044 19064 44056
rect 18012 44016 19064 44044
rect 18012 44004 18018 44016
rect 19058 44004 19064 44016
rect 19116 44004 19122 44056
rect 17770 43936 17776 43988
rect 17828 43976 17834 43988
rect 18414 43976 18420 43988
rect 17828 43948 18420 43976
rect 17828 43936 17834 43948
rect 18414 43936 18420 43948
rect 18472 43936 18478 43988
rect 16850 43636 16856 43648
rect 12406 43608 16856 43636
rect 16850 43596 16856 43608
rect 16908 43596 16914 43648
rect 1104 43546 24723 43568
rect 1104 43494 6814 43546
rect 6866 43494 6878 43546
rect 6930 43494 6942 43546
rect 6994 43494 7006 43546
rect 7058 43494 7070 43546
rect 7122 43494 12679 43546
rect 12731 43494 12743 43546
rect 12795 43494 12807 43546
rect 12859 43494 12871 43546
rect 12923 43494 12935 43546
rect 12987 43494 18544 43546
rect 18596 43494 18608 43546
rect 18660 43494 18672 43546
rect 18724 43494 18736 43546
rect 18788 43494 18800 43546
rect 18852 43494 24409 43546
rect 24461 43494 24473 43546
rect 24525 43494 24537 43546
rect 24589 43494 24601 43546
rect 24653 43494 24665 43546
rect 24717 43494 24723 43546
rect 1104 43472 24723 43494
rect 1578 43392 1584 43444
rect 1636 43392 1642 43444
rect 2317 43435 2375 43441
rect 2317 43401 2329 43435
rect 2363 43432 2375 43435
rect 3142 43432 3148 43444
rect 2363 43404 3148 43432
rect 2363 43401 2375 43404
rect 2317 43395 2375 43401
rect 3142 43392 3148 43404
rect 3200 43392 3206 43444
rect 5626 43432 5632 43444
rect 3528 43404 5632 43432
rect 2682 43324 2688 43376
rect 2740 43324 2746 43376
rect 3053 43367 3111 43373
rect 3053 43333 3065 43367
rect 3099 43364 3111 43367
rect 3528 43364 3556 43404
rect 5626 43392 5632 43404
rect 5684 43392 5690 43444
rect 5902 43392 5908 43444
rect 5960 43392 5966 43444
rect 6089 43435 6147 43441
rect 6089 43401 6101 43435
rect 6135 43432 6147 43435
rect 6730 43432 6736 43444
rect 6135 43404 6736 43432
rect 6135 43401 6147 43404
rect 6089 43395 6147 43401
rect 6730 43392 6736 43404
rect 6788 43392 6794 43444
rect 7190 43392 7196 43444
rect 7248 43392 7254 43444
rect 8205 43435 8263 43441
rect 8205 43401 8217 43435
rect 8251 43432 8263 43435
rect 8665 43435 8723 43441
rect 8251 43404 8524 43432
rect 8251 43401 8263 43404
rect 8205 43395 8263 43401
rect 3099 43336 3556 43364
rect 3605 43367 3663 43373
rect 3099 43333 3111 43336
rect 3053 43327 3111 43333
rect 3605 43333 3617 43367
rect 3651 43364 3663 43367
rect 5920 43364 5948 43392
rect 7742 43364 7748 43376
rect 3651 43336 5948 43364
rect 6288 43336 7748 43364
rect 3651 43333 3663 43336
rect 3605 43327 3663 43333
rect 1394 43256 1400 43308
rect 1452 43256 1458 43308
rect 2041 43299 2099 43305
rect 2041 43265 2053 43299
rect 2087 43296 2099 43299
rect 2958 43296 2964 43308
rect 2087 43268 2964 43296
rect 2087 43265 2099 43268
rect 2041 43259 2099 43265
rect 2958 43256 2964 43268
rect 3016 43256 3022 43308
rect 3234 43256 3240 43308
rect 3292 43256 3298 43308
rect 4063 43299 4121 43305
rect 4063 43265 4075 43299
rect 4109 43296 4121 43299
rect 4706 43296 4712 43308
rect 4109 43268 4712 43296
rect 4109 43265 4121 43268
rect 4063 43259 4121 43265
rect 4706 43256 4712 43268
rect 4764 43256 4770 43308
rect 5261 43299 5319 43305
rect 5261 43265 5273 43299
rect 5307 43296 5319 43299
rect 5718 43296 5724 43308
rect 5307 43268 5724 43296
rect 5307 43265 5319 43268
rect 5261 43259 5319 43265
rect 5718 43256 5724 43268
rect 5776 43256 5782 43308
rect 5813 43299 5871 43305
rect 5813 43265 5825 43299
rect 5859 43296 5871 43299
rect 6288 43296 6316 43336
rect 7742 43324 7748 43336
rect 7800 43324 7806 43376
rect 5859 43268 6316 43296
rect 6365 43299 6423 43305
rect 5859 43265 5871 43268
rect 5813 43259 5871 43265
rect 6365 43265 6377 43299
rect 6411 43265 6423 43299
rect 6365 43259 6423 43265
rect 3326 43188 3332 43240
rect 3384 43228 3390 43240
rect 3789 43231 3847 43237
rect 3789 43228 3801 43231
rect 3384 43200 3801 43228
rect 3384 43188 3390 43200
rect 3789 43197 3801 43200
rect 3835 43197 3847 43231
rect 3789 43191 3847 43197
rect 5534 43188 5540 43240
rect 5592 43188 5598 43240
rect 2498 43120 2504 43172
rect 2556 43160 2562 43172
rect 4801 43163 4859 43169
rect 2556 43132 3832 43160
rect 2556 43120 2562 43132
rect 3804 43092 3832 43132
rect 4801 43129 4813 43163
rect 4847 43129 4859 43163
rect 4801 43123 4859 43129
rect 4816 43092 4844 43123
rect 3804 43064 4844 43092
rect 6380 43092 6408 43259
rect 6638 43256 6644 43308
rect 6696 43296 6702 43308
rect 8496 43305 8524 43404
rect 8665 43401 8677 43435
rect 8711 43432 8723 43435
rect 8938 43432 8944 43444
rect 8711 43404 8944 43432
rect 8711 43401 8723 43404
rect 8665 43395 8723 43401
rect 8938 43392 8944 43404
rect 8996 43392 9002 43444
rect 9125 43435 9183 43441
rect 9125 43401 9137 43435
rect 9171 43432 9183 43435
rect 9490 43432 9496 43444
rect 9171 43404 9496 43432
rect 9171 43401 9183 43404
rect 9125 43395 9183 43401
rect 9490 43392 9496 43404
rect 9548 43392 9554 43444
rect 9677 43435 9735 43441
rect 9677 43401 9689 43435
rect 9723 43432 9735 43435
rect 9766 43432 9772 43444
rect 9723 43404 9772 43432
rect 9723 43401 9735 43404
rect 9677 43395 9735 43401
rect 9766 43392 9772 43404
rect 9824 43392 9830 43444
rect 9858 43392 9864 43444
rect 9916 43432 9922 43444
rect 10045 43435 10103 43441
rect 10045 43432 10057 43435
rect 9916 43404 10057 43432
rect 9916 43392 9922 43404
rect 10045 43401 10057 43404
rect 10091 43401 10103 43435
rect 10045 43395 10103 43401
rect 12158 43392 12164 43444
rect 12216 43432 12222 43444
rect 14277 43435 14335 43441
rect 14277 43432 14289 43435
rect 12216 43404 14289 43432
rect 12216 43392 12222 43404
rect 14277 43401 14289 43404
rect 14323 43401 14335 43435
rect 14277 43395 14335 43401
rect 16114 43392 16120 43444
rect 16172 43432 16178 43444
rect 16172 43404 17172 43432
rect 16172 43392 16178 43404
rect 8772 43336 9812 43364
rect 6917 43299 6975 43305
rect 6917 43296 6929 43299
rect 6696 43268 6929 43296
rect 6696 43256 6702 43268
rect 6917 43265 6929 43268
rect 6963 43265 6975 43299
rect 6917 43259 6975 43265
rect 7469 43299 7527 43305
rect 7469 43265 7481 43299
rect 7515 43296 7527 43299
rect 8481 43299 8539 43305
rect 7515 43268 8432 43296
rect 7515 43265 7527 43268
rect 7469 43259 7527 43265
rect 7558 43188 7564 43240
rect 7616 43188 7622 43240
rect 8404 43228 8432 43268
rect 8481 43265 8493 43299
rect 8527 43296 8539 43299
rect 8772 43296 8800 43336
rect 9784 43308 9812 43336
rect 9968 43336 12204 43364
rect 8527 43268 8800 43296
rect 8941 43299 8999 43305
rect 8527 43265 8539 43268
rect 8481 43259 8539 43265
rect 8941 43265 8953 43299
rect 8987 43296 8999 43299
rect 9401 43299 9459 43305
rect 8987 43268 9352 43296
rect 8987 43265 8999 43268
rect 8941 43259 8999 43265
rect 9122 43228 9128 43240
rect 8404 43200 9128 43228
rect 9122 43188 9128 43200
rect 9180 43188 9186 43240
rect 6549 43163 6607 43169
rect 6549 43129 6561 43163
rect 6595 43160 6607 43163
rect 7576 43160 7604 43188
rect 6595 43132 7604 43160
rect 7745 43163 7803 43169
rect 6595 43129 6607 43132
rect 6549 43123 6607 43129
rect 7745 43129 7757 43163
rect 7791 43160 7803 43163
rect 8662 43160 8668 43172
rect 7791 43132 8668 43160
rect 7791 43129 7803 43132
rect 7745 43123 7803 43129
rect 8662 43120 8668 43132
rect 8720 43120 8726 43172
rect 9324 43160 9352 43268
rect 9401 43265 9413 43299
rect 9447 43296 9459 43299
rect 9582 43296 9588 43308
rect 9447 43268 9588 43296
rect 9447 43265 9459 43268
rect 9401 43259 9459 43265
rect 9582 43256 9588 43268
rect 9640 43256 9646 43308
rect 9766 43256 9772 43308
rect 9824 43256 9830 43308
rect 9968 43305 9996 43336
rect 9953 43299 10011 43305
rect 9953 43265 9965 43299
rect 9999 43265 10011 43299
rect 9953 43259 10011 43265
rect 10226 43256 10232 43308
rect 10284 43296 10290 43308
rect 10413 43299 10471 43305
rect 10413 43296 10425 43299
rect 10284 43268 10425 43296
rect 10284 43256 10290 43268
rect 10413 43265 10425 43268
rect 10459 43265 10471 43299
rect 10413 43259 10471 43265
rect 10962 43256 10968 43308
rect 11020 43256 11026 43308
rect 11146 43256 11152 43308
rect 11204 43296 11210 43308
rect 11517 43299 11575 43305
rect 11517 43296 11529 43299
rect 11204 43268 11529 43296
rect 11204 43256 11210 43268
rect 11517 43265 11529 43268
rect 11563 43265 11575 43299
rect 11517 43259 11575 43265
rect 12066 43256 12072 43308
rect 12124 43256 12130 43308
rect 12176 43296 12204 43336
rect 12250 43324 12256 43376
rect 12308 43364 12314 43376
rect 12437 43367 12495 43373
rect 12437 43364 12449 43367
rect 12308 43336 12449 43364
rect 12308 43324 12314 43336
rect 12437 43333 12449 43336
rect 12483 43333 12495 43367
rect 12437 43327 12495 43333
rect 13170 43324 13176 43376
rect 13228 43324 13234 43376
rect 13538 43324 13544 43376
rect 13596 43324 13602 43376
rect 15286 43324 15292 43376
rect 15344 43364 15350 43376
rect 15841 43367 15899 43373
rect 15841 43364 15853 43367
rect 15344 43336 15853 43364
rect 15344 43324 15350 43336
rect 15841 43333 15853 43336
rect 15887 43333 15899 43367
rect 15841 43327 15899 43333
rect 16022 43324 16028 43376
rect 16080 43364 16086 43376
rect 16761 43367 16819 43373
rect 16761 43364 16773 43367
rect 16080 43336 16773 43364
rect 16080 43324 16086 43336
rect 16761 43333 16773 43336
rect 16807 43333 16819 43367
rect 16761 43327 16819 43333
rect 16850 43324 16856 43376
rect 16908 43364 16914 43376
rect 17144 43373 17172 43404
rect 17310 43392 17316 43444
rect 17368 43432 17374 43444
rect 18325 43435 18383 43441
rect 18325 43432 18337 43435
rect 17368 43404 18337 43432
rect 17368 43392 17374 43404
rect 18325 43401 18337 43404
rect 18371 43401 18383 43435
rect 18325 43395 18383 43401
rect 20254 43392 20260 43444
rect 20312 43432 20318 43444
rect 20349 43435 20407 43441
rect 20349 43432 20361 43435
rect 20312 43404 20361 43432
rect 20312 43392 20318 43404
rect 20349 43401 20361 43404
rect 20395 43401 20407 43435
rect 20349 43395 20407 43401
rect 20530 43392 20536 43444
rect 20588 43432 20594 43444
rect 20717 43435 20775 43441
rect 20717 43432 20729 43435
rect 20588 43404 20729 43432
rect 20588 43392 20594 43404
rect 20717 43401 20729 43404
rect 20763 43401 20775 43435
rect 20717 43395 20775 43401
rect 21358 43392 21364 43444
rect 21416 43432 21422 43444
rect 22373 43435 22431 43441
rect 22373 43432 22385 43435
rect 21416 43404 22385 43432
rect 21416 43392 21422 43404
rect 22373 43401 22385 43404
rect 22419 43401 22431 43435
rect 22373 43395 22431 43401
rect 23750 43392 23756 43444
rect 23808 43392 23814 43444
rect 25498 43392 25504 43444
rect 25556 43392 25562 43444
rect 16945 43367 17003 43373
rect 16945 43364 16957 43367
rect 16908 43336 16957 43364
rect 16908 43324 16914 43336
rect 16945 43333 16957 43336
rect 16991 43333 17003 43367
rect 16945 43327 17003 43333
rect 17129 43367 17187 43373
rect 17129 43333 17141 43367
rect 17175 43333 17187 43367
rect 17129 43327 17187 43333
rect 17218 43324 17224 43376
rect 17276 43364 17282 43376
rect 17276 43336 18276 43364
rect 17276 43324 17282 43336
rect 12342 43296 12348 43308
rect 12176 43268 12348 43296
rect 12342 43256 12348 43268
rect 12400 43256 12406 43308
rect 12805 43299 12863 43305
rect 12805 43265 12817 43299
rect 12851 43296 12863 43299
rect 13078 43296 13084 43308
rect 12851 43268 13084 43296
rect 12851 43265 12863 43268
rect 12805 43259 12863 43265
rect 13078 43256 13084 43268
rect 13136 43256 13142 43308
rect 14090 43256 14096 43308
rect 14148 43256 14154 43308
rect 14458 43256 14464 43308
rect 14516 43256 14522 43308
rect 14826 43256 14832 43308
rect 14884 43256 14890 43308
rect 15562 43256 15568 43308
rect 15620 43296 15626 43308
rect 16117 43299 16175 43305
rect 16117 43296 16129 43299
rect 15620 43268 16129 43296
rect 15620 43256 15626 43268
rect 16117 43265 16129 43268
rect 16163 43265 16175 43299
rect 16117 43259 16175 43265
rect 16390 43256 16396 43308
rect 16448 43296 16454 43308
rect 18248 43305 18276 43336
rect 18414 43324 18420 43376
rect 18472 43364 18478 43376
rect 18472 43336 18828 43364
rect 18472 43324 18478 43336
rect 18800 43305 18828 43336
rect 18874 43324 18880 43376
rect 18932 43364 18938 43376
rect 21637 43367 21695 43373
rect 18932 43336 20024 43364
rect 18932 43324 18938 43336
rect 17405 43299 17463 43305
rect 17405 43296 17417 43299
rect 16448 43268 17417 43296
rect 16448 43256 16454 43268
rect 17405 43265 17417 43268
rect 17451 43265 17463 43299
rect 17405 43259 17463 43265
rect 17957 43299 18015 43305
rect 17957 43265 17969 43299
rect 18003 43265 18015 43299
rect 17957 43259 18015 43265
rect 18233 43299 18291 43305
rect 18233 43265 18245 43299
rect 18279 43265 18291 43299
rect 18233 43259 18291 43265
rect 18509 43299 18567 43305
rect 18509 43265 18521 43299
rect 18555 43265 18567 43299
rect 18509 43259 18567 43265
rect 18785 43299 18843 43305
rect 18785 43265 18797 43299
rect 18831 43265 18843 43299
rect 18785 43259 18843 43265
rect 10502 43188 10508 43240
rect 10560 43228 10566 43240
rect 10597 43231 10655 43237
rect 10597 43228 10609 43231
rect 10560 43200 10609 43228
rect 10560 43188 10566 43200
rect 10597 43197 10609 43200
rect 10643 43197 10655 43231
rect 13170 43228 13176 43240
rect 10597 43191 10655 43197
rect 11164 43200 13176 43228
rect 10410 43160 10416 43172
rect 9324 43132 10416 43160
rect 10410 43120 10416 43132
rect 10468 43120 10474 43172
rect 11164 43169 11192 43200
rect 13170 43188 13176 43200
rect 13228 43188 13234 43240
rect 15010 43188 15016 43240
rect 15068 43228 15074 43240
rect 15105 43231 15163 43237
rect 15105 43228 15117 43231
rect 15068 43200 15117 43228
rect 15068 43188 15074 43200
rect 15105 43197 15117 43200
rect 15151 43197 15163 43231
rect 15105 43191 15163 43197
rect 16666 43188 16672 43240
rect 16724 43228 16730 43240
rect 17972 43228 18000 43259
rect 16724 43200 18000 43228
rect 16724 43188 16730 43200
rect 18046 43188 18052 43240
rect 18104 43228 18110 43240
rect 18524 43228 18552 43259
rect 19058 43256 19064 43308
rect 19116 43256 19122 43308
rect 19150 43256 19156 43308
rect 19208 43296 19214 43308
rect 19996 43305 20024 43336
rect 21637 43333 21649 43367
rect 21683 43364 21695 43367
rect 25516 43364 25544 43392
rect 21683 43336 25544 43364
rect 21683 43333 21695 43336
rect 21637 43327 21695 43333
rect 19429 43299 19487 43305
rect 19429 43296 19441 43299
rect 19208 43268 19441 43296
rect 19208 43256 19214 43268
rect 19429 43265 19441 43268
rect 19475 43265 19487 43299
rect 19429 43259 19487 43265
rect 19705 43299 19763 43305
rect 19705 43265 19717 43299
rect 19751 43265 19763 43299
rect 19705 43259 19763 43265
rect 19981 43299 20039 43305
rect 19981 43265 19993 43299
rect 20027 43265 20039 43299
rect 19981 43259 20039 43265
rect 18104 43200 18552 43228
rect 18104 43188 18110 43200
rect 18690 43188 18696 43240
rect 18748 43228 18754 43240
rect 19720 43228 19748 43259
rect 20162 43256 20168 43308
rect 20220 43256 20226 43308
rect 20625 43299 20683 43305
rect 20625 43296 20637 43299
rect 20272 43268 20637 43296
rect 18748 43200 19748 43228
rect 18748 43188 18754 43200
rect 20070 43188 20076 43240
rect 20128 43228 20134 43240
rect 20272 43228 20300 43268
rect 20625 43265 20637 43268
rect 20671 43265 20683 43299
rect 20625 43259 20683 43265
rect 21266 43256 21272 43308
rect 21324 43256 21330 43308
rect 21821 43299 21879 43305
rect 21821 43265 21833 43299
rect 21867 43296 21879 43299
rect 22281 43299 22339 43305
rect 21867 43268 22048 43296
rect 21867 43265 21879 43268
rect 21821 43259 21879 43265
rect 20128 43200 20300 43228
rect 20128 43188 20134 43200
rect 20806 43188 20812 43240
rect 20864 43188 20870 43240
rect 22020 43228 22048 43268
rect 22281 43265 22293 43299
rect 22327 43296 22339 43299
rect 22370 43296 22376 43308
rect 22327 43268 22376 43296
rect 22327 43265 22339 43268
rect 22281 43259 22339 43265
rect 22370 43256 22376 43268
rect 22428 43256 22434 43308
rect 22830 43256 22836 43308
rect 22888 43256 22894 43308
rect 23477 43299 23535 43305
rect 23477 43265 23489 43299
rect 23523 43265 23535 43299
rect 23477 43259 23535 43265
rect 23492 43228 23520 43259
rect 23658 43256 23664 43308
rect 23716 43256 23722 43308
rect 24210 43228 24216 43240
rect 22020 43200 23336 43228
rect 23492 43200 24216 43228
rect 11149 43163 11207 43169
rect 11149 43129 11161 43163
rect 11195 43129 11207 43163
rect 11149 43123 11207 43129
rect 11882 43120 11888 43172
rect 11940 43160 11946 43172
rect 12989 43163 13047 43169
rect 12989 43160 13001 43163
rect 11940 43132 13001 43160
rect 11940 43120 11946 43132
rect 12989 43129 13001 43132
rect 13035 43129 13047 43163
rect 12989 43123 13047 43129
rect 13354 43120 13360 43172
rect 13412 43120 13418 43172
rect 14182 43120 14188 43172
rect 14240 43160 14246 43172
rect 14240 43132 17264 43160
rect 14240 43120 14246 43132
rect 9674 43092 9680 43104
rect 6380 43064 9680 43092
rect 9674 43052 9680 43064
rect 9732 43052 9738 43104
rect 9766 43052 9772 43104
rect 9824 43092 9830 43104
rect 10870 43092 10876 43104
rect 9824 43064 10876 43092
rect 9824 43052 9830 43064
rect 10870 43052 10876 43064
rect 10928 43052 10934 43104
rect 11701 43095 11759 43101
rect 11701 43061 11713 43095
rect 11747 43092 11759 43095
rect 11790 43092 11796 43104
rect 11747 43064 11796 43092
rect 11747 43061 11759 43064
rect 11701 43055 11759 43061
rect 11790 43052 11796 43064
rect 11848 43052 11854 43104
rect 11974 43052 11980 43104
rect 12032 43092 12038 43104
rect 12253 43095 12311 43101
rect 12253 43092 12265 43095
rect 12032 43064 12265 43092
rect 12032 43052 12038 43064
rect 12253 43061 12265 43064
rect 12299 43061 12311 43095
rect 12253 43055 12311 43061
rect 12526 43052 12532 43104
rect 12584 43052 12590 43104
rect 13630 43052 13636 43104
rect 13688 43052 13694 43104
rect 14642 43052 14648 43104
rect 14700 43052 14706 43104
rect 15470 43052 15476 43104
rect 15528 43092 15534 43104
rect 15933 43095 15991 43101
rect 15933 43092 15945 43095
rect 15528 43064 15945 43092
rect 15528 43052 15534 43064
rect 15933 43061 15945 43064
rect 15979 43061 15991 43095
rect 15933 43055 15991 43061
rect 16298 43052 16304 43104
rect 16356 43052 16362 43104
rect 17236 43101 17264 43132
rect 17862 43120 17868 43172
rect 17920 43160 17926 43172
rect 18877 43163 18935 43169
rect 18877 43160 18889 43163
rect 17920 43132 18889 43160
rect 17920 43120 17926 43132
rect 18877 43129 18889 43132
rect 18923 43129 18935 43163
rect 18877 43123 18935 43129
rect 19610 43120 19616 43172
rect 19668 43160 19674 43172
rect 20530 43160 20536 43172
rect 19668 43132 20536 43160
rect 19668 43120 19674 43132
rect 20530 43120 20536 43132
rect 20588 43120 20594 43172
rect 20824 43160 20852 43188
rect 23308 43169 23336 43200
rect 24210 43188 24216 43200
rect 24268 43188 24274 43240
rect 22005 43163 22063 43169
rect 22005 43160 22017 43163
rect 20824 43132 22017 43160
rect 22005 43129 22017 43132
rect 22051 43129 22063 43163
rect 22005 43123 22063 43129
rect 23293 43163 23351 43169
rect 23293 43129 23305 43163
rect 23339 43129 23351 43163
rect 23293 43123 23351 43129
rect 17221 43095 17279 43101
rect 17221 43061 17233 43095
rect 17267 43061 17279 43095
rect 17221 43055 17279 43061
rect 17586 43052 17592 43104
rect 17644 43052 17650 43104
rect 17770 43052 17776 43104
rect 17828 43052 17834 43104
rect 18046 43052 18052 43104
rect 18104 43052 18110 43104
rect 18598 43052 18604 43104
rect 18656 43052 18662 43104
rect 19242 43052 19248 43104
rect 19300 43052 19306 43104
rect 19426 43052 19432 43104
rect 19484 43092 19490 43104
rect 19521 43095 19579 43101
rect 19521 43092 19533 43095
rect 19484 43064 19533 43092
rect 19484 43052 19490 43064
rect 19521 43061 19533 43064
rect 19567 43061 19579 43095
rect 19521 43055 19579 43061
rect 19794 43052 19800 43104
rect 19852 43052 19858 43104
rect 21910 43052 21916 43104
rect 21968 43092 21974 43104
rect 22925 43095 22983 43101
rect 22925 43092 22937 43095
rect 21968 43064 22937 43092
rect 21968 43052 21974 43064
rect 22925 43061 22937 43064
rect 22971 43061 22983 43095
rect 22925 43055 22983 43061
rect 1104 43002 24564 43024
rect 1104 42950 3882 43002
rect 3934 42950 3946 43002
rect 3998 42950 4010 43002
rect 4062 42950 4074 43002
rect 4126 42950 4138 43002
rect 4190 42950 9747 43002
rect 9799 42950 9811 43002
rect 9863 42950 9875 43002
rect 9927 42950 9939 43002
rect 9991 42950 10003 43002
rect 10055 42950 15612 43002
rect 15664 42950 15676 43002
rect 15728 42950 15740 43002
rect 15792 42950 15804 43002
rect 15856 42950 15868 43002
rect 15920 42950 21477 43002
rect 21529 42950 21541 43002
rect 21593 42950 21605 43002
rect 21657 42950 21669 43002
rect 21721 42950 21733 43002
rect 21785 42950 24564 43002
rect 1104 42928 24564 42950
rect 2961 42891 3019 42897
rect 2961 42857 2973 42891
rect 3007 42888 3019 42891
rect 3050 42888 3056 42900
rect 3007 42860 3056 42888
rect 3007 42857 3019 42860
rect 2961 42851 3019 42857
rect 3050 42848 3056 42860
rect 3108 42848 3114 42900
rect 3712 42860 6132 42888
rect 3234 42780 3240 42832
rect 3292 42820 3298 42832
rect 3510 42820 3516 42832
rect 3292 42792 3516 42820
rect 3292 42780 3298 42792
rect 3510 42780 3516 42792
rect 3568 42780 3574 42832
rect 1857 42755 1915 42761
rect 1857 42721 1869 42755
rect 1903 42752 1915 42755
rect 3418 42752 3424 42764
rect 1903 42724 3424 42752
rect 1903 42721 1915 42724
rect 1857 42715 1915 42721
rect 3418 42712 3424 42724
rect 3476 42712 3482 42764
rect 934 42644 940 42696
rect 992 42684 998 42696
rect 3712 42684 3740 42860
rect 3789 42823 3847 42829
rect 3789 42789 3801 42823
rect 3835 42789 3847 42823
rect 3789 42783 3847 42789
rect 992 42656 3740 42684
rect 992 42644 998 42656
rect 1581 42619 1639 42625
rect 1581 42585 1593 42619
rect 1627 42616 1639 42619
rect 1946 42616 1952 42628
rect 1627 42588 1952 42616
rect 1627 42585 1639 42588
rect 1581 42579 1639 42585
rect 1946 42576 1952 42588
rect 2004 42576 2010 42628
rect 2317 42619 2375 42625
rect 2317 42585 2329 42619
rect 2363 42616 2375 42619
rect 2682 42616 2688 42628
rect 2363 42588 2688 42616
rect 2363 42585 2375 42588
rect 2317 42579 2375 42585
rect 2682 42576 2688 42588
rect 2740 42576 2746 42628
rect 3234 42576 3240 42628
rect 3292 42576 3298 42628
rect 3804 42616 3832 42783
rect 6104 42752 6132 42860
rect 7926 42848 7932 42900
rect 7984 42848 7990 42900
rect 8478 42848 8484 42900
rect 8536 42848 8542 42900
rect 8588 42860 9076 42888
rect 8018 42780 8024 42832
rect 8076 42820 8082 42832
rect 8588 42820 8616 42860
rect 8076 42792 8616 42820
rect 9048 42820 9076 42860
rect 9490 42848 9496 42900
rect 9548 42848 9554 42900
rect 9582 42848 9588 42900
rect 9640 42888 9646 42900
rect 14918 42888 14924 42900
rect 9640 42860 14924 42888
rect 9640 42848 9646 42860
rect 14918 42848 14924 42860
rect 14976 42848 14982 42900
rect 18598 42888 18604 42900
rect 17972 42860 18604 42888
rect 10226 42820 10232 42832
rect 9048 42792 10232 42820
rect 8076 42780 8082 42792
rect 10226 42780 10232 42792
rect 10284 42780 10290 42832
rect 10781 42823 10839 42829
rect 10781 42789 10793 42823
rect 10827 42789 10839 42823
rect 10781 42783 10839 42789
rect 14461 42823 14519 42829
rect 14461 42789 14473 42823
rect 14507 42789 14519 42823
rect 17770 42820 17776 42832
rect 14461 42783 14519 42789
rect 16960 42792 17776 42820
rect 7377 42755 7435 42761
rect 7377 42752 7389 42755
rect 6104 42724 7389 42752
rect 7377 42721 7389 42724
rect 7423 42721 7435 42755
rect 7377 42715 7435 42721
rect 9490 42712 9496 42764
rect 9548 42752 9554 42764
rect 10796 42752 10824 42783
rect 9548 42724 10824 42752
rect 9548 42712 9554 42724
rect 13078 42712 13084 42764
rect 13136 42752 13142 42764
rect 14476 42752 14504 42783
rect 13136 42724 14504 42752
rect 13136 42712 13142 42724
rect 3970 42644 3976 42696
rect 4028 42644 4034 42696
rect 4065 42687 4123 42693
rect 4065 42653 4077 42687
rect 4111 42684 4123 42687
rect 4246 42684 4252 42696
rect 4111 42656 4252 42684
rect 4111 42653 4123 42656
rect 4065 42647 4123 42653
rect 4246 42644 4252 42656
rect 4304 42644 4310 42696
rect 4339 42687 4397 42693
rect 4339 42653 4351 42687
rect 4385 42684 4397 42687
rect 4430 42684 4436 42696
rect 4385 42656 4436 42684
rect 4385 42653 4397 42656
rect 4339 42647 4397 42653
rect 4430 42644 4436 42656
rect 4488 42684 4494 42696
rect 4706 42684 4712 42696
rect 4488 42656 4712 42684
rect 4488 42644 4494 42656
rect 4706 42644 4712 42656
rect 4764 42644 4770 42696
rect 4890 42644 4896 42696
rect 4948 42684 4954 42696
rect 5350 42684 5356 42696
rect 4948 42656 5356 42684
rect 4948 42644 4954 42656
rect 5350 42644 5356 42656
rect 5408 42684 5414 42696
rect 5445 42687 5503 42693
rect 5445 42684 5457 42687
rect 5408 42656 5457 42684
rect 5408 42644 5414 42656
rect 5445 42653 5457 42656
rect 5491 42653 5503 42687
rect 5718 42684 5724 42696
rect 5679 42656 5724 42684
rect 5445 42647 5503 42653
rect 5718 42644 5724 42656
rect 5776 42644 5782 42696
rect 7837 42687 7895 42693
rect 7837 42684 7849 42687
rect 5828 42656 7849 42684
rect 5828 42616 5856 42656
rect 7837 42653 7849 42656
rect 7883 42653 7895 42687
rect 7837 42647 7895 42653
rect 8938 42644 8944 42696
rect 8996 42644 9002 42696
rect 9861 42687 9919 42693
rect 9861 42653 9873 42687
rect 9907 42684 9919 42687
rect 10134 42684 10140 42696
rect 9907 42656 10140 42684
rect 9907 42653 9919 42656
rect 9861 42647 9919 42653
rect 10134 42644 10140 42656
rect 10192 42644 10198 42696
rect 10226 42644 10232 42696
rect 10284 42644 10290 42696
rect 10594 42644 10600 42696
rect 10652 42644 10658 42696
rect 11422 42644 11428 42696
rect 11480 42684 11486 42696
rect 11701 42687 11759 42693
rect 11701 42684 11713 42687
rect 11480 42656 11713 42684
rect 11480 42644 11486 42656
rect 11701 42653 11713 42656
rect 11747 42653 11759 42687
rect 11701 42647 11759 42653
rect 11790 42644 11796 42696
rect 11848 42644 11854 42696
rect 12618 42644 12624 42696
rect 12676 42644 12682 42696
rect 13722 42644 13728 42696
rect 13780 42644 13786 42696
rect 14274 42644 14280 42696
rect 14332 42644 14338 42696
rect 15102 42644 15108 42696
rect 15160 42644 15166 42696
rect 16301 42687 16359 42693
rect 16301 42653 16313 42687
rect 16347 42684 16359 42687
rect 16960 42684 16988 42792
rect 17770 42780 17776 42792
rect 17828 42780 17834 42832
rect 17972 42752 18000 42860
rect 18598 42848 18604 42860
rect 18656 42848 18662 42900
rect 19150 42848 19156 42900
rect 19208 42888 19214 42900
rect 19208 42860 20116 42888
rect 19208 42848 19214 42860
rect 19242 42820 19248 42832
rect 17420 42724 18000 42752
rect 18156 42792 19248 42820
rect 16347 42656 16988 42684
rect 17037 42687 17095 42693
rect 16347 42653 16359 42656
rect 16301 42647 16359 42653
rect 17037 42653 17049 42687
rect 17083 42684 17095 42687
rect 17310 42684 17316 42696
rect 17083 42656 17316 42684
rect 17083 42653 17095 42656
rect 17037 42647 17095 42653
rect 17310 42644 17316 42656
rect 17368 42644 17374 42696
rect 17420 42693 17448 42724
rect 17405 42687 17463 42693
rect 17405 42653 17417 42687
rect 17451 42653 17463 42687
rect 17405 42647 17463 42653
rect 17773 42687 17831 42693
rect 17773 42653 17785 42687
rect 17819 42684 17831 42687
rect 17862 42684 17868 42696
rect 17819 42656 17868 42684
rect 17819 42653 17831 42656
rect 17773 42647 17831 42653
rect 17862 42644 17868 42656
rect 17920 42644 17926 42696
rect 18046 42644 18052 42696
rect 18104 42644 18110 42696
rect 18156 42693 18184 42792
rect 19242 42780 19248 42792
rect 19300 42780 19306 42832
rect 19794 42780 19800 42832
rect 19852 42780 19858 42832
rect 19981 42823 20039 42829
rect 19981 42789 19993 42823
rect 20027 42789 20039 42823
rect 19981 42783 20039 42789
rect 19812 42752 19840 42780
rect 18892 42724 19840 42752
rect 18141 42687 18199 42693
rect 18141 42653 18153 42687
rect 18187 42653 18199 42687
rect 18141 42647 18199 42653
rect 18322 42644 18328 42696
rect 18380 42644 18386 42696
rect 18892 42693 18920 42724
rect 18877 42687 18935 42693
rect 18877 42653 18889 42687
rect 18923 42653 18935 42687
rect 18877 42647 18935 42653
rect 19337 42687 19395 42693
rect 19337 42653 19349 42687
rect 19383 42684 19395 42687
rect 19996 42684 20024 42783
rect 20088 42752 20116 42860
rect 20162 42848 20168 42900
rect 20220 42888 20226 42900
rect 20257 42891 20315 42897
rect 20257 42888 20269 42891
rect 20220 42860 20269 42888
rect 20220 42848 20226 42860
rect 20257 42857 20269 42860
rect 20303 42857 20315 42891
rect 20257 42851 20315 42857
rect 20533 42891 20591 42897
rect 20533 42857 20545 42891
rect 20579 42888 20591 42891
rect 20622 42888 20628 42900
rect 20579 42860 20628 42888
rect 20579 42857 20591 42860
rect 20533 42851 20591 42857
rect 20622 42848 20628 42860
rect 20680 42848 20686 42900
rect 22005 42891 22063 42897
rect 22005 42857 22017 42891
rect 22051 42888 22063 42891
rect 22094 42888 22100 42900
rect 22051 42860 22100 42888
rect 22051 42857 22063 42860
rect 22005 42851 22063 42857
rect 22094 42848 22100 42860
rect 22152 42848 22158 42900
rect 22646 42848 22652 42900
rect 22704 42888 22710 42900
rect 23477 42891 23535 42897
rect 23477 42888 23489 42891
rect 22704 42860 23489 42888
rect 22704 42848 22710 42860
rect 23477 42857 23489 42860
rect 23523 42857 23535 42891
rect 23477 42851 23535 42857
rect 20346 42780 20352 42832
rect 20404 42820 20410 42832
rect 22830 42820 22836 42832
rect 20404 42792 22836 42820
rect 20404 42780 20410 42792
rect 22830 42780 22836 42792
rect 22888 42780 22894 42832
rect 20088 42724 20208 42752
rect 20180 42693 20208 42724
rect 20254 42712 20260 42764
rect 20312 42752 20318 42764
rect 21910 42752 21916 42764
rect 20312 42724 21036 42752
rect 20312 42712 20318 42724
rect 19383 42656 20024 42684
rect 20165 42687 20223 42693
rect 19383 42653 19395 42656
rect 19337 42647 19395 42653
rect 20165 42653 20177 42687
rect 20211 42653 20223 42687
rect 20165 42647 20223 42653
rect 20438 42644 20444 42696
rect 20496 42644 20502 42696
rect 20530 42644 20536 42696
rect 20588 42684 20594 42696
rect 21008 42693 21036 42724
rect 21192 42724 21916 42752
rect 20717 42687 20775 42693
rect 20717 42684 20729 42687
rect 20588 42656 20729 42684
rect 20588 42644 20594 42656
rect 20717 42653 20729 42656
rect 20763 42653 20775 42687
rect 20717 42647 20775 42653
rect 20993 42687 21051 42693
rect 20993 42653 21005 42687
rect 21039 42653 21051 42687
rect 20993 42647 21051 42653
rect 7006 42616 7012 42628
rect 3804 42588 5856 42616
rect 5920 42588 7012 42616
rect 1210 42508 1216 42560
rect 1268 42548 1274 42560
rect 3418 42548 3424 42560
rect 1268 42520 3424 42548
rect 1268 42508 1274 42520
rect 3418 42508 3424 42520
rect 3476 42508 3482 42560
rect 3513 42551 3571 42557
rect 3513 42517 3525 42551
rect 3559 42548 3571 42551
rect 4798 42548 4804 42560
rect 3559 42520 4804 42548
rect 3559 42517 3571 42520
rect 3513 42511 3571 42517
rect 4798 42508 4804 42520
rect 4856 42508 4862 42560
rect 5074 42508 5080 42560
rect 5132 42508 5138 42560
rect 5258 42508 5264 42560
rect 5316 42548 5322 42560
rect 5920 42548 5948 42588
rect 7006 42576 7012 42588
rect 7064 42576 7070 42628
rect 7101 42619 7159 42625
rect 7101 42585 7113 42619
rect 7147 42616 7159 42619
rect 7558 42616 7564 42628
rect 7147 42588 7564 42616
rect 7147 42585 7159 42588
rect 7101 42579 7159 42585
rect 7558 42576 7564 42588
rect 7616 42576 7622 42628
rect 8294 42576 8300 42628
rect 8352 42576 8358 42628
rect 8389 42619 8447 42625
rect 8389 42585 8401 42619
rect 8435 42616 8447 42619
rect 9214 42616 9220 42628
rect 8435 42588 9220 42616
rect 8435 42585 8447 42588
rect 8389 42579 8447 42585
rect 9214 42576 9220 42588
rect 9272 42576 9278 42628
rect 9398 42576 9404 42628
rect 9456 42576 9462 42628
rect 10778 42616 10784 42628
rect 10060 42588 10784 42616
rect 5316 42520 5948 42548
rect 5316 42508 5322 42520
rect 6454 42508 6460 42560
rect 6512 42508 6518 42560
rect 8312 42548 8340 42576
rect 10060 42557 10088 42588
rect 10778 42576 10784 42588
rect 10836 42576 10842 42628
rect 12066 42576 12072 42628
rect 12124 42616 12130 42628
rect 12124 42588 13952 42616
rect 12124 42576 12130 42588
rect 9125 42551 9183 42557
rect 9125 42548 9137 42551
rect 8312 42520 9137 42548
rect 9125 42517 9137 42520
rect 9171 42517 9183 42551
rect 9125 42511 9183 42517
rect 10045 42551 10103 42557
rect 10045 42517 10057 42551
rect 10091 42517 10103 42551
rect 10045 42511 10103 42517
rect 10134 42508 10140 42560
rect 10192 42548 10198 42560
rect 10413 42551 10471 42557
rect 10413 42548 10425 42551
rect 10192 42520 10425 42548
rect 10192 42508 10198 42520
rect 10413 42517 10425 42520
rect 10459 42517 10471 42551
rect 10413 42511 10471 42517
rect 11514 42508 11520 42560
rect 11572 42508 11578 42560
rect 11606 42508 11612 42560
rect 11664 42548 11670 42560
rect 11977 42551 12035 42557
rect 11977 42548 11989 42551
rect 11664 42520 11989 42548
rect 11664 42508 11670 42520
rect 11977 42517 11989 42520
rect 12023 42517 12035 42551
rect 11977 42511 12035 42517
rect 12434 42508 12440 42560
rect 12492 42548 12498 42560
rect 13924 42557 13952 42588
rect 16482 42576 16488 42628
rect 16540 42576 16546 42628
rect 16669 42619 16727 42625
rect 16669 42585 16681 42619
rect 16715 42616 16727 42619
rect 16715 42588 17632 42616
rect 16715 42585 16727 42588
rect 16669 42579 16727 42585
rect 12805 42551 12863 42557
rect 12805 42548 12817 42551
rect 12492 42520 12817 42548
rect 12492 42508 12498 42520
rect 12805 42517 12817 42520
rect 12851 42517 12863 42551
rect 12805 42511 12863 42517
rect 13909 42551 13967 42557
rect 13909 42517 13921 42551
rect 13955 42517 13967 42551
rect 13909 42511 13967 42517
rect 14090 42508 14096 42560
rect 14148 42548 14154 42560
rect 15289 42551 15347 42557
rect 15289 42548 15301 42551
rect 14148 42520 15301 42548
rect 14148 42508 14154 42520
rect 15289 42517 15301 42520
rect 15335 42517 15347 42551
rect 15289 42511 15347 42517
rect 16758 42508 16764 42560
rect 16816 42508 16822 42560
rect 17126 42508 17132 42560
rect 17184 42508 17190 42560
rect 17494 42508 17500 42560
rect 17552 42508 17558 42560
rect 17604 42548 17632 42588
rect 17954 42576 17960 42628
rect 18012 42576 18018 42628
rect 18064 42548 18092 42644
rect 18509 42619 18567 42625
rect 18509 42585 18521 42619
rect 18555 42616 18567 42619
rect 19426 42616 19432 42628
rect 18555 42588 19432 42616
rect 18555 42585 18567 42588
rect 18509 42579 18567 42585
rect 19426 42576 19432 42588
rect 19484 42576 19490 42628
rect 19518 42576 19524 42628
rect 19576 42576 19582 42628
rect 19705 42619 19763 42625
rect 19705 42585 19717 42619
rect 19751 42616 19763 42619
rect 20622 42616 20628 42628
rect 19751 42588 20628 42616
rect 19751 42585 19763 42588
rect 19705 42579 19763 42585
rect 20622 42576 20628 42588
rect 20680 42576 20686 42628
rect 21192 42625 21220 42724
rect 21910 42712 21916 42724
rect 21968 42712 21974 42764
rect 22002 42712 22008 42764
rect 22060 42752 22066 42764
rect 22557 42755 22615 42761
rect 22557 42752 22569 42755
rect 22060 42724 22569 42752
rect 22060 42712 22066 42724
rect 22557 42721 22569 42724
rect 22603 42721 22615 42755
rect 23014 42752 23020 42764
rect 22557 42715 22615 42721
rect 22664 42724 23020 42752
rect 22664 42684 22692 42724
rect 23014 42712 23020 42724
rect 23072 42712 23078 42764
rect 21560 42656 21864 42684
rect 21560 42625 21588 42656
rect 21177 42619 21235 42625
rect 21177 42585 21189 42619
rect 21223 42585 21235 42619
rect 21177 42579 21235 42585
rect 21545 42619 21603 42625
rect 21545 42585 21557 42619
rect 21591 42585 21603 42619
rect 21545 42579 21603 42585
rect 21729 42619 21787 42625
rect 21729 42585 21741 42619
rect 21775 42585 21787 42619
rect 21729 42579 21787 42585
rect 17604 42520 18092 42548
rect 18322 42508 18328 42560
rect 18380 42548 18386 42560
rect 18601 42551 18659 42557
rect 18601 42548 18613 42551
rect 18380 42520 18613 42548
rect 18380 42508 18386 42520
rect 18601 42517 18613 42520
rect 18647 42517 18659 42551
rect 18601 42511 18659 42517
rect 18690 42508 18696 42560
rect 18748 42548 18754 42560
rect 18969 42551 19027 42557
rect 18969 42548 18981 42551
rect 18748 42520 18981 42548
rect 18748 42508 18754 42520
rect 18969 42517 18981 42520
rect 19015 42517 19027 42551
rect 18969 42511 19027 42517
rect 19794 42508 19800 42560
rect 19852 42508 19858 42560
rect 20162 42508 20168 42560
rect 20220 42548 20226 42560
rect 20714 42548 20720 42560
rect 20220 42520 20720 42548
rect 20220 42508 20226 42520
rect 20714 42508 20720 42520
rect 20772 42508 20778 42560
rect 20806 42508 20812 42560
rect 20864 42508 20870 42560
rect 21266 42508 21272 42560
rect 21324 42548 21330 42560
rect 21744 42548 21772 42579
rect 21324 42520 21772 42548
rect 21836 42548 21864 42656
rect 22112 42656 22692 42684
rect 22833 42687 22891 42693
rect 22112 42548 22140 42656
rect 22833 42653 22845 42687
rect 22879 42684 22891 42687
rect 23474 42684 23480 42696
rect 22879 42656 23480 42684
rect 22879 42653 22891 42656
rect 22833 42647 22891 42653
rect 23474 42644 23480 42656
rect 23532 42644 23538 42696
rect 23750 42644 23756 42696
rect 23808 42684 23814 42696
rect 23937 42687 23995 42693
rect 23937 42684 23949 42687
rect 23808 42656 23949 42684
rect 23808 42644 23814 42656
rect 23937 42653 23949 42656
rect 23983 42653 23995 42687
rect 23937 42647 23995 42653
rect 22278 42576 22284 42628
rect 22336 42576 22342 42628
rect 22646 42576 22652 42628
rect 22704 42616 22710 42628
rect 23385 42619 23443 42625
rect 23385 42616 23397 42619
rect 22704 42588 23397 42616
rect 22704 42576 22710 42588
rect 23385 42585 23397 42588
rect 23431 42585 23443 42619
rect 23385 42579 23443 42585
rect 21836 42520 22140 42548
rect 21324 42508 21330 42520
rect 22186 42508 22192 42560
rect 22244 42548 22250 42560
rect 22925 42551 22983 42557
rect 22925 42548 22937 42551
rect 22244 42520 22937 42548
rect 22244 42508 22250 42520
rect 22925 42517 22937 42520
rect 22971 42517 22983 42551
rect 22925 42511 22983 42517
rect 24118 42508 24124 42560
rect 24176 42508 24182 42560
rect 1104 42458 24723 42480
rect 1104 42406 6814 42458
rect 6866 42406 6878 42458
rect 6930 42406 6942 42458
rect 6994 42406 7006 42458
rect 7058 42406 7070 42458
rect 7122 42406 12679 42458
rect 12731 42406 12743 42458
rect 12795 42406 12807 42458
rect 12859 42406 12871 42458
rect 12923 42406 12935 42458
rect 12987 42406 18544 42458
rect 18596 42406 18608 42458
rect 18660 42406 18672 42458
rect 18724 42406 18736 42458
rect 18788 42406 18800 42458
rect 18852 42406 24409 42458
rect 24461 42406 24473 42458
rect 24525 42406 24537 42458
rect 24589 42406 24601 42458
rect 24653 42406 24665 42458
rect 24717 42406 24723 42458
rect 1104 42384 24723 42406
rect 2317 42347 2375 42353
rect 2317 42313 2329 42347
rect 2363 42344 2375 42347
rect 2590 42344 2596 42356
rect 2363 42316 2596 42344
rect 2363 42313 2375 42316
rect 2317 42307 2375 42313
rect 2590 42304 2596 42316
rect 2648 42304 2654 42356
rect 3418 42304 3424 42356
rect 3476 42344 3482 42356
rect 5905 42347 5963 42353
rect 5905 42344 5917 42347
rect 3476 42316 5917 42344
rect 3476 42304 3482 42316
rect 5905 42313 5917 42316
rect 5951 42313 5963 42347
rect 5905 42307 5963 42313
rect 6641 42347 6699 42353
rect 6641 42313 6653 42347
rect 6687 42344 6699 42347
rect 7282 42344 7288 42356
rect 6687 42316 7288 42344
rect 6687 42313 6699 42316
rect 6641 42307 6699 42313
rect 7282 42304 7288 42316
rect 7340 42304 7346 42356
rect 7742 42304 7748 42356
rect 7800 42344 7806 42356
rect 7800 42316 8984 42344
rect 7800 42304 7806 42316
rect 2222 42236 2228 42288
rect 2280 42276 2286 42288
rect 2685 42279 2743 42285
rect 2280 42248 2636 42276
rect 2280 42236 2286 42248
rect 1397 42211 1455 42217
rect 1397 42177 1409 42211
rect 1443 42208 1455 42211
rect 1670 42208 1676 42220
rect 1443 42180 1676 42208
rect 1443 42177 1455 42180
rect 1397 42171 1455 42177
rect 1670 42168 1676 42180
rect 1728 42168 1734 42220
rect 2038 42168 2044 42220
rect 2096 42168 2102 42220
rect 2608 42208 2636 42248
rect 2685 42245 2697 42279
rect 2731 42276 2743 42279
rect 3142 42276 3148 42288
rect 2731 42248 3148 42276
rect 2731 42245 2743 42248
rect 2685 42239 2743 42245
rect 3142 42236 3148 42248
rect 3200 42236 3206 42288
rect 3789 42279 3847 42285
rect 3789 42245 3801 42279
rect 3835 42276 3847 42279
rect 4154 42276 4160 42288
rect 3835 42248 4160 42276
rect 3835 42245 3847 42248
rect 3789 42239 3847 42245
rect 4154 42236 4160 42248
rect 4212 42236 4218 42288
rect 4246 42236 4252 42288
rect 4304 42276 4310 42288
rect 4798 42276 4804 42288
rect 4304 42248 4804 42276
rect 4304 42236 4310 42248
rect 4798 42236 4804 42248
rect 4856 42236 4862 42288
rect 4890 42236 4896 42288
rect 4948 42276 4954 42288
rect 5166 42276 5172 42288
rect 4948 42248 5172 42276
rect 4948 42236 4954 42248
rect 5166 42236 5172 42248
rect 5224 42236 5230 42288
rect 5350 42236 5356 42288
rect 5408 42276 5414 42288
rect 8956 42276 8984 42316
rect 9122 42304 9128 42356
rect 9180 42304 9186 42356
rect 9950 42304 9956 42356
rect 10008 42304 10014 42356
rect 10229 42347 10287 42353
rect 10229 42313 10241 42347
rect 10275 42313 10287 42347
rect 10229 42307 10287 42313
rect 10244 42276 10272 42307
rect 16482 42304 16488 42356
rect 16540 42304 16546 42356
rect 16758 42304 16764 42356
rect 16816 42304 16822 42356
rect 20806 42344 20812 42356
rect 18432 42316 20812 42344
rect 16390 42276 16396 42288
rect 5408 42248 5764 42276
rect 5408 42236 5414 42248
rect 2961 42211 3019 42217
rect 2961 42208 2973 42211
rect 2608 42180 2973 42208
rect 2961 42177 2973 42180
rect 3007 42177 3019 42211
rect 2961 42171 3019 42177
rect 3050 42168 3056 42220
rect 3108 42168 3114 42220
rect 3421 42211 3479 42217
rect 3421 42177 3433 42211
rect 3467 42208 3479 42211
rect 4338 42208 4344 42220
rect 3467 42180 4344 42208
rect 3467 42177 3479 42180
rect 3421 42171 3479 42177
rect 4338 42168 4344 42180
rect 4396 42168 4402 42220
rect 4431 42211 4489 42217
rect 4431 42177 4443 42211
rect 4477 42208 4489 42211
rect 5442 42208 5448 42220
rect 4477 42180 5448 42208
rect 4477 42177 4489 42180
rect 4431 42171 4489 42177
rect 5442 42168 5448 42180
rect 5500 42168 5506 42220
rect 2504 42152 2556 42158
rect 1578 42100 1584 42152
rect 1636 42100 1642 42152
rect 3878 42100 3884 42152
rect 3936 42140 3942 42152
rect 4157 42143 4215 42149
rect 4157 42140 4169 42143
rect 3936 42112 4169 42140
rect 3936 42100 3942 42112
rect 4157 42109 4169 42112
rect 4203 42109 4215 42143
rect 5736 42140 5764 42248
rect 6472 42248 8892 42276
rect 8956 42248 10272 42276
rect 12406 42248 16396 42276
rect 5813 42211 5871 42217
rect 5813 42177 5825 42211
rect 5859 42208 5871 42211
rect 6362 42208 6368 42220
rect 5859 42180 6368 42208
rect 5859 42177 5871 42180
rect 5813 42171 5871 42177
rect 6362 42168 6368 42180
rect 6420 42168 6426 42220
rect 6472 42217 6500 42248
rect 6457 42211 6515 42217
rect 6457 42177 6469 42211
rect 6503 42177 6515 42211
rect 6457 42171 6515 42177
rect 7099 42211 7157 42217
rect 7099 42177 7111 42211
rect 7145 42208 7157 42211
rect 7466 42208 7472 42220
rect 7145 42180 7472 42208
rect 7145 42177 7157 42180
rect 7099 42171 7157 42177
rect 7466 42168 7472 42180
rect 7524 42168 7530 42220
rect 8294 42168 8300 42220
rect 8352 42168 8358 42220
rect 6822 42140 6828 42152
rect 5736 42112 6828 42140
rect 4157 42103 4215 42109
rect 6822 42100 6828 42112
rect 6880 42100 6886 42152
rect 7558 42100 7564 42152
rect 7616 42140 7622 42152
rect 7616 42112 8800 42140
rect 7616 42100 7622 42112
rect 2504 42094 2556 42100
rect 6638 42072 6644 42084
rect 4816 42044 6644 42072
rect 3973 42007 4031 42013
rect 3973 41973 3985 42007
rect 4019 42004 4031 42007
rect 4430 42004 4436 42016
rect 4019 41976 4436 42004
rect 4019 41973 4031 41976
rect 3973 41967 4031 41973
rect 4430 41964 4436 41976
rect 4488 41964 4494 42016
rect 4614 41964 4620 42016
rect 4672 42004 4678 42016
rect 4816 42004 4844 42044
rect 6638 42032 6644 42044
rect 6696 42032 6702 42084
rect 4672 41976 4844 42004
rect 4672 41964 4678 41976
rect 5166 41964 5172 42016
rect 5224 41964 5230 42016
rect 5442 41964 5448 42016
rect 5500 42004 5506 42016
rect 6914 42004 6920 42016
rect 5500 41976 6920 42004
rect 5500 41964 5506 41976
rect 6914 41964 6920 41976
rect 6972 42004 6978 42016
rect 7650 42004 7656 42016
rect 6972 41976 7656 42004
rect 6972 41964 6978 41976
rect 7650 41964 7656 41976
rect 7708 41964 7714 42016
rect 7834 41964 7840 42016
rect 7892 41964 7898 42016
rect 7926 41964 7932 42016
rect 7984 42004 7990 42016
rect 8389 42007 8447 42013
rect 8389 42004 8401 42007
rect 7984 41976 8401 42004
rect 7984 41964 7990 41976
rect 8389 41973 8401 41976
rect 8435 41973 8447 42007
rect 8772 42004 8800 42112
rect 8864 42081 8892 42248
rect 9030 42168 9036 42220
rect 9088 42168 9094 42220
rect 9306 42168 9312 42220
rect 9364 42168 9370 42220
rect 9677 42211 9735 42217
rect 9677 42177 9689 42211
rect 9723 42208 9735 42211
rect 10134 42208 10140 42220
rect 9723 42180 10140 42208
rect 9723 42177 9735 42180
rect 9677 42171 9735 42177
rect 10134 42168 10140 42180
rect 10192 42168 10198 42220
rect 10410 42168 10416 42220
rect 10468 42168 10474 42220
rect 8849 42075 8907 42081
rect 8849 42041 8861 42075
rect 8895 42041 8907 42075
rect 8849 42035 8907 42041
rect 12406 42004 12434 42248
rect 16390 42236 16396 42248
rect 16448 42236 16454 42288
rect 16500 42072 16528 42304
rect 16776 42140 16804 42304
rect 18432 42285 18460 42316
rect 20806 42304 20812 42316
rect 20864 42304 20870 42356
rect 21082 42304 21088 42356
rect 21140 42344 21146 42356
rect 21545 42347 21603 42353
rect 21545 42344 21557 42347
rect 21140 42316 21557 42344
rect 21140 42304 21146 42316
rect 21545 42313 21557 42316
rect 21591 42313 21603 42347
rect 21545 42307 21603 42313
rect 22281 42347 22339 42353
rect 22281 42313 22293 42347
rect 22327 42344 22339 42347
rect 22738 42344 22744 42356
rect 22327 42316 22744 42344
rect 22327 42313 22339 42316
rect 22281 42307 22339 42313
rect 22738 42304 22744 42316
rect 22796 42304 22802 42356
rect 22833 42347 22891 42353
rect 22833 42313 22845 42347
rect 22879 42344 22891 42347
rect 22922 42344 22928 42356
rect 22879 42316 22928 42344
rect 22879 42313 22891 42316
rect 22833 42307 22891 42313
rect 22922 42304 22928 42316
rect 22980 42304 22986 42356
rect 23937 42347 23995 42353
rect 23937 42313 23949 42347
rect 23983 42344 23995 42347
rect 24854 42344 24860 42356
rect 23983 42316 24860 42344
rect 23983 42313 23995 42316
rect 23937 42307 23995 42313
rect 24854 42304 24860 42316
rect 24912 42304 24918 42356
rect 18417 42279 18475 42285
rect 18417 42245 18429 42279
rect 18463 42245 18475 42279
rect 18417 42239 18475 42245
rect 20162 42236 20168 42288
rect 20220 42276 20226 42288
rect 20441 42279 20499 42285
rect 20441 42276 20453 42279
rect 20220 42248 20453 42276
rect 20220 42236 20226 42248
rect 20441 42245 20453 42248
rect 20487 42245 20499 42279
rect 20441 42239 20499 42245
rect 23477 42279 23535 42285
rect 23477 42245 23489 42279
rect 23523 42276 23535 42279
rect 24026 42276 24032 42288
rect 23523 42248 24032 42276
rect 23523 42245 23535 42248
rect 23477 42239 23535 42245
rect 24026 42236 24032 42248
rect 24084 42236 24090 42288
rect 18690 42168 18696 42220
rect 18748 42168 18754 42220
rect 19058 42168 19064 42220
rect 19116 42208 19122 42220
rect 20254 42208 20260 42220
rect 19116 42180 20260 42208
rect 19116 42168 19122 42180
rect 20254 42168 20260 42180
rect 20312 42168 20318 42220
rect 20717 42211 20775 42217
rect 20717 42208 20729 42211
rect 20456 42180 20729 42208
rect 20162 42140 20168 42152
rect 16776 42112 20168 42140
rect 20162 42100 20168 42112
rect 20220 42100 20226 42152
rect 16500 42044 19288 42072
rect 8772 41976 12434 42004
rect 8389 41967 8447 41973
rect 18506 41964 18512 42016
rect 18564 41964 18570 42016
rect 19260 42004 19288 42044
rect 19334 42032 19340 42084
rect 19392 42072 19398 42084
rect 20456 42072 20484 42180
rect 20717 42177 20729 42180
rect 20763 42177 20775 42211
rect 20717 42171 20775 42177
rect 20990 42168 20996 42220
rect 21048 42168 21054 42220
rect 21082 42168 21088 42220
rect 21140 42208 21146 42220
rect 21269 42211 21327 42217
rect 21269 42208 21281 42211
rect 21140 42180 21281 42208
rect 21140 42168 21146 42180
rect 21269 42177 21281 42180
rect 21315 42177 21327 42211
rect 21269 42171 21327 42177
rect 21358 42168 21364 42220
rect 21416 42168 21422 42220
rect 22005 42211 22063 42217
rect 22005 42177 22017 42211
rect 22051 42177 22063 42211
rect 22005 42171 22063 42177
rect 20622 42140 20628 42152
rect 20548 42112 20628 42140
rect 20548 42081 20576 42112
rect 20622 42100 20628 42112
rect 20680 42100 20686 42152
rect 22020 42140 22048 42171
rect 22554 42168 22560 42220
rect 22612 42168 22618 42220
rect 23106 42168 23112 42220
rect 23164 42168 23170 42220
rect 23566 42168 23572 42220
rect 23624 42208 23630 42220
rect 23661 42211 23719 42217
rect 23661 42208 23673 42211
rect 23624 42180 23673 42208
rect 23624 42168 23630 42180
rect 23661 42177 23673 42180
rect 23707 42177 23719 42211
rect 23661 42171 23719 42177
rect 22922 42140 22928 42152
rect 22020 42112 22928 42140
rect 22922 42100 22928 42112
rect 22980 42100 22986 42152
rect 19392 42044 20484 42072
rect 20533 42075 20591 42081
rect 19392 42032 19398 42044
rect 20533 42041 20545 42075
rect 20579 42041 20591 42075
rect 20533 42035 20591 42041
rect 20254 42004 20260 42016
rect 19260 41976 20260 42004
rect 20254 41964 20260 41976
rect 20312 41964 20318 42016
rect 20809 42007 20867 42013
rect 20809 41973 20821 42007
rect 20855 42004 20867 42007
rect 20898 42004 20904 42016
rect 20855 41976 20904 42004
rect 20855 41973 20867 41976
rect 20809 41967 20867 41973
rect 20898 41964 20904 41976
rect 20956 41964 20962 42016
rect 21085 42007 21143 42013
rect 21085 41973 21097 42007
rect 21131 42004 21143 42007
rect 21450 42004 21456 42016
rect 21131 41976 21456 42004
rect 21131 41973 21143 41976
rect 21085 41967 21143 41973
rect 21450 41964 21456 41976
rect 21508 41964 21514 42016
rect 1104 41914 24564 41936
rect 1104 41862 3882 41914
rect 3934 41862 3946 41914
rect 3998 41862 4010 41914
rect 4062 41862 4074 41914
rect 4126 41862 4138 41914
rect 4190 41862 9747 41914
rect 9799 41862 9811 41914
rect 9863 41862 9875 41914
rect 9927 41862 9939 41914
rect 9991 41862 10003 41914
rect 10055 41862 15612 41914
rect 15664 41862 15676 41914
rect 15728 41862 15740 41914
rect 15792 41862 15804 41914
rect 15856 41862 15868 41914
rect 15920 41862 21477 41914
rect 21529 41862 21541 41914
rect 21593 41862 21605 41914
rect 21657 41862 21669 41914
rect 21721 41862 21733 41914
rect 21785 41862 24564 41914
rect 1104 41840 24564 41862
rect 2332 41772 3004 41800
rect 2332 41673 2360 41772
rect 2976 41732 3004 41772
rect 3050 41760 3056 41812
rect 3108 41800 3114 41812
rect 3329 41803 3387 41809
rect 3329 41800 3341 41803
rect 3108 41772 3341 41800
rect 3108 41760 3114 41772
rect 3329 41769 3341 41772
rect 3375 41769 3387 41803
rect 3329 41763 3387 41769
rect 4065 41803 4123 41809
rect 4065 41769 4077 41803
rect 4111 41800 4123 41803
rect 4890 41800 4896 41812
rect 4111 41772 4896 41800
rect 4111 41769 4123 41772
rect 4065 41763 4123 41769
rect 4890 41760 4896 41772
rect 4948 41760 4954 41812
rect 6454 41760 6460 41812
rect 6512 41760 6518 41812
rect 6546 41760 6552 41812
rect 6604 41800 6610 41812
rect 7285 41803 7343 41809
rect 7285 41800 7297 41803
rect 6604 41772 7297 41800
rect 6604 41760 6610 41772
rect 7285 41769 7297 41772
rect 7331 41769 7343 41803
rect 7285 41763 7343 41769
rect 7392 41772 8156 41800
rect 3234 41732 3240 41744
rect 2976 41704 3240 41732
rect 3234 41692 3240 41704
rect 3292 41692 3298 41744
rect 3418 41692 3424 41744
rect 3476 41732 3482 41744
rect 4614 41732 4620 41744
rect 3476 41704 4620 41732
rect 3476 41692 3482 41704
rect 4614 41692 4620 41704
rect 4672 41692 4678 41744
rect 6472 41732 6500 41760
rect 6196 41704 6500 41732
rect 5080 41676 5132 41682
rect 2317 41667 2375 41673
rect 2317 41633 2329 41667
rect 2363 41633 2375 41667
rect 2317 41627 2375 41633
rect 3142 41624 3148 41676
rect 3200 41664 3206 41676
rect 4706 41664 4712 41676
rect 3200 41636 4712 41664
rect 3200 41624 3206 41636
rect 4706 41624 4712 41636
rect 4764 41624 4770 41676
rect 4798 41624 4804 41676
rect 4856 41624 4862 41676
rect 1394 41556 1400 41608
rect 1452 41556 1458 41608
rect 1765 41599 1823 41605
rect 1765 41565 1777 41599
rect 1811 41596 1823 41599
rect 1811 41568 2268 41596
rect 1811 41565 1823 41568
rect 1765 41559 1823 41565
rect 2038 41488 2044 41540
rect 2096 41488 2102 41540
rect 2240 41528 2268 41568
rect 2498 41556 2504 41608
rect 2556 41596 2562 41608
rect 2591 41599 2649 41605
rect 2591 41596 2603 41599
rect 2556 41568 2603 41596
rect 2556 41556 2562 41568
rect 2591 41565 2603 41568
rect 2637 41565 2649 41599
rect 2591 41559 2649 41565
rect 3881 41599 3939 41605
rect 3881 41565 3893 41599
rect 3927 41596 3939 41599
rect 4525 41599 4583 41605
rect 4525 41596 4537 41599
rect 3927 41568 4537 41596
rect 3927 41565 3939 41568
rect 3881 41559 3939 41565
rect 4525 41565 4537 41568
rect 4571 41596 4583 41599
rect 4816 41596 4844 41624
rect 5080 41618 5132 41624
rect 4571 41568 4844 41596
rect 5433 41599 5491 41605
rect 4571 41565 4583 41568
rect 4525 41559 4583 41565
rect 5433 41565 5445 41599
rect 5479 41596 5491 41599
rect 6196 41596 6224 41704
rect 6730 41692 6736 41744
rect 6788 41732 6794 41744
rect 7392 41732 7420 41772
rect 6788 41704 7420 41732
rect 8128 41732 8156 41772
rect 8938 41760 8944 41812
rect 8996 41760 9002 41812
rect 9214 41760 9220 41812
rect 9272 41760 9278 41812
rect 15194 41760 15200 41812
rect 15252 41800 15258 41812
rect 19334 41800 19340 41812
rect 15252 41772 19340 41800
rect 15252 41760 15258 41772
rect 19334 41760 19340 41772
rect 19392 41760 19398 41812
rect 19889 41803 19947 41809
rect 19889 41769 19901 41803
rect 19935 41800 19947 41803
rect 20438 41800 20444 41812
rect 19935 41772 20444 41800
rect 19935 41769 19947 41772
rect 19889 41763 19947 41769
rect 20438 41760 20444 41772
rect 20496 41760 20502 41812
rect 20625 41803 20683 41809
rect 20625 41769 20637 41803
rect 20671 41769 20683 41803
rect 20625 41763 20683 41769
rect 21177 41803 21235 41809
rect 21177 41769 21189 41803
rect 21223 41800 21235 41803
rect 21266 41800 21272 41812
rect 21223 41772 21272 41800
rect 21223 41769 21235 41772
rect 21177 41763 21235 41769
rect 8128 41704 9536 41732
rect 6788 41692 6794 41704
rect 6362 41624 6368 41676
rect 6420 41624 6426 41676
rect 6822 41624 6828 41676
rect 6880 41664 6886 41676
rect 7469 41667 7527 41673
rect 7469 41664 7481 41667
rect 6880 41636 7481 41664
rect 6880 41624 6886 41636
rect 7469 41633 7481 41636
rect 7515 41633 7527 41667
rect 9508 41664 9536 41704
rect 10226 41692 10232 41744
rect 10284 41732 10290 41744
rect 10284 41704 19932 41732
rect 10284 41692 10290 41704
rect 13906 41664 13912 41676
rect 9508 41636 13912 41664
rect 7469 41627 7527 41633
rect 13906 41624 13912 41636
rect 13964 41624 13970 41676
rect 5479 41568 6224 41596
rect 6380 41596 6408 41624
rect 6380 41568 7052 41596
rect 5479 41565 5491 41568
rect 5433 41559 5491 41565
rect 2774 41528 2780 41540
rect 2240 41500 2780 41528
rect 2774 41488 2780 41500
rect 2832 41488 2838 41540
rect 2958 41488 2964 41540
rect 3016 41528 3022 41540
rect 3510 41528 3516 41540
rect 3016 41500 3516 41528
rect 3016 41488 3022 41500
rect 3510 41488 3516 41500
rect 3568 41488 3574 41540
rect 4706 41488 4712 41540
rect 4764 41528 4770 41540
rect 5077 41531 5135 41537
rect 5077 41528 5089 41531
rect 4764 41500 5089 41528
rect 4764 41488 4770 41500
rect 5077 41497 5089 41500
rect 5123 41528 5135 41531
rect 5258 41528 5264 41540
rect 5123 41500 5264 41528
rect 5123 41497 5135 41500
rect 5077 41491 5135 41497
rect 5258 41488 5264 41500
rect 5316 41488 5322 41540
rect 5353 41531 5411 41537
rect 5353 41497 5365 41531
rect 5399 41528 5411 41531
rect 5399 41500 5476 41528
rect 5399 41497 5411 41500
rect 5353 41491 5411 41497
rect 5448 41472 5476 41500
rect 5534 41488 5540 41540
rect 5592 41528 5598 41540
rect 5813 41531 5871 41537
rect 5813 41528 5825 41531
rect 5592 41500 5825 41528
rect 5592 41488 5598 41500
rect 5813 41497 5825 41500
rect 5859 41497 5871 41531
rect 5813 41491 5871 41497
rect 5902 41488 5908 41540
rect 5960 41528 5966 41540
rect 5960 41500 6500 41528
rect 5960 41488 5966 41500
rect 1581 41463 1639 41469
rect 1581 41429 1593 41463
rect 1627 41460 1639 41463
rect 4982 41460 4988 41472
rect 1627 41432 4988 41460
rect 1627 41429 1639 41432
rect 1581 41423 1639 41429
rect 4982 41420 4988 41432
rect 5040 41420 5046 41472
rect 5442 41420 5448 41472
rect 5500 41420 5506 41472
rect 5626 41420 5632 41472
rect 5684 41460 5690 41472
rect 6181 41463 6239 41469
rect 6181 41460 6193 41463
rect 5684 41432 6193 41460
rect 5684 41420 5690 41432
rect 6181 41429 6193 41432
rect 6227 41429 6239 41463
rect 6181 41423 6239 41429
rect 6362 41420 6368 41472
rect 6420 41420 6426 41472
rect 6472 41460 6500 41500
rect 6638 41488 6644 41540
rect 6696 41488 6702 41540
rect 6733 41463 6791 41469
rect 6733 41460 6745 41463
rect 6472 41432 6745 41460
rect 6733 41429 6745 41432
rect 6779 41429 6791 41463
rect 7024 41460 7052 41568
rect 7098 41556 7104 41608
rect 7156 41556 7162 41608
rect 7650 41556 7656 41608
rect 7708 41596 7714 41608
rect 7743 41599 7801 41605
rect 7743 41596 7755 41599
rect 7708 41568 7755 41596
rect 7708 41556 7714 41568
rect 7743 41565 7755 41568
rect 7789 41565 7801 41599
rect 7743 41559 7801 41565
rect 9122 41556 9128 41608
rect 9180 41556 9186 41608
rect 9214 41556 9220 41608
rect 9272 41596 9278 41608
rect 9401 41599 9459 41605
rect 9401 41596 9413 41599
rect 9272 41568 9413 41596
rect 9272 41556 9278 41568
rect 9401 41565 9413 41568
rect 9447 41565 9459 41599
rect 9401 41559 9459 41565
rect 13814 41556 13820 41608
rect 13872 41596 13878 41608
rect 19426 41596 19432 41608
rect 13872 41568 19432 41596
rect 13872 41556 13878 41568
rect 19426 41556 19432 41568
rect 19484 41556 19490 41608
rect 19797 41599 19855 41605
rect 19797 41596 19809 41599
rect 19720 41568 19809 41596
rect 10962 41528 10968 41540
rect 7785 41500 10968 41528
rect 7785 41460 7813 41500
rect 10962 41488 10968 41500
rect 11020 41488 11026 41540
rect 19334 41488 19340 41540
rect 19392 41488 19398 41540
rect 7024 41432 7813 41460
rect 6733 41423 6791 41429
rect 8478 41420 8484 41472
rect 8536 41420 8542 41472
rect 19426 41420 19432 41472
rect 19484 41420 19490 41472
rect 19610 41420 19616 41472
rect 19668 41420 19674 41472
rect 19720 41460 19748 41568
rect 19797 41565 19809 41568
rect 19843 41565 19855 41599
rect 19904 41596 19932 41704
rect 20070 41692 20076 41744
rect 20128 41732 20134 41744
rect 20128 41704 20300 41732
rect 20128 41692 20134 41704
rect 20272 41664 20300 41704
rect 20346 41692 20352 41744
rect 20404 41692 20410 41744
rect 20640 41664 20668 41763
rect 21266 41760 21272 41772
rect 21324 41760 21330 41812
rect 21729 41803 21787 41809
rect 21729 41769 21741 41803
rect 21775 41800 21787 41803
rect 22554 41800 22560 41812
rect 21775 41772 22560 41800
rect 21775 41769 21787 41772
rect 21729 41763 21787 41769
rect 22554 41760 22560 41772
rect 22612 41760 22618 41812
rect 23290 41760 23296 41812
rect 23348 41760 23354 41812
rect 23934 41760 23940 41812
rect 23992 41760 23998 41812
rect 24302 41760 24308 41812
rect 24360 41760 24366 41812
rect 21453 41735 21511 41741
rect 21453 41701 21465 41735
rect 21499 41732 21511 41735
rect 22370 41732 22376 41744
rect 21499 41704 22376 41732
rect 21499 41701 21511 41704
rect 21453 41695 21511 41701
rect 22370 41692 22376 41704
rect 22428 41692 22434 41744
rect 22465 41735 22523 41741
rect 22465 41701 22477 41735
rect 22511 41732 22523 41735
rect 23308 41732 23336 41760
rect 22511 41704 23336 41732
rect 23569 41735 23627 41741
rect 22511 41701 22523 41704
rect 22465 41695 22523 41701
rect 23569 41701 23581 41735
rect 23615 41732 23627 41735
rect 24320 41732 24348 41760
rect 23615 41704 24348 41732
rect 23615 41701 23627 41704
rect 23569 41695 23627 41701
rect 20272 41636 20668 41664
rect 20898 41624 20904 41676
rect 20956 41624 20962 41676
rect 25130 41664 25136 41676
rect 21192 41636 25136 41664
rect 20073 41599 20131 41605
rect 20073 41596 20085 41599
rect 19904 41568 20085 41596
rect 19797 41559 19855 41565
rect 20073 41565 20085 41568
rect 20119 41565 20131 41599
rect 20073 41559 20131 41565
rect 20530 41556 20536 41608
rect 20588 41556 20594 41608
rect 20809 41599 20867 41605
rect 20809 41565 20821 41599
rect 20855 41596 20867 41599
rect 20916 41596 20944 41624
rect 20855 41568 20944 41596
rect 21085 41599 21143 41605
rect 20855 41565 20867 41568
rect 20809 41559 20867 41565
rect 21085 41565 21097 41599
rect 21131 41592 21143 41599
rect 21192 41592 21220 41636
rect 25130 41624 25136 41636
rect 25188 41624 25194 41676
rect 21131 41565 21220 41592
rect 21085 41564 21220 41565
rect 21085 41559 21143 41564
rect 21266 41556 21272 41608
rect 21324 41596 21330 41608
rect 21361 41599 21419 41605
rect 21361 41596 21373 41599
rect 21324 41568 21373 41596
rect 21324 41556 21330 41568
rect 21361 41565 21373 41568
rect 21407 41565 21419 41599
rect 21361 41559 21419 41565
rect 21634 41556 21640 41608
rect 21692 41556 21698 41608
rect 21818 41556 21824 41608
rect 21876 41596 21882 41608
rect 21913 41599 21971 41605
rect 21913 41596 21925 41599
rect 21876 41568 21925 41596
rect 21876 41556 21882 41568
rect 21913 41565 21925 41568
rect 21959 41565 21971 41599
rect 21913 41559 21971 41565
rect 23109 41599 23167 41605
rect 23109 41565 23121 41599
rect 23155 41596 23167 41599
rect 24946 41596 24952 41608
rect 23155 41568 24952 41596
rect 23155 41565 23167 41568
rect 23109 41559 23167 41565
rect 24946 41556 24952 41568
rect 25004 41556 25010 41608
rect 22094 41528 22100 41540
rect 20916 41500 22100 41528
rect 20622 41460 20628 41472
rect 19720 41432 20628 41460
rect 20622 41420 20628 41432
rect 20680 41420 20686 41472
rect 20916 41469 20944 41500
rect 22094 41488 22100 41500
rect 22152 41488 22158 41540
rect 22186 41488 22192 41540
rect 22244 41488 22250 41540
rect 22741 41531 22799 41537
rect 22741 41497 22753 41531
rect 22787 41497 22799 41531
rect 22741 41491 22799 41497
rect 20901 41463 20959 41469
rect 20901 41429 20913 41463
rect 20947 41429 20959 41463
rect 20901 41423 20959 41429
rect 21542 41420 21548 41472
rect 21600 41460 21606 41472
rect 22370 41460 22376 41472
rect 21600 41432 22376 41460
rect 21600 41420 21606 41432
rect 22370 41420 22376 41432
rect 22428 41420 22434 41472
rect 22756 41460 22784 41491
rect 23290 41488 23296 41540
rect 23348 41488 23354 41540
rect 23842 41488 23848 41540
rect 23900 41488 23906 41540
rect 24026 41460 24032 41472
rect 22756 41432 24032 41460
rect 24026 41420 24032 41432
rect 24084 41420 24090 41472
rect 1104 41370 24723 41392
rect 1104 41318 6814 41370
rect 6866 41318 6878 41370
rect 6930 41318 6942 41370
rect 6994 41318 7006 41370
rect 7058 41318 7070 41370
rect 7122 41318 12679 41370
rect 12731 41318 12743 41370
rect 12795 41318 12807 41370
rect 12859 41318 12871 41370
rect 12923 41318 12935 41370
rect 12987 41318 18544 41370
rect 18596 41318 18608 41370
rect 18660 41318 18672 41370
rect 18724 41318 18736 41370
rect 18788 41318 18800 41370
rect 18852 41318 24409 41370
rect 24461 41318 24473 41370
rect 24525 41318 24537 41370
rect 24589 41318 24601 41370
rect 24653 41318 24665 41370
rect 24717 41318 24723 41370
rect 1104 41296 24723 41318
rect 2777 41259 2835 41265
rect 2777 41225 2789 41259
rect 2823 41256 2835 41259
rect 3694 41256 3700 41268
rect 2823 41228 3700 41256
rect 2823 41225 2835 41228
rect 2777 41219 2835 41225
rect 3694 41216 3700 41228
rect 3752 41216 3758 41268
rect 4430 41256 4436 41268
rect 3804 41228 4436 41256
rect 2406 41148 2412 41200
rect 2464 41188 2470 41200
rect 3804 41188 3832 41228
rect 4430 41216 4436 41228
rect 4488 41216 4494 41268
rect 4525 41259 4583 41265
rect 4525 41225 4537 41259
rect 4571 41256 4583 41259
rect 4706 41256 4712 41268
rect 4571 41228 4712 41256
rect 4571 41225 4583 41228
rect 4525 41219 4583 41225
rect 4706 41216 4712 41228
rect 4764 41216 4770 41268
rect 5813 41259 5871 41265
rect 5813 41256 5825 41259
rect 4816 41228 5825 41256
rect 2464 41160 3832 41188
rect 2464 41148 2470 41160
rect 4338 41148 4344 41200
rect 4396 41188 4402 41200
rect 4816 41188 4844 41228
rect 5813 41225 5825 41228
rect 5859 41225 5871 41259
rect 5813 41219 5871 41225
rect 4396 41160 4844 41188
rect 4893 41191 4951 41197
rect 4396 41148 4402 41160
rect 4893 41157 4905 41191
rect 4939 41188 4951 41191
rect 5166 41188 5172 41200
rect 4939 41160 5172 41188
rect 4939 41157 4951 41160
rect 4893 41151 4951 41157
rect 5166 41148 5172 41160
rect 5224 41148 5230 41200
rect 5261 41191 5319 41197
rect 5261 41157 5273 41191
rect 5307 41188 5319 41191
rect 5534 41188 5540 41200
rect 5307 41160 5540 41188
rect 5307 41157 5319 41160
rect 5261 41151 5319 41157
rect 5534 41148 5540 41160
rect 5592 41148 5598 41200
rect 5626 41148 5632 41200
rect 5684 41148 5690 41200
rect 5828 41188 5856 41219
rect 5994 41216 6000 41268
rect 6052 41216 6058 41268
rect 7650 41256 7656 41268
rect 7208 41228 7656 41256
rect 7208 41188 7236 41228
rect 7650 41216 7656 41228
rect 7708 41216 7714 41268
rect 8665 41259 8723 41265
rect 8665 41225 8677 41259
rect 8711 41225 8723 41259
rect 8665 41219 8723 41225
rect 20349 41259 20407 41265
rect 20349 41225 20361 41259
rect 20395 41256 20407 41259
rect 20901 41259 20959 41265
rect 20395 41228 20852 41256
rect 20395 41225 20407 41228
rect 20349 41219 20407 41225
rect 5828 41160 7236 41188
rect 7300 41160 7512 41188
rect 1394 41080 1400 41132
rect 1452 41080 1458 41132
rect 2498 41080 2504 41132
rect 2556 41080 2562 41132
rect 3235 41123 3293 41129
rect 3235 41089 3247 41123
rect 3281 41120 3293 41123
rect 4430 41120 4436 41132
rect 3281 41092 4436 41120
rect 3281 41089 3293 41092
rect 3235 41083 3293 41089
rect 4430 41080 4436 41092
rect 4488 41080 4494 41132
rect 4801 41123 4859 41129
rect 4801 41089 4813 41123
rect 4847 41120 4859 41123
rect 5074 41120 5080 41132
rect 4847 41092 5080 41120
rect 4847 41089 4859 41092
rect 4801 41083 4859 41089
rect 5074 41080 5080 41092
rect 5132 41120 5138 41132
rect 5442 41120 5448 41132
rect 5132 41092 5448 41120
rect 5132 41080 5138 41092
rect 5442 41080 5448 41092
rect 5500 41080 5506 41132
rect 842 41012 848 41064
rect 900 41052 906 41064
rect 2133 41055 2191 41061
rect 2133 41052 2145 41055
rect 900 41024 2145 41052
rect 900 41012 906 41024
rect 2133 41021 2145 41024
rect 2179 41052 2191 41055
rect 2314 41052 2320 41064
rect 2179 41024 2320 41052
rect 2179 41021 2191 41024
rect 2133 41015 2191 41021
rect 2314 41012 2320 41024
rect 2372 41012 2378 41064
rect 2958 41012 2964 41064
rect 3016 41012 3022 41064
rect 3973 40987 4031 40993
rect 3973 40953 3985 40987
rect 4019 40984 4031 40987
rect 4356 40984 4384 41038
rect 4019 40956 4384 40984
rect 5644 40984 5672 41148
rect 5810 41080 5816 41132
rect 5868 41120 5874 41132
rect 7300 41129 7328 41160
rect 6181 41123 6239 41129
rect 6181 41120 6193 41123
rect 5868 41092 6193 41120
rect 5868 41080 5874 41092
rect 6181 41089 6193 41092
rect 6227 41089 6239 41123
rect 6181 41083 6239 41089
rect 6457 41123 6515 41129
rect 6457 41089 6469 41123
rect 6503 41089 6515 41123
rect 6457 41083 6515 41089
rect 7285 41123 7343 41129
rect 7285 41089 7297 41123
rect 7331 41089 7343 41123
rect 7484 41120 7512 41160
rect 7558 41148 7564 41200
rect 7616 41148 7622 41200
rect 7929 41191 7987 41197
rect 7929 41157 7941 41191
rect 7975 41188 7987 41191
rect 8478 41188 8484 41200
rect 7975 41160 8484 41188
rect 7975 41157 7987 41160
rect 7929 41151 7987 41157
rect 8478 41148 8484 41160
rect 8536 41148 8542 41200
rect 8680 41132 8708 41219
rect 13906 41148 13912 41200
rect 13964 41188 13970 41200
rect 20824 41188 20852 41228
rect 20901 41225 20913 41259
rect 20947 41256 20959 41259
rect 21082 41256 21088 41268
rect 20947 41228 21088 41256
rect 20947 41225 20959 41228
rect 20901 41219 20959 41225
rect 21082 41216 21088 41228
rect 21140 41216 21146 41268
rect 21177 41259 21235 41265
rect 21177 41225 21189 41259
rect 21223 41225 21235 41259
rect 21177 41219 21235 41225
rect 21453 41259 21511 41265
rect 21453 41225 21465 41259
rect 21499 41256 21511 41259
rect 22186 41256 22192 41268
rect 21499 41228 22192 41256
rect 21499 41225 21511 41228
rect 21453 41219 21511 41225
rect 20990 41188 20996 41200
rect 13964 41160 19380 41188
rect 20824 41160 20996 41188
rect 13964 41148 13970 41160
rect 7837 41123 7895 41129
rect 7837 41120 7849 41123
rect 7484 41092 7849 41120
rect 7285 41083 7343 41089
rect 7837 41089 7849 41092
rect 7883 41089 7895 41123
rect 7837 41083 7895 41089
rect 5718 41012 5724 41064
rect 5776 41052 5782 41064
rect 6472 41052 6500 41083
rect 8110 41080 8116 41132
rect 8168 41120 8174 41132
rect 8297 41123 8355 41129
rect 8297 41120 8309 41123
rect 8168 41092 8309 41120
rect 8168 41080 8174 41092
rect 8297 41089 8309 41092
rect 8343 41089 8355 41123
rect 8297 41083 8355 41089
rect 8662 41080 8668 41132
rect 8720 41080 8726 41132
rect 19242 41080 19248 41132
rect 19300 41080 19306 41132
rect 19352 41120 19380 41160
rect 20990 41148 20996 41160
rect 21048 41148 21054 41200
rect 21192 41188 21220 41219
rect 22186 41216 22192 41228
rect 22244 41216 22250 41268
rect 22281 41259 22339 41265
rect 22281 41225 22293 41259
rect 22327 41256 22339 41259
rect 22646 41256 22652 41268
rect 22327 41228 22652 41256
rect 22327 41225 22339 41228
rect 22281 41219 22339 41225
rect 22646 41216 22652 41228
rect 22704 41216 22710 41268
rect 23106 41216 23112 41268
rect 23164 41216 23170 41268
rect 23382 41216 23388 41268
rect 23440 41216 23446 41268
rect 23474 41216 23480 41268
rect 23532 41256 23538 41268
rect 23842 41256 23848 41268
rect 23532 41228 23848 41256
rect 23532 41216 23538 41228
rect 23842 41216 23848 41228
rect 23900 41216 23906 41268
rect 23937 41259 23995 41265
rect 23937 41225 23949 41259
rect 23983 41256 23995 41259
rect 24762 41256 24768 41268
rect 23983 41228 24768 41256
rect 23983 41225 23995 41228
rect 23937 41219 23995 41225
rect 24762 41216 24768 41228
rect 24820 41216 24826 41268
rect 23124 41188 23152 41216
rect 21192 41160 23152 41188
rect 20533 41123 20591 41129
rect 20533 41120 20545 41123
rect 19352 41092 20545 41120
rect 20533 41089 20545 41092
rect 20579 41089 20591 41123
rect 20809 41123 20867 41129
rect 20809 41120 20821 41123
rect 20533 41083 20591 41089
rect 20640 41092 20821 41120
rect 5776 41024 6500 41052
rect 5776 41012 5782 41024
rect 7742 41012 7748 41064
rect 7800 41012 7806 41064
rect 16206 41012 16212 41064
rect 16264 41052 16270 41064
rect 20640 41052 20668 41092
rect 20809 41089 20821 41092
rect 20855 41089 20867 41123
rect 21085 41123 21143 41129
rect 21085 41120 21097 41123
rect 20809 41083 20867 41089
rect 20916 41092 21097 41120
rect 16264 41024 20668 41052
rect 16264 41012 16270 41024
rect 5994 40984 6000 40996
rect 5644 40956 6000 40984
rect 4019 40953 4031 40956
rect 3973 40947 4031 40953
rect 5994 40944 6000 40956
rect 6052 40944 6058 40996
rect 20625 40987 20683 40993
rect 20625 40953 20637 40987
rect 20671 40984 20683 40987
rect 20916 40984 20944 41092
rect 21085 41089 21097 41092
rect 21131 41089 21143 41123
rect 21085 41083 21143 41089
rect 21266 41080 21272 41132
rect 21324 41120 21330 41132
rect 21361 41123 21419 41129
rect 21361 41120 21373 41123
rect 21324 41092 21373 41120
rect 21324 41080 21330 41092
rect 21361 41089 21373 41092
rect 21407 41089 21419 41123
rect 21361 41083 21419 41089
rect 21450 41080 21456 41132
rect 21508 41120 21514 41132
rect 21637 41123 21695 41129
rect 21637 41120 21649 41123
rect 21508 41092 21649 41120
rect 21508 41080 21514 41092
rect 21637 41089 21649 41092
rect 21683 41089 21695 41123
rect 21637 41083 21695 41089
rect 22002 41080 22008 41132
rect 22060 41120 22066 41132
rect 22060 41080 22094 41120
rect 22186 41080 22192 41132
rect 22244 41080 22250 41132
rect 22462 41080 22468 41132
rect 22520 41080 22526 41132
rect 22649 41123 22707 41129
rect 22649 41089 22661 41123
rect 22695 41089 22707 41123
rect 22649 41083 22707 41089
rect 21910 41012 21916 41064
rect 21968 41012 21974 41064
rect 22066 41052 22094 41080
rect 22664 41052 22692 41083
rect 23106 41080 23112 41132
rect 23164 41080 23170 41132
rect 23661 41123 23719 41129
rect 23661 41089 23673 41123
rect 23707 41120 23719 41123
rect 23842 41120 23848 41132
rect 23707 41092 23848 41120
rect 23707 41089 23719 41092
rect 23661 41083 23719 41089
rect 23842 41080 23848 41092
rect 23900 41080 23906 41132
rect 22066 41024 22692 41052
rect 21928 40984 21956 41012
rect 22005 40987 22063 40993
rect 22005 40984 22017 40987
rect 20671 40956 20944 40984
rect 21100 40956 21312 40984
rect 21928 40956 22017 40984
rect 20671 40953 20683 40956
rect 20625 40947 20683 40953
rect 2130 40876 2136 40928
rect 2188 40916 2194 40928
rect 2682 40916 2688 40928
rect 2188 40888 2688 40916
rect 2188 40876 2194 40888
rect 2682 40876 2688 40888
rect 2740 40876 2746 40928
rect 3234 40876 3240 40928
rect 3292 40916 3298 40928
rect 4338 40916 4344 40928
rect 3292 40888 4344 40916
rect 3292 40876 3298 40888
rect 4338 40876 4344 40888
rect 4396 40876 4402 40928
rect 6546 40876 6552 40928
rect 6604 40876 6610 40928
rect 8849 40919 8907 40925
rect 8849 40885 8861 40919
rect 8895 40916 8907 40919
rect 17034 40916 17040 40928
rect 8895 40888 17040 40916
rect 8895 40885 8907 40888
rect 8849 40879 8907 40885
rect 17034 40876 17040 40888
rect 17092 40876 17098 40928
rect 19061 40919 19119 40925
rect 19061 40885 19073 40919
rect 19107 40916 19119 40919
rect 21100 40916 21128 40956
rect 19107 40888 21128 40916
rect 21284 40916 21312 40956
rect 22005 40953 22017 40956
rect 22051 40953 22063 40987
rect 22005 40947 22063 40953
rect 22756 40956 23796 40984
rect 22756 40916 22784 40956
rect 23768 40928 23796 40956
rect 21284 40888 22784 40916
rect 22833 40919 22891 40925
rect 19107 40885 19119 40888
rect 19061 40879 19119 40885
rect 22833 40885 22845 40919
rect 22879 40916 22891 40919
rect 23658 40916 23664 40928
rect 22879 40888 23664 40916
rect 22879 40885 22891 40888
rect 22833 40879 22891 40885
rect 23658 40876 23664 40888
rect 23716 40876 23722 40928
rect 23750 40876 23756 40928
rect 23808 40876 23814 40928
rect 1104 40826 24564 40848
rect 1104 40774 3882 40826
rect 3934 40774 3946 40826
rect 3998 40774 4010 40826
rect 4062 40774 4074 40826
rect 4126 40774 4138 40826
rect 4190 40774 9747 40826
rect 9799 40774 9811 40826
rect 9863 40774 9875 40826
rect 9927 40774 9939 40826
rect 9991 40774 10003 40826
rect 10055 40774 15612 40826
rect 15664 40774 15676 40826
rect 15728 40774 15740 40826
rect 15792 40774 15804 40826
rect 15856 40774 15868 40826
rect 15920 40774 21477 40826
rect 21529 40774 21541 40826
rect 21593 40774 21605 40826
rect 21657 40774 21669 40826
rect 21721 40774 21733 40826
rect 21785 40774 24564 40826
rect 1104 40752 24564 40774
rect 2682 40672 2688 40724
rect 2740 40712 2746 40724
rect 2740 40684 3280 40712
rect 2740 40672 2746 40684
rect 3252 40644 3280 40684
rect 3418 40672 3424 40724
rect 3476 40672 3482 40724
rect 3973 40715 4031 40721
rect 3973 40681 3985 40715
rect 4019 40681 4031 40715
rect 3973 40675 4031 40681
rect 3988 40644 4016 40675
rect 4062 40672 4068 40724
rect 4120 40712 4126 40724
rect 4525 40715 4583 40721
rect 4525 40712 4537 40715
rect 4120 40684 4537 40712
rect 4120 40672 4126 40684
rect 4525 40681 4537 40684
rect 4571 40681 4583 40715
rect 4525 40675 4583 40681
rect 4706 40672 4712 40724
rect 4764 40712 4770 40724
rect 5629 40715 5687 40721
rect 5629 40712 5641 40715
rect 4764 40684 5641 40712
rect 4764 40672 4770 40684
rect 5629 40681 5641 40684
rect 5675 40681 5687 40715
rect 5629 40675 5687 40681
rect 5718 40672 5724 40724
rect 5776 40672 5782 40724
rect 5902 40672 5908 40724
rect 5960 40672 5966 40724
rect 5997 40715 6055 40721
rect 5997 40681 6009 40715
rect 6043 40712 6055 40715
rect 6086 40712 6092 40724
rect 6043 40684 6092 40712
rect 6043 40681 6055 40684
rect 5997 40675 6055 40681
rect 6086 40672 6092 40684
rect 6144 40672 6150 40724
rect 7190 40672 7196 40724
rect 7248 40672 7254 40724
rect 18417 40715 18475 40721
rect 18417 40681 18429 40715
rect 18463 40712 18475 40715
rect 19242 40712 19248 40724
rect 18463 40684 19248 40712
rect 18463 40681 18475 40684
rect 18417 40675 18475 40681
rect 19242 40672 19248 40684
rect 19300 40672 19306 40724
rect 19978 40672 19984 40724
rect 20036 40712 20042 40724
rect 21545 40715 21603 40721
rect 21545 40712 21557 40715
rect 20036 40684 21557 40712
rect 20036 40672 20042 40684
rect 21545 40681 21557 40684
rect 21591 40681 21603 40715
rect 21545 40675 21603 40681
rect 21637 40715 21695 40721
rect 21637 40681 21649 40715
rect 21683 40712 21695 40715
rect 21818 40712 21824 40724
rect 21683 40684 21824 40712
rect 21683 40681 21695 40684
rect 21637 40675 21695 40681
rect 21818 40672 21824 40684
rect 21876 40672 21882 40724
rect 21910 40672 21916 40724
rect 21968 40672 21974 40724
rect 22189 40715 22247 40721
rect 22189 40681 22201 40715
rect 22235 40712 22247 40715
rect 22462 40712 22468 40724
rect 22235 40684 22468 40712
rect 22235 40681 22247 40684
rect 22189 40675 22247 40681
rect 22462 40672 22468 40684
rect 22520 40672 22526 40724
rect 23109 40715 23167 40721
rect 23109 40681 23121 40715
rect 23155 40712 23167 40715
rect 23290 40712 23296 40724
rect 23155 40684 23296 40712
rect 23155 40681 23167 40684
rect 23109 40675 23167 40681
rect 23290 40672 23296 40684
rect 23348 40672 23354 40724
rect 24121 40715 24179 40721
rect 24121 40681 24133 40715
rect 24167 40712 24179 40715
rect 25222 40712 25228 40724
rect 24167 40684 25228 40712
rect 24167 40681 24179 40684
rect 24121 40675 24179 40681
rect 25222 40672 25228 40684
rect 25280 40672 25286 40724
rect 3252 40616 4016 40644
rect 2130 40536 2136 40588
rect 2188 40536 2194 40588
rect 2406 40536 2412 40588
rect 2464 40536 2470 40588
rect 2547 40579 2605 40585
rect 2547 40545 2559 40579
rect 2593 40576 2605 40579
rect 3234 40576 3240 40588
rect 2593 40548 3240 40576
rect 2593 40545 2605 40548
rect 2547 40539 2605 40545
rect 3234 40536 3240 40548
rect 3292 40536 3298 40588
rect 3329 40579 3387 40585
rect 3329 40545 3341 40579
rect 3375 40576 3387 40579
rect 5736 40576 5764 40672
rect 5920 40644 5948 40672
rect 6917 40647 6975 40653
rect 6917 40644 6929 40647
rect 5920 40616 6929 40644
rect 6917 40613 6929 40616
rect 6963 40613 6975 40647
rect 6917 40607 6975 40613
rect 7466 40604 7472 40656
rect 7524 40644 7530 40656
rect 7834 40644 7840 40656
rect 7524 40616 7840 40644
rect 7524 40604 7530 40616
rect 7834 40604 7840 40616
rect 7892 40604 7898 40656
rect 21082 40604 21088 40656
rect 21140 40604 21146 40656
rect 22370 40604 22376 40656
rect 22428 40644 22434 40656
rect 23014 40644 23020 40656
rect 22428 40616 23020 40644
rect 22428 40604 22434 40616
rect 23014 40604 23020 40616
rect 23072 40604 23078 40656
rect 23569 40647 23627 40653
rect 23569 40613 23581 40647
rect 23615 40644 23627 40647
rect 24946 40644 24952 40656
rect 23615 40616 24952 40644
rect 23615 40613 23627 40616
rect 23569 40607 23627 40613
rect 24946 40604 24952 40616
rect 25004 40604 25010 40656
rect 3375 40548 5764 40576
rect 3375 40545 3387 40548
rect 3329 40539 3387 40545
rect 6270 40536 6276 40588
rect 6328 40576 6334 40588
rect 9490 40576 9496 40588
rect 6328 40548 9496 40576
rect 6328 40536 6334 40548
rect 9490 40536 9496 40548
rect 9548 40536 9554 40588
rect 20806 40536 20812 40588
rect 20864 40576 20870 40588
rect 20864 40548 21404 40576
rect 20864 40536 20870 40548
rect 1489 40511 1547 40517
rect 1489 40477 1501 40511
rect 1535 40477 1547 40511
rect 1489 40471 1547 40477
rect 1504 40372 1532 40471
rect 1670 40468 1676 40520
rect 1728 40468 1734 40520
rect 2682 40468 2688 40520
rect 2740 40468 2746 40520
rect 3602 40468 3608 40520
rect 3660 40468 3666 40520
rect 4246 40468 4252 40520
rect 4304 40508 4310 40520
rect 4304 40480 5028 40508
rect 4304 40468 4310 40480
rect 3234 40400 3240 40452
rect 3292 40440 3298 40452
rect 3881 40443 3939 40449
rect 3881 40440 3893 40443
rect 3292 40412 3893 40440
rect 3292 40400 3298 40412
rect 3881 40409 3893 40412
rect 3927 40409 3939 40443
rect 3881 40403 3939 40409
rect 4430 40400 4436 40452
rect 4488 40400 4494 40452
rect 5000 40449 5028 40480
rect 6178 40468 6184 40520
rect 6236 40468 6242 40520
rect 7101 40511 7159 40517
rect 7101 40508 7113 40511
rect 6564 40480 7113 40508
rect 4985 40443 5043 40449
rect 4985 40409 4997 40443
rect 5031 40409 5043 40443
rect 4985 40403 5043 40409
rect 5534 40400 5540 40452
rect 5592 40400 5598 40452
rect 5626 40400 5632 40452
rect 5684 40440 5690 40452
rect 5902 40440 5908 40452
rect 5684 40412 5908 40440
rect 5684 40400 5690 40412
rect 5902 40400 5908 40412
rect 5960 40400 5966 40452
rect 2314 40372 2320 40384
rect 1504 40344 2320 40372
rect 2314 40332 2320 40344
rect 2372 40332 2378 40384
rect 2958 40332 2964 40384
rect 3016 40372 3022 40384
rect 5077 40375 5135 40381
rect 5077 40372 5089 40375
rect 3016 40344 5089 40372
rect 3016 40332 3022 40344
rect 5077 40341 5089 40344
rect 5123 40341 5135 40375
rect 5077 40335 5135 40341
rect 5718 40332 5724 40384
rect 5776 40372 5782 40384
rect 6564 40381 6592 40480
rect 7101 40477 7113 40480
rect 7147 40477 7159 40511
rect 7101 40471 7159 40477
rect 7190 40468 7196 40520
rect 7248 40508 7254 40520
rect 7377 40511 7435 40517
rect 7377 40508 7389 40511
rect 7248 40480 7389 40508
rect 7248 40468 7254 40480
rect 7377 40477 7389 40480
rect 7423 40477 7435 40511
rect 7377 40471 7435 40477
rect 10502 40468 10508 40520
rect 10560 40508 10566 40520
rect 21376 40517 21404 40548
rect 21910 40536 21916 40588
rect 21968 40576 21974 40588
rect 23658 40576 23664 40588
rect 21968 40548 23664 40576
rect 21968 40536 21974 40548
rect 23658 40536 23664 40548
rect 23716 40536 23722 40588
rect 18601 40511 18659 40517
rect 18601 40508 18613 40511
rect 10560 40480 18613 40508
rect 10560 40468 10566 40480
rect 18601 40477 18613 40480
rect 18647 40477 18659 40511
rect 21269 40511 21327 40517
rect 21269 40508 21281 40511
rect 18601 40471 18659 40477
rect 18708 40480 21281 40508
rect 13538 40400 13544 40452
rect 13596 40440 13602 40452
rect 18708 40440 18736 40480
rect 21269 40477 21281 40480
rect 21315 40477 21327 40511
rect 21269 40471 21327 40477
rect 21361 40511 21419 40517
rect 21361 40477 21373 40511
rect 21407 40477 21419 40511
rect 21361 40471 21419 40477
rect 21821 40511 21879 40517
rect 21821 40477 21833 40511
rect 21867 40477 21879 40511
rect 21821 40471 21879 40477
rect 13596 40412 18736 40440
rect 13596 40400 13602 40412
rect 20806 40400 20812 40452
rect 20864 40440 20870 40452
rect 21836 40440 21864 40471
rect 22094 40468 22100 40520
rect 22152 40468 22158 40520
rect 22373 40511 22431 40517
rect 22373 40477 22385 40511
rect 22419 40477 22431 40511
rect 22373 40471 22431 40477
rect 22388 40440 22416 40471
rect 22462 40468 22468 40520
rect 22520 40508 22526 40520
rect 22833 40511 22891 40517
rect 22833 40508 22845 40511
rect 22520 40480 22845 40508
rect 22520 40468 22526 40480
rect 22833 40477 22845 40480
rect 22879 40477 22891 40511
rect 22833 40471 22891 40477
rect 23290 40468 23296 40520
rect 23348 40468 23354 40520
rect 23385 40511 23443 40517
rect 23385 40477 23397 40511
rect 23431 40477 23443 40511
rect 23385 40471 23443 40477
rect 20864 40412 21864 40440
rect 22066 40412 22416 40440
rect 20864 40400 20870 40412
rect 6549 40375 6607 40381
rect 6549 40372 6561 40375
rect 5776 40344 6561 40372
rect 5776 40332 5782 40344
rect 6549 40341 6561 40344
rect 6595 40341 6607 40375
rect 6549 40335 6607 40341
rect 19702 40332 19708 40384
rect 19760 40372 19766 40384
rect 22066 40372 22094 40412
rect 23198 40400 23204 40452
rect 23256 40440 23262 40452
rect 23400 40440 23428 40471
rect 23256 40412 23428 40440
rect 23256 40400 23262 40412
rect 23750 40400 23756 40452
rect 23808 40440 23814 40452
rect 23845 40443 23903 40449
rect 23845 40440 23857 40443
rect 23808 40412 23857 40440
rect 23808 40400 23814 40412
rect 23845 40409 23857 40412
rect 23891 40409 23903 40443
rect 23845 40403 23903 40409
rect 19760 40344 22094 40372
rect 19760 40332 19766 40344
rect 22646 40332 22652 40384
rect 22704 40332 22710 40384
rect 1104 40282 24723 40304
rect 1104 40230 6814 40282
rect 6866 40230 6878 40282
rect 6930 40230 6942 40282
rect 6994 40230 7006 40282
rect 7058 40230 7070 40282
rect 7122 40230 12679 40282
rect 12731 40230 12743 40282
rect 12795 40230 12807 40282
rect 12859 40230 12871 40282
rect 12923 40230 12935 40282
rect 12987 40230 18544 40282
rect 18596 40230 18608 40282
rect 18660 40230 18672 40282
rect 18724 40230 18736 40282
rect 18788 40230 18800 40282
rect 18852 40230 24409 40282
rect 24461 40230 24473 40282
rect 24525 40230 24537 40282
rect 24589 40230 24601 40282
rect 24653 40230 24665 40282
rect 24717 40230 24723 40282
rect 1104 40208 24723 40230
rect 2593 40171 2651 40177
rect 2593 40137 2605 40171
rect 2639 40168 2651 40171
rect 2682 40168 2688 40180
rect 2639 40140 2688 40168
rect 2639 40137 2651 40140
rect 2593 40131 2651 40137
rect 2682 40128 2688 40140
rect 2740 40128 2746 40180
rect 6546 40168 6552 40180
rect 2884 40140 6552 40168
rect 382 40060 388 40112
rect 440 40100 446 40112
rect 2884 40100 2912 40140
rect 6546 40128 6552 40140
rect 6604 40128 6610 40180
rect 19334 40128 19340 40180
rect 19392 40168 19398 40180
rect 21453 40171 21511 40177
rect 21453 40168 21465 40171
rect 19392 40140 21465 40168
rect 19392 40128 19398 40140
rect 21453 40137 21465 40140
rect 21499 40137 21511 40171
rect 21453 40131 21511 40137
rect 22002 40128 22008 40180
rect 22060 40128 22066 40180
rect 22281 40171 22339 40177
rect 22281 40137 22293 40171
rect 22327 40137 22339 40171
rect 22281 40131 22339 40137
rect 440 40072 2912 40100
rect 440 40060 446 40072
rect 2958 40060 2964 40112
rect 3016 40060 3022 40112
rect 3510 40060 3516 40112
rect 3568 40100 3574 40112
rect 5905 40103 5963 40109
rect 5905 40100 5917 40103
rect 3568 40072 5917 40100
rect 3568 40060 3574 40072
rect 5905 40069 5917 40072
rect 5951 40100 5963 40103
rect 6454 40100 6460 40112
rect 5951 40072 6460 40100
rect 5951 40069 5963 40072
rect 5905 40063 5963 40069
rect 6454 40060 6460 40072
rect 6512 40060 6518 40112
rect 6564 40072 6868 40100
rect 1855 40035 1913 40041
rect 1855 40001 1867 40035
rect 1901 40032 1913 40035
rect 2314 40032 2320 40044
rect 1901 40004 2320 40032
rect 1901 40001 1913 40004
rect 1855 39995 1913 40001
rect 2314 39992 2320 40004
rect 2372 39992 2378 40044
rect 3418 39992 3424 40044
rect 3476 40032 3482 40044
rect 4215 40035 4273 40041
rect 4215 40032 4227 40035
rect 3476 40004 4227 40032
rect 3476 39992 3482 40004
rect 4215 40001 4227 40004
rect 4261 40001 4273 40035
rect 4215 39995 4273 40001
rect 4798 39992 4804 40044
rect 4856 40032 4862 40044
rect 6564 40032 6592 40072
rect 4856 40004 6592 40032
rect 6639 40035 6697 40041
rect 4856 39992 4862 40004
rect 6639 40001 6651 40035
rect 6685 40032 6697 40035
rect 6730 40032 6736 40044
rect 6685 40004 6736 40032
rect 6685 40001 6697 40004
rect 6639 39995 6697 40001
rect 6730 39992 6736 40004
rect 6788 39992 6794 40044
rect 6840 40032 6868 40072
rect 19886 40060 19892 40112
rect 19944 40100 19950 40112
rect 22296 40100 22324 40131
rect 22646 40128 22652 40180
rect 22704 40128 22710 40180
rect 22922 40128 22928 40180
rect 22980 40128 22986 40180
rect 23201 40171 23259 40177
rect 23201 40137 23213 40171
rect 23247 40168 23259 40171
rect 23566 40168 23572 40180
rect 23247 40140 23572 40168
rect 23247 40137 23259 40140
rect 23201 40131 23259 40137
rect 23566 40128 23572 40140
rect 23624 40128 23630 40180
rect 23658 40128 23664 40180
rect 23716 40128 23722 40180
rect 19944 40072 21220 40100
rect 19944 40060 19950 40072
rect 10502 40032 10508 40044
rect 6840 40004 10508 40032
rect 10502 39992 10508 40004
rect 10560 39992 10566 40044
rect 10962 39992 10968 40044
rect 11020 40032 11026 40044
rect 16574 40032 16580 40044
rect 11020 40004 16580 40032
rect 11020 39992 11026 40004
rect 16574 39992 16580 40004
rect 16632 39992 16638 40044
rect 21192 40032 21220 40072
rect 22204 40072 22324 40100
rect 22664 40100 22692 40128
rect 23676 40100 23704 40128
rect 23845 40103 23903 40109
rect 23845 40100 23857 40103
rect 22664 40072 23428 40100
rect 23676 40072 23857 40100
rect 22204 40041 22232 40072
rect 21637 40035 21695 40041
rect 21637 40032 21649 40035
rect 21192 40004 21649 40032
rect 21637 40001 21649 40004
rect 21683 40001 21695 40035
rect 21637 39995 21695 40001
rect 22189 40035 22247 40041
rect 22189 40001 22201 40035
rect 22235 40001 22247 40035
rect 22189 39995 22247 40001
rect 22370 39992 22376 40044
rect 22428 40032 22434 40044
rect 22465 40035 22523 40041
rect 22465 40032 22477 40035
rect 22428 40004 22477 40032
rect 22428 39992 22434 40004
rect 22465 40001 22477 40004
rect 22511 40032 22523 40035
rect 22741 40035 22799 40041
rect 22741 40032 22753 40035
rect 22511 40004 22753 40032
rect 22511 40001 22523 40004
rect 22465 39995 22523 40001
rect 22741 40001 22753 40004
rect 22787 40001 22799 40035
rect 22741 39995 22799 40001
rect 23014 39992 23020 40044
rect 23072 40032 23078 40044
rect 23400 40041 23428 40072
rect 23845 40069 23857 40072
rect 23891 40069 23903 40103
rect 25498 40100 25504 40112
rect 23845 40063 23903 40069
rect 23952 40072 25504 40100
rect 23109 40035 23167 40041
rect 23109 40032 23121 40035
rect 23072 40004 23121 40032
rect 23072 39992 23078 40004
rect 23109 40001 23121 40004
rect 23155 40001 23167 40035
rect 23109 39995 23167 40001
rect 23385 40035 23443 40041
rect 23385 40001 23397 40035
rect 23431 40001 23443 40035
rect 23385 39995 23443 40001
rect 23661 40035 23719 40041
rect 23661 40001 23673 40035
rect 23707 40032 23719 40035
rect 23952 40032 23980 40072
rect 25498 40060 25504 40072
rect 25556 40060 25562 40112
rect 23707 40004 23980 40032
rect 23707 40001 23719 40004
rect 23661 39995 23719 40001
rect 1578 39924 1584 39976
rect 1636 39924 1642 39976
rect 3694 39924 3700 39976
rect 3752 39924 3758 39976
rect 3786 39924 3792 39976
rect 3844 39924 3850 39976
rect 3970 39924 3976 39976
rect 4028 39924 4034 39976
rect 6365 39967 6423 39973
rect 6365 39933 6377 39967
rect 6411 39933 6423 39967
rect 6365 39927 6423 39933
rect 3712 39896 3740 39924
rect 3988 39896 4016 39924
rect 3712 39868 4016 39896
rect 4632 39868 5120 39896
rect 3510 39788 3516 39840
rect 3568 39828 3574 39840
rect 4632 39828 4660 39868
rect 3568 39800 4660 39828
rect 3568 39788 3574 39800
rect 4982 39788 4988 39840
rect 5040 39788 5046 39840
rect 5092 39828 5120 39868
rect 5626 39856 5632 39908
rect 5684 39856 5690 39908
rect 6178 39856 6184 39908
rect 6236 39896 6242 39908
rect 6380 39896 6408 39927
rect 7650 39924 7656 39976
rect 7708 39964 7714 39976
rect 7708 39936 10824 39964
rect 7708 39924 7714 39936
rect 6236 39868 6408 39896
rect 7024 39868 8340 39896
rect 6236 39856 6242 39868
rect 7024 39828 7052 39868
rect 8312 39840 8340 39868
rect 10796 39840 10824 39936
rect 22066 39936 23612 39964
rect 13630 39856 13636 39908
rect 13688 39896 13694 39908
rect 22066 39896 22094 39936
rect 23477 39899 23535 39905
rect 23477 39896 23489 39899
rect 13688 39868 22094 39896
rect 22296 39868 23489 39896
rect 13688 39856 13694 39868
rect 5092 39800 7052 39828
rect 7374 39788 7380 39840
rect 7432 39788 7438 39840
rect 8294 39788 8300 39840
rect 8352 39788 8358 39840
rect 10778 39788 10784 39840
rect 10836 39788 10842 39840
rect 21266 39788 21272 39840
rect 21324 39828 21330 39840
rect 22296 39828 22324 39868
rect 23477 39865 23489 39868
rect 23523 39865 23535 39899
rect 23477 39859 23535 39865
rect 23584 39840 23612 39936
rect 21324 39800 22324 39828
rect 21324 39788 21330 39800
rect 23566 39788 23572 39840
rect 23624 39788 23630 39840
rect 24118 39788 24124 39840
rect 24176 39788 24182 39840
rect 1104 39738 24564 39760
rect 1104 39686 3882 39738
rect 3934 39686 3946 39738
rect 3998 39686 4010 39738
rect 4062 39686 4074 39738
rect 4126 39686 4138 39738
rect 4190 39686 9747 39738
rect 9799 39686 9811 39738
rect 9863 39686 9875 39738
rect 9927 39686 9939 39738
rect 9991 39686 10003 39738
rect 10055 39686 15612 39738
rect 15664 39686 15676 39738
rect 15728 39686 15740 39738
rect 15792 39686 15804 39738
rect 15856 39686 15868 39738
rect 15920 39686 21477 39738
rect 21529 39686 21541 39738
rect 21593 39686 21605 39738
rect 21657 39686 21669 39738
rect 21721 39686 21733 39738
rect 21785 39686 24564 39738
rect 1104 39664 24564 39686
rect 1673 39627 1731 39633
rect 1673 39593 1685 39627
rect 1719 39624 1731 39627
rect 2222 39624 2228 39636
rect 1719 39596 2228 39624
rect 1719 39593 1731 39596
rect 1673 39587 1731 39593
rect 2222 39584 2228 39596
rect 2280 39584 2286 39636
rect 2590 39584 2596 39636
rect 2648 39624 2654 39636
rect 4341 39627 4399 39633
rect 4341 39624 4353 39627
rect 2648 39596 4353 39624
rect 2648 39584 2654 39596
rect 4341 39593 4353 39596
rect 4387 39593 4399 39627
rect 8202 39624 8208 39636
rect 4341 39587 4399 39593
rect 6104 39596 8208 39624
rect 1486 39516 1492 39568
rect 1544 39556 1550 39568
rect 2041 39559 2099 39565
rect 2041 39556 2053 39559
rect 1544 39528 2053 39556
rect 1544 39516 1550 39528
rect 2041 39525 2053 39528
rect 2087 39525 2099 39559
rect 2041 39519 2099 39525
rect 3973 39491 4031 39497
rect 3973 39488 3985 39491
rect 3712 39460 3985 39488
rect 2317 39423 2375 39429
rect 2317 39389 2329 39423
rect 2363 39389 2375 39423
rect 2317 39383 2375 39389
rect 1854 39312 1860 39364
rect 1912 39312 1918 39364
rect 2332 39352 2360 39383
rect 2498 39380 2504 39432
rect 2556 39420 2562 39432
rect 2591 39423 2649 39429
rect 2591 39420 2603 39423
rect 2556 39392 2603 39420
rect 2556 39380 2562 39392
rect 2591 39389 2603 39392
rect 2637 39389 2649 39423
rect 2591 39383 2649 39389
rect 2682 39380 2688 39432
rect 2740 39420 2746 39432
rect 3712 39420 3740 39460
rect 3973 39457 3985 39460
rect 4019 39457 4031 39491
rect 3973 39451 4031 39457
rect 2740 39392 3740 39420
rect 2740 39380 2746 39392
rect 3786 39380 3792 39432
rect 3844 39380 3850 39432
rect 3050 39352 3056 39364
rect 2332 39324 3056 39352
rect 3050 39312 3056 39324
rect 3108 39312 3114 39364
rect 3988 39352 4016 39451
rect 4982 39448 4988 39500
rect 5040 39448 5046 39500
rect 4522 39380 4528 39432
rect 4580 39380 4586 39432
rect 4706 39380 4712 39432
rect 4764 39420 4770 39432
rect 5537 39423 5595 39429
rect 4764 39392 5488 39420
rect 4764 39380 4770 39392
rect 3988 39324 5028 39352
rect 3326 39244 3332 39296
rect 3384 39244 3390 39296
rect 4801 39287 4859 39293
rect 4801 39253 4813 39287
rect 4847 39284 4859 39287
rect 4890 39284 4896 39296
rect 4847 39256 4896 39284
rect 4847 39253 4859 39256
rect 4801 39247 4859 39253
rect 4890 39244 4896 39256
rect 4948 39244 4954 39296
rect 5000 39284 5028 39324
rect 5074 39312 5080 39364
rect 5132 39312 5138 39364
rect 5166 39312 5172 39364
rect 5224 39312 5230 39364
rect 5460 39352 5488 39392
rect 5537 39389 5549 39423
rect 5583 39420 5595 39423
rect 5902 39420 5908 39432
rect 5583 39392 5908 39420
rect 5583 39389 5595 39392
rect 5537 39383 5595 39389
rect 5902 39380 5908 39392
rect 5960 39380 5966 39432
rect 6104 39352 6132 39596
rect 8202 39584 8208 39596
rect 8260 39584 8266 39636
rect 9125 39627 9183 39633
rect 9125 39593 9137 39627
rect 9171 39624 9183 39627
rect 9398 39624 9404 39636
rect 9171 39596 9404 39624
rect 9171 39593 9183 39596
rect 9125 39587 9183 39593
rect 9398 39584 9404 39596
rect 9456 39584 9462 39636
rect 10226 39624 10232 39636
rect 9876 39596 10232 39624
rect 9033 39559 9091 39565
rect 9033 39525 9045 39559
rect 9079 39556 9091 39559
rect 9677 39559 9735 39565
rect 9677 39556 9689 39559
rect 9079 39528 9689 39556
rect 9079 39525 9091 39528
rect 9033 39519 9091 39525
rect 9677 39525 9689 39528
rect 9723 39525 9735 39559
rect 9677 39519 9735 39525
rect 9876 39497 9904 39596
rect 10226 39584 10232 39596
rect 10284 39584 10290 39636
rect 21358 39584 21364 39636
rect 21416 39624 21422 39636
rect 22833 39627 22891 39633
rect 22833 39624 22845 39627
rect 21416 39596 22845 39624
rect 21416 39584 21422 39596
rect 22833 39593 22845 39596
rect 22879 39593 22891 39627
rect 22833 39587 22891 39593
rect 23198 39584 23204 39636
rect 23256 39584 23262 39636
rect 23290 39584 23296 39636
rect 23348 39624 23354 39636
rect 23661 39627 23719 39633
rect 23661 39624 23673 39627
rect 23348 39596 23673 39624
rect 23348 39584 23354 39596
rect 23661 39593 23673 39596
rect 23707 39593 23719 39627
rect 23661 39587 23719 39593
rect 19337 39559 19395 39565
rect 19337 39525 19349 39559
rect 19383 39556 19395 39559
rect 21910 39556 21916 39568
rect 19383 39528 21916 39556
rect 19383 39525 19395 39528
rect 19337 39519 19395 39525
rect 21910 39516 21916 39528
rect 21968 39516 21974 39568
rect 22373 39559 22431 39565
rect 22373 39525 22385 39559
rect 22419 39556 22431 39559
rect 23216 39556 23244 39584
rect 22419 39528 23244 39556
rect 23385 39559 23443 39565
rect 22419 39525 22431 39528
rect 22373 39519 22431 39525
rect 23385 39525 23397 39559
rect 23431 39525 23443 39559
rect 23385 39519 23443 39525
rect 9217 39491 9275 39497
rect 9217 39457 9229 39491
rect 9263 39488 9275 39491
rect 9401 39491 9459 39497
rect 9401 39488 9413 39491
rect 9263 39460 9413 39488
rect 9263 39457 9275 39460
rect 9217 39451 9275 39457
rect 9401 39457 9413 39460
rect 9447 39457 9459 39491
rect 9401 39451 9459 39457
rect 9861 39491 9919 39497
rect 9861 39457 9873 39491
rect 9907 39457 9919 39491
rect 9861 39451 9919 39457
rect 20346 39448 20352 39500
rect 20404 39488 20410 39500
rect 20404 39460 22094 39488
rect 20404 39448 20410 39460
rect 6178 39380 6184 39432
rect 6236 39420 6242 39432
rect 6825 39423 6883 39429
rect 6825 39420 6837 39423
rect 6236 39392 6837 39420
rect 6236 39380 6242 39392
rect 6825 39389 6837 39392
rect 6871 39389 6883 39423
rect 6825 39383 6883 39389
rect 7099 39423 7157 39429
rect 7099 39389 7111 39423
rect 7145 39420 7157 39423
rect 8110 39420 8116 39432
rect 7145 39392 8116 39420
rect 7145 39389 7157 39392
rect 7099 39383 7157 39389
rect 5460 39324 6132 39352
rect 6840 39352 6868 39383
rect 8110 39380 8116 39392
rect 8168 39380 8174 39432
rect 8941 39423 8999 39429
rect 8941 39389 8953 39423
rect 8987 39420 8999 39423
rect 9309 39423 9367 39429
rect 9309 39420 9321 39423
rect 8987 39392 9321 39420
rect 8987 39389 8999 39392
rect 8941 39383 8999 39389
rect 9309 39389 9321 39392
rect 9355 39420 9367 39423
rect 9355 39392 9444 39420
rect 9355 39389 9367 39392
rect 9309 39383 9367 39389
rect 7282 39352 7288 39364
rect 6840 39324 7288 39352
rect 7282 39312 7288 39324
rect 7340 39312 7346 39364
rect 7392 39324 9260 39352
rect 5626 39284 5632 39296
rect 5000 39256 5632 39284
rect 5626 39244 5632 39256
rect 5684 39244 5690 39296
rect 5905 39287 5963 39293
rect 5905 39253 5917 39287
rect 5951 39284 5963 39287
rect 5994 39284 6000 39296
rect 5951 39256 6000 39284
rect 5951 39253 5963 39256
rect 5905 39247 5963 39253
rect 5994 39244 6000 39256
rect 6052 39244 6058 39296
rect 6086 39244 6092 39296
rect 6144 39244 6150 39296
rect 6454 39244 6460 39296
rect 6512 39284 6518 39296
rect 7392 39284 7420 39324
rect 6512 39256 7420 39284
rect 6512 39244 6518 39256
rect 7466 39244 7472 39296
rect 7524 39284 7530 39296
rect 7837 39287 7895 39293
rect 7837 39284 7849 39287
rect 7524 39256 7849 39284
rect 7524 39244 7530 39256
rect 7837 39253 7849 39256
rect 7883 39284 7895 39287
rect 7926 39284 7932 39296
rect 7883 39256 7932 39284
rect 7883 39253 7895 39256
rect 7837 39247 7895 39253
rect 7926 39244 7932 39256
rect 7984 39244 7990 39296
rect 9232 39284 9260 39324
rect 9416 39296 9444 39392
rect 9490 39380 9496 39432
rect 9548 39380 9554 39432
rect 9582 39380 9588 39432
rect 9640 39380 9646 39432
rect 10135 39423 10193 39429
rect 10135 39420 10147 39423
rect 9692 39392 10147 39420
rect 9306 39284 9312 39296
rect 9232 39256 9312 39284
rect 9306 39244 9312 39256
rect 9364 39244 9370 39296
rect 9398 39244 9404 39296
rect 9456 39244 9462 39296
rect 9490 39244 9496 39296
rect 9548 39284 9554 39296
rect 9692 39284 9720 39392
rect 10135 39389 10147 39392
rect 10181 39420 10193 39423
rect 12434 39420 12440 39432
rect 10181 39392 12440 39420
rect 10181 39389 10193 39392
rect 10135 39383 10193 39389
rect 12434 39380 12440 39392
rect 12492 39380 12498 39432
rect 19518 39380 19524 39432
rect 19576 39380 19582 39432
rect 9766 39312 9772 39364
rect 9824 39352 9830 39364
rect 22066 39352 22094 39460
rect 22554 39380 22560 39432
rect 22612 39380 22618 39432
rect 23017 39423 23075 39429
rect 23017 39389 23029 39423
rect 23063 39420 23075 39423
rect 23198 39420 23204 39432
rect 23063 39392 23204 39420
rect 23063 39389 23075 39392
rect 23017 39383 23075 39389
rect 23198 39380 23204 39392
rect 23256 39380 23262 39432
rect 23293 39423 23351 39429
rect 23293 39389 23305 39423
rect 23339 39420 23351 39423
rect 23400 39420 23428 39519
rect 25222 39488 25228 39500
rect 23860 39460 25228 39488
rect 23339 39392 23428 39420
rect 23339 39389 23351 39392
rect 23293 39383 23351 39389
rect 23566 39380 23572 39432
rect 23624 39380 23630 39432
rect 23860 39429 23888 39460
rect 25222 39448 25228 39460
rect 25280 39448 25286 39500
rect 23845 39423 23903 39429
rect 23845 39389 23857 39423
rect 23891 39389 23903 39423
rect 23845 39383 23903 39389
rect 23937 39423 23995 39429
rect 23937 39389 23949 39423
rect 23983 39389 23995 39423
rect 23937 39383 23995 39389
rect 23952 39352 23980 39383
rect 9824 39324 12112 39352
rect 22066 39324 23980 39352
rect 9824 39312 9830 39324
rect 12084 39296 12112 39324
rect 9548 39256 9720 39284
rect 9548 39244 9554 39256
rect 10410 39244 10416 39296
rect 10468 39284 10474 39296
rect 10873 39287 10931 39293
rect 10873 39284 10885 39287
rect 10468 39256 10885 39284
rect 10468 39244 10474 39256
rect 10873 39253 10885 39256
rect 10919 39253 10931 39287
rect 10873 39247 10931 39253
rect 12066 39244 12072 39296
rect 12124 39244 12130 39296
rect 23109 39287 23167 39293
rect 23109 39253 23121 39287
rect 23155 39284 23167 39287
rect 23474 39284 23480 39296
rect 23155 39256 23480 39284
rect 23155 39253 23167 39256
rect 23109 39247 23167 39253
rect 23474 39244 23480 39256
rect 23532 39244 23538 39296
rect 24121 39287 24179 39293
rect 24121 39253 24133 39287
rect 24167 39284 24179 39287
rect 24854 39284 24860 39296
rect 24167 39256 24860 39284
rect 24167 39253 24179 39256
rect 24121 39247 24179 39253
rect 24854 39244 24860 39256
rect 24912 39244 24918 39296
rect 1104 39194 24723 39216
rect 1104 39142 6814 39194
rect 6866 39142 6878 39194
rect 6930 39142 6942 39194
rect 6994 39142 7006 39194
rect 7058 39142 7070 39194
rect 7122 39142 12679 39194
rect 12731 39142 12743 39194
rect 12795 39142 12807 39194
rect 12859 39142 12871 39194
rect 12923 39142 12935 39194
rect 12987 39142 18544 39194
rect 18596 39142 18608 39194
rect 18660 39142 18672 39194
rect 18724 39142 18736 39194
rect 18788 39142 18800 39194
rect 18852 39142 24409 39194
rect 24461 39142 24473 39194
rect 24525 39142 24537 39194
rect 24589 39142 24601 39194
rect 24653 39142 24665 39194
rect 24717 39142 24723 39194
rect 1104 39120 24723 39142
rect 3418 39080 3424 39092
rect 1688 39052 3424 39080
rect 1688 38983 1716 39052
rect 3418 39040 3424 39052
rect 3476 39040 3482 39092
rect 5166 39040 5172 39092
rect 5224 39080 5230 39092
rect 5905 39083 5963 39089
rect 5905 39080 5917 39083
rect 5224 39052 5917 39080
rect 5224 39040 5230 39052
rect 5905 39049 5917 39052
rect 5951 39049 5963 39083
rect 8757 39083 8815 39089
rect 5905 39043 5963 39049
rect 6012 39052 8432 39080
rect 1655 38977 1716 38983
rect 1655 38943 1667 38977
rect 1701 38946 1716 38977
rect 2314 38972 2320 39024
rect 2372 39012 2378 39024
rect 6012 39012 6040 39052
rect 2372 38984 5120 39012
rect 2372 38972 2378 38984
rect 1701 38943 1713 38946
rect 1655 38937 1713 38943
rect 2038 38904 2044 38956
rect 2096 38944 2102 38956
rect 2682 38944 2688 38956
rect 2096 38916 2688 38944
rect 2096 38904 2102 38916
rect 2682 38904 2688 38916
rect 2740 38904 2746 38956
rect 2774 38904 2780 38956
rect 2832 38904 2838 38956
rect 3050 38904 3056 38956
rect 3108 38944 3114 38956
rect 3789 38947 3847 38953
rect 3789 38944 3801 38947
rect 3108 38916 3801 38944
rect 3108 38904 3114 38916
rect 3789 38913 3801 38916
rect 3835 38913 3847 38947
rect 3789 38907 3847 38913
rect 3970 38904 3976 38956
rect 4028 38944 4034 38956
rect 4065 38947 4123 38953
rect 4065 38944 4077 38947
rect 4028 38916 4077 38944
rect 4028 38904 4034 38916
rect 4065 38913 4077 38916
rect 4111 38913 4123 38947
rect 4065 38907 4123 38913
rect 4338 38904 4344 38956
rect 4396 38904 4402 38956
rect 5092 38954 5120 38984
rect 5276 38984 6040 39012
rect 8404 39012 8432 39052
rect 8757 39049 8769 39083
rect 8803 39080 8815 39083
rect 9582 39080 9588 39092
rect 8803 39052 9588 39080
rect 8803 39049 8815 39052
rect 8757 39043 8815 39049
rect 9582 39040 9588 39052
rect 9640 39040 9646 39092
rect 9766 39040 9772 39092
rect 9824 39040 9830 39092
rect 10410 39080 10416 39092
rect 10336 39052 10416 39080
rect 9490 39012 9496 39024
rect 8404 38984 9496 39012
rect 5167 38957 5225 38963
rect 5167 38954 5179 38957
rect 4893 38947 4951 38953
rect 4893 38944 4905 38947
rect 4540 38916 4905 38944
rect 4540 38888 4568 38916
rect 4893 38913 4905 38916
rect 4939 38913 4951 38947
rect 5092 38926 5179 38954
rect 5167 38923 5179 38926
rect 5213 38954 5225 38957
rect 5276 38954 5304 38984
rect 9490 38972 9496 38984
rect 9548 38972 9554 39024
rect 10042 38972 10048 39024
rect 10100 38972 10106 39024
rect 10137 39015 10195 39021
rect 10137 38981 10149 39015
rect 10183 39012 10195 39015
rect 10336 39012 10364 39052
rect 10410 39040 10416 39052
rect 10468 39040 10474 39092
rect 20346 39040 20352 39092
rect 20404 39040 20410 39092
rect 21821 39083 21879 39089
rect 21821 39049 21833 39083
rect 21867 39080 21879 39083
rect 22554 39080 22560 39092
rect 21867 39052 22560 39080
rect 21867 39049 21879 39052
rect 21821 39043 21879 39049
rect 22554 39040 22560 39052
rect 22612 39040 22618 39092
rect 22925 39083 22983 39089
rect 22925 39049 22937 39083
rect 22971 39080 22983 39083
rect 23934 39080 23940 39092
rect 22971 39052 23940 39080
rect 22971 39049 22983 39052
rect 22925 39043 22983 39049
rect 23934 39040 23940 39052
rect 23992 39040 23998 39092
rect 10183 38984 10364 39012
rect 10183 38981 10195 38984
rect 10137 38975 10195 38981
rect 10686 38972 10692 39024
rect 10744 39012 10750 39024
rect 10873 39015 10931 39021
rect 10873 39012 10885 39015
rect 10744 38984 10885 39012
rect 10744 38972 10750 38984
rect 10873 38981 10885 38984
rect 10919 38981 10931 39015
rect 10873 38975 10931 38981
rect 10962 38972 10968 39024
rect 11020 38972 11026 39024
rect 21082 38972 21088 39024
rect 21140 39012 21146 39024
rect 21140 38984 23152 39012
rect 21140 38972 21146 38984
rect 5213 38926 5304 38954
rect 6917 38947 6975 38953
rect 6917 38944 6929 38947
rect 5213 38923 5225 38926
rect 5167 38917 5225 38923
rect 4893 38907 4951 38913
rect 6564 38916 6929 38944
rect 6564 38888 6592 38916
rect 6917 38913 6929 38916
rect 6963 38913 6975 38947
rect 6917 38907 6975 38913
rect 7650 38904 7656 38956
rect 7708 38904 7714 38956
rect 7742 38904 7748 38956
rect 7800 38953 7806 38956
rect 7800 38947 7828 38953
rect 7816 38913 7828 38947
rect 7800 38907 7828 38913
rect 7800 38904 7806 38907
rect 7926 38904 7932 38956
rect 7984 38904 7990 38956
rect 8938 38904 8944 38956
rect 8996 38904 9002 38956
rect 9309 38947 9367 38953
rect 9309 38913 9321 38947
rect 9355 38944 9367 38947
rect 10505 38947 10563 38953
rect 10505 38944 10517 38947
rect 9355 38916 10517 38944
rect 9355 38913 9367 38916
rect 9309 38907 9367 38913
rect 10505 38913 10517 38916
rect 10551 38944 10563 38947
rect 10980 38944 11008 38972
rect 10551 38916 11008 38944
rect 11517 38947 11575 38953
rect 10551 38913 10563 38916
rect 10505 38907 10563 38913
rect 11517 38913 11529 38947
rect 11563 38944 11575 38947
rect 12066 38944 12072 38956
rect 11563 38916 12072 38944
rect 11563 38913 11575 38916
rect 11517 38907 11575 38913
rect 12066 38904 12072 38916
rect 12124 38904 12130 38956
rect 20530 38904 20536 38956
rect 20588 38904 20594 38956
rect 22002 38904 22008 38956
rect 22060 38904 22066 38956
rect 23124 38953 23152 38984
rect 23198 38972 23204 39024
rect 23256 39012 23262 39024
rect 23845 39015 23903 39021
rect 23845 39012 23857 39015
rect 23256 38984 23857 39012
rect 23256 38972 23262 38984
rect 23845 38981 23857 38984
rect 23891 38981 23903 39015
rect 23845 38975 23903 38981
rect 23109 38947 23167 38953
rect 23109 38913 23121 38947
rect 23155 38913 23167 38947
rect 23109 38907 23167 38913
rect 23385 38947 23443 38953
rect 23385 38913 23397 38947
rect 23431 38913 23443 38947
rect 23385 38907 23443 38913
rect 1397 38879 1455 38885
rect 1397 38845 1409 38879
rect 1443 38845 1455 38879
rect 1397 38839 1455 38845
rect 1412 38808 1440 38839
rect 3602 38836 3608 38888
rect 3660 38836 3666 38888
rect 3694 38836 3700 38888
rect 3752 38876 3758 38888
rect 4522 38876 4528 38888
rect 3752 38848 4528 38876
rect 3752 38836 3758 38848
rect 4522 38836 4528 38848
rect 4580 38836 4586 38888
rect 4617 38879 4675 38885
rect 4617 38845 4629 38879
rect 4663 38876 4675 38879
rect 4706 38876 4712 38888
rect 4663 38848 4712 38876
rect 4663 38845 4675 38848
rect 4617 38839 4675 38845
rect 4706 38836 4712 38848
rect 4764 38836 4770 38888
rect 6362 38836 6368 38888
rect 6420 38836 6426 38888
rect 6546 38836 6552 38888
rect 6604 38836 6610 38888
rect 6733 38879 6791 38885
rect 6733 38845 6745 38879
rect 6779 38845 6791 38879
rect 6733 38839 6791 38845
rect 1412 38780 1532 38808
rect 1504 38752 1532 38780
rect 2130 38768 2136 38820
rect 2188 38808 2194 38820
rect 2409 38811 2467 38817
rect 2409 38808 2421 38811
rect 2188 38780 2421 38808
rect 2188 38768 2194 38780
rect 2409 38777 2421 38780
rect 2455 38777 2467 38811
rect 2409 38771 2467 38777
rect 2498 38768 2504 38820
rect 2556 38808 2562 38820
rect 4798 38808 4804 38820
rect 2556 38780 4804 38808
rect 2556 38768 2562 38780
rect 4798 38768 4804 38780
rect 4856 38768 4862 38820
rect 6380 38808 6408 38836
rect 6748 38808 6776 38839
rect 7374 38836 7380 38888
rect 7432 38836 7438 38888
rect 10226 38836 10232 38888
rect 10284 38836 10290 38888
rect 20990 38836 20996 38888
rect 21048 38876 21054 38888
rect 23400 38876 23428 38907
rect 21048 38848 23428 38876
rect 21048 38836 21054 38848
rect 6380 38780 6776 38808
rect 14642 38768 14648 38820
rect 14700 38808 14706 38820
rect 14700 38780 22094 38808
rect 14700 38768 14706 38780
rect 1486 38700 1492 38752
rect 1544 38700 1550 38752
rect 3418 38700 3424 38752
rect 3476 38740 3482 38752
rect 3602 38740 3608 38752
rect 3476 38712 3608 38740
rect 3476 38700 3482 38712
rect 3602 38700 3608 38712
rect 3660 38700 3666 38752
rect 3694 38700 3700 38752
rect 3752 38740 3758 38752
rect 8018 38740 8024 38752
rect 3752 38712 8024 38740
rect 3752 38700 3758 38712
rect 8018 38700 8024 38712
rect 8076 38700 8082 38752
rect 8570 38700 8576 38752
rect 8628 38700 8634 38752
rect 10962 38700 10968 38752
rect 11020 38740 11026 38752
rect 11057 38743 11115 38749
rect 11057 38740 11069 38743
rect 11020 38712 11069 38740
rect 11020 38700 11026 38712
rect 11057 38709 11069 38712
rect 11103 38709 11115 38743
rect 11057 38703 11115 38709
rect 11698 38700 11704 38752
rect 11756 38700 11762 38752
rect 22066 38740 22094 38780
rect 23106 38768 23112 38820
rect 23164 38808 23170 38820
rect 23201 38811 23259 38817
rect 23201 38808 23213 38811
rect 23164 38780 23213 38808
rect 23164 38768 23170 38780
rect 23201 38777 23213 38780
rect 23247 38777 23259 38811
rect 24302 38808 24308 38820
rect 23201 38771 23259 38777
rect 23308 38780 24308 38808
rect 23308 38740 23336 38780
rect 24302 38768 24308 38780
rect 24360 38768 24366 38820
rect 22066 38712 23336 38740
rect 24118 38700 24124 38752
rect 24176 38700 24182 38752
rect 1104 38650 24564 38672
rect 1104 38598 3882 38650
rect 3934 38598 3946 38650
rect 3998 38598 4010 38650
rect 4062 38598 4074 38650
rect 4126 38598 4138 38650
rect 4190 38598 9747 38650
rect 9799 38598 9811 38650
rect 9863 38598 9875 38650
rect 9927 38598 9939 38650
rect 9991 38598 10003 38650
rect 10055 38598 15612 38650
rect 15664 38598 15676 38650
rect 15728 38598 15740 38650
rect 15792 38598 15804 38650
rect 15856 38598 15868 38650
rect 15920 38598 21477 38650
rect 21529 38598 21541 38650
rect 21593 38598 21605 38650
rect 21657 38598 21669 38650
rect 21721 38598 21733 38650
rect 21785 38598 24564 38650
rect 1104 38576 24564 38598
rect 1026 38496 1032 38548
rect 1084 38536 1090 38548
rect 5718 38536 5724 38548
rect 1084 38508 5724 38536
rect 1084 38496 1090 38508
rect 5718 38496 5724 38508
rect 5776 38496 5782 38548
rect 7374 38536 7380 38548
rect 7116 38508 7380 38536
rect 3694 38468 3700 38480
rect 2240 38440 3700 38468
rect 2240 38409 2268 38440
rect 3694 38428 3700 38440
rect 3752 38428 3758 38480
rect 4706 38428 4712 38480
rect 4764 38468 4770 38480
rect 4801 38471 4859 38477
rect 4801 38468 4813 38471
rect 4764 38440 4813 38468
rect 4764 38428 4770 38440
rect 4801 38437 4813 38440
rect 4847 38437 4859 38471
rect 4801 38431 4859 38437
rect 5442 38428 5448 38480
rect 5500 38468 5506 38480
rect 7116 38477 7144 38508
rect 7374 38496 7380 38508
rect 7432 38496 7438 38548
rect 7466 38496 7472 38548
rect 7524 38536 7530 38548
rect 8297 38539 8355 38545
rect 7524 38508 8064 38536
rect 7524 38496 7530 38508
rect 7101 38471 7159 38477
rect 5500 38440 5764 38468
rect 5500 38428 5506 38440
rect 2225 38403 2283 38409
rect 2225 38369 2237 38403
rect 2271 38369 2283 38403
rect 2225 38363 2283 38369
rect 3234 38360 3240 38412
rect 3292 38400 3298 38412
rect 3789 38403 3847 38409
rect 3789 38400 3801 38403
rect 3292 38372 3801 38400
rect 3292 38360 3298 38372
rect 3789 38369 3801 38372
rect 3835 38369 3847 38403
rect 3789 38363 3847 38369
rect 2409 38335 2467 38341
rect 2409 38301 2421 38335
rect 2455 38332 2467 38335
rect 2774 38332 2780 38344
rect 2455 38304 2780 38332
rect 2455 38301 2467 38304
rect 2409 38295 2467 38301
rect 2774 38292 2780 38304
rect 2832 38292 2838 38344
rect 2958 38292 2964 38344
rect 3016 38292 3022 38344
rect 4062 38292 4068 38344
rect 4120 38332 4126 38344
rect 4120 38304 4163 38332
rect 4120 38292 4126 38304
rect 4982 38292 4988 38344
rect 5040 38332 5046 38344
rect 5169 38335 5227 38341
rect 5169 38332 5181 38335
rect 5040 38304 5181 38332
rect 5040 38292 5046 38304
rect 5169 38301 5181 38304
rect 5215 38301 5227 38335
rect 5169 38295 5227 38301
rect 750 38224 756 38276
rect 808 38264 814 38276
rect 1397 38267 1455 38273
rect 1397 38264 1409 38267
rect 808 38236 1409 38264
rect 808 38224 814 38236
rect 1397 38233 1409 38236
rect 1443 38233 1455 38267
rect 1397 38227 1455 38233
rect 2590 38224 2596 38276
rect 2648 38264 2654 38276
rect 2685 38267 2743 38273
rect 2685 38264 2697 38267
rect 2648 38236 2697 38264
rect 2648 38224 2654 38236
rect 2685 38233 2697 38236
rect 2731 38233 2743 38267
rect 2685 38227 2743 38233
rect 2700 38196 2728 38227
rect 2866 38224 2872 38276
rect 2924 38264 2930 38276
rect 3237 38267 3295 38273
rect 3237 38264 3249 38267
rect 2924 38236 3249 38264
rect 2924 38224 2930 38236
rect 3237 38233 3249 38236
rect 3283 38233 3295 38267
rect 3237 38227 3295 38233
rect 4154 38224 4160 38276
rect 4212 38264 4218 38276
rect 5258 38264 5264 38276
rect 4212 38236 5264 38264
rect 4212 38224 4218 38236
rect 5258 38224 5264 38236
rect 5316 38224 5322 38276
rect 5442 38224 5448 38276
rect 5500 38224 5506 38276
rect 5736 38264 5764 38440
rect 7101 38437 7113 38471
rect 7147 38437 7159 38471
rect 7101 38431 7159 38437
rect 5810 38360 5816 38412
rect 5868 38400 5874 38412
rect 6086 38400 6092 38412
rect 5868 38372 6092 38400
rect 5868 38360 5874 38372
rect 6086 38360 6092 38372
rect 6144 38400 6150 38412
rect 7377 38403 7435 38409
rect 7377 38400 7389 38403
rect 6144 38372 7389 38400
rect 6144 38360 6150 38372
rect 7377 38369 7389 38372
rect 7423 38369 7435 38403
rect 7377 38363 7435 38369
rect 7653 38403 7711 38409
rect 7653 38369 7665 38403
rect 7699 38400 7711 38403
rect 8036 38400 8064 38508
rect 8297 38505 8309 38539
rect 8343 38536 8355 38539
rect 8938 38536 8944 38548
rect 8343 38508 8944 38536
rect 8343 38505 8355 38508
rect 8297 38499 8355 38505
rect 8938 38496 8944 38508
rect 8996 38496 9002 38548
rect 10134 38536 10140 38548
rect 9232 38508 10140 38536
rect 9232 38409 9260 38508
rect 10134 38496 10140 38508
rect 10192 38496 10198 38548
rect 10226 38496 10232 38548
rect 10284 38496 10290 38548
rect 18601 38539 18659 38545
rect 18601 38505 18613 38539
rect 18647 38536 18659 38539
rect 19518 38536 19524 38548
rect 18647 38508 19524 38536
rect 18647 38505 18659 38508
rect 18601 38499 18659 38505
rect 19518 38496 19524 38508
rect 19576 38496 19582 38548
rect 19705 38539 19763 38545
rect 19705 38505 19717 38539
rect 19751 38536 19763 38539
rect 20530 38536 20536 38548
rect 19751 38508 20536 38536
rect 19751 38505 19763 38508
rect 19705 38499 19763 38505
rect 20530 38496 20536 38508
rect 20588 38496 20594 38548
rect 22649 38539 22707 38545
rect 22649 38505 22661 38539
rect 22695 38536 22707 38539
rect 23198 38536 23204 38548
rect 22695 38508 23204 38536
rect 22695 38505 22707 38508
rect 22649 38499 22707 38505
rect 23198 38496 23204 38508
rect 23256 38496 23262 38548
rect 10152 38468 10180 38496
rect 10410 38468 10416 38480
rect 10152 38440 10416 38468
rect 10410 38428 10416 38440
rect 10468 38428 10474 38480
rect 10778 38428 10784 38480
rect 10836 38468 10842 38480
rect 10962 38468 10968 38480
rect 10836 38440 10968 38468
rect 10836 38428 10842 38440
rect 10962 38428 10968 38440
rect 11020 38428 11026 38480
rect 7699 38372 8064 38400
rect 9217 38403 9275 38409
rect 7699 38369 7711 38372
rect 7653 38363 7711 38369
rect 9217 38369 9229 38403
rect 9263 38369 9275 38403
rect 9217 38363 9275 38369
rect 10226 38360 10232 38412
rect 10284 38400 10290 38412
rect 22002 38400 22008 38412
rect 10284 38372 22008 38400
rect 10284 38360 10290 38372
rect 22002 38360 22008 38372
rect 22060 38360 22066 38412
rect 6454 38292 6460 38344
rect 6512 38292 6518 38344
rect 6641 38335 6699 38341
rect 6641 38301 6653 38335
rect 6687 38301 6699 38335
rect 6641 38295 6699 38301
rect 6656 38264 6684 38295
rect 7466 38292 7472 38344
rect 7524 38341 7530 38344
rect 7524 38335 7552 38341
rect 7540 38301 7552 38335
rect 7524 38295 7552 38301
rect 7524 38292 7530 38295
rect 8570 38292 8576 38344
rect 8628 38332 8634 38344
rect 9125 38335 9183 38341
rect 9125 38332 9137 38335
rect 8628 38304 9137 38332
rect 8628 38292 8634 38304
rect 9125 38301 9137 38304
rect 9171 38301 9183 38335
rect 9490 38332 9496 38344
rect 9451 38304 9496 38332
rect 9125 38295 9183 38301
rect 9490 38292 9496 38304
rect 9548 38292 9554 38344
rect 18785 38335 18843 38341
rect 18785 38332 18797 38335
rect 9646 38304 18797 38332
rect 5736 38236 6684 38264
rect 8202 38224 8208 38276
rect 8260 38264 8266 38276
rect 8260 38236 9444 38264
rect 8260 38224 8266 38236
rect 3602 38196 3608 38208
rect 2700 38168 3608 38196
rect 3602 38156 3608 38168
rect 3660 38156 3666 38208
rect 3970 38156 3976 38208
rect 4028 38196 4034 38208
rect 7190 38196 7196 38208
rect 4028 38168 7196 38196
rect 4028 38156 4034 38168
rect 7190 38156 7196 38168
rect 7248 38156 7254 38208
rect 8941 38199 8999 38205
rect 8941 38165 8953 38199
rect 8987 38196 8999 38199
rect 9214 38196 9220 38208
rect 8987 38168 9220 38196
rect 8987 38165 8999 38168
rect 8941 38159 8999 38165
rect 9214 38156 9220 38168
rect 9272 38156 9278 38208
rect 9416 38196 9444 38236
rect 9646 38196 9674 38304
rect 18785 38301 18797 38304
rect 18831 38301 18843 38335
rect 18785 38295 18843 38301
rect 19889 38335 19947 38341
rect 19889 38301 19901 38335
rect 19935 38301 19947 38335
rect 19889 38295 19947 38301
rect 15470 38224 15476 38276
rect 15528 38264 15534 38276
rect 19904 38264 19932 38295
rect 22830 38292 22836 38344
rect 22888 38292 22894 38344
rect 23934 38292 23940 38344
rect 23992 38292 23998 38344
rect 15528 38236 19932 38264
rect 15528 38224 15534 38236
rect 9416 38168 9674 38196
rect 24121 38199 24179 38205
rect 24121 38165 24133 38199
rect 24167 38196 24179 38199
rect 24854 38196 24860 38208
rect 24167 38168 24860 38196
rect 24167 38165 24179 38168
rect 24121 38159 24179 38165
rect 24854 38156 24860 38168
rect 24912 38156 24918 38208
rect 1104 38106 24723 38128
rect 1104 38054 6814 38106
rect 6866 38054 6878 38106
rect 6930 38054 6942 38106
rect 6994 38054 7006 38106
rect 7058 38054 7070 38106
rect 7122 38054 12679 38106
rect 12731 38054 12743 38106
rect 12795 38054 12807 38106
rect 12859 38054 12871 38106
rect 12923 38054 12935 38106
rect 12987 38054 18544 38106
rect 18596 38054 18608 38106
rect 18660 38054 18672 38106
rect 18724 38054 18736 38106
rect 18788 38054 18800 38106
rect 18852 38054 24409 38106
rect 24461 38054 24473 38106
rect 24525 38054 24537 38106
rect 24589 38054 24601 38106
rect 24653 38054 24665 38106
rect 24717 38054 24723 38106
rect 1104 38032 24723 38054
rect 14 37952 20 38004
rect 72 37992 78 38004
rect 3970 37992 3976 38004
rect 72 37964 3976 37992
rect 72 37952 78 37964
rect 3970 37952 3976 37964
rect 4028 37952 4034 38004
rect 4062 37952 4068 38004
rect 4120 37992 4126 38004
rect 4120 37964 5580 37992
rect 4120 37952 4126 37964
rect 2314 37884 2320 37936
rect 2372 37924 2378 37936
rect 2372 37896 3556 37924
rect 2372 37884 2378 37896
rect 1763 37859 1821 37865
rect 1763 37825 1775 37859
rect 1809 37856 1821 37859
rect 2590 37856 2596 37868
rect 1809 37828 2596 37856
rect 1809 37825 1821 37828
rect 1763 37819 1821 37825
rect 2590 37816 2596 37828
rect 2648 37816 2654 37868
rect 3142 37816 3148 37868
rect 3200 37856 3206 37868
rect 3235 37859 3293 37865
rect 3235 37856 3247 37859
rect 3200 37828 3247 37856
rect 3200 37816 3206 37828
rect 3235 37825 3247 37828
rect 3281 37825 3293 37859
rect 3528 37856 3556 37896
rect 3602 37884 3608 37936
rect 3660 37924 3666 37936
rect 5166 37924 5172 37936
rect 3660 37896 5172 37924
rect 3660 37884 3666 37896
rect 5166 37884 5172 37896
rect 5224 37884 5230 37936
rect 4341 37859 4399 37865
rect 3528 37828 4108 37856
rect 3235 37819 3293 37825
rect 1486 37748 1492 37800
rect 1544 37748 1550 37800
rect 2961 37791 3019 37797
rect 2961 37757 2973 37791
rect 3007 37757 3019 37791
rect 2961 37751 3019 37757
rect 2501 37655 2559 37661
rect 2501 37621 2513 37655
rect 2547 37652 2559 37655
rect 2590 37652 2596 37664
rect 2547 37624 2596 37652
rect 2547 37621 2559 37624
rect 2501 37615 2559 37621
rect 2590 37612 2596 37624
rect 2648 37612 2654 37664
rect 2976 37652 3004 37751
rect 3234 37652 3240 37664
rect 2976 37624 3240 37652
rect 3234 37612 3240 37624
rect 3292 37612 3298 37664
rect 3418 37612 3424 37664
rect 3476 37652 3482 37664
rect 3973 37655 4031 37661
rect 3973 37652 3985 37655
rect 3476 37624 3985 37652
rect 3476 37612 3482 37624
rect 3973 37621 3985 37624
rect 4019 37621 4031 37655
rect 4080 37652 4108 37828
rect 4341 37825 4353 37859
rect 4387 37856 4399 37859
rect 4522 37856 4528 37868
rect 4387 37828 4528 37856
rect 4387 37825 4399 37828
rect 4341 37819 4399 37825
rect 4522 37816 4528 37828
rect 4580 37816 4586 37868
rect 4615 37859 4673 37865
rect 4615 37825 4627 37859
rect 4661 37856 4673 37859
rect 5552 37856 5580 37964
rect 5626 37952 5632 38004
rect 5684 37952 5690 38004
rect 9398 37952 9404 38004
rect 9456 37952 9462 38004
rect 21913 37995 21971 38001
rect 21913 37961 21925 37995
rect 21959 37992 21971 37995
rect 22830 37992 22836 38004
rect 21959 37964 22836 37992
rect 21959 37961 21971 37964
rect 21913 37955 21971 37961
rect 22830 37952 22836 37964
rect 22888 37952 22894 38004
rect 23382 37952 23388 38004
rect 23440 37952 23446 38004
rect 23661 37995 23719 38001
rect 23661 37961 23673 37995
rect 23707 37992 23719 37995
rect 23934 37992 23940 38004
rect 23707 37964 23940 37992
rect 23707 37961 23719 37964
rect 23661 37955 23719 37961
rect 23934 37952 23940 37964
rect 23992 37952 23998 38004
rect 5644 37924 5672 37952
rect 5644 37896 11818 37924
rect 8631 37859 8689 37865
rect 8631 37856 8643 37859
rect 4661 37828 5488 37856
rect 5552 37828 8643 37856
rect 4661 37825 4673 37828
rect 4615 37819 4673 37825
rect 5460 37788 5488 37828
rect 8631 37825 8643 37828
rect 8677 37856 8689 37859
rect 11330 37856 11336 37868
rect 8677 37828 11336 37856
rect 8677 37825 8689 37828
rect 8631 37819 8689 37825
rect 11330 37816 11336 37828
rect 11388 37816 11394 37868
rect 11790 37865 11818 37896
rect 11790 37859 11849 37865
rect 11790 37828 11803 37859
rect 11791 37825 11803 37828
rect 11837 37856 11849 37859
rect 15470 37856 15476 37868
rect 11837 37828 15476 37856
rect 11837 37825 11849 37828
rect 11791 37819 11849 37825
rect 15470 37816 15476 37828
rect 15528 37816 15534 37868
rect 22097 37859 22155 37865
rect 22097 37825 22109 37859
rect 22143 37825 22155 37859
rect 22097 37819 22155 37825
rect 5718 37788 5724 37800
rect 5460 37760 5724 37788
rect 5718 37748 5724 37760
rect 5776 37748 5782 37800
rect 7650 37748 7656 37800
rect 7708 37748 7714 37800
rect 8389 37791 8447 37797
rect 8389 37757 8401 37791
rect 8435 37757 8447 37791
rect 8389 37751 8447 37757
rect 11517 37791 11575 37797
rect 11517 37757 11529 37791
rect 11563 37757 11575 37791
rect 11517 37751 11575 37757
rect 7668 37720 7696 37748
rect 5000 37692 7696 37720
rect 5000 37652 5028 37692
rect 4080 37624 5028 37652
rect 3973 37615 4031 37621
rect 5350 37612 5356 37664
rect 5408 37612 5414 37664
rect 5442 37612 5448 37664
rect 5500 37652 5506 37664
rect 7650 37652 7656 37664
rect 5500 37624 7656 37652
rect 5500 37612 5506 37624
rect 7650 37612 7656 37624
rect 7708 37612 7714 37664
rect 8404 37652 8432 37751
rect 11532 37664 11560 37751
rect 13538 37748 13544 37800
rect 13596 37748 13602 37800
rect 13814 37748 13820 37800
rect 13872 37788 13878 37800
rect 22112 37788 22140 37819
rect 23566 37816 23572 37868
rect 23624 37816 23630 37868
rect 23845 37859 23903 37865
rect 23845 37825 23857 37859
rect 23891 37825 23903 37859
rect 23845 37819 23903 37825
rect 23937 37859 23995 37865
rect 23937 37825 23949 37859
rect 23983 37825 23995 37859
rect 23937 37819 23995 37825
rect 13872 37760 22140 37788
rect 13872 37748 13878 37760
rect 23382 37748 23388 37800
rect 23440 37788 23446 37800
rect 23860 37788 23888 37819
rect 23440 37760 23888 37788
rect 23440 37748 23446 37760
rect 13556 37720 13584 37748
rect 12176 37692 13584 37720
rect 9122 37652 9128 37664
rect 8404 37624 9128 37652
rect 9122 37612 9128 37624
rect 9180 37612 9186 37664
rect 11514 37612 11520 37664
rect 11572 37652 11578 37664
rect 12176 37652 12204 37692
rect 23014 37680 23020 37732
rect 23072 37720 23078 37732
rect 23952 37720 23980 37819
rect 23072 37692 23980 37720
rect 23072 37680 23078 37692
rect 11572 37624 12204 37652
rect 11572 37612 11578 37624
rect 12526 37612 12532 37664
rect 12584 37612 12590 37664
rect 24118 37612 24124 37664
rect 24176 37612 24182 37664
rect 1104 37562 24564 37584
rect 1104 37510 3882 37562
rect 3934 37510 3946 37562
rect 3998 37510 4010 37562
rect 4062 37510 4074 37562
rect 4126 37510 4138 37562
rect 4190 37510 9747 37562
rect 9799 37510 9811 37562
rect 9863 37510 9875 37562
rect 9927 37510 9939 37562
rect 9991 37510 10003 37562
rect 10055 37510 15612 37562
rect 15664 37510 15676 37562
rect 15728 37510 15740 37562
rect 15792 37510 15804 37562
rect 15856 37510 15868 37562
rect 15920 37510 21477 37562
rect 21529 37510 21541 37562
rect 21593 37510 21605 37562
rect 21657 37510 21669 37562
rect 21721 37510 21733 37562
rect 21785 37510 24564 37562
rect 1104 37488 24564 37510
rect 1854 37408 1860 37460
rect 1912 37448 1918 37460
rect 3237 37451 3295 37457
rect 3237 37448 3249 37451
rect 1912 37420 3249 37448
rect 1912 37408 1918 37420
rect 3237 37417 3249 37420
rect 3283 37417 3295 37451
rect 3237 37411 3295 37417
rect 4522 37408 4528 37460
rect 4580 37448 4586 37460
rect 4982 37448 4988 37460
rect 4580 37420 4988 37448
rect 4580 37408 4586 37420
rect 4982 37408 4988 37420
rect 5040 37408 5046 37460
rect 6178 37408 6184 37460
rect 6236 37448 6242 37460
rect 10502 37448 10508 37460
rect 6236 37420 10508 37448
rect 6236 37408 6242 37420
rect 10502 37408 10508 37420
rect 10560 37408 10566 37460
rect 23382 37408 23388 37460
rect 23440 37408 23446 37460
rect 23566 37408 23572 37460
rect 23624 37448 23630 37460
rect 23661 37451 23719 37457
rect 23661 37448 23673 37451
rect 23624 37420 23673 37448
rect 23624 37408 23630 37420
rect 23661 37417 23673 37420
rect 23707 37417 23719 37451
rect 23661 37411 23719 37417
rect 6273 37383 6331 37389
rect 6273 37349 6285 37383
rect 6319 37380 6331 37383
rect 6546 37380 6552 37392
rect 6319 37352 6552 37380
rect 6319 37349 6331 37352
rect 6273 37343 6331 37349
rect 6546 37340 6552 37352
rect 6604 37340 6610 37392
rect 7650 37340 7656 37392
rect 7708 37380 7714 37392
rect 10226 37380 10232 37392
rect 7708 37352 10232 37380
rect 7708 37340 7714 37352
rect 10226 37340 10232 37352
rect 10284 37340 10290 37392
rect 11977 37383 12035 37389
rect 11977 37349 11989 37383
rect 12023 37380 12035 37383
rect 12158 37380 12164 37392
rect 12023 37352 12164 37380
rect 12023 37349 12035 37352
rect 11977 37343 12035 37349
rect 12158 37340 12164 37352
rect 12216 37340 12222 37392
rect 21729 37383 21787 37389
rect 21729 37349 21741 37383
rect 21775 37349 21787 37383
rect 21729 37343 21787 37349
rect 1320 37284 1532 37312
rect 658 37204 664 37256
rect 716 37244 722 37256
rect 1320 37244 1348 37284
rect 716 37216 1348 37244
rect 1397 37247 1455 37253
rect 716 37204 722 37216
rect 1397 37213 1409 37247
rect 1443 37213 1455 37247
rect 1504 37244 1532 37284
rect 2038 37272 2044 37324
rect 2096 37272 2102 37324
rect 2314 37272 2320 37324
rect 2372 37272 2378 37324
rect 2406 37272 2412 37324
rect 2464 37321 2470 37324
rect 2464 37315 2492 37321
rect 2480 37281 2492 37315
rect 2464 37275 2492 37281
rect 2464 37272 2470 37275
rect 2590 37272 2596 37324
rect 2648 37272 2654 37324
rect 5442 37272 5448 37324
rect 5500 37272 5506 37324
rect 10962 37272 10968 37324
rect 11020 37272 11026 37324
rect 21744 37312 21772 37343
rect 21744 37284 22048 37312
rect 1581 37247 1639 37253
rect 1581 37244 1593 37247
rect 1504 37216 1593 37244
rect 1397 37207 1455 37213
rect 1581 37213 1593 37216
rect 1627 37213 1639 37247
rect 1581 37207 1639 37213
rect 1412 37108 1440 37207
rect 3234 37204 3240 37256
rect 3292 37244 3298 37256
rect 3789 37247 3847 37253
rect 3789 37244 3801 37247
rect 3292 37216 3801 37244
rect 3292 37204 3298 37216
rect 3789 37213 3801 37216
rect 3835 37213 3847 37247
rect 3789 37207 3847 37213
rect 5074 37204 5080 37256
rect 5132 37244 5138 37256
rect 5261 37247 5319 37253
rect 5261 37244 5273 37247
rect 5132 37216 5273 37244
rect 5132 37204 5138 37216
rect 5261 37213 5273 37216
rect 5307 37244 5319 37247
rect 5307 37216 6040 37244
rect 5307 37213 5319 37216
rect 5261 37207 5319 37213
rect 6012 37188 6040 37216
rect 6914 37204 6920 37256
rect 6972 37204 6978 37256
rect 7191 37247 7249 37253
rect 7191 37244 7203 37247
rect 7022 37216 7203 37244
rect 3970 37136 3976 37188
rect 4028 37176 4034 37188
rect 4065 37179 4123 37185
rect 4065 37176 4077 37179
rect 4028 37148 4077 37176
rect 4028 37136 4034 37148
rect 4065 37145 4077 37148
rect 4111 37145 4123 37179
rect 4065 37139 4123 37145
rect 4890 37136 4896 37188
rect 4948 37176 4954 37188
rect 4985 37179 5043 37185
rect 4985 37176 4997 37179
rect 4948 37148 4997 37176
rect 4948 37136 4954 37148
rect 4985 37145 4997 37148
rect 5031 37145 5043 37179
rect 4985 37139 5043 37145
rect 5350 37136 5356 37188
rect 5408 37136 5414 37188
rect 5626 37136 5632 37188
rect 5684 37176 5690 37188
rect 5721 37179 5779 37185
rect 5721 37176 5733 37179
rect 5684 37148 5733 37176
rect 5684 37136 5690 37148
rect 5721 37145 5733 37148
rect 5767 37176 5779 37179
rect 5902 37176 5908 37188
rect 5767 37148 5908 37176
rect 5767 37145 5779 37148
rect 5721 37139 5779 37145
rect 5902 37136 5908 37148
rect 5960 37136 5966 37188
rect 5994 37136 6000 37188
rect 6052 37136 6058 37188
rect 6086 37136 6092 37188
rect 6144 37136 6150 37188
rect 2498 37108 2504 37120
rect 1412 37080 2504 37108
rect 2498 37068 2504 37080
rect 2556 37068 2562 37120
rect 2590 37068 2596 37120
rect 2648 37108 2654 37120
rect 3878 37108 3884 37120
rect 2648 37080 3884 37108
rect 2648 37068 2654 37080
rect 3878 37068 3884 37080
rect 3936 37068 3942 37120
rect 5258 37068 5264 37120
rect 5316 37108 5322 37120
rect 7022 37108 7050 37216
rect 7191 37213 7203 37216
rect 7237 37244 7249 37247
rect 8846 37244 8852 37256
rect 7237 37216 8852 37244
rect 7237 37213 7249 37216
rect 7191 37207 7249 37213
rect 8846 37204 8852 37216
rect 8904 37204 8910 37256
rect 9214 37204 9220 37256
rect 9272 37244 9278 37256
rect 10226 37244 10232 37256
rect 9272 37216 10232 37244
rect 9272 37204 9278 37216
rect 10226 37204 10232 37216
rect 10284 37204 10290 37256
rect 11057 37247 11115 37253
rect 11057 37213 11069 37247
rect 11103 37244 11115 37247
rect 12526 37244 12532 37256
rect 11103 37216 12532 37244
rect 11103 37213 11115 37216
rect 7466 37136 7472 37188
rect 7524 37176 7530 37188
rect 7742 37176 7748 37188
rect 7524 37148 7748 37176
rect 7524 37136 7530 37148
rect 7742 37136 7748 37148
rect 7800 37136 7806 37188
rect 8018 37136 8024 37188
rect 8076 37176 8082 37188
rect 9398 37176 9404 37188
rect 8076 37148 9404 37176
rect 8076 37136 8082 37148
rect 9398 37136 9404 37148
rect 9456 37136 9462 37188
rect 10612 37185 10730 37210
rect 11057 37207 11115 37213
rect 12526 37204 12532 37216
rect 12584 37204 12590 37256
rect 20990 37204 20996 37256
rect 21048 37204 21054 37256
rect 21910 37204 21916 37256
rect 21968 37204 21974 37256
rect 10612 37182 10747 37185
rect 10612 37176 10640 37182
rect 9646 37148 10640 37176
rect 10689 37179 10747 37182
rect 5316 37080 7050 37108
rect 5316 37068 5322 37080
rect 7926 37068 7932 37120
rect 7984 37068 7990 37120
rect 8202 37068 8208 37120
rect 8260 37108 8266 37120
rect 9646 37108 9674 37148
rect 10689 37145 10701 37179
rect 10735 37145 10747 37179
rect 10689 37139 10747 37145
rect 10778 37136 10784 37188
rect 10836 37176 10842 37188
rect 10965 37179 11023 37185
rect 10965 37176 10977 37179
rect 10836 37148 10977 37176
rect 10836 37136 10842 37148
rect 10965 37145 10977 37148
rect 11011 37145 11023 37179
rect 10965 37139 11023 37145
rect 11422 37136 11428 37188
rect 11480 37136 11486 37188
rect 11793 37179 11851 37185
rect 11793 37145 11805 37179
rect 11839 37145 11851 37179
rect 22020 37176 22048 37284
rect 23860 37284 24072 37312
rect 23566 37204 23572 37256
rect 23624 37204 23630 37256
rect 23860 37253 23888 37284
rect 23845 37247 23903 37253
rect 23845 37213 23857 37247
rect 23891 37213 23903 37247
rect 23845 37207 23903 37213
rect 23937 37247 23995 37253
rect 23937 37213 23949 37247
rect 23983 37213 23995 37247
rect 24044 37244 24072 37284
rect 25590 37244 25596 37256
rect 24044 37216 25596 37244
rect 23937 37207 23995 37213
rect 23952 37176 23980 37207
rect 25590 37204 25596 37216
rect 25648 37204 25654 37256
rect 11793 37139 11851 37145
rect 20824 37148 21864 37176
rect 22020 37148 23980 37176
rect 8260 37080 9674 37108
rect 8260 37068 8266 37080
rect 10502 37068 10508 37120
rect 10560 37108 10566 37120
rect 11808 37108 11836 37139
rect 20824 37117 20852 37148
rect 10560 37080 11836 37108
rect 20809 37111 20867 37117
rect 10560 37068 10566 37080
rect 20809 37077 20821 37111
rect 20855 37077 20867 37111
rect 21836 37108 21864 37148
rect 23014 37108 23020 37120
rect 21836 37080 23020 37108
rect 20809 37071 20867 37077
rect 23014 37068 23020 37080
rect 23072 37068 23078 37120
rect 24121 37111 24179 37117
rect 24121 37077 24133 37111
rect 24167 37108 24179 37111
rect 24854 37108 24860 37120
rect 24167 37080 24860 37108
rect 24167 37077 24179 37080
rect 24121 37071 24179 37077
rect 24854 37068 24860 37080
rect 24912 37068 24918 37120
rect 1104 37018 24723 37040
rect 1104 36966 6814 37018
rect 6866 36966 6878 37018
rect 6930 36966 6942 37018
rect 6994 36966 7006 37018
rect 7058 36966 7070 37018
rect 7122 36966 12679 37018
rect 12731 36966 12743 37018
rect 12795 36966 12807 37018
rect 12859 36966 12871 37018
rect 12923 36966 12935 37018
rect 12987 36966 18544 37018
rect 18596 36966 18608 37018
rect 18660 36966 18672 37018
rect 18724 36966 18736 37018
rect 18788 36966 18800 37018
rect 18852 36966 24409 37018
rect 24461 36966 24473 37018
rect 24525 36966 24537 37018
rect 24589 36966 24601 37018
rect 24653 36966 24665 37018
rect 24717 36966 24723 37018
rect 1104 36944 24723 36966
rect 2038 36864 2044 36916
rect 2096 36904 2102 36916
rect 2409 36907 2467 36913
rect 2409 36904 2421 36907
rect 2096 36876 2421 36904
rect 2096 36864 2102 36876
rect 2409 36873 2421 36876
rect 2455 36873 2467 36907
rect 2409 36867 2467 36873
rect 3050 36864 3056 36916
rect 3108 36864 3114 36916
rect 4890 36864 4896 36916
rect 4948 36904 4954 36916
rect 5258 36904 5264 36916
rect 4948 36876 5264 36904
rect 4948 36864 4954 36876
rect 5258 36864 5264 36876
rect 5316 36864 5322 36916
rect 5350 36864 5356 36916
rect 5408 36904 5414 36916
rect 5905 36907 5963 36913
rect 5905 36904 5917 36907
rect 5408 36876 5917 36904
rect 5408 36864 5414 36876
rect 5905 36873 5917 36876
rect 5951 36873 5963 36907
rect 5905 36867 5963 36873
rect 6270 36864 6276 36916
rect 6328 36904 6334 36916
rect 10502 36904 10508 36916
rect 6328 36876 10508 36904
rect 6328 36864 6334 36876
rect 10502 36864 10508 36876
rect 10560 36864 10566 36916
rect 10962 36864 10968 36916
rect 11020 36864 11026 36916
rect 20165 36907 20223 36913
rect 20165 36873 20177 36907
rect 20211 36904 20223 36907
rect 20990 36904 20996 36916
rect 20211 36876 20996 36904
rect 20211 36873 20223 36876
rect 20165 36867 20223 36873
rect 20990 36864 20996 36876
rect 21048 36864 21054 36916
rect 21910 36864 21916 36916
rect 21968 36864 21974 36916
rect 23566 36904 23572 36916
rect 22066 36876 23572 36904
rect 3068 36836 3096 36864
rect 1686 36808 3096 36836
rect 1686 36777 1714 36808
rect 4154 36796 4160 36848
rect 4212 36796 4218 36848
rect 4430 36796 4436 36848
rect 4488 36836 4494 36848
rect 5074 36836 5080 36848
rect 4488 36808 5080 36836
rect 4488 36796 4494 36808
rect 5074 36796 5080 36808
rect 5132 36796 5138 36848
rect 7098 36796 7104 36848
rect 7156 36836 7162 36848
rect 7466 36836 7472 36848
rect 7156 36808 7472 36836
rect 7156 36796 7162 36808
rect 7466 36796 7472 36808
rect 7524 36796 7530 36848
rect 7558 36796 7564 36848
rect 7616 36836 7622 36848
rect 7745 36839 7803 36845
rect 7745 36836 7757 36839
rect 7616 36808 7757 36836
rect 7616 36796 7622 36808
rect 7745 36805 7757 36808
rect 7791 36805 7803 36839
rect 7745 36799 7803 36805
rect 7837 36839 7895 36845
rect 7837 36805 7849 36839
rect 7883 36836 7895 36839
rect 8386 36836 8392 36848
rect 7883 36808 8392 36836
rect 7883 36805 7895 36808
rect 7837 36799 7895 36805
rect 8386 36796 8392 36808
rect 8444 36796 8450 36848
rect 8573 36839 8631 36845
rect 8573 36805 8585 36839
rect 8619 36836 8631 36839
rect 8662 36836 8668 36848
rect 8619 36808 8668 36836
rect 8619 36805 8631 36808
rect 8573 36799 8631 36805
rect 8662 36796 8668 36808
rect 8720 36796 8726 36848
rect 11514 36836 11520 36848
rect 9968 36808 11520 36836
rect 1671 36771 1729 36777
rect 1671 36737 1683 36771
rect 1717 36737 1729 36771
rect 1671 36731 1729 36737
rect 2774 36728 2780 36780
rect 2832 36728 2838 36780
rect 3050 36728 3056 36780
rect 3108 36768 3114 36780
rect 3329 36771 3387 36777
rect 3329 36768 3341 36771
rect 3108 36740 3341 36768
rect 3108 36728 3114 36740
rect 3329 36737 3341 36740
rect 3375 36737 3387 36771
rect 3329 36731 3387 36737
rect 3602 36728 3608 36780
rect 3660 36768 3666 36780
rect 3881 36771 3939 36777
rect 3881 36768 3893 36771
rect 3660 36740 3893 36768
rect 3660 36728 3666 36740
rect 3881 36737 3893 36740
rect 3927 36737 3939 36771
rect 5166 36768 5172 36780
rect 5127 36740 5172 36768
rect 3881 36731 3939 36737
rect 5166 36728 5172 36740
rect 5224 36728 5230 36780
rect 7374 36728 7380 36780
rect 7432 36768 7438 36780
rect 8202 36768 8208 36780
rect 7432 36740 8208 36768
rect 7432 36728 7438 36740
rect 8202 36728 8208 36740
rect 8260 36728 8266 36780
rect 9122 36728 9128 36780
rect 9180 36768 9186 36780
rect 9968 36777 9996 36808
rect 11514 36796 11520 36808
rect 11572 36796 11578 36848
rect 13814 36796 13820 36848
rect 13872 36796 13878 36848
rect 9953 36771 10011 36777
rect 9953 36768 9965 36771
rect 9180 36740 9965 36768
rect 9180 36728 9186 36740
rect 9953 36737 9965 36740
rect 9999 36737 10011 36771
rect 9953 36731 10011 36737
rect 10134 36728 10140 36780
rect 10192 36768 10198 36780
rect 10227 36771 10285 36777
rect 10227 36768 10239 36771
rect 10192 36740 10239 36768
rect 10192 36728 10198 36740
rect 10227 36737 10239 36740
rect 10273 36768 10285 36771
rect 13832 36768 13860 36796
rect 14182 36768 14188 36780
rect 10273 36740 14188 36768
rect 10273 36737 10285 36740
rect 10227 36731 10285 36737
rect 14182 36728 14188 36740
rect 14240 36728 14246 36780
rect 20346 36728 20352 36780
rect 20404 36728 20410 36780
rect 21177 36771 21235 36777
rect 21177 36737 21189 36771
rect 21223 36737 21235 36771
rect 21177 36731 21235 36737
rect 1394 36660 1400 36712
rect 1452 36660 1458 36712
rect 2961 36703 3019 36709
rect 2961 36669 2973 36703
rect 3007 36669 3019 36703
rect 2961 36663 3019 36669
rect 3513 36703 3571 36709
rect 3513 36669 3525 36703
rect 3559 36669 3571 36703
rect 3513 36663 3571 36669
rect 2590 36632 2596 36644
rect 2424 36604 2596 36632
rect 658 36524 664 36576
rect 716 36564 722 36576
rect 2424 36564 2452 36604
rect 2590 36592 2596 36604
rect 2648 36592 2654 36644
rect 716 36536 2452 36564
rect 2976 36564 3004 36663
rect 3528 36632 3556 36663
rect 3694 36660 3700 36712
rect 3752 36700 3758 36712
rect 3970 36700 3976 36712
rect 3752 36672 3976 36700
rect 3752 36660 3758 36672
rect 3970 36660 3976 36672
rect 4028 36660 4034 36712
rect 4430 36660 4436 36712
rect 4488 36700 4494 36712
rect 4617 36703 4675 36709
rect 4617 36700 4629 36703
rect 4488 36672 4629 36700
rect 4488 36660 4494 36672
rect 4617 36669 4629 36672
rect 4663 36669 4675 36703
rect 4617 36663 4675 36669
rect 4706 36660 4712 36712
rect 4764 36700 4770 36712
rect 4893 36703 4951 36709
rect 4893 36700 4905 36703
rect 4764 36672 4905 36700
rect 4764 36660 4770 36672
rect 4893 36669 4905 36672
rect 4939 36669 4951 36703
rect 4893 36663 4951 36669
rect 7926 36660 7932 36712
rect 7984 36660 7990 36712
rect 18138 36660 18144 36712
rect 18196 36700 18202 36712
rect 21192 36700 21220 36731
rect 18196 36672 21220 36700
rect 18196 36660 18202 36672
rect 3528 36604 5028 36632
rect 4890 36564 4896 36576
rect 2976 36536 4896 36564
rect 716 36524 722 36536
rect 4890 36524 4896 36536
rect 4948 36524 4954 36576
rect 5000 36564 5028 36604
rect 10686 36592 10692 36644
rect 10744 36632 10750 36644
rect 10962 36632 10968 36644
rect 10744 36604 10968 36632
rect 10744 36592 10750 36604
rect 10962 36592 10968 36604
rect 11020 36592 11026 36644
rect 20993 36635 21051 36641
rect 20993 36601 21005 36635
rect 21039 36632 21051 36635
rect 21928 36632 21956 36864
rect 21039 36604 21956 36632
rect 21039 36601 21051 36604
rect 20993 36595 21051 36601
rect 7282 36564 7288 36576
rect 5000 36536 7288 36564
rect 7282 36524 7288 36536
rect 7340 36524 7346 36576
rect 8757 36567 8815 36573
rect 8757 36533 8769 36567
rect 8803 36564 8815 36567
rect 8938 36564 8944 36576
rect 8803 36536 8944 36564
rect 8803 36533 8815 36536
rect 8757 36527 8815 36533
rect 8938 36524 8944 36536
rect 8996 36524 9002 36576
rect 9030 36524 9036 36576
rect 9088 36564 9094 36576
rect 10226 36564 10232 36576
rect 9088 36536 10232 36564
rect 9088 36524 9094 36536
rect 10226 36524 10232 36536
rect 10284 36524 10290 36576
rect 13262 36524 13268 36576
rect 13320 36564 13326 36576
rect 13538 36564 13544 36576
rect 13320 36536 13544 36564
rect 13320 36524 13326 36536
rect 13538 36524 13544 36536
rect 13596 36524 13602 36576
rect 19334 36524 19340 36576
rect 19392 36564 19398 36576
rect 22066 36564 22094 36876
rect 23566 36864 23572 36876
rect 23624 36864 23630 36916
rect 23658 36728 23664 36780
rect 23716 36728 23722 36780
rect 23934 36728 23940 36780
rect 23992 36728 23998 36780
rect 24026 36660 24032 36712
rect 24084 36660 24090 36712
rect 23477 36635 23535 36641
rect 23477 36601 23489 36635
rect 23523 36632 23535 36635
rect 24044 36632 24072 36660
rect 23523 36604 24072 36632
rect 23523 36601 23535 36604
rect 23477 36595 23535 36601
rect 24946 36592 24952 36644
rect 25004 36632 25010 36644
rect 25222 36632 25228 36644
rect 25004 36604 25228 36632
rect 25004 36592 25010 36604
rect 25222 36592 25228 36604
rect 25280 36592 25286 36644
rect 19392 36536 22094 36564
rect 19392 36524 19398 36536
rect 24118 36524 24124 36576
rect 24176 36524 24182 36576
rect 1104 36474 24564 36496
rect 1104 36422 3882 36474
rect 3934 36422 3946 36474
rect 3998 36422 4010 36474
rect 4062 36422 4074 36474
rect 4126 36422 4138 36474
rect 4190 36422 9747 36474
rect 9799 36422 9811 36474
rect 9863 36422 9875 36474
rect 9927 36422 9939 36474
rect 9991 36422 10003 36474
rect 10055 36422 15612 36474
rect 15664 36422 15676 36474
rect 15728 36422 15740 36474
rect 15792 36422 15804 36474
rect 15856 36422 15868 36474
rect 15920 36422 21477 36474
rect 21529 36422 21541 36474
rect 21593 36422 21605 36474
rect 21657 36422 21669 36474
rect 21721 36422 21733 36474
rect 21785 36422 24564 36474
rect 1104 36400 24564 36422
rect 2590 36360 2596 36372
rect 2332 36332 2596 36360
rect 1673 36227 1731 36233
rect 1673 36193 1685 36227
rect 1719 36224 1731 36227
rect 2130 36224 2136 36236
rect 1719 36196 2136 36224
rect 1719 36193 1731 36196
rect 1673 36187 1731 36193
rect 2130 36184 2136 36196
rect 2188 36184 2194 36236
rect 2332 36233 2360 36332
rect 2590 36320 2596 36332
rect 2648 36360 2654 36372
rect 3142 36360 3148 36372
rect 2648 36332 3148 36360
rect 2648 36320 2654 36332
rect 3142 36320 3148 36332
rect 3200 36320 3206 36372
rect 7190 36320 7196 36372
rect 7248 36360 7254 36372
rect 9122 36360 9128 36372
rect 7248 36332 9128 36360
rect 7248 36320 7254 36332
rect 3329 36295 3387 36301
rect 3329 36261 3341 36295
rect 3375 36292 3387 36295
rect 3375 36264 3832 36292
rect 3375 36261 3387 36264
rect 3329 36255 3387 36261
rect 2317 36227 2375 36233
rect 2317 36193 2329 36227
rect 2363 36193 2375 36227
rect 3804 36210 3832 36264
rect 2317 36187 2375 36193
rect 7374 36184 7380 36236
rect 7432 36224 7438 36236
rect 7484 36233 7512 36332
rect 9048 36233 9076 36332
rect 9122 36320 9128 36332
rect 9180 36320 9186 36372
rect 9398 36320 9404 36372
rect 9456 36360 9462 36372
rect 21269 36363 21327 36369
rect 9456 36332 11192 36360
rect 9456 36320 9462 36332
rect 7469 36227 7527 36233
rect 7469 36224 7481 36227
rect 7432 36196 7481 36224
rect 7432 36184 7438 36196
rect 7469 36193 7481 36196
rect 7515 36193 7527 36227
rect 7469 36187 7527 36193
rect 9033 36227 9091 36233
rect 9033 36193 9045 36227
rect 9079 36193 9091 36227
rect 9033 36187 9091 36193
rect 10226 36184 10232 36236
rect 10284 36224 10290 36236
rect 10413 36227 10471 36233
rect 10413 36224 10425 36227
rect 10284 36196 10425 36224
rect 10284 36184 10290 36196
rect 10413 36193 10425 36196
rect 10459 36193 10471 36227
rect 10413 36187 10471 36193
rect 11164 36224 11192 36332
rect 21269 36329 21281 36363
rect 21315 36360 21327 36363
rect 23934 36360 23940 36372
rect 21315 36332 23940 36360
rect 21315 36329 21327 36332
rect 21269 36323 21327 36329
rect 23934 36320 23940 36332
rect 23992 36320 23998 36372
rect 23385 36295 23443 36301
rect 23385 36261 23397 36295
rect 23431 36292 23443 36295
rect 23842 36292 23848 36304
rect 23431 36264 23848 36292
rect 23431 36261 23443 36264
rect 23385 36255 23443 36261
rect 23842 36252 23848 36264
rect 23900 36252 23906 36304
rect 11422 36224 11428 36236
rect 11164 36196 11428 36224
rect 1394 36116 1400 36168
rect 1452 36116 1458 36168
rect 4341 36159 4399 36165
rect 2575 36129 2633 36135
rect 2575 36126 2587 36129
rect 2314 36048 2320 36100
rect 2372 36088 2378 36100
rect 2516 36098 2587 36126
rect 2516 36088 2544 36098
rect 2575 36095 2587 36098
rect 2621 36095 2633 36129
rect 4341 36125 4353 36159
rect 4387 36156 4399 36159
rect 4387 36128 4568 36156
rect 4387 36125 4399 36128
rect 4341 36119 4399 36125
rect 2575 36089 2633 36095
rect 4249 36091 4307 36097
rect 2372 36060 2544 36088
rect 2372 36048 2378 36060
rect 4249 36057 4261 36091
rect 4295 36088 4307 36091
rect 4295 36060 4476 36088
rect 4295 36057 4307 36060
rect 4249 36051 4307 36057
rect 4448 36032 4476 36060
rect 4540 36032 4568 36128
rect 4724 36097 4844 36122
rect 5442 36116 5448 36168
rect 5500 36116 5506 36168
rect 6638 36116 6644 36168
rect 6696 36156 6702 36168
rect 7742 36165 7748 36168
rect 7711 36159 7748 36165
rect 7711 36156 7723 36159
rect 6696 36128 7723 36156
rect 6696 36116 6702 36128
rect 7711 36125 7723 36128
rect 7711 36119 7748 36125
rect 7742 36116 7748 36119
rect 7800 36116 7806 36168
rect 8294 36116 8300 36168
rect 8352 36156 8358 36168
rect 9275 36159 9333 36165
rect 9275 36156 9287 36159
rect 8352 36128 9287 36156
rect 8352 36116 8358 36128
rect 9275 36125 9287 36128
rect 9321 36156 9333 36159
rect 10687 36159 10745 36165
rect 9321 36128 10640 36156
rect 9321 36125 9333 36128
rect 9275 36119 9333 36125
rect 4709 36094 4844 36097
rect 4709 36091 4767 36094
rect 4709 36057 4721 36091
rect 4755 36057 4767 36091
rect 4709 36051 4767 36057
rect 3142 35980 3148 36032
rect 3200 36020 3206 36032
rect 3973 36023 4031 36029
rect 3973 36020 3985 36023
rect 3200 35992 3985 36020
rect 3200 35980 3206 35992
rect 3973 35989 3985 35992
rect 4019 35989 4031 36023
rect 3973 35983 4031 35989
rect 4062 35980 4068 36032
rect 4120 36020 4126 36032
rect 4430 36020 4436 36032
rect 4120 35992 4436 36020
rect 4120 35980 4126 35992
rect 4430 35980 4436 35992
rect 4488 35980 4494 36032
rect 4522 35980 4528 36032
rect 4580 35980 4586 36032
rect 4816 36020 4844 36094
rect 5718 36048 5724 36100
rect 5776 36088 5782 36100
rect 10612 36088 10640 36128
rect 10687 36125 10699 36159
rect 10733 36156 10745 36159
rect 11164 36156 11192 36196
rect 11422 36184 11428 36196
rect 11480 36184 11486 36236
rect 19978 36224 19984 36236
rect 19306 36196 19984 36224
rect 10733 36128 11192 36156
rect 10733 36125 10745 36128
rect 10687 36119 10745 36125
rect 14550 36116 14556 36168
rect 14608 36116 14614 36168
rect 14737 36159 14795 36165
rect 14737 36125 14749 36159
rect 14783 36156 14795 36159
rect 15010 36156 15016 36168
rect 14783 36128 15016 36156
rect 14783 36125 14795 36128
rect 14737 36119 14795 36125
rect 15010 36116 15016 36128
rect 15068 36116 15074 36168
rect 10778 36088 10784 36100
rect 5776 36060 10548 36088
rect 10612 36060 10784 36088
rect 5776 36048 5782 36060
rect 4890 36020 4896 36032
rect 4816 35992 4896 36020
rect 4890 35980 4896 35992
rect 4948 35980 4954 36032
rect 5074 35980 5080 36032
rect 5132 35980 5138 36032
rect 5261 36023 5319 36029
rect 5261 35989 5273 36023
rect 5307 36020 5319 36023
rect 5442 36020 5448 36032
rect 5307 35992 5448 36020
rect 5307 35989 5319 35992
rect 5261 35983 5319 35989
rect 5442 35980 5448 35992
rect 5500 35980 5506 36032
rect 8478 35980 8484 36032
rect 8536 35980 8542 36032
rect 9766 35980 9772 36032
rect 9824 36020 9830 36032
rect 10045 36023 10103 36029
rect 10045 36020 10057 36023
rect 9824 35992 10057 36020
rect 9824 35980 9830 35992
rect 10045 35989 10057 35992
rect 10091 35989 10103 36023
rect 10520 36020 10548 36060
rect 10778 36048 10784 36060
rect 10836 36048 10842 36100
rect 13170 36088 13176 36100
rect 10888 36060 13176 36088
rect 10888 36020 10916 36060
rect 13170 36048 13176 36060
rect 13228 36088 13234 36100
rect 19306 36088 19334 36196
rect 19978 36184 19984 36196
rect 20036 36224 20042 36236
rect 20036 36196 20668 36224
rect 20036 36184 20042 36196
rect 20640 36165 20668 36196
rect 20625 36159 20683 36165
rect 20625 36125 20637 36159
rect 20671 36125 20683 36159
rect 20625 36119 20683 36125
rect 21453 36159 21511 36165
rect 21453 36125 21465 36159
rect 21499 36125 21511 36159
rect 21453 36119 21511 36125
rect 21468 36088 21496 36119
rect 23290 36116 23296 36168
rect 23348 36116 23354 36168
rect 23566 36116 23572 36168
rect 23624 36116 23630 36168
rect 23845 36091 23903 36097
rect 23845 36088 23857 36091
rect 13228 36060 19334 36088
rect 20456 36060 21496 36088
rect 23124 36060 23857 36088
rect 13228 36048 13234 36060
rect 10520 35992 10916 36020
rect 11425 36023 11483 36029
rect 10045 35983 10103 35989
rect 11425 35989 11437 36023
rect 11471 36020 11483 36023
rect 11790 36020 11796 36032
rect 11471 35992 11796 36020
rect 11471 35989 11483 35992
rect 11425 35983 11483 35989
rect 11790 35980 11796 35992
rect 11848 35980 11854 36032
rect 12434 35980 12440 36032
rect 12492 36020 12498 36032
rect 13814 36020 13820 36032
rect 12492 35992 13820 36020
rect 12492 35980 12498 35992
rect 13814 35980 13820 35992
rect 13872 35980 13878 36032
rect 14734 35980 14740 36032
rect 14792 35980 14798 36032
rect 20456 36029 20484 36060
rect 23124 36029 23152 36060
rect 23845 36057 23857 36060
rect 23891 36057 23903 36091
rect 23845 36051 23903 36057
rect 24213 36091 24271 36097
rect 24213 36057 24225 36091
rect 24259 36088 24271 36091
rect 24946 36088 24952 36100
rect 24259 36060 24952 36088
rect 24259 36057 24271 36060
rect 24213 36051 24271 36057
rect 24946 36048 24952 36060
rect 25004 36048 25010 36100
rect 20441 36023 20499 36029
rect 20441 35989 20453 36023
rect 20487 35989 20499 36023
rect 20441 35983 20499 35989
rect 23109 36023 23167 36029
rect 23109 35989 23121 36023
rect 23155 35989 23167 36023
rect 23109 35983 23167 35989
rect 1104 35930 24723 35952
rect 1104 35878 6814 35930
rect 6866 35878 6878 35930
rect 6930 35878 6942 35930
rect 6994 35878 7006 35930
rect 7058 35878 7070 35930
rect 7122 35878 12679 35930
rect 12731 35878 12743 35930
rect 12795 35878 12807 35930
rect 12859 35878 12871 35930
rect 12923 35878 12935 35930
rect 12987 35878 18544 35930
rect 18596 35878 18608 35930
rect 18660 35878 18672 35930
rect 18724 35878 18736 35930
rect 18788 35878 18800 35930
rect 18852 35878 24409 35930
rect 24461 35878 24473 35930
rect 24525 35878 24537 35930
rect 24589 35878 24601 35930
rect 24653 35878 24665 35930
rect 24717 35878 24723 35930
rect 1104 35856 24723 35878
rect 2038 35776 2044 35828
rect 2096 35816 2102 35828
rect 2958 35816 2964 35828
rect 2096 35788 2964 35816
rect 2096 35776 2102 35788
rect 2958 35776 2964 35788
rect 3016 35776 3022 35828
rect 3053 35819 3111 35825
rect 3053 35785 3065 35819
rect 3099 35816 3111 35819
rect 3142 35816 3148 35828
rect 3099 35788 3148 35816
rect 3099 35785 3111 35788
rect 3053 35779 3111 35785
rect 3142 35776 3148 35788
rect 3200 35776 3206 35828
rect 3970 35816 3976 35828
rect 3344 35788 3976 35816
rect 1762 35708 1768 35760
rect 1820 35748 1826 35760
rect 2406 35748 2412 35760
rect 1820 35720 2412 35748
rect 1820 35708 1826 35720
rect 2406 35708 2412 35720
rect 2464 35708 2470 35760
rect 3344 35757 3372 35788
rect 3970 35776 3976 35788
rect 4028 35776 4034 35828
rect 6178 35776 6184 35828
rect 6236 35816 6242 35828
rect 6730 35816 6736 35828
rect 6236 35788 6736 35816
rect 6236 35776 6242 35788
rect 6730 35776 6736 35788
rect 6788 35776 6794 35828
rect 8386 35776 8392 35828
rect 8444 35776 8450 35828
rect 8496 35788 11560 35816
rect 3329 35751 3387 35757
rect 3329 35717 3341 35751
rect 3375 35717 3387 35751
rect 3329 35711 3387 35717
rect 3418 35708 3424 35760
rect 3476 35708 3482 35760
rect 3789 35751 3847 35757
rect 3789 35717 3801 35751
rect 3835 35748 3847 35751
rect 4982 35748 4988 35760
rect 3835 35720 4988 35748
rect 3835 35717 3847 35720
rect 3789 35711 3847 35717
rect 4982 35708 4988 35720
rect 5040 35748 5046 35760
rect 8496 35748 8524 35788
rect 5040 35720 8524 35748
rect 5040 35708 5046 35720
rect 8938 35708 8944 35760
rect 8996 35708 9002 35760
rect 9309 35751 9367 35757
rect 9309 35717 9321 35751
rect 9355 35748 9367 35751
rect 9766 35748 9772 35760
rect 9355 35720 9772 35748
rect 9355 35717 9367 35720
rect 9309 35711 9367 35717
rect 9766 35708 9772 35720
rect 9824 35708 9830 35760
rect 10042 35708 10048 35760
rect 10100 35748 10106 35760
rect 10100 35720 11466 35748
rect 10100 35708 10106 35720
rect 1671 35683 1729 35689
rect 1671 35649 1683 35683
rect 1717 35680 1729 35683
rect 2958 35680 2964 35692
rect 1717 35652 2964 35680
rect 1717 35649 1729 35652
rect 1671 35643 1729 35649
rect 2958 35640 2964 35652
rect 3016 35640 3022 35692
rect 4181 35683 4239 35689
rect 4181 35649 4193 35683
rect 4227 35680 4239 35683
rect 5074 35680 5080 35692
rect 4227 35652 5080 35680
rect 4227 35649 4239 35652
rect 4181 35643 4239 35649
rect 5074 35640 5080 35652
rect 5132 35640 5138 35692
rect 5167 35683 5225 35689
rect 5167 35649 5179 35683
rect 5213 35680 5225 35683
rect 5258 35680 5264 35692
rect 5213 35652 5264 35680
rect 5213 35649 5225 35652
rect 5167 35643 5225 35649
rect 5258 35640 5264 35652
rect 5316 35640 5322 35692
rect 7282 35640 7288 35692
rect 7340 35680 7346 35692
rect 7650 35689 7656 35692
rect 7619 35683 7656 35689
rect 7619 35680 7631 35683
rect 7340 35652 7631 35680
rect 7340 35640 7346 35652
rect 7619 35649 7631 35652
rect 7619 35643 7656 35649
rect 7650 35640 7656 35643
rect 7708 35640 7714 35692
rect 9214 35680 9220 35692
rect 8036 35652 9220 35680
rect 1397 35615 1455 35621
rect 1397 35581 1409 35615
rect 1443 35581 1455 35615
rect 1397 35575 1455 35581
rect 1412 35544 1440 35575
rect 3326 35572 3332 35624
rect 3384 35572 3390 35624
rect 4798 35572 4804 35624
rect 4856 35612 4862 35624
rect 4893 35615 4951 35621
rect 4893 35612 4905 35615
rect 4856 35584 4905 35612
rect 4856 35572 4862 35584
rect 4893 35581 4905 35584
rect 4939 35581 4951 35615
rect 4893 35575 4951 35581
rect 7374 35572 7380 35624
rect 7432 35572 7438 35624
rect 1412 35516 1532 35544
rect 1504 35488 1532 35516
rect 5828 35516 7512 35544
rect 1486 35436 1492 35488
rect 1544 35436 1550 35488
rect 2406 35436 2412 35488
rect 2464 35436 2470 35488
rect 4338 35436 4344 35488
rect 4396 35476 4402 35488
rect 5828 35476 5856 35516
rect 4396 35448 5856 35476
rect 4396 35436 4402 35448
rect 5902 35436 5908 35488
rect 5960 35436 5966 35488
rect 7484 35476 7512 35516
rect 8036 35476 8064 35652
rect 9214 35640 9220 35652
rect 9272 35640 9278 35692
rect 9677 35683 9735 35689
rect 9677 35649 9689 35683
rect 9723 35680 9735 35683
rect 10134 35680 10140 35692
rect 9723 35652 10140 35680
rect 9723 35649 9735 35652
rect 9677 35643 9735 35649
rect 10134 35640 10140 35652
rect 10192 35640 10198 35692
rect 10226 35640 10232 35692
rect 10284 35680 10290 35692
rect 10686 35680 10692 35692
rect 10284 35652 10692 35680
rect 10284 35640 10290 35652
rect 10686 35640 10692 35652
rect 10744 35640 10750 35692
rect 8478 35572 8484 35624
rect 8536 35612 8542 35624
rect 11333 35615 11391 35621
rect 8536 35584 8786 35612
rect 8536 35572 8542 35584
rect 11333 35581 11345 35615
rect 11379 35581 11391 35615
rect 11438 35612 11466 35720
rect 11532 35689 11560 35788
rect 13630 35776 13636 35828
rect 13688 35776 13694 35828
rect 14461 35819 14519 35825
rect 14461 35785 14473 35819
rect 14507 35816 14519 35819
rect 14550 35816 14556 35828
rect 14507 35788 14556 35816
rect 14507 35785 14519 35788
rect 14461 35779 14519 35785
rect 14550 35776 14556 35788
rect 14608 35776 14614 35828
rect 14918 35776 14924 35828
rect 14976 35816 14982 35828
rect 15105 35819 15163 35825
rect 15105 35816 15117 35819
rect 14976 35788 15117 35816
rect 14976 35776 14982 35788
rect 15105 35785 15117 35788
rect 15151 35785 15163 35819
rect 15105 35779 15163 35785
rect 21821 35819 21879 35825
rect 21821 35785 21833 35819
rect 21867 35816 21879 35819
rect 22554 35816 22560 35828
rect 21867 35788 22560 35816
rect 21867 35785 21879 35788
rect 21821 35779 21879 35785
rect 22554 35776 22560 35788
rect 22612 35776 22618 35828
rect 22649 35819 22707 35825
rect 22649 35785 22661 35819
rect 22695 35816 22707 35819
rect 23290 35816 23296 35828
rect 22695 35788 23296 35816
rect 22695 35785 22707 35788
rect 22649 35779 22707 35785
rect 23290 35776 23296 35788
rect 23348 35776 23354 35828
rect 23658 35776 23664 35828
rect 23716 35776 23722 35828
rect 24210 35816 24216 35828
rect 23768 35788 24216 35816
rect 11517 35683 11575 35689
rect 11517 35649 11529 35683
rect 11563 35649 11575 35683
rect 11517 35643 11575 35649
rect 13449 35683 13507 35689
rect 13449 35649 13461 35683
rect 13495 35680 13507 35683
rect 13648 35680 13676 35776
rect 13814 35748 13820 35760
rect 13740 35720 13820 35748
rect 13740 35719 13768 35720
rect 13495 35652 13676 35680
rect 13707 35713 13768 35719
rect 13707 35679 13719 35713
rect 13753 35682 13768 35713
rect 13814 35708 13820 35720
rect 13872 35708 13878 35760
rect 13753 35679 13765 35682
rect 13707 35673 13765 35679
rect 14568 35680 14596 35776
rect 23768 35748 23796 35788
rect 24210 35776 24216 35788
rect 24268 35776 24274 35828
rect 22940 35720 23796 35748
rect 23860 35720 24072 35748
rect 14829 35683 14887 35689
rect 14829 35680 14841 35683
rect 14568 35652 14841 35680
rect 13495 35649 13507 35652
rect 13449 35643 13507 35649
rect 14829 35649 14841 35652
rect 14875 35649 14887 35683
rect 14829 35643 14887 35649
rect 14918 35640 14924 35692
rect 14976 35680 14982 35692
rect 15197 35683 15255 35689
rect 15197 35680 15209 35683
rect 14976 35652 15209 35680
rect 14976 35640 14982 35652
rect 15197 35649 15209 35652
rect 15243 35649 15255 35683
rect 15197 35643 15255 35649
rect 19334 35640 19340 35692
rect 19392 35680 19398 35692
rect 20533 35683 20591 35689
rect 20533 35680 20545 35683
rect 19392 35652 20545 35680
rect 19392 35640 19398 35652
rect 20533 35649 20545 35652
rect 20579 35649 20591 35683
rect 20533 35643 20591 35649
rect 22005 35683 22063 35689
rect 22005 35649 22017 35683
rect 22051 35649 22063 35683
rect 22005 35643 22063 35649
rect 11701 35615 11759 35621
rect 11701 35612 11713 35615
rect 11438 35584 11713 35612
rect 11333 35575 11391 35581
rect 11701 35581 11713 35584
rect 11747 35581 11759 35615
rect 11701 35575 11759 35581
rect 10226 35504 10232 35556
rect 10284 35504 10290 35556
rect 11348 35544 11376 35575
rect 11790 35572 11796 35624
rect 11848 35612 11854 35624
rect 12161 35615 12219 35621
rect 12161 35612 12173 35615
rect 11848 35584 12173 35612
rect 11848 35572 11854 35584
rect 12161 35581 12173 35584
rect 12207 35581 12219 35615
rect 12437 35615 12495 35621
rect 12437 35612 12449 35615
rect 12161 35575 12219 35581
rect 12268 35584 12449 35612
rect 12268 35544 12296 35584
rect 12437 35581 12449 35584
rect 12483 35581 12495 35615
rect 12437 35575 12495 35581
rect 12526 35572 12532 35624
rect 12584 35621 12590 35624
rect 12584 35615 12612 35621
rect 12600 35581 12612 35615
rect 12584 35575 12612 35581
rect 12584 35572 12590 35575
rect 12710 35572 12716 35624
rect 12768 35572 12774 35624
rect 14734 35572 14740 35624
rect 14792 35612 14798 35624
rect 15105 35615 15163 35621
rect 15105 35612 15117 35615
rect 14792 35584 15117 35612
rect 14792 35572 14798 35584
rect 15105 35581 15117 35584
rect 15151 35581 15163 35615
rect 15105 35575 15163 35581
rect 17218 35572 17224 35624
rect 17276 35612 17282 35624
rect 22020 35612 22048 35643
rect 22554 35640 22560 35692
rect 22612 35640 22618 35692
rect 22830 35640 22836 35692
rect 22888 35640 22894 35692
rect 22940 35612 22968 35720
rect 23198 35640 23204 35692
rect 23256 35680 23262 35692
rect 23860 35689 23888 35720
rect 23569 35683 23627 35689
rect 23569 35680 23581 35683
rect 23256 35652 23581 35680
rect 23256 35640 23262 35652
rect 23569 35649 23581 35652
rect 23615 35649 23627 35683
rect 23569 35643 23627 35649
rect 23845 35683 23903 35689
rect 23845 35649 23857 35683
rect 23891 35649 23903 35683
rect 23845 35643 23903 35649
rect 23937 35683 23995 35689
rect 23937 35649 23949 35683
rect 23983 35649 23995 35683
rect 23937 35643 23995 35649
rect 23952 35612 23980 35643
rect 17276 35584 22048 35612
rect 22296 35584 22968 35612
rect 23124 35584 23980 35612
rect 17276 35572 17282 35584
rect 11348 35516 12296 35544
rect 14921 35547 14979 35553
rect 14921 35513 14933 35547
rect 14967 35544 14979 35547
rect 15289 35547 15347 35553
rect 15289 35544 15301 35547
rect 14967 35516 15301 35544
rect 14967 35513 14979 35516
rect 14921 35507 14979 35513
rect 15289 35513 15301 35516
rect 15335 35513 15347 35547
rect 15289 35507 15347 35513
rect 20364 35516 21956 35544
rect 7484 35448 8064 35476
rect 13357 35479 13415 35485
rect 13357 35445 13369 35479
rect 13403 35476 13415 35479
rect 17310 35476 17316 35488
rect 13403 35448 17316 35476
rect 13403 35445 13415 35448
rect 13357 35439 13415 35445
rect 17310 35436 17316 35448
rect 17368 35436 17374 35488
rect 20364 35485 20392 35516
rect 20349 35479 20407 35485
rect 20349 35445 20361 35479
rect 20395 35445 20407 35479
rect 21928 35476 21956 35516
rect 22296 35476 22324 35584
rect 21928 35448 22324 35476
rect 22373 35479 22431 35485
rect 20349 35439 20407 35445
rect 22373 35445 22385 35479
rect 22419 35476 22431 35479
rect 23124 35476 23152 35584
rect 24044 35544 24072 35720
rect 23308 35516 24072 35544
rect 23308 35488 23336 35516
rect 22419 35448 23152 35476
rect 22419 35445 22431 35448
rect 22373 35439 22431 35445
rect 23290 35436 23296 35488
rect 23348 35436 23354 35488
rect 23382 35436 23388 35488
rect 23440 35436 23446 35488
rect 24118 35436 24124 35488
rect 24176 35436 24182 35488
rect 1104 35386 24564 35408
rect 1104 35334 3882 35386
rect 3934 35334 3946 35386
rect 3998 35334 4010 35386
rect 4062 35334 4074 35386
rect 4126 35334 4138 35386
rect 4190 35334 9747 35386
rect 9799 35334 9811 35386
rect 9863 35334 9875 35386
rect 9927 35334 9939 35386
rect 9991 35334 10003 35386
rect 10055 35334 15612 35386
rect 15664 35334 15676 35386
rect 15728 35334 15740 35386
rect 15792 35334 15804 35386
rect 15856 35334 15868 35386
rect 15920 35334 21477 35386
rect 21529 35334 21541 35386
rect 21593 35334 21605 35386
rect 21657 35334 21669 35386
rect 21721 35334 21733 35386
rect 21785 35334 24564 35386
rect 1104 35312 24564 35334
rect 2406 35232 2412 35284
rect 2464 35232 2470 35284
rect 2958 35232 2964 35284
rect 3016 35272 3022 35284
rect 3326 35272 3332 35284
rect 3016 35244 3332 35272
rect 3016 35232 3022 35244
rect 3326 35232 3332 35244
rect 3384 35272 3390 35284
rect 3602 35272 3608 35284
rect 3384 35244 3608 35272
rect 3384 35232 3390 35244
rect 3602 35232 3608 35244
rect 3660 35232 3666 35284
rect 11514 35272 11520 35284
rect 6564 35244 8984 35272
rect 2317 35207 2375 35213
rect 2317 35173 2329 35207
rect 2363 35204 2375 35207
rect 2424 35204 2452 35232
rect 2363 35176 2452 35204
rect 2363 35173 2375 35176
rect 2317 35167 2375 35173
rect 2406 35096 2412 35148
rect 2464 35136 2470 35148
rect 2593 35139 2651 35145
rect 2593 35136 2605 35139
rect 2464 35108 2605 35136
rect 2464 35096 2470 35108
rect 2593 35105 2605 35108
rect 2639 35105 2651 35139
rect 2593 35099 2651 35105
rect 2710 35139 2768 35145
rect 2710 35105 2722 35139
rect 2756 35136 2768 35139
rect 2756 35108 5028 35136
rect 2756 35105 2768 35108
rect 2710 35099 2768 35105
rect 1673 35071 1731 35077
rect 1673 35037 1685 35071
rect 1719 35068 1731 35071
rect 1762 35068 1768 35080
rect 1719 35040 1768 35068
rect 1719 35037 1731 35040
rect 1673 35031 1731 35037
rect 1762 35028 1768 35040
rect 1820 35028 1826 35080
rect 1857 35071 1915 35077
rect 1857 35037 1869 35071
rect 1903 35037 1915 35071
rect 1857 35031 1915 35037
rect 1872 34932 1900 35031
rect 2866 35028 2872 35080
rect 2924 35028 2930 35080
rect 3510 35028 3516 35080
rect 3568 35028 3574 35080
rect 3602 35028 3608 35080
rect 3660 35028 3666 35080
rect 3786 35028 3792 35080
rect 3844 35028 3850 35080
rect 3878 35028 3884 35080
rect 3936 35068 3942 35080
rect 4341 35071 4399 35077
rect 4341 35068 4353 35071
rect 3936 35040 4353 35068
rect 3936 35028 3942 35040
rect 4341 35037 4353 35040
rect 4387 35037 4399 35071
rect 5000 35068 5028 35108
rect 5718 35096 5724 35148
rect 5776 35096 5782 35148
rect 5629 35071 5687 35077
rect 5000 35040 5488 35068
rect 4341 35031 4399 35037
rect 3620 35000 3648 35028
rect 5460 35012 5488 35040
rect 5629 35037 5641 35071
rect 5675 35068 5687 35071
rect 5902 35068 5908 35080
rect 5675 35040 5908 35068
rect 5675 35037 5687 35040
rect 5629 35031 5687 35037
rect 5902 35028 5908 35040
rect 5960 35028 5966 35080
rect 5994 35028 6000 35080
rect 6052 35028 6058 35080
rect 6564 35068 6592 35244
rect 8956 35216 8984 35244
rect 11164 35244 11520 35272
rect 7834 35204 7840 35216
rect 7668 35176 7840 35204
rect 6472 35040 6592 35068
rect 4065 35003 4123 35009
rect 4065 35000 4077 35003
rect 3620 34972 4077 35000
rect 4065 34969 4077 34972
rect 4111 34969 4123 35003
rect 4065 34963 4123 34969
rect 4614 34960 4620 35012
rect 4672 34960 4678 35012
rect 5442 34960 5448 35012
rect 5500 35000 5506 35012
rect 5537 35003 5595 35009
rect 5537 35000 5549 35003
rect 5500 34972 5549 35000
rect 5500 34960 5506 34972
rect 5537 34969 5549 34972
rect 5583 35000 5595 35003
rect 6472 35000 6500 35040
rect 6638 35028 6644 35080
rect 6696 35068 6702 35080
rect 6733 35071 6791 35077
rect 6733 35068 6745 35071
rect 6696 35040 6745 35068
rect 6696 35028 6702 35040
rect 6733 35037 6745 35040
rect 6779 35037 6791 35071
rect 6733 35031 6791 35037
rect 7007 35071 7065 35077
rect 7007 35037 7019 35071
rect 7053 35068 7065 35071
rect 7668 35068 7696 35176
rect 7834 35164 7840 35176
rect 7892 35164 7898 35216
rect 8938 35164 8944 35216
rect 8996 35164 9002 35216
rect 10686 35096 10692 35148
rect 10744 35136 10750 35148
rect 11164 35145 11192 35244
rect 11514 35232 11520 35244
rect 11572 35232 11578 35284
rect 12161 35275 12219 35281
rect 12161 35241 12173 35275
rect 12207 35272 12219 35275
rect 12710 35272 12716 35284
rect 12207 35244 12716 35272
rect 12207 35241 12219 35244
rect 12161 35235 12219 35241
rect 12710 35232 12716 35244
rect 12768 35232 12774 35284
rect 14737 35275 14795 35281
rect 14737 35241 14749 35275
rect 14783 35272 14795 35275
rect 14918 35272 14924 35284
rect 14783 35244 14924 35272
rect 14783 35241 14795 35244
rect 14737 35235 14795 35241
rect 14918 35232 14924 35244
rect 14976 35232 14982 35284
rect 15010 35232 15016 35284
rect 15068 35232 15074 35284
rect 17218 35232 17224 35284
rect 17276 35232 17282 35284
rect 19242 35232 19248 35284
rect 19300 35272 19306 35284
rect 22833 35275 22891 35281
rect 19300 35244 22094 35272
rect 19300 35232 19306 35244
rect 11149 35139 11207 35145
rect 11149 35136 11161 35139
rect 10744 35108 11161 35136
rect 10744 35096 10750 35108
rect 11149 35105 11161 35108
rect 11195 35105 11207 35139
rect 17236 35136 17264 35232
rect 19337 35207 19395 35213
rect 19337 35173 19349 35207
rect 19383 35204 19395 35207
rect 19383 35176 20024 35204
rect 19383 35173 19395 35176
rect 19337 35167 19395 35173
rect 11149 35099 11207 35105
rect 12406 35108 17264 35136
rect 7053 35040 7696 35068
rect 7053 35037 7065 35040
rect 7007 35031 7065 35037
rect 7742 35028 7748 35080
rect 7800 35068 7806 35080
rect 7800 35040 9674 35068
rect 7800 35028 7806 35040
rect 7466 35000 7472 35012
rect 5583 34972 6500 35000
rect 6564 34972 7472 35000
rect 5583 34969 5595 34972
rect 5537 34963 5595 34969
rect 3418 34932 3424 34944
rect 1872 34904 3424 34932
rect 3418 34892 3424 34904
rect 3476 34892 3482 34944
rect 4522 34892 4528 34944
rect 4580 34932 4586 34944
rect 4890 34932 4896 34944
rect 4580 34904 4896 34932
rect 4580 34892 4586 34904
rect 4890 34892 4896 34904
rect 4948 34892 4954 34944
rect 4982 34892 4988 34944
rect 5040 34932 5046 34944
rect 5166 34932 5172 34944
rect 5040 34904 5172 34932
rect 5040 34892 5046 34904
rect 5166 34892 5172 34904
rect 5224 34892 5230 34944
rect 5258 34892 5264 34944
rect 5316 34892 5322 34944
rect 5626 34892 5632 34944
rect 5684 34932 5690 34944
rect 6270 34932 6276 34944
rect 5684 34904 6276 34932
rect 5684 34892 5690 34904
rect 6270 34892 6276 34904
rect 6328 34932 6334 34944
rect 6564 34941 6592 34972
rect 7466 34960 7472 34972
rect 7524 34960 7530 35012
rect 9646 35000 9674 35040
rect 11330 35028 11336 35080
rect 11388 35068 11394 35080
rect 11423 35071 11481 35077
rect 11423 35068 11435 35071
rect 11388 35040 11435 35068
rect 11388 35028 11394 35040
rect 11423 35037 11435 35040
rect 11469 35068 11481 35071
rect 11790 35068 11796 35080
rect 11469 35040 11796 35068
rect 11469 35037 11481 35040
rect 11423 35031 11481 35037
rect 11790 35028 11796 35040
rect 11848 35028 11854 35080
rect 12406 35000 12434 35108
rect 14918 35028 14924 35080
rect 14976 35028 14982 35080
rect 15194 35028 15200 35080
rect 15252 35028 15258 35080
rect 17310 35028 17316 35080
rect 17368 35068 17374 35080
rect 19150 35068 19156 35080
rect 17368 35040 19156 35068
rect 17368 35028 17374 35040
rect 19150 35028 19156 35040
rect 19208 35068 19214 35080
rect 19996 35077 20024 35176
rect 19521 35071 19579 35077
rect 19521 35068 19533 35071
rect 19208 35040 19533 35068
rect 19208 35028 19214 35040
rect 19521 35037 19533 35040
rect 19567 35037 19579 35071
rect 19521 35031 19579 35037
rect 19981 35071 20039 35077
rect 19981 35037 19993 35071
rect 20027 35037 20039 35071
rect 19981 35031 20039 35037
rect 20254 35028 20260 35080
rect 20312 35068 20318 35080
rect 20533 35071 20591 35077
rect 20533 35068 20545 35071
rect 20312 35040 20545 35068
rect 20312 35028 20318 35040
rect 20533 35037 20545 35040
rect 20579 35037 20591 35071
rect 22066 35068 22094 35244
rect 22833 35241 22845 35275
rect 22879 35272 22891 35275
rect 23198 35272 23204 35284
rect 22879 35244 23204 35272
rect 22879 35241 22891 35244
rect 22833 35235 22891 35241
rect 23198 35232 23204 35244
rect 23256 35232 23262 35284
rect 23382 35232 23388 35284
rect 23440 35232 23446 35284
rect 23566 35232 23572 35284
rect 23624 35272 23630 35284
rect 23661 35275 23719 35281
rect 23661 35272 23673 35275
rect 23624 35244 23673 35272
rect 23624 35232 23630 35244
rect 23661 35241 23673 35244
rect 23707 35241 23719 35275
rect 23661 35235 23719 35241
rect 23400 35136 23428 35232
rect 23400 35108 23980 35136
rect 23952 35077 23980 35108
rect 23017 35071 23075 35077
rect 23017 35068 23029 35071
rect 22066 35040 23029 35068
rect 20533 35031 20591 35037
rect 23017 35037 23029 35040
rect 23063 35037 23075 35071
rect 23845 35071 23903 35077
rect 23845 35068 23857 35071
rect 23017 35031 23075 35037
rect 23308 35040 23857 35068
rect 9646 34972 12434 35000
rect 19996 34972 21772 35000
rect 6365 34935 6423 34941
rect 6365 34932 6377 34935
rect 6328 34904 6377 34932
rect 6328 34892 6334 34904
rect 6365 34901 6377 34904
rect 6411 34901 6423 34935
rect 6365 34895 6423 34901
rect 6549 34935 6607 34941
rect 6549 34901 6561 34935
rect 6595 34901 6607 34935
rect 6549 34895 6607 34901
rect 6730 34892 6736 34944
rect 6788 34932 6794 34944
rect 7745 34935 7803 34941
rect 7745 34932 7757 34935
rect 6788 34904 7757 34932
rect 6788 34892 6794 34904
rect 7745 34901 7757 34904
rect 7791 34901 7803 34935
rect 7745 34895 7803 34901
rect 15102 34892 15108 34944
rect 15160 34932 15166 34944
rect 16482 34932 16488 34944
rect 15160 34904 16488 34932
rect 15160 34892 15166 34904
rect 16482 34892 16488 34904
rect 16540 34932 16546 34944
rect 19996 34932 20024 34972
rect 21744 34944 21772 34972
rect 16540 34904 20024 34932
rect 16540 34892 16546 34904
rect 20070 34892 20076 34944
rect 20128 34892 20134 34944
rect 20346 34892 20352 34944
rect 20404 34892 20410 34944
rect 21726 34892 21732 34944
rect 21784 34892 21790 34944
rect 22922 34892 22928 34944
rect 22980 34932 22986 34944
rect 23308 34941 23336 35040
rect 23845 35037 23857 35040
rect 23891 35037 23903 35071
rect 23845 35031 23903 35037
rect 23937 35071 23995 35077
rect 23937 35037 23949 35071
rect 23983 35037 23995 35071
rect 23937 35031 23995 35037
rect 23293 34935 23351 34941
rect 23293 34932 23305 34935
rect 22980 34904 23305 34932
rect 22980 34892 22986 34904
rect 23293 34901 23305 34904
rect 23339 34901 23351 34935
rect 23293 34895 23351 34901
rect 24121 34935 24179 34941
rect 24121 34901 24133 34935
rect 24167 34932 24179 34935
rect 24854 34932 24860 34944
rect 24167 34904 24860 34932
rect 24167 34901 24179 34904
rect 24121 34895 24179 34901
rect 24854 34892 24860 34904
rect 24912 34892 24918 34944
rect 1104 34842 24723 34864
rect 1104 34790 6814 34842
rect 6866 34790 6878 34842
rect 6930 34790 6942 34842
rect 6994 34790 7006 34842
rect 7058 34790 7070 34842
rect 7122 34790 12679 34842
rect 12731 34790 12743 34842
rect 12795 34790 12807 34842
rect 12859 34790 12871 34842
rect 12923 34790 12935 34842
rect 12987 34790 18544 34842
rect 18596 34790 18608 34842
rect 18660 34790 18672 34842
rect 18724 34790 18736 34842
rect 18788 34790 18800 34842
rect 18852 34790 24409 34842
rect 24461 34790 24473 34842
rect 24525 34790 24537 34842
rect 24589 34790 24601 34842
rect 24653 34790 24665 34842
rect 24717 34790 24723 34842
rect 1104 34768 24723 34790
rect 2774 34688 2780 34740
rect 2832 34688 2838 34740
rect 2884 34700 4660 34728
rect 2884 34660 2912 34700
rect 4632 34672 4660 34700
rect 4982 34688 4988 34740
rect 5040 34688 5046 34740
rect 5718 34688 5724 34740
rect 5776 34688 5782 34740
rect 7466 34688 7472 34740
rect 7524 34728 7530 34740
rect 9582 34728 9588 34740
rect 7524 34700 9588 34728
rect 7524 34688 7530 34700
rect 9582 34688 9588 34700
rect 9640 34688 9646 34740
rect 9861 34731 9919 34737
rect 9861 34697 9873 34731
rect 9907 34728 9919 34731
rect 10318 34728 10324 34740
rect 9907 34700 10324 34728
rect 9907 34697 9919 34700
rect 9861 34691 9919 34697
rect 10318 34688 10324 34700
rect 10376 34688 10382 34740
rect 10778 34688 10784 34740
rect 10836 34728 10842 34740
rect 12250 34728 12256 34740
rect 10836 34700 12256 34728
rect 10836 34688 10842 34700
rect 12250 34688 12256 34700
rect 12308 34688 12314 34740
rect 12526 34728 12532 34740
rect 12406 34700 12532 34728
rect 2054 34632 2912 34660
rect 2054 34631 2082 34632
rect 2023 34625 2082 34631
rect 2023 34591 2035 34625
rect 2069 34594 2082 34625
rect 3403 34625 3461 34631
rect 2069 34591 2081 34594
rect 3403 34592 3415 34625
rect 2023 34585 2081 34591
rect 3068 34591 3415 34592
rect 3449 34622 3461 34625
rect 3449 34591 3464 34622
rect 4614 34620 4620 34672
rect 4672 34620 4678 34672
rect 4798 34660 4804 34672
rect 4724 34632 4804 34660
rect 4724 34601 4752 34632
rect 4798 34620 4804 34632
rect 4856 34660 4862 34672
rect 5000 34660 5028 34688
rect 4856 34632 5028 34660
rect 4856 34620 4862 34632
rect 9214 34620 9220 34672
rect 9272 34660 9278 34672
rect 12406 34660 12434 34700
rect 12526 34688 12532 34700
rect 12584 34688 12590 34740
rect 20070 34688 20076 34740
rect 20128 34688 20134 34740
rect 20254 34688 20260 34740
rect 20312 34688 20318 34740
rect 20346 34688 20352 34740
rect 20404 34728 20410 34740
rect 20404 34700 21220 34728
rect 20404 34688 20410 34700
rect 19150 34669 19156 34672
rect 19144 34660 19156 34669
rect 9272 34632 12434 34660
rect 19111 34632 19156 34660
rect 9272 34620 9278 34632
rect 19144 34623 19156 34632
rect 19150 34620 19156 34623
rect 19208 34620 19214 34672
rect 3068 34564 3464 34591
rect 4709 34595 4767 34601
rect 1486 34484 1492 34536
rect 1544 34524 1550 34536
rect 1765 34527 1823 34533
rect 1765 34524 1777 34527
rect 1544 34496 1777 34524
rect 1544 34484 1550 34496
rect 1765 34493 1777 34496
rect 1811 34493 1823 34527
rect 1765 34487 1823 34493
rect 2958 34484 2964 34536
rect 3016 34524 3022 34536
rect 3068 34524 3096 34564
rect 4709 34561 4721 34595
rect 4755 34561 4767 34595
rect 4709 34555 4767 34561
rect 4890 34552 4896 34604
rect 4948 34592 4954 34604
rect 4983 34595 5041 34601
rect 4983 34592 4995 34595
rect 4948 34564 4995 34592
rect 4948 34552 4954 34564
rect 4983 34561 4995 34564
rect 5029 34561 5041 34595
rect 4983 34555 5041 34561
rect 5902 34552 5908 34604
rect 5960 34592 5966 34604
rect 6178 34592 6184 34604
rect 5960 34564 6184 34592
rect 5960 34552 5966 34564
rect 6178 34552 6184 34564
rect 6236 34592 6242 34604
rect 6883 34595 6941 34601
rect 6883 34592 6895 34595
rect 6236 34564 6895 34592
rect 6236 34552 6242 34564
rect 6883 34561 6895 34564
rect 6929 34561 6941 34595
rect 6883 34555 6941 34561
rect 9585 34595 9643 34601
rect 9585 34561 9597 34595
rect 9631 34592 9643 34595
rect 10318 34592 10324 34604
rect 9631 34564 10324 34592
rect 9631 34561 9643 34564
rect 9585 34555 9643 34561
rect 10318 34552 10324 34564
rect 10376 34552 10382 34604
rect 12250 34552 12256 34604
rect 12308 34552 12314 34604
rect 13814 34552 13820 34604
rect 13872 34592 13878 34604
rect 16666 34592 16672 34604
rect 13872 34564 16672 34592
rect 13872 34552 13878 34564
rect 16666 34552 16672 34564
rect 16724 34552 16730 34604
rect 18874 34552 18880 34604
rect 18932 34552 18938 34604
rect 20088 34592 20116 34688
rect 20901 34663 20959 34669
rect 20901 34629 20913 34663
rect 20947 34660 20959 34663
rect 21085 34663 21143 34669
rect 21085 34660 21097 34663
rect 20947 34632 21097 34660
rect 20947 34629 20959 34632
rect 20901 34623 20959 34629
rect 21085 34629 21097 34632
rect 21131 34629 21143 34663
rect 21085 34623 21143 34629
rect 20533 34595 20591 34601
rect 20533 34592 20545 34595
rect 18984 34564 20024 34592
rect 20088 34564 20545 34592
rect 3016 34496 3096 34524
rect 3145 34527 3203 34533
rect 3016 34484 3022 34496
rect 3145 34493 3157 34527
rect 3191 34493 3203 34527
rect 3145 34487 3203 34493
rect 3160 34388 3188 34487
rect 6086 34484 6092 34536
rect 6144 34524 6150 34536
rect 6638 34524 6644 34536
rect 6144 34496 6644 34524
rect 6144 34484 6150 34496
rect 6638 34484 6644 34496
rect 6696 34484 6702 34536
rect 9861 34527 9919 34533
rect 9861 34493 9873 34527
rect 9907 34524 9919 34527
rect 10778 34524 10784 34536
rect 9907 34496 10784 34524
rect 9907 34493 9919 34496
rect 9861 34487 9919 34493
rect 10778 34484 10784 34496
rect 10836 34484 10842 34536
rect 12268 34524 12296 34552
rect 18984 34524 19012 34564
rect 12268 34496 19012 34524
rect 19996 34524 20024 34564
rect 20533 34561 20545 34564
rect 20579 34561 20591 34595
rect 20533 34555 20591 34561
rect 20622 34552 20628 34604
rect 20680 34592 20686 34604
rect 21192 34601 21220 34700
rect 21818 34688 21824 34740
rect 21876 34688 21882 34740
rect 22649 34731 22707 34737
rect 22649 34697 22661 34731
rect 22695 34697 22707 34731
rect 22649 34691 22707 34697
rect 23385 34731 23443 34737
rect 23385 34697 23397 34731
rect 23431 34697 23443 34731
rect 23385 34691 23443 34697
rect 22664 34660 22692 34691
rect 23400 34660 23428 34691
rect 23845 34663 23903 34669
rect 23845 34660 23857 34663
rect 22664 34632 23152 34660
rect 23400 34632 23857 34660
rect 20717 34595 20775 34601
rect 20717 34592 20729 34595
rect 20680 34564 20729 34592
rect 20680 34552 20686 34564
rect 20717 34561 20729 34564
rect 20763 34592 20775 34595
rect 20993 34595 21051 34601
rect 20993 34592 21005 34595
rect 20763 34564 21005 34592
rect 20763 34561 20775 34564
rect 20717 34555 20775 34561
rect 20993 34561 21005 34564
rect 21039 34561 21051 34595
rect 20993 34555 21051 34561
rect 21177 34595 21235 34601
rect 21177 34561 21189 34595
rect 21223 34561 21235 34595
rect 21177 34555 21235 34561
rect 22002 34552 22008 34604
rect 22060 34552 22066 34604
rect 22833 34595 22891 34601
rect 22833 34561 22845 34595
rect 22879 34561 22891 34595
rect 23124 34592 23152 34632
rect 23845 34629 23857 34632
rect 23891 34629 23903 34663
rect 23845 34623 23903 34629
rect 23569 34595 23627 34601
rect 23569 34592 23581 34595
rect 23124 34564 23581 34592
rect 22833 34555 22891 34561
rect 23569 34561 23581 34564
rect 23615 34561 23627 34595
rect 23569 34555 23627 34561
rect 22848 34524 22876 34555
rect 19996 34496 21404 34524
rect 7300 34428 17264 34456
rect 3602 34388 3608 34400
rect 3160 34360 3608 34388
rect 3602 34348 3608 34360
rect 3660 34348 3666 34400
rect 4157 34391 4215 34397
rect 4157 34357 4169 34391
rect 4203 34388 4215 34391
rect 4246 34388 4252 34400
rect 4203 34360 4252 34388
rect 4203 34357 4215 34360
rect 4157 34351 4215 34357
rect 4246 34348 4252 34360
rect 4304 34348 4310 34400
rect 4614 34348 4620 34400
rect 4672 34388 4678 34400
rect 5442 34388 5448 34400
rect 4672 34360 5448 34388
rect 4672 34348 4678 34360
rect 5442 34348 5448 34360
rect 5500 34388 5506 34400
rect 7300 34388 7328 34428
rect 17236 34400 17264 34428
rect 20530 34416 20536 34468
rect 20588 34416 20594 34468
rect 21376 34400 21404 34496
rect 22020 34496 22876 34524
rect 21726 34416 21732 34468
rect 21784 34456 21790 34468
rect 22020 34456 22048 34496
rect 24118 34484 24124 34536
rect 24176 34484 24182 34536
rect 21784 34428 22048 34456
rect 21784 34416 21790 34428
rect 5500 34360 7328 34388
rect 5500 34348 5506 34360
rect 7650 34348 7656 34400
rect 7708 34348 7714 34400
rect 8662 34348 8668 34400
rect 8720 34388 8726 34400
rect 9677 34391 9735 34397
rect 9677 34388 9689 34391
rect 8720 34360 9689 34388
rect 8720 34348 8726 34360
rect 9677 34357 9689 34360
rect 9723 34357 9735 34391
rect 9677 34351 9735 34357
rect 11330 34348 11336 34400
rect 11388 34388 11394 34400
rect 15102 34388 15108 34400
rect 11388 34360 15108 34388
rect 11388 34348 11394 34360
rect 15102 34348 15108 34360
rect 15160 34348 15166 34400
rect 17218 34348 17224 34400
rect 17276 34348 17282 34400
rect 21358 34348 21364 34400
rect 21416 34388 21422 34400
rect 22830 34388 22836 34400
rect 21416 34360 22836 34388
rect 21416 34348 21422 34360
rect 22830 34348 22836 34360
rect 22888 34348 22894 34400
rect 1104 34298 24564 34320
rect 1104 34246 3882 34298
rect 3934 34246 3946 34298
rect 3998 34246 4010 34298
rect 4062 34246 4074 34298
rect 4126 34246 4138 34298
rect 4190 34246 9747 34298
rect 9799 34246 9811 34298
rect 9863 34246 9875 34298
rect 9927 34246 9939 34298
rect 9991 34246 10003 34298
rect 10055 34246 15612 34298
rect 15664 34246 15676 34298
rect 15728 34246 15740 34298
rect 15792 34246 15804 34298
rect 15856 34246 15868 34298
rect 15920 34246 21477 34298
rect 21529 34246 21541 34298
rect 21593 34246 21605 34298
rect 21657 34246 21669 34298
rect 21721 34246 21733 34298
rect 21785 34246 24564 34298
rect 1104 34224 24564 34246
rect 3602 34144 3608 34196
rect 3660 34184 3666 34196
rect 4062 34184 4068 34196
rect 3660 34156 4068 34184
rect 3660 34144 3666 34156
rect 4062 34144 4068 34156
rect 4120 34144 4126 34196
rect 5258 34144 5264 34196
rect 5316 34184 5322 34196
rect 5353 34187 5411 34193
rect 5353 34184 5365 34187
rect 5316 34156 5365 34184
rect 5316 34144 5322 34156
rect 5353 34153 5365 34156
rect 5399 34153 5411 34187
rect 5353 34147 5411 34153
rect 8662 34144 8668 34196
rect 8720 34144 8726 34196
rect 9398 34184 9404 34196
rect 8956 34156 9404 34184
rect 7834 34076 7840 34128
rect 7892 34116 7898 34128
rect 8956 34116 8984 34156
rect 9398 34144 9404 34156
rect 9456 34184 9462 34196
rect 9456 34156 10272 34184
rect 9456 34144 9462 34156
rect 7892 34088 8984 34116
rect 9033 34119 9091 34125
rect 7892 34076 7898 34088
rect 9033 34085 9045 34119
rect 9079 34085 9091 34119
rect 10244 34116 10272 34156
rect 10318 34144 10324 34196
rect 10376 34144 10382 34196
rect 10778 34144 10784 34196
rect 10836 34144 10842 34196
rect 13262 34184 13268 34196
rect 10888 34156 13268 34184
rect 10888 34116 10916 34156
rect 13262 34144 13268 34156
rect 13320 34144 13326 34196
rect 19702 34184 19708 34196
rect 14752 34156 15976 34184
rect 10244 34088 10916 34116
rect 9033 34079 9091 34085
rect 1302 34008 1308 34060
rect 1360 34048 1366 34060
rect 3329 34051 3387 34057
rect 1360 34020 2774 34048
rect 1360 34008 1366 34020
rect 1394 33940 1400 33992
rect 1452 33940 1458 33992
rect 1946 33940 1952 33992
rect 2004 33940 2010 33992
rect 2501 33983 2559 33989
rect 2501 33949 2513 33983
rect 2547 33949 2559 33983
rect 2746 33980 2774 34020
rect 3329 34017 3341 34051
rect 3375 34048 3387 34051
rect 3694 34048 3700 34060
rect 3375 34020 3700 34048
rect 3375 34017 3387 34020
rect 3329 34011 3387 34017
rect 3694 34008 3700 34020
rect 3752 34008 3758 34060
rect 4246 34008 4252 34060
rect 4304 34008 4310 34060
rect 6730 34008 6736 34060
rect 6788 34008 6794 34060
rect 3053 33983 3111 33989
rect 3053 33980 3065 33983
rect 2746 33952 3065 33980
rect 2501 33943 2559 33949
rect 3053 33949 3065 33952
rect 3099 33949 3111 33983
rect 6270 33980 6276 33992
rect 3053 33943 3111 33949
rect 3528 33952 6276 33980
rect 1670 33872 1676 33924
rect 1728 33872 1734 33924
rect 2222 33872 2228 33924
rect 2280 33872 2286 33924
rect 1118 33804 1124 33856
rect 1176 33844 1182 33856
rect 2516 33844 2544 33943
rect 2777 33915 2835 33921
rect 2777 33881 2789 33915
rect 2823 33912 2835 33915
rect 3528 33912 3556 33952
rect 6270 33940 6276 33952
rect 6328 33940 6334 33992
rect 6454 33940 6460 33992
rect 6512 33940 6518 33992
rect 6638 33940 6644 33992
rect 6696 33980 6702 33992
rect 6825 33983 6883 33989
rect 6825 33980 6837 33983
rect 6696 33952 6837 33980
rect 6696 33940 6702 33952
rect 6825 33949 6837 33952
rect 6871 33949 6883 33983
rect 6825 33943 6883 33949
rect 6917 33983 6975 33989
rect 6917 33949 6929 33983
rect 6963 33980 6975 33983
rect 7650 33980 7656 33992
rect 6963 33952 7656 33980
rect 6963 33949 6975 33952
rect 6917 33943 6975 33949
rect 7650 33940 7656 33952
rect 7708 33940 7714 33992
rect 8573 33983 8631 33989
rect 8573 33949 8585 33983
rect 8619 33980 8631 33983
rect 9048 33980 9076 34079
rect 12158 34076 12164 34128
rect 12216 34116 12222 34128
rect 12342 34116 12348 34128
rect 12216 34088 12348 34116
rect 12216 34076 12222 34088
rect 12342 34076 12348 34088
rect 12400 34076 12406 34128
rect 10318 34008 10324 34060
rect 10376 34008 10382 34060
rect 10410 34008 10416 34060
rect 10468 34048 10474 34060
rect 11241 34051 11299 34057
rect 11241 34048 11253 34051
rect 10468 34020 11253 34048
rect 10468 34008 10474 34020
rect 11241 34017 11253 34020
rect 11287 34017 11299 34051
rect 11241 34011 11299 34017
rect 8619 33952 9076 33980
rect 8619 33949 8631 33952
rect 8573 33943 8631 33949
rect 9122 33940 9128 33992
rect 9180 33980 9186 33992
rect 9217 33983 9275 33989
rect 9217 33980 9229 33983
rect 9180 33952 9229 33980
rect 9180 33940 9186 33952
rect 9217 33949 9229 33952
rect 9263 33949 9275 33983
rect 9217 33943 9275 33949
rect 9306 33940 9312 33992
rect 9364 33940 9370 33992
rect 9490 33940 9496 33992
rect 9548 33980 9554 33992
rect 9583 33983 9641 33989
rect 9583 33980 9595 33983
rect 9548 33952 9595 33980
rect 9548 33940 9554 33952
rect 9583 33949 9595 33952
rect 9629 33949 9641 33983
rect 10336 33980 10364 34008
rect 10689 33983 10747 33989
rect 10689 33980 10701 33983
rect 10336 33952 10701 33980
rect 9583 33943 9641 33949
rect 10689 33949 10701 33952
rect 10735 33949 10747 33983
rect 10689 33943 10747 33949
rect 10778 33940 10784 33992
rect 10836 33980 10842 33992
rect 10873 33983 10931 33989
rect 10873 33980 10885 33983
rect 10836 33952 10885 33980
rect 10836 33940 10842 33952
rect 10873 33949 10885 33952
rect 10919 33949 10931 33983
rect 11515 33983 11573 33989
rect 11515 33980 11527 33983
rect 10873 33943 10931 33949
rect 11498 33949 11527 33980
rect 11561 33980 11573 33983
rect 14752 33980 14780 34156
rect 15948 34060 15976 34156
rect 19444 34156 19708 34184
rect 15930 34008 15936 34060
rect 15988 34008 15994 34060
rect 19444 34057 19472 34156
rect 19702 34144 19708 34156
rect 19760 34144 19766 34196
rect 20441 34187 20499 34193
rect 20441 34153 20453 34187
rect 20487 34184 20499 34187
rect 20622 34184 20628 34196
rect 20487 34156 20628 34184
rect 20487 34153 20499 34156
rect 20441 34147 20499 34153
rect 20622 34144 20628 34156
rect 20680 34144 20686 34196
rect 21453 34187 21511 34193
rect 21453 34153 21465 34187
rect 21499 34184 21511 34187
rect 22002 34184 22008 34196
rect 21499 34156 22008 34184
rect 21499 34153 21511 34156
rect 21453 34147 21511 34153
rect 22002 34144 22008 34156
rect 22060 34144 22066 34196
rect 23661 34119 23719 34125
rect 23661 34085 23673 34119
rect 23707 34085 23719 34119
rect 23661 34079 23719 34085
rect 19429 34051 19487 34057
rect 19429 34017 19441 34051
rect 19475 34017 19487 34051
rect 23676 34048 23704 34079
rect 23676 34020 23980 34048
rect 19429 34011 19487 34017
rect 11561 33952 14780 33980
rect 14829 33983 14887 33989
rect 11561 33949 11573 33952
rect 11498 33943 11573 33949
rect 14829 33949 14841 33983
rect 14875 33980 14887 33983
rect 15010 33980 15016 33992
rect 14875 33952 15016 33980
rect 14875 33949 14887 33952
rect 14829 33943 14887 33949
rect 2823 33884 3556 33912
rect 2823 33881 2835 33884
rect 2777 33875 2835 33881
rect 3602 33872 3608 33924
rect 3660 33912 3666 33924
rect 4338 33912 4344 33924
rect 3660 33884 4344 33912
rect 3660 33872 3666 33884
rect 4338 33872 4344 33884
rect 4396 33872 4402 33924
rect 4433 33915 4491 33921
rect 4433 33881 4445 33915
rect 4479 33881 4491 33915
rect 4433 33875 4491 33881
rect 1176 33816 2544 33844
rect 1176 33804 1182 33816
rect 3234 33804 3240 33856
rect 3292 33844 3298 33856
rect 4065 33847 4123 33853
rect 4065 33844 4077 33847
rect 3292 33816 4077 33844
rect 3292 33804 3298 33816
rect 4065 33813 4077 33816
rect 4111 33813 4123 33847
rect 4065 33807 4123 33813
rect 4154 33804 4160 33856
rect 4212 33844 4218 33856
rect 4448 33844 4476 33875
rect 4706 33872 4712 33924
rect 4764 33912 4770 33924
rect 4801 33915 4859 33921
rect 4801 33912 4813 33915
rect 4764 33884 4813 33912
rect 4764 33872 4770 33884
rect 4801 33881 4813 33884
rect 4847 33881 4859 33915
rect 6472 33912 6500 33940
rect 6472 33884 6868 33912
rect 4801 33875 4859 33881
rect 4212 33816 4476 33844
rect 4212 33804 4218 33816
rect 4614 33804 4620 33856
rect 4672 33844 4678 33856
rect 5074 33844 5080 33856
rect 4672 33816 5080 33844
rect 4672 33804 4678 33816
rect 5074 33804 5080 33816
rect 5132 33844 5138 33856
rect 5169 33847 5227 33853
rect 5169 33844 5181 33847
rect 5132 33816 5181 33844
rect 5132 33804 5138 33816
rect 5169 33813 5181 33816
rect 5215 33813 5227 33847
rect 5169 33807 5227 33813
rect 6178 33804 6184 33856
rect 6236 33844 6242 33856
rect 6549 33847 6607 33853
rect 6549 33844 6561 33847
rect 6236 33816 6561 33844
rect 6236 33804 6242 33816
rect 6549 33813 6561 33816
rect 6595 33813 6607 33847
rect 6840 33844 6868 33884
rect 7282 33872 7288 33924
rect 7340 33872 7346 33924
rect 10318 33912 10324 33924
rect 7852 33884 10324 33912
rect 7852 33853 7880 33884
rect 10318 33872 10324 33884
rect 10376 33872 10382 33924
rect 7653 33847 7711 33853
rect 7653 33844 7665 33847
rect 6840 33816 7665 33844
rect 6549 33807 6607 33813
rect 7653 33813 7665 33816
rect 7699 33813 7711 33847
rect 7653 33807 7711 33813
rect 7837 33847 7895 33853
rect 7837 33813 7849 33847
rect 7883 33813 7895 33847
rect 7837 33807 7895 33813
rect 7926 33804 7932 33856
rect 7984 33844 7990 33856
rect 11498 33844 11526 33943
rect 15010 33940 15016 33952
rect 15068 33940 15074 33992
rect 15102 33940 15108 33992
rect 15160 33980 15166 33992
rect 15160 33952 15203 33980
rect 15160 33940 15166 33952
rect 19610 33940 19616 33992
rect 19668 33980 19674 33992
rect 19703 33983 19761 33989
rect 19703 33980 19715 33983
rect 19668 33952 19715 33980
rect 19668 33940 19674 33952
rect 19703 33949 19715 33952
rect 19749 33980 19761 33983
rect 20070 33980 20076 33992
rect 19749 33952 20076 33980
rect 19749 33949 19761 33952
rect 19703 33943 19761 33949
rect 20070 33940 20076 33952
rect 20128 33940 20134 33992
rect 21637 33983 21695 33989
rect 21637 33949 21649 33983
rect 21683 33949 21695 33983
rect 21637 33943 21695 33949
rect 13078 33872 13084 33924
rect 13136 33912 13142 33924
rect 17954 33912 17960 33924
rect 13136 33884 17960 33912
rect 13136 33872 13142 33884
rect 17954 33872 17960 33884
rect 18012 33872 18018 33924
rect 18046 33872 18052 33924
rect 18104 33912 18110 33924
rect 21652 33912 21680 33943
rect 23842 33940 23848 33992
rect 23900 33940 23906 33992
rect 23952 33989 23980 34020
rect 23937 33983 23995 33989
rect 23937 33949 23949 33983
rect 23983 33949 23995 33983
rect 23937 33943 23995 33949
rect 18104 33884 21680 33912
rect 18104 33872 18110 33884
rect 7984 33816 11526 33844
rect 7984 33804 7990 33816
rect 12250 33804 12256 33856
rect 12308 33804 12314 33856
rect 15378 33804 15384 33856
rect 15436 33844 15442 33856
rect 15841 33847 15899 33853
rect 15841 33844 15853 33847
rect 15436 33816 15853 33844
rect 15436 33804 15442 33816
rect 15841 33813 15853 33816
rect 15887 33813 15899 33847
rect 15841 33807 15899 33813
rect 17218 33804 17224 33856
rect 17276 33844 17282 33856
rect 22738 33844 22744 33856
rect 17276 33816 22744 33844
rect 17276 33804 17282 33816
rect 22738 33804 22744 33816
rect 22796 33804 22802 33856
rect 24121 33847 24179 33853
rect 24121 33813 24133 33847
rect 24167 33844 24179 33847
rect 24854 33844 24860 33856
rect 24167 33816 24860 33844
rect 24167 33813 24179 33816
rect 24121 33807 24179 33813
rect 24854 33804 24860 33816
rect 24912 33804 24918 33856
rect 1104 33754 24723 33776
rect 1104 33702 6814 33754
rect 6866 33702 6878 33754
rect 6930 33702 6942 33754
rect 6994 33702 7006 33754
rect 7058 33702 7070 33754
rect 7122 33702 12679 33754
rect 12731 33702 12743 33754
rect 12795 33702 12807 33754
rect 12859 33702 12871 33754
rect 12923 33702 12935 33754
rect 12987 33702 18544 33754
rect 18596 33702 18608 33754
rect 18660 33702 18672 33754
rect 18724 33702 18736 33754
rect 18788 33702 18800 33754
rect 18852 33702 24409 33754
rect 24461 33702 24473 33754
rect 24525 33702 24537 33754
rect 24589 33702 24601 33754
rect 24653 33702 24665 33754
rect 24717 33702 24723 33754
rect 1104 33680 24723 33702
rect 4157 33643 4215 33649
rect 4157 33609 4169 33643
rect 4203 33640 4215 33643
rect 4338 33640 4344 33652
rect 4203 33612 4344 33640
rect 4203 33609 4215 33612
rect 4157 33603 4215 33609
rect 4338 33600 4344 33612
rect 4396 33600 4402 33652
rect 4890 33600 4896 33652
rect 4948 33640 4954 33652
rect 5261 33643 5319 33649
rect 5261 33640 5273 33643
rect 4948 33612 5273 33640
rect 4948 33600 4954 33612
rect 5261 33609 5273 33612
rect 5307 33609 5319 33643
rect 5261 33603 5319 33609
rect 5626 33600 5632 33652
rect 5684 33640 5690 33652
rect 6362 33640 6368 33652
rect 5684 33612 6368 33640
rect 5684 33600 5690 33612
rect 6362 33600 6368 33612
rect 6420 33640 6426 33652
rect 6638 33640 6644 33652
rect 6420 33612 6644 33640
rect 6420 33600 6426 33612
rect 6638 33600 6644 33612
rect 6696 33600 6702 33652
rect 7006 33600 7012 33652
rect 7064 33640 7070 33652
rect 7466 33640 7472 33652
rect 7064 33612 7472 33640
rect 7064 33600 7070 33612
rect 7466 33600 7472 33612
rect 7524 33600 7530 33652
rect 7650 33600 7656 33652
rect 7708 33640 7714 33652
rect 9306 33640 9312 33652
rect 7708 33612 9312 33640
rect 7708 33600 7714 33612
rect 9306 33600 9312 33612
rect 9364 33600 9370 33652
rect 9677 33643 9735 33649
rect 9677 33609 9689 33643
rect 9723 33640 9735 33643
rect 10778 33640 10784 33652
rect 9723 33612 10784 33640
rect 9723 33609 9735 33612
rect 9677 33603 9735 33609
rect 10778 33600 10784 33612
rect 10836 33600 10842 33652
rect 11698 33600 11704 33652
rect 11756 33600 11762 33652
rect 12250 33600 12256 33652
rect 12308 33600 12314 33652
rect 13078 33640 13084 33652
rect 12406 33612 13084 33640
rect 1302 33532 1308 33584
rect 1360 33572 1366 33584
rect 1360 33544 2820 33572
rect 1360 33532 1366 33544
rect 1578 33464 1584 33516
rect 1636 33504 1642 33516
rect 1671 33507 1729 33513
rect 1671 33504 1683 33507
rect 1636 33476 1683 33504
rect 1636 33464 1642 33476
rect 1671 33473 1683 33476
rect 1717 33473 1729 33507
rect 1671 33467 1729 33473
rect 2130 33464 2136 33516
rect 2188 33504 2194 33516
rect 2590 33504 2596 33516
rect 2188 33476 2596 33504
rect 2188 33464 2194 33476
rect 2590 33464 2596 33476
rect 2648 33464 2654 33516
rect 2792 33513 2820 33544
rect 5994 33532 6000 33584
rect 6052 33532 6058 33584
rect 6178 33532 6184 33584
rect 6236 33572 6242 33584
rect 8202 33572 8208 33584
rect 6236 33544 8208 33572
rect 6236 33532 6242 33544
rect 8202 33532 8208 33544
rect 8260 33532 8266 33584
rect 11330 33572 11336 33584
rect 10334 33544 11336 33572
rect 4491 33517 4549 33523
rect 4491 33516 4503 33517
rect 2777 33507 2835 33513
rect 2777 33473 2789 33507
rect 2823 33473 2835 33507
rect 2777 33467 2835 33473
rect 3970 33464 3976 33516
rect 4028 33464 4034 33516
rect 4062 33464 4068 33516
rect 4120 33504 4126 33516
rect 4249 33507 4307 33513
rect 4249 33504 4261 33507
rect 4120 33476 4261 33504
rect 4120 33464 4126 33476
rect 4249 33473 4261 33476
rect 4295 33473 4307 33507
rect 4249 33467 4307 33473
rect 4430 33464 4436 33516
rect 4488 33483 4503 33516
rect 4537 33483 4549 33517
rect 4488 33477 4549 33483
rect 6012 33504 6040 33532
rect 7926 33513 7932 33516
rect 7895 33507 7932 33513
rect 7895 33504 7907 33507
rect 4488 33464 4494 33477
rect 6012 33476 7907 33504
rect 7895 33473 7907 33476
rect 7895 33467 7932 33473
rect 7926 33464 7932 33467
rect 7984 33464 7990 33516
rect 9398 33464 9404 33516
rect 9456 33504 9462 33516
rect 10334 33513 10362 33544
rect 11330 33532 11336 33544
rect 11388 33532 11394 33584
rect 11974 33532 11980 33584
rect 12032 33532 12038 33584
rect 12069 33575 12127 33581
rect 12069 33541 12081 33575
rect 12115 33572 12127 33575
rect 12268 33572 12296 33600
rect 12406 33572 12434 33612
rect 13078 33600 13084 33612
rect 13136 33600 13142 33652
rect 13630 33640 13636 33652
rect 13188 33612 13636 33640
rect 12115 33544 12296 33572
rect 12360 33544 12434 33572
rect 12115 33541 12127 33544
rect 12069 33535 12127 33541
rect 9861 33507 9919 33513
rect 9861 33504 9873 33507
rect 9456 33476 9873 33504
rect 9456 33464 9462 33476
rect 9861 33473 9873 33476
rect 9907 33473 9919 33507
rect 10319 33507 10377 33513
rect 10319 33504 10331 33507
rect 9861 33467 9919 33473
rect 9968 33476 10331 33504
rect 842 33396 848 33448
rect 900 33436 906 33448
rect 1118 33436 1124 33448
rect 900 33408 1124 33436
rect 900 33396 906 33408
rect 1118 33396 1124 33408
rect 1176 33396 1182 33448
rect 1397 33439 1455 33445
rect 1397 33405 1409 33439
rect 1443 33405 1455 33439
rect 1397 33399 1455 33405
rect 3053 33439 3111 33445
rect 3053 33405 3065 33439
rect 3099 33405 3111 33439
rect 3053 33399 3111 33405
rect 1412 33368 1440 33399
rect 1412 33340 1532 33368
rect 1504 33312 1532 33340
rect 1486 33260 1492 33312
rect 1544 33260 1550 33312
rect 2130 33260 2136 33312
rect 2188 33300 2194 33312
rect 2409 33303 2467 33309
rect 2409 33300 2421 33303
rect 2188 33272 2421 33300
rect 2188 33260 2194 33272
rect 2409 33269 2421 33272
rect 2455 33269 2467 33303
rect 3068 33300 3096 33399
rect 3786 33396 3792 33448
rect 3844 33436 3850 33448
rect 4080 33436 4108 33464
rect 3844 33408 4108 33436
rect 3844 33396 3850 33408
rect 7466 33396 7472 33448
rect 7524 33436 7530 33448
rect 7650 33436 7656 33448
rect 7524 33408 7656 33436
rect 7524 33396 7530 33408
rect 7650 33396 7656 33408
rect 7708 33396 7714 33448
rect 8846 33396 8852 33448
rect 8904 33436 8910 33448
rect 9968 33436 9996 33476
rect 10319 33473 10331 33476
rect 10365 33473 10377 33507
rect 12360 33504 12388 33544
rect 12802 33532 12808 33584
rect 12860 33532 12866 33584
rect 10319 33467 10377 33473
rect 10704 33476 12388 33504
rect 8904 33408 9996 33436
rect 8904 33396 8910 33408
rect 10042 33396 10048 33448
rect 10100 33396 10106 33448
rect 3326 33328 3332 33380
rect 3384 33368 3390 33380
rect 4246 33368 4252 33380
rect 3384 33340 4252 33368
rect 3384 33328 3390 33340
rect 4246 33328 4252 33340
rect 4304 33328 4310 33380
rect 5534 33328 5540 33380
rect 5592 33368 5598 33380
rect 7282 33368 7288 33380
rect 5592 33340 7288 33368
rect 5592 33328 5598 33340
rect 7282 33328 7288 33340
rect 7340 33328 7346 33380
rect 9490 33368 9496 33380
rect 8588 33340 9496 33368
rect 8588 33300 8616 33340
rect 9490 33328 9496 33340
rect 9548 33328 9554 33380
rect 3068 33272 8616 33300
rect 8665 33303 8723 33309
rect 2409 33263 2467 33269
rect 8665 33269 8677 33303
rect 8711 33300 8723 33303
rect 8754 33300 8760 33312
rect 8711 33272 8760 33300
rect 8711 33269 8723 33272
rect 8665 33263 8723 33269
rect 8754 33260 8760 33272
rect 8812 33260 8818 33312
rect 8846 33260 8852 33312
rect 8904 33300 8910 33312
rect 10704 33300 10732 33476
rect 12434 33464 12440 33516
rect 12492 33464 12498 33516
rect 12526 33464 12532 33516
rect 12584 33504 12590 33516
rect 13188 33504 13216 33612
rect 13630 33600 13636 33612
rect 13688 33600 13694 33652
rect 14200 33612 16342 33640
rect 13262 33532 13268 33584
rect 13320 33532 13326 33584
rect 12584 33476 13216 33504
rect 13280 33504 13308 33532
rect 13539 33507 13597 33513
rect 13539 33504 13551 33507
rect 13280 33476 13551 33504
rect 12584 33464 12590 33476
rect 13188 33436 13216 33476
rect 13539 33473 13551 33476
rect 13585 33504 13597 33507
rect 14200 33504 14228 33612
rect 16314 33572 16342 33612
rect 16390 33600 16396 33652
rect 16448 33640 16454 33652
rect 16485 33643 16543 33649
rect 16485 33640 16497 33643
rect 16448 33612 16497 33640
rect 16448 33600 16454 33612
rect 16485 33609 16497 33612
rect 16531 33609 16543 33643
rect 16485 33603 16543 33609
rect 21637 33643 21695 33649
rect 21637 33609 21649 33643
rect 21683 33640 21695 33643
rect 23201 33643 23259 33649
rect 21683 33612 22600 33640
rect 21683 33609 21695 33612
rect 21637 33603 21695 33609
rect 16314 33544 16436 33572
rect 13585 33476 14228 33504
rect 13585 33473 13597 33476
rect 13539 33467 13597 33473
rect 15562 33464 15568 33516
rect 15620 33464 15626 33516
rect 16408 33504 16436 33544
rect 16758 33532 16764 33584
rect 16816 33572 16822 33584
rect 20502 33575 20560 33581
rect 20502 33572 20514 33575
rect 16816 33544 20514 33572
rect 16816 33532 16822 33544
rect 20502 33541 20514 33544
rect 20548 33572 20560 33575
rect 20548 33541 20576 33572
rect 20502 33535 20576 33541
rect 16850 33504 16856 33516
rect 16408 33476 16856 33504
rect 16850 33464 16856 33476
rect 16908 33464 16914 33516
rect 17954 33464 17960 33516
rect 18012 33464 18018 33516
rect 18874 33464 18880 33516
rect 18932 33504 18938 33516
rect 20257 33507 20315 33513
rect 20257 33504 20269 33507
rect 18932 33476 20269 33504
rect 18932 33464 18938 33476
rect 20257 33473 20269 33476
rect 20303 33473 20315 33507
rect 20548 33504 20576 33535
rect 22572 33513 22600 33612
rect 23201 33609 23213 33643
rect 23247 33640 23259 33643
rect 23842 33640 23848 33652
rect 23247 33612 23848 33640
rect 23247 33609 23259 33612
rect 23201 33603 23259 33609
rect 23842 33600 23848 33612
rect 23900 33600 23906 33652
rect 22756 33544 23428 33572
rect 22756 33516 22784 33544
rect 22005 33507 22063 33513
rect 22005 33504 22017 33507
rect 20548 33476 22017 33504
rect 20257 33467 20315 33473
rect 22005 33473 22017 33476
rect 22051 33473 22063 33507
rect 22005 33467 22063 33473
rect 22097 33507 22155 33513
rect 22097 33473 22109 33507
rect 22143 33473 22155 33507
rect 22097 33467 22155 33473
rect 22557 33507 22615 33513
rect 22557 33473 22569 33507
rect 22603 33473 22615 33507
rect 22557 33467 22615 33473
rect 13265 33439 13323 33445
rect 13265 33436 13277 33439
rect 11057 33371 11115 33377
rect 11057 33337 11069 33371
rect 11103 33368 11115 33371
rect 11532 33368 11560 33422
rect 13188 33408 13277 33436
rect 13265 33405 13277 33408
rect 13311 33405 13323 33439
rect 13265 33399 13323 33405
rect 14642 33396 14648 33448
rect 14700 33396 14706 33448
rect 14826 33436 14832 33448
rect 14752 33408 14832 33436
rect 14752 33368 14780 33408
rect 14826 33396 14832 33408
rect 14884 33396 14890 33448
rect 15286 33396 15292 33448
rect 15344 33396 15350 33448
rect 15682 33439 15740 33445
rect 15682 33436 15694 33439
rect 15396 33408 15694 33436
rect 11103 33340 11560 33368
rect 14200 33340 14780 33368
rect 11103 33337 11115 33340
rect 11057 33331 11115 33337
rect 8904 33272 10732 33300
rect 12989 33303 13047 33309
rect 8904 33260 8910 33272
rect 12989 33269 13001 33303
rect 13035 33300 13047 33303
rect 13078 33300 13084 33312
rect 13035 33272 13084 33300
rect 13035 33269 13047 33272
rect 12989 33263 13047 33269
rect 13078 33260 13084 33272
rect 13136 33260 13142 33312
rect 13262 33260 13268 33312
rect 13320 33300 13326 33312
rect 14200 33300 14228 33340
rect 13320 33272 14228 33300
rect 14277 33303 14335 33309
rect 13320 33260 13326 33272
rect 14277 33269 14289 33303
rect 14323 33300 14335 33303
rect 14366 33300 14372 33312
rect 14323 33272 14372 33300
rect 14323 33269 14335 33272
rect 14277 33263 14335 33269
rect 14366 33260 14372 33272
rect 14424 33260 14430 33312
rect 15102 33260 15108 33312
rect 15160 33300 15166 33312
rect 15396 33300 15424 33408
rect 15682 33405 15694 33408
rect 15728 33405 15740 33439
rect 15682 33399 15740 33405
rect 15841 33439 15899 33445
rect 15841 33405 15853 33439
rect 15887 33436 15899 33439
rect 16482 33436 16488 33448
rect 15887 33408 16488 33436
rect 15887 33405 15899 33408
rect 15841 33399 15899 33405
rect 16482 33396 16488 33408
rect 16540 33396 16546 33448
rect 15160 33272 15424 33300
rect 17972 33300 18000 33464
rect 22112 33436 22140 33467
rect 22738 33464 22744 33516
rect 22796 33464 22802 33516
rect 23400 33513 23428 33544
rect 23109 33507 23167 33513
rect 23109 33473 23121 33507
rect 23155 33473 23167 33507
rect 23109 33467 23167 33473
rect 23385 33507 23443 33513
rect 23385 33473 23397 33507
rect 23431 33473 23443 33507
rect 23753 33507 23811 33513
rect 23753 33504 23765 33507
rect 23385 33467 23443 33473
rect 23492 33476 23765 33504
rect 23124 33436 23152 33467
rect 21836 33408 22140 33436
rect 22204 33408 23152 33436
rect 21836 33377 21864 33408
rect 21821 33371 21879 33377
rect 21821 33337 21833 33371
rect 21867 33337 21879 33371
rect 22204 33368 22232 33408
rect 21821 33331 21879 33337
rect 22066 33340 22232 33368
rect 22925 33371 22983 33377
rect 21266 33300 21272 33312
rect 17972 33272 21272 33300
rect 15160 33260 15166 33272
rect 21266 33260 21272 33272
rect 21324 33300 21330 33312
rect 22066 33300 22094 33340
rect 22925 33337 22937 33371
rect 22971 33368 22983 33371
rect 23492 33368 23520 33476
rect 23753 33473 23765 33476
rect 23799 33473 23811 33507
rect 23753 33467 23811 33473
rect 23937 33507 23995 33513
rect 23937 33473 23949 33507
rect 23983 33473 23995 33507
rect 23937 33467 23995 33473
rect 23952 33436 23980 33467
rect 23584 33408 23980 33436
rect 23584 33377 23612 33408
rect 22971 33340 23520 33368
rect 23569 33371 23627 33377
rect 22971 33337 22983 33340
rect 22925 33331 22983 33337
rect 23569 33337 23581 33371
rect 23615 33337 23627 33371
rect 23569 33331 23627 33337
rect 21324 33272 22094 33300
rect 21324 33260 21330 33272
rect 22186 33260 22192 33312
rect 22244 33260 22250 33312
rect 22373 33303 22431 33309
rect 22373 33269 22385 33303
rect 22419 33300 22431 33303
rect 23014 33300 23020 33312
rect 22419 33272 23020 33300
rect 22419 33269 22431 33272
rect 22373 33263 22431 33269
rect 23014 33260 23020 33272
rect 23072 33260 23078 33312
rect 24118 33260 24124 33312
rect 24176 33260 24182 33312
rect 1104 33210 24564 33232
rect 1104 33158 3882 33210
rect 3934 33158 3946 33210
rect 3998 33158 4010 33210
rect 4062 33158 4074 33210
rect 4126 33158 4138 33210
rect 4190 33158 9747 33210
rect 9799 33158 9811 33210
rect 9863 33158 9875 33210
rect 9927 33158 9939 33210
rect 9991 33158 10003 33210
rect 10055 33158 15612 33210
rect 15664 33158 15676 33210
rect 15728 33158 15740 33210
rect 15792 33158 15804 33210
rect 15856 33158 15868 33210
rect 15920 33158 21477 33210
rect 21529 33158 21541 33210
rect 21593 33158 21605 33210
rect 21657 33158 21669 33210
rect 21721 33158 21733 33210
rect 21785 33158 24564 33210
rect 1104 33136 24564 33158
rect 3145 33099 3203 33105
rect 3145 33065 3157 33099
rect 3191 33096 3203 33099
rect 6178 33096 6184 33108
rect 3191 33068 6184 33096
rect 3191 33065 3203 33068
rect 3145 33059 3203 33065
rect 6178 33056 6184 33068
rect 6236 33056 6242 33108
rect 6730 33056 6736 33108
rect 6788 33096 6794 33108
rect 13541 33099 13599 33105
rect 6788 33068 13492 33096
rect 6788 33056 6794 33068
rect 3418 32988 3424 33040
rect 3476 33028 3482 33040
rect 7006 33028 7012 33040
rect 3476 33000 7012 33028
rect 3476 32988 3482 33000
rect 7006 32988 7012 33000
rect 7064 32988 7070 33040
rect 8294 32988 8300 33040
rect 8352 33028 8358 33040
rect 9214 33028 9220 33040
rect 8352 33000 9220 33028
rect 8352 32988 8358 33000
rect 9214 32988 9220 33000
rect 9272 32988 9278 33040
rect 10686 32988 10692 33040
rect 10744 33028 10750 33040
rect 11882 33028 11888 33040
rect 10744 33000 11888 33028
rect 10744 32988 10750 33000
rect 11882 32988 11888 33000
rect 11940 32988 11946 33040
rect 3326 32960 3332 32972
rect 2884 32932 3332 32960
rect 1486 32852 1492 32904
rect 1544 32892 1550 32904
rect 1581 32895 1639 32901
rect 1581 32892 1593 32895
rect 1544 32864 1593 32892
rect 1544 32852 1550 32864
rect 1581 32861 1593 32864
rect 1627 32861 1639 32895
rect 2884 32892 2912 32932
rect 3326 32920 3332 32932
rect 3384 32920 3390 32972
rect 7098 32920 7104 32972
rect 7156 32920 7162 32972
rect 12526 32920 12532 32972
rect 12584 32920 12590 32972
rect 13464 32960 13492 33068
rect 13541 33065 13553 33099
rect 13587 33096 13599 33099
rect 13814 33096 13820 33108
rect 13587 33068 13820 33096
rect 13587 33065 13599 33068
rect 13541 33059 13599 33065
rect 13814 33056 13820 33068
rect 13872 33096 13878 33108
rect 13872 33068 14780 33096
rect 13872 33056 13878 33068
rect 13630 32988 13636 33040
rect 13688 33028 13694 33040
rect 14752 33037 14780 33068
rect 15194 33056 15200 33108
rect 15252 33096 15258 33108
rect 15933 33099 15991 33105
rect 15933 33096 15945 33099
rect 15252 33068 15945 33096
rect 15252 33056 15258 33068
rect 15933 33065 15945 33068
rect 15979 33065 15991 33099
rect 15933 33059 15991 33065
rect 16482 33056 16488 33108
rect 16540 33096 16546 33108
rect 17037 33099 17095 33105
rect 17037 33096 17049 33099
rect 16540 33068 17049 33096
rect 16540 33056 16546 33068
rect 17037 33065 17049 33068
rect 17083 33065 17095 33099
rect 17037 33059 17095 33065
rect 17218 33056 17224 33108
rect 17276 33096 17282 33108
rect 19058 33096 19064 33108
rect 17276 33068 19064 33096
rect 17276 33056 17282 33068
rect 19058 33056 19064 33068
rect 19116 33096 19122 33108
rect 19702 33096 19708 33108
rect 19116 33068 19708 33096
rect 19116 33056 19122 33068
rect 19702 33056 19708 33068
rect 19760 33056 19766 33108
rect 22186 33056 22192 33108
rect 22244 33096 22250 33108
rect 22557 33099 22615 33105
rect 22557 33096 22569 33099
rect 22244 33068 22569 33096
rect 22244 33056 22250 33068
rect 22557 33065 22569 33068
rect 22603 33065 22615 33099
rect 22557 33059 22615 33065
rect 22649 33099 22707 33105
rect 22649 33065 22661 33099
rect 22695 33096 22707 33099
rect 25590 33096 25596 33108
rect 22695 33068 25596 33096
rect 22695 33065 22707 33068
rect 22649 33059 22707 33065
rect 25590 33056 25596 33068
rect 25648 33056 25654 33108
rect 14737 33031 14795 33037
rect 13688 33000 14486 33028
rect 13688 32988 13694 33000
rect 14458 32960 14486 33000
rect 14737 32997 14749 33031
rect 14783 32997 14795 33031
rect 14737 32991 14795 32997
rect 22097 33031 22155 33037
rect 22097 32997 22109 33031
rect 22143 32997 22155 33031
rect 22097 32991 22155 32997
rect 23661 33031 23719 33037
rect 23661 32997 23673 33031
rect 23707 32997 23719 33031
rect 23661 32991 23719 32997
rect 15013 32963 15071 32969
rect 15013 32960 15025 32963
rect 13464 32932 14412 32960
rect 14458 32932 15025 32960
rect 1581 32855 1639 32861
rect 1839 32865 1897 32871
rect 1839 32831 1851 32865
rect 1885 32862 1897 32865
rect 2056 32864 2912 32892
rect 2961 32895 3019 32901
rect 1885 32831 1898 32862
rect 2056 32836 2084 32864
rect 2961 32861 2973 32895
rect 3007 32892 3019 32895
rect 4617 32895 4675 32901
rect 3007 32864 3096 32892
rect 3007 32861 3019 32864
rect 2961 32855 3019 32861
rect 1839 32825 1898 32831
rect 1870 32824 1898 32825
rect 2038 32824 2044 32836
rect 1870 32796 2044 32824
rect 2038 32784 2044 32796
rect 2096 32784 2102 32836
rect 3068 32768 3096 32864
rect 4617 32861 4629 32895
rect 4663 32892 4675 32895
rect 7343 32895 7401 32901
rect 7343 32892 7355 32895
rect 4663 32864 7355 32892
rect 4663 32861 4675 32864
rect 4617 32855 4675 32861
rect 7343 32861 7355 32864
rect 7389 32892 7401 32895
rect 7742 32892 7748 32904
rect 7389 32864 7748 32892
rect 7389 32861 7401 32864
rect 7343 32855 7401 32861
rect 7742 32852 7748 32864
rect 7800 32852 7806 32904
rect 11698 32852 11704 32904
rect 11756 32892 11762 32904
rect 12069 32895 12127 32901
rect 12069 32892 12081 32895
rect 11756 32864 12081 32892
rect 11756 32852 11762 32864
rect 12069 32861 12081 32864
rect 12115 32861 12127 32895
rect 12069 32855 12127 32861
rect 12342 32852 12348 32904
rect 12400 32892 12406 32904
rect 12544 32892 12572 32920
rect 12787 32895 12845 32901
rect 12787 32892 12799 32895
rect 12400 32864 12572 32892
rect 12728 32864 12799 32892
rect 12400 32852 12406 32864
rect 3142 32784 3148 32836
rect 3200 32824 3206 32836
rect 3789 32827 3847 32833
rect 3789 32824 3801 32827
rect 3200 32796 3801 32824
rect 3200 32784 3206 32796
rect 3789 32793 3801 32796
rect 3835 32793 3847 32827
rect 3789 32787 3847 32793
rect 5166 32784 5172 32836
rect 5224 32824 5230 32836
rect 6178 32824 6184 32836
rect 5224 32796 6184 32824
rect 5224 32784 5230 32796
rect 6178 32784 6184 32796
rect 6236 32784 6242 32836
rect 6270 32784 6276 32836
rect 6328 32824 6334 32836
rect 6328 32796 12434 32824
rect 6328 32784 6334 32796
rect 2590 32716 2596 32768
rect 2648 32716 2654 32768
rect 3050 32716 3056 32768
rect 3108 32716 3114 32768
rect 5350 32716 5356 32768
rect 5408 32756 5414 32768
rect 5994 32756 6000 32768
rect 5408 32728 6000 32756
rect 5408 32716 5414 32728
rect 5994 32716 6000 32728
rect 6052 32716 6058 32768
rect 8110 32716 8116 32768
rect 8168 32716 8174 32768
rect 9306 32716 9312 32768
rect 9364 32756 9370 32768
rect 9674 32756 9680 32768
rect 9364 32728 9680 32756
rect 9364 32716 9370 32728
rect 9674 32716 9680 32728
rect 9732 32716 9738 32768
rect 11698 32716 11704 32768
rect 11756 32756 11762 32768
rect 12161 32759 12219 32765
rect 12161 32756 12173 32759
rect 11756 32728 12173 32756
rect 11756 32716 11762 32728
rect 12161 32725 12173 32728
rect 12207 32725 12219 32759
rect 12406 32756 12434 32796
rect 12728 32756 12756 32864
rect 12787 32861 12799 32864
rect 12833 32861 12845 32895
rect 12787 32855 12845 32861
rect 14093 32895 14151 32901
rect 14093 32861 14105 32895
rect 14139 32861 14151 32895
rect 14093 32855 14151 32861
rect 13078 32784 13084 32836
rect 13136 32824 13142 32836
rect 13630 32824 13636 32836
rect 13136 32796 13636 32824
rect 13136 32784 13142 32796
rect 13630 32784 13636 32796
rect 13688 32784 13694 32836
rect 13998 32756 14004 32768
rect 12406 32728 14004 32756
rect 12161 32719 12219 32725
rect 13998 32716 14004 32728
rect 14056 32716 14062 32768
rect 14108 32756 14136 32855
rect 14274 32852 14280 32904
rect 14332 32852 14338 32904
rect 14384 32892 14412 32932
rect 15013 32929 15025 32932
rect 15059 32929 15071 32963
rect 15013 32923 15071 32929
rect 15102 32920 15108 32972
rect 15160 32969 15166 32972
rect 15160 32963 15188 32969
rect 15176 32929 15188 32963
rect 15160 32923 15188 32929
rect 15160 32920 15166 32923
rect 15838 32920 15844 32972
rect 15896 32960 15902 32972
rect 16025 32963 16083 32969
rect 16025 32960 16037 32963
rect 15896 32932 16037 32960
rect 15896 32920 15902 32932
rect 16025 32929 16037 32932
rect 16071 32929 16083 32963
rect 16025 32923 16083 32929
rect 20714 32920 20720 32972
rect 20772 32960 20778 32972
rect 20990 32960 20996 32972
rect 20772 32932 20996 32960
rect 20772 32920 20778 32932
rect 20990 32920 20996 32932
rect 21048 32960 21054 32972
rect 21085 32963 21143 32969
rect 21085 32960 21097 32963
rect 21048 32932 21097 32960
rect 21048 32920 21054 32932
rect 21085 32929 21097 32932
rect 21131 32929 21143 32963
rect 21085 32923 21143 32929
rect 14458 32892 14464 32904
rect 14384 32864 14464 32892
rect 14458 32852 14464 32864
rect 14516 32852 14522 32904
rect 15286 32852 15292 32904
rect 15344 32852 15350 32904
rect 15930 32852 15936 32904
rect 15988 32892 15994 32904
rect 16299 32895 16357 32901
rect 16299 32892 16311 32895
rect 15988 32864 16311 32892
rect 15988 32852 15994 32864
rect 16299 32861 16311 32864
rect 16345 32892 16357 32895
rect 19242 32892 19248 32904
rect 16345 32864 19248 32892
rect 16345 32861 16357 32864
rect 16299 32855 16357 32861
rect 19242 32852 19248 32864
rect 19300 32852 19306 32904
rect 21358 32892 21364 32904
rect 21319 32864 21364 32892
rect 21358 32852 21364 32864
rect 21416 32852 21422 32904
rect 22112 32892 22140 32991
rect 22741 32963 22799 32969
rect 22741 32929 22753 32963
rect 22787 32960 22799 32963
rect 22925 32963 22983 32969
rect 22925 32960 22937 32963
rect 22787 32932 22937 32960
rect 22787 32929 22799 32932
rect 22741 32923 22799 32929
rect 22925 32929 22937 32932
rect 22971 32929 22983 32963
rect 23676 32960 23704 32991
rect 23676 32932 23980 32960
rect 22925 32923 22983 32929
rect 22465 32895 22523 32901
rect 22465 32892 22477 32895
rect 22112 32864 22477 32892
rect 22465 32861 22477 32864
rect 22511 32892 22523 32895
rect 22833 32895 22891 32901
rect 22833 32892 22845 32895
rect 22511 32864 22845 32892
rect 22511 32861 22523 32864
rect 22465 32855 22523 32861
rect 22833 32861 22845 32864
rect 22879 32861 22891 32895
rect 22833 32855 22891 32861
rect 23014 32852 23020 32904
rect 23072 32852 23078 32904
rect 23952 32901 23980 32932
rect 23293 32895 23351 32901
rect 23293 32892 23305 32895
rect 23124 32864 23305 32892
rect 23124 32824 23152 32864
rect 23293 32861 23305 32864
rect 23339 32861 23351 32895
rect 23845 32895 23903 32901
rect 23845 32892 23857 32895
rect 23293 32855 23351 32861
rect 23492 32864 23857 32892
rect 22066 32796 23152 32824
rect 16114 32756 16120 32768
rect 14108 32728 16120 32756
rect 16114 32716 16120 32728
rect 16172 32716 16178 32768
rect 16666 32716 16672 32768
rect 16724 32756 16730 32768
rect 17218 32756 17224 32768
rect 16724 32728 17224 32756
rect 16724 32716 16730 32728
rect 17218 32716 17224 32728
rect 17276 32756 17282 32768
rect 22066 32756 22094 32796
rect 17276 32728 22094 32756
rect 23109 32759 23167 32765
rect 17276 32716 17282 32728
rect 23109 32725 23121 32759
rect 23155 32756 23167 32759
rect 23492 32756 23520 32864
rect 23845 32861 23857 32864
rect 23891 32861 23903 32895
rect 23845 32855 23903 32861
rect 23937 32895 23995 32901
rect 23937 32861 23949 32895
rect 23983 32861 23995 32895
rect 23937 32855 23995 32861
rect 23155 32728 23520 32756
rect 24121 32759 24179 32765
rect 23155 32725 23167 32728
rect 23109 32719 23167 32725
rect 24121 32725 24133 32759
rect 24167 32756 24179 32759
rect 24854 32756 24860 32768
rect 24167 32728 24860 32756
rect 24167 32725 24179 32728
rect 24121 32719 24179 32725
rect 24854 32716 24860 32728
rect 24912 32716 24918 32768
rect 1104 32666 24723 32688
rect 1104 32614 6814 32666
rect 6866 32614 6878 32666
rect 6930 32614 6942 32666
rect 6994 32614 7006 32666
rect 7058 32614 7070 32666
rect 7122 32614 12679 32666
rect 12731 32614 12743 32666
rect 12795 32614 12807 32666
rect 12859 32614 12871 32666
rect 12923 32614 12935 32666
rect 12987 32614 18544 32666
rect 18596 32614 18608 32666
rect 18660 32614 18672 32666
rect 18724 32614 18736 32666
rect 18788 32614 18800 32666
rect 18852 32614 24409 32666
rect 24461 32614 24473 32666
rect 24525 32614 24537 32666
rect 24589 32614 24601 32666
rect 24653 32614 24665 32666
rect 24717 32614 24723 32666
rect 1104 32592 24723 32614
rect 2314 32512 2320 32564
rect 2372 32552 2378 32564
rect 5166 32552 5172 32564
rect 2372 32524 5172 32552
rect 2372 32512 2378 32524
rect 5166 32512 5172 32524
rect 5224 32512 5230 32564
rect 5258 32512 5264 32564
rect 5316 32552 5322 32564
rect 5316 32524 6316 32552
rect 5316 32512 5322 32524
rect 3602 32444 3608 32496
rect 3660 32444 3666 32496
rect 5994 32444 6000 32496
rect 6052 32484 6058 32496
rect 6052 32456 6224 32484
rect 6052 32444 6058 32456
rect 6196 32428 6224 32456
rect 1578 32376 1584 32428
rect 1636 32376 1642 32428
rect 2314 32376 2320 32428
rect 2372 32376 2378 32428
rect 2590 32376 2596 32428
rect 2648 32376 2654 32428
rect 3329 32419 3387 32425
rect 3329 32385 3341 32419
rect 3375 32385 3387 32419
rect 3329 32379 3387 32385
rect 1394 32308 1400 32360
rect 1452 32308 1458 32360
rect 2041 32351 2099 32357
rect 2041 32317 2053 32351
rect 2087 32348 2099 32351
rect 2130 32348 2136 32360
rect 2087 32320 2136 32348
rect 2087 32317 2099 32320
rect 2041 32311 2099 32317
rect 2130 32308 2136 32320
rect 2188 32308 2194 32360
rect 2455 32351 2513 32357
rect 2455 32317 2467 32351
rect 2501 32348 2513 32351
rect 2774 32348 2780 32360
rect 2501 32320 2780 32348
rect 2501 32317 2513 32320
rect 2455 32311 2513 32317
rect 2774 32308 2780 32320
rect 2832 32308 2838 32360
rect 3344 32280 3372 32379
rect 3418 32376 3424 32428
rect 3476 32416 3482 32428
rect 3881 32419 3939 32425
rect 3881 32416 3893 32419
rect 3476 32388 3893 32416
rect 3476 32376 3482 32388
rect 3881 32385 3893 32388
rect 3927 32385 3939 32419
rect 3881 32379 3939 32385
rect 4338 32376 4344 32428
rect 4396 32416 4402 32428
rect 5135 32419 5193 32425
rect 5135 32416 5147 32419
rect 4396 32388 5147 32416
rect 4396 32376 4402 32388
rect 5135 32385 5147 32388
rect 5181 32385 5193 32419
rect 5135 32379 5193 32385
rect 6178 32376 6184 32428
rect 6236 32376 6242 32428
rect 6288 32416 6316 32524
rect 9398 32512 9404 32564
rect 9456 32512 9462 32564
rect 14918 32512 14924 32564
rect 14976 32552 14982 32564
rect 15013 32555 15071 32561
rect 15013 32552 15025 32555
rect 14976 32524 15025 32552
rect 14976 32512 14982 32524
rect 15013 32521 15025 32524
rect 15059 32521 15071 32555
rect 15013 32515 15071 32521
rect 17402 32512 17408 32564
rect 17460 32552 17466 32564
rect 19334 32552 19340 32564
rect 17460 32524 19340 32552
rect 17460 32512 17466 32524
rect 19334 32512 19340 32524
rect 19392 32512 19398 32564
rect 22557 32555 22615 32561
rect 22557 32521 22569 32555
rect 22603 32521 22615 32555
rect 22557 32515 22615 32521
rect 23201 32555 23259 32561
rect 23201 32521 23213 32555
rect 23247 32552 23259 32555
rect 23247 32524 23980 32552
rect 23247 32521 23259 32524
rect 23201 32515 23259 32521
rect 20714 32484 20720 32496
rect 16132 32456 20720 32484
rect 6914 32416 6920 32428
rect 6288 32388 6920 32416
rect 6914 32376 6920 32388
rect 6972 32416 6978 32428
rect 7561 32419 7619 32425
rect 7561 32416 7573 32419
rect 6972 32388 7573 32416
rect 6972 32376 6978 32388
rect 7561 32385 7573 32388
rect 7607 32385 7619 32419
rect 7561 32379 7619 32385
rect 8754 32376 8760 32428
rect 8812 32376 8818 32428
rect 13262 32376 13268 32428
rect 13320 32416 13326 32428
rect 13357 32419 13415 32425
rect 13357 32416 13369 32419
rect 13320 32388 13369 32416
rect 13320 32376 13326 32388
rect 13357 32385 13369 32388
rect 13403 32385 13415 32419
rect 13357 32379 13415 32385
rect 14366 32376 14372 32428
rect 14424 32376 14430 32428
rect 3602 32308 3608 32360
rect 3660 32348 3666 32360
rect 3786 32348 3792 32360
rect 3660 32320 3792 32348
rect 3660 32308 3666 32320
rect 3786 32308 3792 32320
rect 3844 32308 3850 32360
rect 4798 32308 4804 32360
rect 4856 32308 4862 32360
rect 4890 32308 4896 32360
rect 4948 32308 4954 32360
rect 7650 32308 7656 32360
rect 7708 32348 7714 32360
rect 7745 32351 7803 32357
rect 7745 32348 7757 32351
rect 7708 32320 7757 32348
rect 7708 32308 7714 32320
rect 7745 32317 7757 32320
rect 7791 32317 7803 32351
rect 7745 32311 7803 32317
rect 8110 32308 8116 32360
rect 8168 32348 8174 32360
rect 8205 32351 8263 32357
rect 8205 32348 8217 32351
rect 8168 32320 8217 32348
rect 8168 32308 8174 32320
rect 8205 32317 8217 32320
rect 8251 32317 8263 32351
rect 8481 32351 8539 32357
rect 8481 32348 8493 32351
rect 8205 32311 8263 32317
rect 8312 32320 8493 32348
rect 4816 32280 4844 32308
rect 6270 32280 6276 32292
rect 3068 32252 3372 32280
rect 3988 32252 4844 32280
rect 5828 32252 6276 32280
rect 1302 32172 1308 32224
rect 1360 32212 1366 32224
rect 3068 32212 3096 32252
rect 1360 32184 3096 32212
rect 3237 32215 3295 32221
rect 1360 32172 1366 32184
rect 3237 32181 3249 32215
rect 3283 32212 3295 32215
rect 3988 32212 4016 32252
rect 3283 32184 4016 32212
rect 4065 32215 4123 32221
rect 3283 32181 3295 32184
rect 3237 32175 3295 32181
rect 4065 32181 4077 32215
rect 4111 32212 4123 32215
rect 5828 32212 5856 32252
rect 6270 32240 6276 32252
rect 6328 32280 6334 32292
rect 8018 32280 8024 32292
rect 6328 32252 8024 32280
rect 6328 32240 6334 32252
rect 8018 32240 8024 32252
rect 8076 32240 8082 32292
rect 4111 32184 5856 32212
rect 4111 32181 4123 32184
rect 4065 32175 4123 32181
rect 5902 32172 5908 32224
rect 5960 32172 5966 32224
rect 6362 32172 6368 32224
rect 6420 32212 6426 32224
rect 8312 32212 8340 32320
rect 8481 32317 8493 32320
rect 8527 32317 8539 32351
rect 8481 32311 8539 32317
rect 8619 32351 8677 32357
rect 8619 32317 8631 32351
rect 8665 32348 8677 32351
rect 8938 32348 8944 32360
rect 8665 32320 8944 32348
rect 8665 32317 8677 32320
rect 8619 32311 8677 32317
rect 8938 32308 8944 32320
rect 8996 32348 9002 32360
rect 9398 32348 9404 32360
rect 8996 32320 9404 32348
rect 8996 32308 9002 32320
rect 9398 32308 9404 32320
rect 9456 32308 9462 32360
rect 13173 32351 13231 32357
rect 13173 32317 13185 32351
rect 13219 32317 13231 32351
rect 13173 32311 13231 32317
rect 8478 32212 8484 32224
rect 6420 32184 8484 32212
rect 6420 32172 6426 32184
rect 8478 32172 8484 32184
rect 8536 32172 8542 32224
rect 8754 32172 8760 32224
rect 8812 32212 8818 32224
rect 11330 32212 11336 32224
rect 8812 32184 11336 32212
rect 8812 32172 8818 32184
rect 11330 32172 11336 32184
rect 11388 32172 11394 32224
rect 13188 32212 13216 32311
rect 13814 32308 13820 32360
rect 13872 32308 13878 32360
rect 14093 32351 14151 32357
rect 14093 32348 14105 32351
rect 13924 32320 14105 32348
rect 13630 32240 13636 32292
rect 13688 32280 13694 32292
rect 13924 32280 13952 32320
rect 14093 32317 14105 32320
rect 14139 32317 14151 32351
rect 14093 32311 14151 32317
rect 14182 32308 14188 32360
rect 14240 32357 14246 32360
rect 14240 32351 14268 32357
rect 14256 32317 14268 32351
rect 14240 32311 14268 32317
rect 14240 32308 14246 32311
rect 16132 32280 16160 32456
rect 20714 32444 20720 32456
rect 20772 32444 20778 32496
rect 22572 32484 22600 32515
rect 22572 32456 23428 32484
rect 17034 32376 17040 32428
rect 17092 32376 17098 32428
rect 18874 32376 18880 32428
rect 18932 32376 18938 32428
rect 19150 32425 19156 32428
rect 19133 32419 19156 32425
rect 19133 32416 19145 32419
rect 18984 32388 19145 32416
rect 17052 32348 17080 32376
rect 18984 32348 19012 32388
rect 19133 32385 19145 32388
rect 19133 32379 19156 32385
rect 19150 32376 19156 32379
rect 19208 32376 19214 32428
rect 22646 32416 22652 32428
rect 22066 32388 22652 32416
rect 17052 32320 19012 32348
rect 22066 32280 22094 32388
rect 22646 32376 22652 32388
rect 22704 32416 22710 32428
rect 23400 32425 23428 32456
rect 22741 32419 22799 32425
rect 22741 32416 22753 32419
rect 22704 32388 22753 32416
rect 22704 32376 22710 32388
rect 22741 32385 22753 32388
rect 22787 32385 22799 32419
rect 22741 32379 22799 32385
rect 23385 32419 23443 32425
rect 23385 32385 23397 32419
rect 23431 32385 23443 32419
rect 23385 32379 23443 32385
rect 23658 32376 23664 32428
rect 23716 32376 23722 32428
rect 23952 32425 23980 32524
rect 23937 32419 23995 32425
rect 23937 32385 23949 32419
rect 23983 32385 23995 32419
rect 23937 32379 23995 32385
rect 13688 32252 13952 32280
rect 15304 32252 16160 32280
rect 19812 32252 22094 32280
rect 13688 32240 13694 32252
rect 14274 32212 14280 32224
rect 13188 32184 14280 32212
rect 14274 32172 14280 32184
rect 14332 32172 14338 32224
rect 14734 32172 14740 32224
rect 14792 32212 14798 32224
rect 15304 32212 15332 32252
rect 14792 32184 15332 32212
rect 14792 32172 14798 32184
rect 16850 32172 16856 32224
rect 16908 32212 16914 32224
rect 19812 32212 19840 32252
rect 23750 32240 23756 32292
rect 23808 32280 23814 32292
rect 23845 32283 23903 32289
rect 23845 32280 23857 32283
rect 23808 32252 23857 32280
rect 23808 32240 23814 32252
rect 23845 32249 23857 32252
rect 23891 32249 23903 32283
rect 23845 32243 23903 32249
rect 16908 32184 19840 32212
rect 16908 32172 16914 32184
rect 20254 32172 20260 32224
rect 20312 32172 20318 32224
rect 24118 32172 24124 32224
rect 24176 32172 24182 32224
rect 1104 32122 24564 32144
rect 1104 32070 3882 32122
rect 3934 32070 3946 32122
rect 3998 32070 4010 32122
rect 4062 32070 4074 32122
rect 4126 32070 4138 32122
rect 4190 32070 9747 32122
rect 9799 32070 9811 32122
rect 9863 32070 9875 32122
rect 9927 32070 9939 32122
rect 9991 32070 10003 32122
rect 10055 32070 15612 32122
rect 15664 32070 15676 32122
rect 15728 32070 15740 32122
rect 15792 32070 15804 32122
rect 15856 32070 15868 32122
rect 15920 32070 21477 32122
rect 21529 32070 21541 32122
rect 21593 32070 21605 32122
rect 21657 32070 21669 32122
rect 21721 32070 21733 32122
rect 21785 32070 24564 32122
rect 1104 32048 24564 32070
rect 3694 32008 3700 32020
rect 2240 31980 3700 32008
rect 2240 31949 2268 31980
rect 3694 31968 3700 31980
rect 3752 31968 3758 32020
rect 3786 31968 3792 32020
rect 3844 32008 3850 32020
rect 3844 31980 4844 32008
rect 3844 31968 3850 31980
rect 4816 31949 4844 31980
rect 5166 31968 5172 32020
rect 5224 32008 5230 32020
rect 5442 32008 5448 32020
rect 5224 31980 5448 32008
rect 5224 31968 5230 31980
rect 5442 31968 5448 31980
rect 5500 31968 5506 32020
rect 6730 31968 6736 32020
rect 6788 31968 6794 32020
rect 8110 32008 8116 32020
rect 7576 31980 8116 32008
rect 2225 31943 2283 31949
rect 2225 31909 2237 31943
rect 2271 31909 2283 31943
rect 2225 31903 2283 31909
rect 4801 31943 4859 31949
rect 4801 31909 4813 31943
rect 4847 31909 4859 31943
rect 5350 31940 5356 31952
rect 4801 31903 4859 31909
rect 5000 31912 5356 31940
rect 3602 31872 3608 31884
rect 3252 31844 3608 31872
rect 1394 31764 1400 31816
rect 1452 31764 1458 31816
rect 1670 31764 1676 31816
rect 1728 31764 1734 31816
rect 2038 31764 2044 31816
rect 2096 31764 2102 31816
rect 2317 31807 2375 31813
rect 2317 31773 2329 31807
rect 2363 31773 2375 31807
rect 2590 31804 2596 31816
rect 2551 31776 2596 31804
rect 2317 31767 2375 31773
rect 1486 31696 1492 31748
rect 1544 31696 1550 31748
rect 2332 31736 2360 31767
rect 2590 31764 2596 31776
rect 2648 31764 2654 31816
rect 3142 31804 3148 31816
rect 2700 31776 3148 31804
rect 2700 31736 2728 31776
rect 3142 31764 3148 31776
rect 3200 31804 3206 31816
rect 3252 31804 3280 31844
rect 3602 31832 3608 31844
rect 3660 31872 3666 31884
rect 3789 31875 3847 31881
rect 3789 31872 3801 31875
rect 3660 31844 3801 31872
rect 3660 31832 3666 31844
rect 3789 31841 3801 31844
rect 3835 31841 3847 31875
rect 3789 31835 3847 31841
rect 5000 31816 5028 31912
rect 5350 31900 5356 31912
rect 5408 31900 5414 31952
rect 7576 31949 7604 31980
rect 8110 31968 8116 31980
rect 8168 31968 8174 32020
rect 8478 31968 8484 32020
rect 8536 31968 8542 32020
rect 8757 32011 8815 32017
rect 8757 31977 8769 32011
rect 8803 32008 8815 32011
rect 9122 32008 9128 32020
rect 8803 31980 9128 32008
rect 8803 31977 8815 31980
rect 8757 31971 8815 31977
rect 9122 31968 9128 31980
rect 9180 31968 9186 32020
rect 12618 32008 12624 32020
rect 10428 31980 12624 32008
rect 7561 31943 7619 31949
rect 7561 31909 7573 31943
rect 7607 31909 7619 31943
rect 8496 31940 8524 31968
rect 10428 31949 10456 31980
rect 12618 31968 12624 31980
rect 12676 31968 12682 32020
rect 13630 31968 13636 32020
rect 13688 32008 13694 32020
rect 16022 32008 16028 32020
rect 13688 31980 16028 32008
rect 13688 31968 13694 31980
rect 16022 31968 16028 31980
rect 16080 31968 16086 32020
rect 17402 32008 17408 32020
rect 16316 31980 17408 32008
rect 10413 31943 10471 31949
rect 8496 31912 8892 31940
rect 7561 31903 7619 31909
rect 5902 31832 5908 31884
rect 5960 31832 5966 31884
rect 7190 31872 7196 31884
rect 6840 31844 7196 31872
rect 3200 31776 3280 31804
rect 3200 31764 3206 31776
rect 3326 31764 3332 31816
rect 3384 31804 3390 31816
rect 4031 31807 4089 31813
rect 4031 31804 4043 31807
rect 3384 31776 4043 31804
rect 3384 31764 3390 31776
rect 4031 31773 4043 31776
rect 4077 31804 4089 31807
rect 4982 31804 4988 31816
rect 4077 31776 4988 31804
rect 4077 31773 4089 31776
rect 4031 31767 4089 31773
rect 4982 31764 4988 31776
rect 5040 31764 5046 31816
rect 5718 31764 5724 31816
rect 5776 31764 5782 31816
rect 5813 31807 5871 31813
rect 5813 31773 5825 31807
rect 5859 31804 5871 31807
rect 6840 31804 6868 31844
rect 7190 31832 7196 31844
rect 7248 31832 7254 31884
rect 8113 31875 8171 31881
rect 8113 31841 8125 31875
rect 8159 31872 8171 31875
rect 8662 31872 8668 31884
rect 8159 31844 8668 31872
rect 8159 31841 8171 31844
rect 8113 31835 8171 31841
rect 8662 31832 8668 31844
rect 8720 31832 8726 31884
rect 5859 31776 6868 31804
rect 6917 31807 6975 31813
rect 5859 31773 5871 31776
rect 5813 31767 5871 31773
rect 6917 31773 6929 31807
rect 6963 31804 6975 31807
rect 6963 31776 7052 31804
rect 6963 31773 6975 31776
rect 6917 31767 6975 31773
rect 5350 31736 5356 31748
rect 2332 31708 2728 31736
rect 3252 31708 5356 31736
rect 1504 31668 1532 31696
rect 1670 31668 1676 31680
rect 1504 31640 1676 31668
rect 1670 31628 1676 31640
rect 1728 31628 1734 31680
rect 2314 31628 2320 31680
rect 2372 31668 2378 31680
rect 3252 31668 3280 31708
rect 5350 31696 5356 31708
rect 5408 31736 5414 31748
rect 5445 31739 5503 31745
rect 5445 31736 5457 31739
rect 5408 31708 5457 31736
rect 5408 31696 5414 31708
rect 5445 31705 5457 31708
rect 5491 31705 5503 31739
rect 5445 31699 5503 31705
rect 2372 31640 3280 31668
rect 2372 31628 2378 31640
rect 3326 31628 3332 31680
rect 3384 31628 3390 31680
rect 3694 31628 3700 31680
rect 3752 31668 3758 31680
rect 5258 31668 5264 31680
rect 3752 31640 5264 31668
rect 3752 31628 3758 31640
rect 5258 31628 5264 31640
rect 5316 31628 5322 31680
rect 5736 31668 5764 31764
rect 5902 31696 5908 31748
rect 5960 31736 5966 31748
rect 6181 31739 6239 31745
rect 6181 31736 6193 31739
rect 5960 31708 6193 31736
rect 5960 31696 5966 31708
rect 6181 31705 6193 31708
rect 6227 31705 6239 31739
rect 6181 31699 6239 31705
rect 6454 31696 6460 31748
rect 6512 31736 6518 31748
rect 6549 31739 6607 31745
rect 6549 31736 6561 31739
rect 6512 31708 6561 31736
rect 6512 31696 6518 31708
rect 6549 31705 6561 31708
rect 6595 31705 6607 31739
rect 6549 31699 6607 31705
rect 5810 31668 5816 31680
rect 5736 31640 5816 31668
rect 5810 31628 5816 31640
rect 5868 31628 5874 31680
rect 6638 31628 6644 31680
rect 6696 31668 6702 31680
rect 6914 31668 6920 31680
rect 6696 31640 6920 31668
rect 6696 31628 6702 31640
rect 6914 31628 6920 31640
rect 6972 31628 6978 31680
rect 7024 31668 7052 31776
rect 7098 31764 7104 31816
rect 7156 31764 7162 31816
rect 7834 31764 7840 31816
rect 7892 31764 7898 31816
rect 8018 31813 8024 31816
rect 7975 31807 8024 31813
rect 7975 31773 7987 31807
rect 8021 31773 8024 31807
rect 7975 31767 8024 31773
rect 8018 31764 8024 31767
rect 8076 31764 8082 31816
rect 8864 31794 8892 31912
rect 10413 31909 10425 31943
rect 10459 31909 10471 31943
rect 10413 31903 10471 31909
rect 14182 31900 14188 31952
rect 14240 31940 14246 31952
rect 14918 31940 14924 31952
rect 14240 31912 14924 31940
rect 14240 31900 14246 31912
rect 14918 31900 14924 31912
rect 14976 31900 14982 31952
rect 8944 31884 8996 31890
rect 12342 31832 12348 31884
rect 12400 31832 12406 31884
rect 13998 31832 14004 31884
rect 14056 31872 14062 31884
rect 14734 31872 14740 31884
rect 14056 31844 14740 31872
rect 14056 31832 14062 31844
rect 14734 31832 14740 31844
rect 14792 31832 14798 31884
rect 16316 31881 16344 31980
rect 17402 31968 17408 31980
rect 17460 31968 17466 32020
rect 17954 31968 17960 32020
rect 18012 32008 18018 32020
rect 18874 32008 18880 32020
rect 18012 31980 18880 32008
rect 18012 31968 18018 31980
rect 18874 31968 18880 31980
rect 18932 31968 18938 32020
rect 19794 32008 19800 32020
rect 19260 31980 19800 32008
rect 17681 31943 17739 31949
rect 17681 31909 17693 31943
rect 17727 31940 17739 31943
rect 18785 31943 18843 31949
rect 17727 31912 18368 31940
rect 17727 31909 17739 31912
rect 17681 31903 17739 31909
rect 16301 31875 16359 31881
rect 16301 31841 16313 31875
rect 16347 31841 16359 31875
rect 16301 31835 16359 31841
rect 8944 31826 8996 31832
rect 9401 31807 9459 31813
rect 9401 31804 9413 31807
rect 9048 31794 9413 31804
rect 8864 31776 9413 31794
rect 8864 31766 9076 31776
rect 9401 31773 9413 31776
rect 9447 31773 9459 31807
rect 9401 31767 9459 31773
rect 9858 31764 9864 31816
rect 9916 31764 9922 31816
rect 11330 31764 11336 31816
rect 11388 31804 11394 31816
rect 12587 31807 12645 31813
rect 12587 31804 12599 31807
rect 11388 31776 12599 31804
rect 11388 31764 11394 31776
rect 12587 31773 12599 31776
rect 12633 31773 12645 31807
rect 12587 31767 12645 31773
rect 13170 31764 13176 31816
rect 13228 31804 13234 31816
rect 13630 31804 13636 31816
rect 13228 31776 13636 31804
rect 13228 31764 13234 31776
rect 13630 31764 13636 31776
rect 13688 31764 13694 31816
rect 14366 31764 14372 31816
rect 14424 31804 14430 31816
rect 14921 31807 14979 31813
rect 14921 31804 14933 31807
rect 14424 31776 14933 31804
rect 14424 31764 14430 31776
rect 14921 31773 14933 31776
rect 14967 31804 14979 31807
rect 14967 31776 15148 31804
rect 14967 31773 14979 31776
rect 14921 31767 14979 31773
rect 9490 31696 9496 31748
rect 9548 31696 9554 31748
rect 10778 31696 10784 31748
rect 10836 31736 10842 31748
rect 10836 31708 14504 31736
rect 10836 31696 10842 31708
rect 14476 31680 14504 31708
rect 7282 31668 7288 31680
rect 7024 31640 7288 31668
rect 7282 31628 7288 31640
rect 7340 31628 7346 31680
rect 7374 31628 7380 31680
rect 7432 31668 7438 31680
rect 7926 31668 7932 31680
rect 7432 31640 7932 31668
rect 7432 31628 7438 31640
rect 7926 31628 7932 31640
rect 7984 31628 7990 31680
rect 8018 31628 8024 31680
rect 8076 31668 8082 31680
rect 9125 31671 9183 31677
rect 9125 31668 9137 31671
rect 8076 31640 9137 31668
rect 8076 31628 8082 31640
rect 9125 31637 9137 31640
rect 9171 31668 9183 31671
rect 10134 31668 10140 31680
rect 9171 31640 10140 31668
rect 9171 31637 9183 31640
rect 9125 31631 9183 31637
rect 10134 31628 10140 31640
rect 10192 31628 10198 31680
rect 10226 31628 10232 31680
rect 10284 31628 10290 31680
rect 13170 31628 13176 31680
rect 13228 31668 13234 31680
rect 13357 31671 13415 31677
rect 13357 31668 13369 31671
rect 13228 31640 13369 31668
rect 13228 31628 13234 31640
rect 13357 31637 13369 31640
rect 13403 31637 13415 31671
rect 13357 31631 13415 31637
rect 14458 31628 14464 31680
rect 14516 31628 14522 31680
rect 15120 31668 15148 31776
rect 15194 31764 15200 31816
rect 15252 31804 15258 31816
rect 16316 31804 16344 31835
rect 15252 31776 15295 31804
rect 15488 31776 16344 31804
rect 16575 31807 16633 31813
rect 15252 31764 15258 31776
rect 15488 31668 15516 31776
rect 16575 31773 16587 31807
rect 16621 31804 16633 31807
rect 16666 31804 16672 31816
rect 16621 31776 16672 31804
rect 16621 31773 16633 31776
rect 16575 31767 16633 31773
rect 16666 31764 16672 31776
rect 16724 31804 16730 31816
rect 17402 31804 17408 31816
rect 16724 31776 17408 31804
rect 16724 31764 16730 31776
rect 17402 31764 17408 31776
rect 17460 31764 17466 31816
rect 18340 31813 18368 31912
rect 18785 31909 18797 31943
rect 18831 31940 18843 31943
rect 19260 31940 19288 31980
rect 19794 31968 19800 31980
rect 19852 31968 19858 32020
rect 20254 31968 20260 32020
rect 20312 32008 20318 32020
rect 23201 32011 23259 32017
rect 20312 31980 21220 32008
rect 20312 31968 20318 31980
rect 18831 31912 19288 31940
rect 19337 31943 19395 31949
rect 18831 31909 18843 31912
rect 18785 31903 18843 31909
rect 19337 31909 19349 31943
rect 19383 31909 19395 31943
rect 19337 31903 19395 31909
rect 19150 31832 19156 31884
rect 19208 31832 19214 31884
rect 19352 31872 19380 31903
rect 20346 31900 20352 31952
rect 20404 31900 20410 31952
rect 21085 31943 21143 31949
rect 21085 31909 21097 31943
rect 21131 31909 21143 31943
rect 21085 31903 21143 31909
rect 19981 31875 20039 31881
rect 19352 31844 19932 31872
rect 17865 31807 17923 31813
rect 17865 31804 17877 31807
rect 17512 31776 17877 31804
rect 17512 31680 17540 31776
rect 17865 31773 17877 31776
rect 17911 31773 17923 31807
rect 17865 31767 17923 31773
rect 18325 31807 18383 31813
rect 18325 31773 18337 31807
rect 18371 31773 18383 31807
rect 18325 31767 18383 31773
rect 18417 31807 18475 31813
rect 18417 31773 18429 31807
rect 18463 31804 18475 31807
rect 18782 31804 18788 31816
rect 18463 31776 18788 31804
rect 18463 31773 18475 31776
rect 18417 31767 18475 31773
rect 18782 31764 18788 31776
rect 18840 31764 18846 31816
rect 18966 31764 18972 31816
rect 19024 31764 19030 31816
rect 19168 31804 19196 31832
rect 19904 31813 19932 31844
rect 19981 31841 19993 31875
rect 20027 31872 20039 31875
rect 20901 31875 20959 31881
rect 20901 31872 20913 31875
rect 20027 31844 20392 31872
rect 20027 31841 20039 31844
rect 19981 31835 20039 31841
rect 19521 31807 19579 31813
rect 19521 31804 19533 31807
rect 19168 31776 19533 31804
rect 19521 31773 19533 31776
rect 19567 31773 19579 31807
rect 19521 31767 19579 31773
rect 19889 31807 19947 31813
rect 19889 31773 19901 31807
rect 19935 31773 19947 31807
rect 19889 31767 19947 31773
rect 20162 31764 20168 31816
rect 20220 31764 20226 31816
rect 20364 31813 20392 31844
rect 20732 31844 20913 31872
rect 20732 31813 20760 31844
rect 20901 31841 20913 31844
rect 20947 31841 20959 31875
rect 20901 31835 20959 31841
rect 20349 31807 20407 31813
rect 20349 31773 20361 31807
rect 20395 31773 20407 31807
rect 20349 31767 20407 31773
rect 20717 31807 20775 31813
rect 20717 31773 20729 31807
rect 20763 31773 20775 31807
rect 20717 31767 20775 31773
rect 20809 31807 20867 31813
rect 20809 31773 20821 31807
rect 20855 31804 20867 31807
rect 20993 31807 21051 31813
rect 20855 31776 20889 31804
rect 20855 31773 20867 31776
rect 20809 31767 20867 31773
rect 20993 31773 21005 31807
rect 21039 31804 21051 31807
rect 21100 31804 21128 31903
rect 21039 31776 21128 31804
rect 21192 31804 21220 31980
rect 23201 31977 23213 32011
rect 23247 32008 23259 32011
rect 23658 32008 23664 32020
rect 23247 31980 23664 32008
rect 23247 31977 23259 31980
rect 23201 31971 23259 31977
rect 23658 31968 23664 31980
rect 23716 31968 23722 32020
rect 22741 31943 22799 31949
rect 22741 31909 22753 31943
rect 22787 31909 22799 31943
rect 22741 31903 22799 31909
rect 23477 31943 23535 31949
rect 23477 31909 23489 31943
rect 23523 31909 23535 31943
rect 23477 31903 23535 31909
rect 22756 31872 22784 31903
rect 23492 31872 23520 31903
rect 22756 31844 23336 31872
rect 23492 31844 23888 31872
rect 21269 31807 21327 31813
rect 21269 31804 21281 31807
rect 21192 31776 21281 31804
rect 21039 31773 21051 31776
rect 20993 31767 21051 31773
rect 21269 31773 21281 31776
rect 21315 31773 21327 31807
rect 22925 31807 22983 31813
rect 22925 31804 22937 31807
rect 21269 31767 21327 31773
rect 21836 31776 22937 31804
rect 20180 31736 20208 31764
rect 20824 31736 20852 31767
rect 20180 31708 20852 31736
rect 21836 31680 21864 31776
rect 22925 31773 22937 31776
rect 22971 31773 22983 31807
rect 22925 31767 22983 31773
rect 23308 31736 23336 31844
rect 23382 31764 23388 31816
rect 23440 31764 23446 31816
rect 23860 31813 23888 31844
rect 23661 31807 23719 31813
rect 23661 31804 23673 31807
rect 23492 31776 23673 31804
rect 23492 31736 23520 31776
rect 23661 31773 23673 31776
rect 23707 31773 23719 31807
rect 23661 31767 23719 31773
rect 23845 31807 23903 31813
rect 23845 31773 23857 31807
rect 23891 31773 23903 31807
rect 23845 31767 23903 31773
rect 24213 31807 24271 31813
rect 24213 31773 24225 31807
rect 24259 31804 24271 31807
rect 25038 31804 25044 31816
rect 24259 31776 25044 31804
rect 24259 31773 24271 31776
rect 24213 31767 24271 31773
rect 25038 31764 25044 31776
rect 25096 31764 25102 31816
rect 23308 31708 23520 31736
rect 15120 31640 15516 31668
rect 15930 31628 15936 31680
rect 15988 31628 15994 31680
rect 17310 31628 17316 31680
rect 17368 31628 17374 31680
rect 17494 31628 17500 31680
rect 17552 31628 17558 31680
rect 20714 31628 20720 31680
rect 20772 31668 20778 31680
rect 21818 31668 21824 31680
rect 20772 31640 21824 31668
rect 20772 31628 20778 31640
rect 21818 31628 21824 31640
rect 21876 31628 21882 31680
rect 1104 31578 24723 31600
rect 1104 31526 6814 31578
rect 6866 31526 6878 31578
rect 6930 31526 6942 31578
rect 6994 31526 7006 31578
rect 7058 31526 7070 31578
rect 7122 31526 12679 31578
rect 12731 31526 12743 31578
rect 12795 31526 12807 31578
rect 12859 31526 12871 31578
rect 12923 31526 12935 31578
rect 12987 31526 18544 31578
rect 18596 31526 18608 31578
rect 18660 31526 18672 31578
rect 18724 31526 18736 31578
rect 18788 31526 18800 31578
rect 18852 31526 24409 31578
rect 24461 31526 24473 31578
rect 24525 31526 24537 31578
rect 24589 31526 24601 31578
rect 24653 31526 24665 31578
rect 24717 31526 24723 31578
rect 1104 31504 24723 31526
rect 3145 31467 3203 31473
rect 3145 31433 3157 31467
rect 3191 31464 3203 31467
rect 4430 31464 4436 31476
rect 3191 31436 4436 31464
rect 3191 31433 3203 31436
rect 3145 31427 3203 31433
rect 4430 31424 4436 31436
rect 4488 31424 4494 31476
rect 4522 31424 4528 31476
rect 4580 31424 4586 31476
rect 4709 31467 4767 31473
rect 4709 31433 4721 31467
rect 4755 31464 4767 31467
rect 7742 31464 7748 31476
rect 4755 31436 7748 31464
rect 4755 31433 4767 31436
rect 4709 31427 4767 31433
rect 7742 31424 7748 31436
rect 7800 31424 7806 31476
rect 8481 31467 8539 31473
rect 8481 31433 8493 31467
rect 8527 31464 8539 31467
rect 8754 31464 8760 31476
rect 8527 31436 8760 31464
rect 8527 31433 8539 31436
rect 8481 31427 8539 31433
rect 8754 31424 8760 31436
rect 8812 31424 8818 31476
rect 9490 31424 9496 31476
rect 9548 31464 9554 31476
rect 9766 31464 9772 31476
rect 9548 31436 9772 31464
rect 9548 31424 9554 31436
rect 9766 31424 9772 31436
rect 9824 31424 9830 31476
rect 9950 31424 9956 31476
rect 10008 31464 10014 31476
rect 10413 31467 10471 31473
rect 10413 31464 10425 31467
rect 10008 31436 10425 31464
rect 10008 31424 10014 31436
rect 10413 31433 10425 31436
rect 10459 31433 10471 31467
rect 10413 31427 10471 31433
rect 11698 31424 11704 31476
rect 11756 31464 11762 31476
rect 12066 31464 12072 31476
rect 11756 31436 12072 31464
rect 11756 31424 11762 31436
rect 12066 31424 12072 31436
rect 12124 31424 12130 31476
rect 13262 31424 13268 31476
rect 13320 31464 13326 31476
rect 13722 31464 13728 31476
rect 13320 31436 13728 31464
rect 13320 31424 13326 31436
rect 13722 31424 13728 31436
rect 13780 31424 13786 31476
rect 14458 31424 14464 31476
rect 14516 31464 14522 31476
rect 18601 31467 18659 31473
rect 14516 31436 18184 31464
rect 14516 31424 14522 31436
rect 1394 31356 1400 31408
rect 1452 31356 1458 31408
rect 2685 31399 2743 31405
rect 2685 31365 2697 31399
rect 2731 31396 2743 31399
rect 2731 31365 2753 31396
rect 2685 31362 2753 31365
rect 2792 31368 3188 31396
rect 2792 31362 2820 31368
rect 2685 31359 2820 31362
rect 1302 31288 1308 31340
rect 1360 31328 1366 31340
rect 2409 31331 2467 31337
rect 2725 31334 2820 31359
rect 2409 31328 2421 31331
rect 1360 31300 2421 31328
rect 1360 31288 1366 31300
rect 2409 31297 2421 31300
rect 2455 31297 2467 31331
rect 2961 31331 3019 31337
rect 2961 31328 2973 31331
rect 2409 31291 2467 31297
rect 2884 31300 2973 31328
rect 2884 31272 2912 31300
rect 2961 31297 2973 31300
rect 3007 31297 3019 31331
rect 3160 31328 3188 31368
rect 3234 31356 3240 31408
rect 3292 31396 3298 31408
rect 3421 31399 3479 31405
rect 3421 31396 3433 31399
rect 3292 31368 3433 31396
rect 3292 31356 3298 31368
rect 3421 31365 3433 31368
rect 3467 31365 3479 31399
rect 3421 31359 3479 31365
rect 3528 31368 4752 31396
rect 3528 31328 3556 31368
rect 3160 31300 3556 31328
rect 2961 31291 3019 31297
rect 3602 31288 3608 31340
rect 3660 31328 3666 31340
rect 3697 31331 3755 31337
rect 3697 31328 3709 31331
rect 3660 31300 3709 31328
rect 3660 31288 3666 31300
rect 3697 31297 3709 31300
rect 3743 31297 3755 31331
rect 3697 31291 3755 31297
rect 3789 31331 3847 31337
rect 3789 31297 3801 31331
rect 3835 31328 3847 31331
rect 3970 31328 3976 31340
rect 3835 31300 3976 31328
rect 3835 31297 3847 31300
rect 3789 31291 3847 31297
rect 3970 31288 3976 31300
rect 4028 31288 4034 31340
rect 4157 31331 4215 31337
rect 4157 31297 4169 31331
rect 4203 31328 4215 31331
rect 4614 31328 4620 31340
rect 4203 31300 4620 31328
rect 4203 31297 4215 31300
rect 4157 31291 4215 31297
rect 4614 31288 4620 31300
rect 4672 31288 4678 31340
rect 1762 31220 1768 31272
rect 1820 31260 1826 31272
rect 2133 31263 2191 31269
rect 2133 31260 2145 31263
rect 1820 31232 2145 31260
rect 1820 31220 1826 31232
rect 2133 31229 2145 31232
rect 2179 31260 2191 31263
rect 2222 31260 2228 31272
rect 2179 31232 2228 31260
rect 2179 31229 2191 31232
rect 2133 31223 2191 31229
rect 2222 31220 2228 31232
rect 2280 31220 2286 31272
rect 2866 31220 2872 31272
rect 2924 31220 2930 31272
rect 3326 31220 3332 31272
rect 3384 31220 3390 31272
rect 4724 31124 4752 31368
rect 4798 31356 4804 31408
rect 4856 31396 4862 31408
rect 5442 31396 5448 31408
rect 4856 31368 5448 31396
rect 4856 31356 4862 31368
rect 5442 31356 5448 31368
rect 5500 31396 5506 31408
rect 5994 31396 6000 31408
rect 5500 31368 6000 31396
rect 5500 31356 5506 31368
rect 5994 31356 6000 31368
rect 6052 31356 6058 31408
rect 7668 31368 8708 31396
rect 5166 31328 5172 31340
rect 5127 31300 5172 31328
rect 5166 31288 5172 31300
rect 5224 31288 5230 31340
rect 5258 31288 5264 31340
rect 5316 31328 5322 31340
rect 5316 31300 7218 31328
rect 5316 31288 5322 31300
rect 4893 31263 4951 31269
rect 4893 31229 4905 31263
rect 4939 31229 4951 31263
rect 4893 31223 4951 31229
rect 4798 31152 4804 31204
rect 4856 31192 4862 31204
rect 4908 31192 4936 31223
rect 7098 31192 7104 31204
rect 4856 31164 4936 31192
rect 5828 31164 7104 31192
rect 4856 31152 4862 31164
rect 5828 31124 5856 31164
rect 7098 31152 7104 31164
rect 7156 31152 7162 31204
rect 4724 31096 5856 31124
rect 5902 31084 5908 31136
rect 5960 31084 5966 31136
rect 7190 31124 7218 31300
rect 7466 31288 7472 31340
rect 7524 31328 7530 31340
rect 7668 31328 7696 31368
rect 7524 31300 7696 31328
rect 7743 31331 7801 31337
rect 7524 31288 7530 31300
rect 7743 31297 7755 31331
rect 7789 31328 7801 31331
rect 8202 31328 8208 31340
rect 7789 31300 8208 31328
rect 7789 31297 7801 31300
rect 7743 31291 7801 31297
rect 8202 31288 8208 31300
rect 8260 31328 8266 31340
rect 8570 31328 8576 31340
rect 8260 31300 8576 31328
rect 8260 31288 8266 31300
rect 8570 31288 8576 31300
rect 8628 31288 8634 31340
rect 8680 31260 8708 31368
rect 9122 31356 9128 31408
rect 9180 31396 9186 31408
rect 9180 31368 12480 31396
rect 9180 31356 9186 31368
rect 9030 31288 9036 31340
rect 9088 31328 9094 31340
rect 9674 31337 9680 31340
rect 9643 31331 9680 31337
rect 9643 31328 9655 31331
rect 9088 31300 9655 31328
rect 9088 31288 9094 31300
rect 9643 31297 9655 31300
rect 9643 31291 9680 31297
rect 9674 31288 9680 31291
rect 9732 31288 9738 31340
rect 10318 31288 10324 31340
rect 10376 31328 10382 31340
rect 10962 31328 10968 31340
rect 10376 31300 10968 31328
rect 10376 31288 10382 31300
rect 10962 31288 10968 31300
rect 11020 31288 11026 31340
rect 11698 31328 11704 31340
rect 11072 31300 11704 31328
rect 9401 31263 9459 31269
rect 9401 31260 9413 31263
rect 8680 31232 9413 31260
rect 9401 31229 9413 31232
rect 9447 31229 9459 31263
rect 9401 31223 9459 31229
rect 11072 31204 11100 31300
rect 11698 31288 11704 31300
rect 11756 31288 11762 31340
rect 12342 31288 12348 31340
rect 12400 31288 12406 31340
rect 12452 31328 12480 31368
rect 13630 31356 13636 31408
rect 13688 31356 13694 31408
rect 14458 31367 14486 31424
rect 18156 31408 18184 31436
rect 18601 31433 18613 31467
rect 18647 31464 18659 31467
rect 18966 31464 18972 31476
rect 18647 31436 18972 31464
rect 18647 31433 18659 31436
rect 18601 31427 18659 31433
rect 18966 31424 18972 31436
rect 19024 31424 19030 31476
rect 19889 31467 19947 31473
rect 19889 31433 19901 31467
rect 19935 31464 19947 31467
rect 20162 31464 20168 31476
rect 19935 31436 20168 31464
rect 19935 31433 19947 31436
rect 19889 31427 19947 31433
rect 20162 31424 20168 31436
rect 20220 31424 20226 31476
rect 23385 31467 23443 31473
rect 23385 31433 23397 31467
rect 23431 31433 23443 31467
rect 23385 31427 23443 31433
rect 14443 31361 14501 31367
rect 13079 31331 13137 31337
rect 13079 31328 13091 31331
rect 12452 31300 13091 31328
rect 13079 31297 13091 31300
rect 13125 31328 13137 31331
rect 13648 31328 13676 31356
rect 13125 31300 13676 31328
rect 14185 31331 14243 31337
rect 13125 31297 13137 31300
rect 13079 31291 13137 31297
rect 14185 31297 14197 31331
rect 14231 31297 14243 31331
rect 14443 31327 14455 31361
rect 14489 31327 14501 31361
rect 14550 31356 14556 31408
rect 14608 31356 14614 31408
rect 17236 31368 18000 31396
rect 14443 31321 14501 31327
rect 14568 31328 14596 31356
rect 17236 31337 17264 31368
rect 17972 31340 18000 31368
rect 18138 31356 18144 31408
rect 18196 31356 18202 31408
rect 18874 31356 18880 31408
rect 18932 31396 18938 31408
rect 23400 31396 23428 31427
rect 18932 31368 20300 31396
rect 23400 31368 23980 31396
rect 18932 31356 18938 31368
rect 17494 31337 17500 31340
rect 17221 31331 17279 31337
rect 14568 31300 17172 31328
rect 14185 31291 14243 31297
rect 12066 31220 12072 31272
rect 12124 31260 12130 31272
rect 12360 31260 12388 31288
rect 12802 31260 12808 31272
rect 12124 31232 12808 31260
rect 12124 31220 12130 31232
rect 12802 31220 12808 31232
rect 12860 31220 12866 31272
rect 14090 31220 14096 31272
rect 14148 31260 14154 31272
rect 14200 31260 14228 31291
rect 14148 31232 14228 31260
rect 14148 31220 14154 31232
rect 8956 31164 9534 31192
rect 8956 31124 8984 31164
rect 7190 31096 8984 31124
rect 9030 31084 9036 31136
rect 9088 31084 9094 31136
rect 9506 31124 9534 31164
rect 11054 31152 11060 31204
rect 11112 31152 11118 31204
rect 11882 31152 11888 31204
rect 11940 31152 11946 31204
rect 12250 31124 12256 31136
rect 9506 31096 12256 31124
rect 12250 31084 12256 31096
rect 12308 31124 12314 31136
rect 13630 31124 13636 31136
rect 12308 31096 13636 31124
rect 12308 31084 12314 31096
rect 13630 31084 13636 31096
rect 13688 31084 13694 31136
rect 13814 31084 13820 31136
rect 13872 31084 13878 31136
rect 14458 31084 14464 31136
rect 14516 31124 14522 31136
rect 15197 31127 15255 31133
rect 15197 31124 15209 31127
rect 14516 31096 15209 31124
rect 14516 31084 14522 31096
rect 15197 31093 15209 31096
rect 15243 31093 15255 31127
rect 17144 31124 17172 31300
rect 17221 31297 17233 31331
rect 17267 31297 17279 31331
rect 17488 31328 17500 31337
rect 17455 31300 17500 31328
rect 17221 31291 17279 31297
rect 17488 31291 17500 31300
rect 17494 31288 17500 31291
rect 17552 31288 17558 31340
rect 17954 31288 17960 31340
rect 18012 31288 18018 31340
rect 19058 31328 19064 31340
rect 18892 31300 19064 31328
rect 18414 31220 18420 31272
rect 18472 31260 18478 31272
rect 18892 31269 18920 31300
rect 19058 31288 19064 31300
rect 19116 31288 19122 31340
rect 19151 31331 19209 31337
rect 19151 31297 19163 31331
rect 19197 31328 19209 31331
rect 19242 31328 19248 31340
rect 19197 31300 19248 31328
rect 19197 31297 19209 31300
rect 19151 31291 19209 31297
rect 19242 31288 19248 31300
rect 19300 31288 19306 31340
rect 20272 31337 20300 31368
rect 20257 31331 20315 31337
rect 20257 31297 20269 31331
rect 20303 31297 20315 31331
rect 20513 31331 20571 31337
rect 20513 31328 20525 31331
rect 20257 31291 20315 31297
rect 20364 31300 20525 31328
rect 18877 31263 18935 31269
rect 18877 31260 18889 31263
rect 18472 31232 18889 31260
rect 18472 31220 18478 31232
rect 18877 31229 18889 31232
rect 18923 31229 18935 31263
rect 20364 31260 20392 31300
rect 20513 31297 20525 31300
rect 20559 31297 20571 31331
rect 20513 31291 20571 31297
rect 23566 31288 23572 31340
rect 23624 31288 23630 31340
rect 23842 31288 23848 31340
rect 23900 31288 23906 31340
rect 23952 31337 23980 31368
rect 23937 31331 23995 31337
rect 23937 31297 23949 31331
rect 23983 31297 23995 31331
rect 23937 31291 23995 31297
rect 18877 31223 18935 31229
rect 20272 31232 20392 31260
rect 20272 31124 20300 31232
rect 20438 31124 20444 31136
rect 17144 31096 20444 31124
rect 15197 31087 15255 31093
rect 20438 31084 20444 31096
rect 20496 31084 20502 31136
rect 21637 31127 21695 31133
rect 21637 31093 21649 31127
rect 21683 31124 21695 31127
rect 23198 31124 23204 31136
rect 21683 31096 23204 31124
rect 21683 31093 21695 31096
rect 21637 31087 21695 31093
rect 23198 31084 23204 31096
rect 23256 31084 23262 31136
rect 23658 31084 23664 31136
rect 23716 31084 23722 31136
rect 24118 31084 24124 31136
rect 24176 31084 24182 31136
rect 1104 31034 24564 31056
rect 1104 30982 3882 31034
rect 3934 30982 3946 31034
rect 3998 30982 4010 31034
rect 4062 30982 4074 31034
rect 4126 30982 4138 31034
rect 4190 30982 9747 31034
rect 9799 30982 9811 31034
rect 9863 30982 9875 31034
rect 9927 30982 9939 31034
rect 9991 30982 10003 31034
rect 10055 30982 15612 31034
rect 15664 30982 15676 31034
rect 15728 30982 15740 31034
rect 15792 30982 15804 31034
rect 15856 30982 15868 31034
rect 15920 30982 21477 31034
rect 21529 30982 21541 31034
rect 21593 30982 21605 31034
rect 21657 30982 21669 31034
rect 21721 30982 21733 31034
rect 21785 30982 24564 31034
rect 1104 30960 24564 30982
rect 1670 30920 1676 30932
rect 1412 30892 1676 30920
rect 1412 30796 1440 30892
rect 1670 30880 1676 30892
rect 1728 30880 1734 30932
rect 2866 30880 2872 30932
rect 2924 30920 2930 30932
rect 3970 30920 3976 30932
rect 2924 30892 3976 30920
rect 2924 30880 2930 30892
rect 3970 30880 3976 30892
rect 4028 30920 4034 30932
rect 4430 30920 4436 30932
rect 4028 30892 4436 30920
rect 4028 30880 4034 30892
rect 4430 30880 4436 30892
rect 4488 30880 4494 30932
rect 5902 30880 5908 30932
rect 5960 30880 5966 30932
rect 5994 30880 6000 30932
rect 6052 30880 6058 30932
rect 7190 30880 7196 30932
rect 7248 30920 7254 30932
rect 7377 30923 7435 30929
rect 7377 30920 7389 30923
rect 7248 30892 7389 30920
rect 7248 30880 7254 30892
rect 7377 30889 7389 30892
rect 7423 30889 7435 30923
rect 10778 30920 10784 30932
rect 7377 30883 7435 30889
rect 9646 30892 10784 30920
rect 1394 30744 1400 30796
rect 1452 30744 1458 30796
rect 3053 30787 3111 30793
rect 3053 30753 3065 30787
rect 3099 30784 3111 30787
rect 3099 30756 4384 30784
rect 3099 30753 3111 30756
rect 3053 30747 3111 30753
rect 1671 30719 1729 30725
rect 1671 30685 1683 30719
rect 1717 30716 1729 30719
rect 2406 30716 2412 30728
rect 1717 30688 2412 30716
rect 1717 30685 1729 30688
rect 1671 30679 1729 30685
rect 2406 30676 2412 30688
rect 2464 30676 2470 30728
rect 2774 30676 2780 30728
rect 2832 30676 2838 30728
rect 2038 30540 2044 30592
rect 2096 30580 2102 30592
rect 2409 30583 2467 30589
rect 2409 30580 2421 30583
rect 2096 30552 2421 30580
rect 2096 30540 2102 30552
rect 2409 30549 2421 30552
rect 2455 30549 2467 30583
rect 2409 30543 2467 30549
rect 4154 30540 4160 30592
rect 4212 30540 4218 30592
rect 4356 30580 4384 30756
rect 4890 30744 4896 30796
rect 4948 30744 4954 30796
rect 4985 30719 5043 30725
rect 4985 30685 4997 30719
rect 5031 30716 5043 30719
rect 5920 30716 5948 30880
rect 6012 30784 6040 30880
rect 7466 30812 7472 30864
rect 7524 30852 7530 30864
rect 9646 30852 9674 30892
rect 10778 30880 10784 30892
rect 10836 30880 10842 30932
rect 17037 30923 17095 30929
rect 17037 30889 17049 30923
rect 17083 30920 17095 30923
rect 17494 30920 17500 30932
rect 17083 30892 17500 30920
rect 17083 30889 17095 30892
rect 17037 30883 17095 30889
rect 17494 30880 17500 30892
rect 17552 30880 17558 30932
rect 19334 30880 19340 30932
rect 19392 30880 19398 30932
rect 19429 30923 19487 30929
rect 19429 30889 19441 30923
rect 19475 30920 19487 30923
rect 23293 30923 23351 30929
rect 19475 30892 23152 30920
rect 19475 30889 19487 30892
rect 19429 30883 19487 30889
rect 7524 30824 9674 30852
rect 7524 30812 7530 30824
rect 10226 30812 10232 30864
rect 10284 30852 10290 30864
rect 10284 30824 10732 30852
rect 10284 30812 10290 30824
rect 6365 30787 6423 30793
rect 6365 30784 6377 30787
rect 6012 30756 6377 30784
rect 6365 30753 6377 30756
rect 6411 30753 6423 30787
rect 6365 30747 6423 30753
rect 7098 30744 7104 30796
rect 7156 30784 7162 30796
rect 10502 30784 10508 30796
rect 7156 30756 10508 30784
rect 7156 30744 7162 30756
rect 10502 30744 10508 30756
rect 10560 30744 10566 30796
rect 10704 30793 10732 30824
rect 14826 30812 14832 30864
rect 14884 30852 14890 30864
rect 15102 30852 15108 30864
rect 14884 30824 15108 30852
rect 14884 30812 14890 30824
rect 15102 30812 15108 30824
rect 15160 30812 15166 30864
rect 15194 30812 15200 30864
rect 15252 30852 15258 30864
rect 15562 30852 15568 30864
rect 15252 30824 15568 30852
rect 15252 30812 15258 30824
rect 15562 30812 15568 30824
rect 15620 30812 15626 30864
rect 15841 30855 15899 30861
rect 15841 30821 15853 30855
rect 15887 30852 15899 30855
rect 15930 30852 15936 30864
rect 15887 30824 15936 30852
rect 15887 30821 15899 30824
rect 15841 30815 15899 30821
rect 15930 30812 15936 30824
rect 15988 30812 15994 30864
rect 18785 30855 18843 30861
rect 18785 30821 18797 30855
rect 18831 30821 18843 30855
rect 18785 30815 18843 30821
rect 10689 30787 10747 30793
rect 10689 30753 10701 30787
rect 10735 30753 10747 30787
rect 10689 30747 10747 30753
rect 5031 30688 5948 30716
rect 5031 30685 5043 30688
rect 4985 30679 5043 30685
rect 6178 30676 6184 30728
rect 6236 30716 6242 30728
rect 6607 30719 6665 30725
rect 6607 30716 6619 30719
rect 6236 30688 6619 30716
rect 6236 30676 6242 30688
rect 6607 30685 6619 30688
rect 6653 30716 6665 30719
rect 7374 30716 7380 30728
rect 6653 30688 7380 30716
rect 6653 30685 6665 30688
rect 6607 30679 6665 30685
rect 7374 30676 7380 30688
rect 7432 30676 7438 30728
rect 8110 30676 8116 30728
rect 8168 30716 8174 30728
rect 10042 30716 10048 30728
rect 8168 30688 10048 30716
rect 8168 30676 8174 30688
rect 10042 30676 10048 30688
rect 10100 30716 10106 30728
rect 10704 30716 10732 30747
rect 13078 30744 13084 30796
rect 13136 30744 13142 30796
rect 16234 30787 16292 30793
rect 16234 30784 16246 30787
rect 14936 30756 16246 30784
rect 14936 30728 14964 30756
rect 16234 30753 16246 30756
rect 16280 30753 16292 30787
rect 16234 30747 16292 30753
rect 16393 30787 16451 30793
rect 16393 30753 16405 30787
rect 16439 30784 16451 30787
rect 17310 30784 17316 30796
rect 16439 30756 17316 30784
rect 16439 30753 16451 30756
rect 16393 30747 16451 30753
rect 17310 30744 17316 30756
rect 17368 30744 17374 30796
rect 10962 30725 10968 30728
rect 10100 30688 10732 30716
rect 10931 30719 10968 30725
rect 10100 30676 10106 30688
rect 10931 30685 10943 30719
rect 10931 30679 10968 30685
rect 10962 30676 10968 30679
rect 11020 30676 11026 30728
rect 12066 30676 12072 30728
rect 12124 30676 12130 30728
rect 12713 30719 12771 30725
rect 12713 30685 12725 30719
rect 12759 30716 12771 30719
rect 13170 30716 13176 30728
rect 12759 30688 13176 30716
rect 12759 30685 12771 30688
rect 12713 30679 12771 30685
rect 13170 30676 13176 30688
rect 13228 30676 13234 30728
rect 13630 30676 13636 30728
rect 13688 30716 13694 30728
rect 14918 30716 14924 30728
rect 13688 30688 14924 30716
rect 13688 30676 13694 30688
rect 14918 30676 14924 30688
rect 14976 30676 14982 30728
rect 15194 30676 15200 30728
rect 15252 30676 15258 30728
rect 15381 30719 15439 30725
rect 15381 30685 15393 30719
rect 15427 30685 15439 30719
rect 15381 30679 15439 30685
rect 4893 30651 4951 30657
rect 4893 30617 4905 30651
rect 4939 30648 4951 30651
rect 5258 30648 5264 30660
rect 4939 30620 5264 30648
rect 4939 30617 4951 30620
rect 4893 30611 4951 30617
rect 5258 30608 5264 30620
rect 5316 30608 5322 30660
rect 5353 30651 5411 30657
rect 5353 30617 5365 30651
rect 5399 30617 5411 30651
rect 5353 30611 5411 30617
rect 4430 30580 4436 30592
rect 4356 30552 4436 30580
rect 4430 30540 4436 30552
rect 4488 30540 4494 30592
rect 4614 30540 4620 30592
rect 4672 30540 4678 30592
rect 4798 30540 4804 30592
rect 4856 30580 4862 30592
rect 5368 30580 5396 30611
rect 5718 30608 5724 30660
rect 5776 30648 5782 30660
rect 12084 30648 12112 30676
rect 5776 30620 9628 30648
rect 5776 30608 5782 30620
rect 9600 30592 9628 30620
rect 11532 30620 12112 30648
rect 11532 30592 11560 30620
rect 12250 30608 12256 30660
rect 12308 30648 12314 30660
rect 12345 30651 12403 30657
rect 12345 30648 12357 30651
rect 12308 30620 12357 30648
rect 12308 30608 12314 30620
rect 12345 30617 12357 30620
rect 12391 30617 12403 30651
rect 12621 30651 12679 30657
rect 12621 30648 12633 30651
rect 12345 30611 12403 30617
rect 12452 30620 12633 30648
rect 4856 30552 5396 30580
rect 4856 30540 4862 30552
rect 5902 30540 5908 30592
rect 5960 30580 5966 30592
rect 6362 30580 6368 30592
rect 5960 30552 6368 30580
rect 5960 30540 5966 30552
rect 6362 30540 6368 30552
rect 6420 30540 6426 30592
rect 7558 30540 7564 30592
rect 7616 30580 7622 30592
rect 7926 30580 7932 30592
rect 7616 30552 7932 30580
rect 7616 30540 7622 30552
rect 7926 30540 7932 30552
rect 7984 30540 7990 30592
rect 9582 30540 9588 30592
rect 9640 30540 9646 30592
rect 11146 30540 11152 30592
rect 11204 30580 11210 30592
rect 11330 30580 11336 30592
rect 11204 30552 11336 30580
rect 11204 30540 11210 30552
rect 11330 30540 11336 30552
rect 11388 30540 11394 30592
rect 11514 30540 11520 30592
rect 11572 30540 11578 30592
rect 11698 30540 11704 30592
rect 11756 30540 11762 30592
rect 12066 30540 12072 30592
rect 12124 30580 12130 30592
rect 12452 30580 12480 30620
rect 12621 30617 12633 30620
rect 12667 30648 12679 30651
rect 12986 30648 12992 30660
rect 12667 30620 12992 30648
rect 12667 30617 12679 30620
rect 12621 30611 12679 30617
rect 12986 30608 12992 30620
rect 13044 30608 13050 30660
rect 13081 30651 13139 30657
rect 13081 30617 13093 30651
rect 13127 30617 13139 30651
rect 13081 30611 13139 30617
rect 12124 30552 12480 30580
rect 12124 30540 12130 30552
rect 12526 30540 12532 30592
rect 12584 30580 12590 30592
rect 13096 30580 13124 30611
rect 12584 30552 13124 30580
rect 12584 30540 12590 30552
rect 13446 30540 13452 30592
rect 13504 30540 13510 30592
rect 13630 30540 13636 30592
rect 13688 30540 13694 30592
rect 14274 30540 14280 30592
rect 14332 30580 14338 30592
rect 14826 30580 14832 30592
rect 14332 30552 14832 30580
rect 14332 30540 14338 30552
rect 14826 30540 14832 30552
rect 14884 30580 14890 30592
rect 15396 30580 15424 30679
rect 16114 30676 16120 30728
rect 16172 30676 16178 30728
rect 17773 30719 17831 30725
rect 17773 30685 17785 30719
rect 17819 30685 17831 30719
rect 17773 30679 17831 30685
rect 18047 30719 18105 30725
rect 18047 30685 18059 30719
rect 18093 30716 18105 30719
rect 18138 30716 18144 30728
rect 18093 30688 18144 30716
rect 18093 30685 18105 30688
rect 18047 30679 18105 30685
rect 17494 30608 17500 30660
rect 17552 30648 17558 30660
rect 17788 30648 17816 30679
rect 18138 30676 18144 30688
rect 18196 30676 18202 30728
rect 18800 30716 18828 30815
rect 20438 30812 20444 30864
rect 20496 30812 20502 30864
rect 23017 30855 23075 30861
rect 23017 30821 23029 30855
rect 23063 30821 23075 30855
rect 23017 30815 23075 30821
rect 19521 30787 19579 30793
rect 19521 30753 19533 30787
rect 19567 30784 19579 30787
rect 19705 30787 19763 30793
rect 19705 30784 19717 30787
rect 19567 30756 19717 30784
rect 19567 30753 19579 30756
rect 19521 30747 19579 30753
rect 19705 30753 19717 30756
rect 19751 30753 19763 30787
rect 19705 30747 19763 30753
rect 19245 30719 19303 30725
rect 19245 30716 19257 30719
rect 18800 30688 19257 30716
rect 19245 30685 19257 30688
rect 19291 30716 19303 30719
rect 19613 30719 19671 30725
rect 19613 30716 19625 30719
rect 19291 30688 19625 30716
rect 19291 30685 19303 30688
rect 19245 30679 19303 30685
rect 19613 30685 19625 30688
rect 19659 30685 19671 30719
rect 19613 30679 19671 30685
rect 19794 30676 19800 30728
rect 19852 30676 19858 30728
rect 20456 30716 20484 30812
rect 20990 30744 20996 30796
rect 21048 30784 21054 30796
rect 21361 30787 21419 30793
rect 21361 30784 21373 30787
rect 21048 30756 21373 30784
rect 21048 30744 21054 30756
rect 21361 30753 21373 30756
rect 21407 30753 21419 30787
rect 21361 30747 21419 30753
rect 21269 30719 21327 30725
rect 21269 30716 21281 30719
rect 20456 30688 21281 30716
rect 21269 30685 21281 30688
rect 21315 30685 21327 30719
rect 21269 30679 21327 30685
rect 21376 30648 21404 30747
rect 22741 30719 22799 30725
rect 21619 30689 21677 30695
rect 21619 30655 21631 30689
rect 21665 30686 21677 30689
rect 21665 30655 21680 30686
rect 22741 30685 22753 30719
rect 22787 30685 22799 30719
rect 22741 30679 22799 30685
rect 22925 30719 22983 30725
rect 22925 30685 22937 30719
rect 22971 30716 22983 30719
rect 23032 30716 23060 30815
rect 22971 30688 23060 30716
rect 22971 30685 22983 30688
rect 22925 30679 22983 30685
rect 21619 30649 21680 30655
rect 17552 30620 21404 30648
rect 21652 30648 21680 30649
rect 21818 30648 21824 30660
rect 21652 30620 21824 30648
rect 17552 30608 17558 30620
rect 21818 30608 21824 30620
rect 21876 30608 21882 30660
rect 14884 30552 15424 30580
rect 14884 30540 14890 30552
rect 21082 30540 21088 30592
rect 21140 30540 21146 30592
rect 22186 30540 22192 30592
rect 22244 30580 22250 30592
rect 22373 30583 22431 30589
rect 22373 30580 22385 30583
rect 22244 30552 22385 30580
rect 22244 30540 22250 30552
rect 22373 30549 22385 30552
rect 22419 30580 22431 30583
rect 22756 30580 22784 30679
rect 22419 30552 22784 30580
rect 22419 30549 22431 30552
rect 22373 30543 22431 30549
rect 22830 30540 22836 30592
rect 22888 30540 22894 30592
rect 23124 30580 23152 30892
rect 23293 30889 23305 30923
rect 23339 30920 23351 30923
rect 23566 30920 23572 30932
rect 23339 30892 23572 30920
rect 23339 30889 23351 30892
rect 23293 30883 23351 30889
rect 23566 30880 23572 30892
rect 23624 30880 23630 30932
rect 23658 30880 23664 30932
rect 23716 30880 23722 30932
rect 23198 30676 23204 30728
rect 23256 30676 23262 30728
rect 23477 30719 23535 30725
rect 23477 30685 23489 30719
rect 23523 30685 23535 30719
rect 23676 30716 23704 30880
rect 23845 30719 23903 30725
rect 23845 30716 23857 30719
rect 23676 30688 23857 30716
rect 23477 30679 23535 30685
rect 23845 30685 23857 30688
rect 23891 30685 23903 30719
rect 23845 30679 23903 30685
rect 23492 30648 23520 30679
rect 24026 30648 24032 30660
rect 23492 30620 24032 30648
rect 24026 30608 24032 30620
rect 24084 30608 24090 30660
rect 24213 30651 24271 30657
rect 24213 30617 24225 30651
rect 24259 30648 24271 30651
rect 24854 30648 24860 30660
rect 24259 30620 24860 30648
rect 24259 30617 24271 30620
rect 24213 30611 24271 30617
rect 24854 30608 24860 30620
rect 24912 30608 24918 30660
rect 25498 30580 25504 30592
rect 23124 30552 25504 30580
rect 25498 30540 25504 30552
rect 25556 30540 25562 30592
rect 1104 30490 24723 30512
rect 1104 30438 6814 30490
rect 6866 30438 6878 30490
rect 6930 30438 6942 30490
rect 6994 30438 7006 30490
rect 7058 30438 7070 30490
rect 7122 30438 12679 30490
rect 12731 30438 12743 30490
rect 12795 30438 12807 30490
rect 12859 30438 12871 30490
rect 12923 30438 12935 30490
rect 12987 30438 18544 30490
rect 18596 30438 18608 30490
rect 18660 30438 18672 30490
rect 18724 30438 18736 30490
rect 18788 30438 18800 30490
rect 18852 30438 24409 30490
rect 24461 30438 24473 30490
rect 24525 30438 24537 30490
rect 24589 30438 24601 30490
rect 24653 30438 24665 30490
rect 24717 30438 24723 30490
rect 1104 30416 24723 30438
rect 1688 30348 4380 30376
rect 1688 30249 1716 30348
rect 1673 30243 1731 30249
rect 1673 30209 1685 30243
rect 1719 30209 1731 30243
rect 1673 30203 1731 30209
rect 2590 30200 2596 30252
rect 2648 30200 2654 30252
rect 2710 30243 2768 30249
rect 2710 30240 2722 30243
rect 2700 30209 2722 30240
rect 2756 30209 2768 30243
rect 2700 30203 2768 30209
rect 1854 30132 1860 30184
rect 1912 30132 1918 30184
rect 2038 30132 2044 30184
rect 2096 30172 2102 30184
rect 2317 30175 2375 30181
rect 2317 30172 2329 30175
rect 2096 30144 2329 30172
rect 2096 30132 2102 30144
rect 2317 30141 2329 30144
rect 2363 30141 2375 30175
rect 2700 30172 2728 30203
rect 2317 30135 2375 30141
rect 2424 30144 2728 30172
rect 2222 30064 2228 30116
rect 2280 30104 2286 30116
rect 2424 30104 2452 30144
rect 2866 30132 2872 30184
rect 2924 30132 2930 30184
rect 3050 30132 3056 30184
rect 3108 30172 3114 30184
rect 3436 30172 3464 30348
rect 3510 30268 3516 30320
rect 3568 30268 3574 30320
rect 4352 30308 4380 30348
rect 4890 30336 4896 30388
rect 4948 30376 4954 30388
rect 4985 30379 5043 30385
rect 4985 30376 4997 30379
rect 4948 30348 4997 30376
rect 4948 30336 4954 30348
rect 4985 30345 4997 30348
rect 5031 30345 5043 30379
rect 4985 30339 5043 30345
rect 5534 30336 5540 30388
rect 5592 30376 5598 30388
rect 5902 30376 5908 30388
rect 5592 30348 5908 30376
rect 5592 30336 5598 30348
rect 5902 30336 5908 30348
rect 5960 30336 5966 30388
rect 6638 30336 6644 30388
rect 6696 30376 6702 30388
rect 13446 30376 13452 30388
rect 6696 30348 13452 30376
rect 6696 30336 6702 30348
rect 13446 30336 13452 30348
rect 13504 30336 13510 30388
rect 14093 30379 14151 30385
rect 14093 30345 14105 30379
rect 14139 30376 14151 30379
rect 15010 30376 15016 30388
rect 14139 30348 15016 30376
rect 14139 30345 14151 30348
rect 14093 30339 14151 30345
rect 14292 30320 14320 30348
rect 15010 30336 15016 30348
rect 15068 30336 15074 30388
rect 15102 30336 15108 30388
rect 15160 30376 15166 30388
rect 15197 30379 15255 30385
rect 15197 30376 15209 30379
rect 15160 30348 15209 30376
rect 15160 30336 15166 30348
rect 15197 30345 15209 30348
rect 15243 30376 15255 30379
rect 16850 30376 16856 30388
rect 15243 30348 16856 30376
rect 15243 30345 15255 30348
rect 15197 30339 15255 30345
rect 16850 30336 16856 30348
rect 16908 30336 16914 30388
rect 22741 30379 22799 30385
rect 22741 30345 22753 30379
rect 22787 30376 22799 30379
rect 23842 30376 23848 30388
rect 22787 30348 23848 30376
rect 22787 30345 22799 30348
rect 22741 30339 22799 30345
rect 23842 30336 23848 30348
rect 23900 30336 23906 30388
rect 10778 30308 10784 30320
rect 4352 30280 10784 30308
rect 10778 30268 10784 30280
rect 10836 30268 10842 30320
rect 10962 30268 10968 30320
rect 11020 30308 11026 30320
rect 11020 30280 12020 30308
rect 11020 30268 11026 30280
rect 4247 30253 4305 30259
rect 4247 30252 4259 30253
rect 4293 30252 4305 30253
rect 3697 30243 3755 30249
rect 3697 30209 3709 30243
rect 3743 30209 3755 30243
rect 3697 30203 3755 30209
rect 3108 30144 3464 30172
rect 3108 30132 3114 30144
rect 3712 30104 3740 30203
rect 4246 30200 4252 30252
rect 4304 30200 4310 30252
rect 4798 30200 4804 30252
rect 4856 30240 4862 30252
rect 5074 30240 5080 30252
rect 4856 30212 5080 30240
rect 4856 30200 4862 30212
rect 5074 30200 5080 30212
rect 5132 30200 5138 30252
rect 5350 30200 5356 30252
rect 5408 30200 5414 30252
rect 5902 30200 5908 30252
rect 5960 30200 5966 30252
rect 7650 30240 7656 30252
rect 7611 30212 7656 30240
rect 7650 30200 7656 30212
rect 7708 30200 7714 30252
rect 10042 30200 10048 30252
rect 10100 30200 10106 30252
rect 10226 30200 10232 30252
rect 10284 30240 10290 30252
rect 10319 30243 10377 30249
rect 10319 30240 10331 30243
rect 10284 30212 10331 30240
rect 10284 30200 10290 30212
rect 10319 30209 10331 30212
rect 10365 30240 10377 30243
rect 10365 30212 10732 30240
rect 10365 30209 10377 30212
rect 10319 30203 10377 30209
rect 3970 30132 3976 30184
rect 4028 30132 4034 30184
rect 5629 30175 5687 30181
rect 5629 30141 5641 30175
rect 5675 30172 5687 30175
rect 6822 30172 6828 30184
rect 5675 30144 6828 30172
rect 5675 30141 5687 30144
rect 5629 30135 5687 30141
rect 6822 30132 6828 30144
rect 6880 30132 6886 30184
rect 7374 30132 7380 30184
rect 7432 30132 7438 30184
rect 2280 30076 2452 30104
rect 3252 30076 3740 30104
rect 6089 30107 6147 30113
rect 2280 30064 2286 30076
rect 1302 29996 1308 30048
rect 1360 30036 1366 30048
rect 3252 30036 3280 30076
rect 6089 30073 6101 30107
rect 6135 30073 6147 30107
rect 10704 30104 10732 30212
rect 11514 30200 11520 30252
rect 11572 30240 11578 30252
rect 11882 30240 11888 30252
rect 11572 30212 11888 30240
rect 11572 30200 11578 30212
rect 11882 30200 11888 30212
rect 11940 30200 11946 30252
rect 11992 30240 12020 30280
rect 12143 30273 12201 30279
rect 12143 30240 12155 30273
rect 11992 30239 12155 30240
rect 12189 30239 12201 30273
rect 12434 30268 12440 30320
rect 12492 30308 12498 30320
rect 13170 30308 13176 30320
rect 12492 30280 13176 30308
rect 12492 30268 12498 30280
rect 13170 30268 13176 30280
rect 13228 30268 13234 30320
rect 13262 30268 13268 30320
rect 13320 30308 13326 30320
rect 13357 30311 13415 30317
rect 13357 30308 13369 30311
rect 13320 30280 13369 30308
rect 13320 30268 13326 30280
rect 13357 30277 13369 30280
rect 13403 30277 13415 30311
rect 13357 30271 13415 30277
rect 14274 30268 14280 30320
rect 14332 30268 14338 30320
rect 14458 30268 14464 30320
rect 14516 30268 14522 30320
rect 22278 30308 22284 30320
rect 14752 30280 15148 30308
rect 11992 30233 12201 30239
rect 14369 30243 14427 30249
rect 11992 30212 12186 30233
rect 14369 30209 14381 30243
rect 14415 30240 14427 30243
rect 14752 30240 14780 30280
rect 14415 30212 14780 30240
rect 14829 30243 14887 30249
rect 14415 30209 14427 30212
rect 14369 30203 14427 30209
rect 14829 30209 14841 30243
rect 14875 30240 14887 30243
rect 14918 30240 14924 30252
rect 14875 30212 14924 30240
rect 14875 30209 14887 30212
rect 14829 30203 14887 30209
rect 14918 30200 14924 30212
rect 14976 30200 14982 30252
rect 15120 30240 15148 30280
rect 16960 30280 22284 30308
rect 15378 30240 15384 30252
rect 15120 30212 15384 30240
rect 15378 30200 15384 30212
rect 15436 30200 15442 30252
rect 13814 30132 13820 30184
rect 13872 30172 13878 30184
rect 13872 30144 13938 30172
rect 13872 30132 13878 30144
rect 15930 30132 15936 30184
rect 15988 30172 15994 30184
rect 16960 30172 16988 30280
rect 22278 30268 22284 30280
rect 22336 30268 22342 30320
rect 22370 30268 22376 30320
rect 22428 30308 22434 30320
rect 22428 30280 23520 30308
rect 22428 30268 22434 30280
rect 21082 30200 21088 30252
rect 21140 30240 21146 30252
rect 21821 30243 21879 30249
rect 21821 30240 21833 30243
rect 21140 30212 21833 30240
rect 21140 30200 21146 30212
rect 21821 30209 21833 30212
rect 21867 30209 21879 30243
rect 21821 30203 21879 30209
rect 22186 30200 22192 30252
rect 22244 30200 22250 30252
rect 22830 30240 22836 30252
rect 22572 30212 22836 30240
rect 22476 30186 22534 30192
rect 15988 30144 16988 30172
rect 15988 30132 15994 30144
rect 17402 30132 17408 30184
rect 17460 30172 17466 30184
rect 17460 30144 22416 30172
rect 22476 30152 22488 30186
rect 22522 30183 22534 30186
rect 22572 30183 22600 30212
rect 22830 30200 22836 30212
rect 22888 30200 22894 30252
rect 23492 30249 23520 30280
rect 22925 30243 22983 30249
rect 22925 30209 22937 30243
rect 22971 30209 22983 30243
rect 22925 30203 22983 30209
rect 23201 30243 23259 30249
rect 23201 30209 23213 30243
rect 23247 30240 23259 30243
rect 23477 30243 23535 30249
rect 23247 30212 23336 30240
rect 23247 30209 23259 30212
rect 23201 30203 23259 30209
rect 22522 30155 22600 30183
rect 22522 30152 22534 30155
rect 22476 30146 22534 30152
rect 17460 30132 17466 30144
rect 10962 30104 10968 30116
rect 6089 30067 6147 30073
rect 8312 30076 9674 30104
rect 10704 30076 10968 30104
rect 1360 30008 3280 30036
rect 1360 29996 1366 30008
rect 3510 29996 3516 30048
rect 3568 30036 3574 30048
rect 3789 30039 3847 30045
rect 3789 30036 3801 30039
rect 3568 30008 3801 30036
rect 3568 29996 3574 30008
rect 3789 30005 3801 30008
rect 3835 30005 3847 30039
rect 3789 29999 3847 30005
rect 4062 29996 4068 30048
rect 4120 30036 4126 30048
rect 6104 30036 6132 30067
rect 4120 30008 6132 30036
rect 4120 29996 4126 30008
rect 6362 29996 6368 30048
rect 6420 30036 6426 30048
rect 8312 30036 8340 30076
rect 6420 30008 8340 30036
rect 6420 29996 6426 30008
rect 8386 29996 8392 30048
rect 8444 29996 8450 30048
rect 9646 30036 9674 30076
rect 10962 30064 10968 30076
rect 11020 30104 11026 30116
rect 11238 30104 11244 30116
rect 11020 30076 11244 30104
rect 11020 30064 11026 30076
rect 11238 30064 11244 30076
rect 11296 30064 11302 30116
rect 12897 30107 12955 30113
rect 12897 30073 12909 30107
rect 12943 30104 12955 30107
rect 13078 30104 13084 30116
rect 12943 30076 13084 30104
rect 12943 30073 12955 30076
rect 12897 30067 12955 30073
rect 13078 30064 13084 30076
rect 13136 30064 13142 30116
rect 22388 30104 22416 30144
rect 22940 30104 22968 30203
rect 23308 30113 23336 30212
rect 23477 30209 23489 30243
rect 23523 30209 23535 30243
rect 23477 30203 23535 30209
rect 23566 30200 23572 30252
rect 23624 30240 23630 30252
rect 23845 30243 23903 30249
rect 23845 30240 23857 30243
rect 23624 30212 23857 30240
rect 23624 30200 23630 30212
rect 23845 30209 23857 30212
rect 23891 30209 23903 30243
rect 23845 30203 23903 30209
rect 23937 30243 23995 30249
rect 23937 30209 23949 30243
rect 23983 30209 23995 30243
rect 23937 30203 23995 30209
rect 23952 30172 23980 30203
rect 23584 30144 23980 30172
rect 22388 30076 22968 30104
rect 23293 30107 23351 30113
rect 23293 30073 23305 30107
rect 23339 30073 23351 30107
rect 23293 30067 23351 30073
rect 10778 30036 10784 30048
rect 9646 30008 10784 30036
rect 10778 29996 10784 30008
rect 10836 29996 10842 30048
rect 11054 29996 11060 30048
rect 11112 29996 11118 30048
rect 11422 29996 11428 30048
rect 11480 30036 11486 30048
rect 12342 30036 12348 30048
rect 11480 30008 12348 30036
rect 11480 29996 11486 30008
rect 12342 29996 12348 30008
rect 12400 29996 12406 30048
rect 13446 29996 13452 30048
rect 13504 29996 13510 30048
rect 15381 30039 15439 30045
rect 15381 30005 15393 30039
rect 15427 30036 15439 30039
rect 16482 30036 16488 30048
rect 15427 30008 16488 30036
rect 15427 30005 15439 30008
rect 15381 29999 15439 30005
rect 16482 29996 16488 30008
rect 16540 29996 16546 30048
rect 16666 29996 16672 30048
rect 16724 30036 16730 30048
rect 20898 30036 20904 30048
rect 16724 30008 20904 30036
rect 16724 29996 16730 30008
rect 20898 29996 20904 30008
rect 20956 29996 20962 30048
rect 21913 30039 21971 30045
rect 21913 30005 21925 30039
rect 21959 30036 21971 30039
rect 22281 30039 22339 30045
rect 22281 30036 22293 30039
rect 21959 30008 22293 30036
rect 21959 30005 21971 30008
rect 21913 29999 21971 30005
rect 22281 30005 22293 30008
rect 22327 30005 22339 30039
rect 22281 29999 22339 30005
rect 22373 30039 22431 30045
rect 22373 30005 22385 30039
rect 22419 30036 22431 30039
rect 22922 30036 22928 30048
rect 22419 30008 22928 30036
rect 22419 30005 22431 30008
rect 22373 29999 22431 30005
rect 22922 29996 22928 30008
rect 22980 29996 22986 30048
rect 23017 30039 23075 30045
rect 23017 30005 23029 30039
rect 23063 30036 23075 30039
rect 23584 30036 23612 30144
rect 23063 30008 23612 30036
rect 23063 30005 23075 30008
rect 23017 29999 23075 30005
rect 23658 29996 23664 30048
rect 23716 29996 23722 30048
rect 24118 29996 24124 30048
rect 24176 29996 24182 30048
rect 1104 29946 24564 29968
rect 1104 29894 3882 29946
rect 3934 29894 3946 29946
rect 3998 29894 4010 29946
rect 4062 29894 4074 29946
rect 4126 29894 4138 29946
rect 4190 29894 9747 29946
rect 9799 29894 9811 29946
rect 9863 29894 9875 29946
rect 9927 29894 9939 29946
rect 9991 29894 10003 29946
rect 10055 29894 15612 29946
rect 15664 29894 15676 29946
rect 15728 29894 15740 29946
rect 15792 29894 15804 29946
rect 15856 29894 15868 29946
rect 15920 29894 21477 29946
rect 21529 29894 21541 29946
rect 21593 29894 21605 29946
rect 21657 29894 21669 29946
rect 21721 29894 21733 29946
rect 21785 29894 24564 29946
rect 1104 29872 24564 29894
rect 2866 29792 2872 29844
rect 2924 29792 2930 29844
rect 6362 29832 6368 29844
rect 4448 29804 6368 29832
rect 4448 29776 4476 29804
rect 6362 29792 6368 29804
rect 6420 29792 6426 29844
rect 9950 29792 9956 29844
rect 10008 29832 10014 29844
rect 10226 29832 10232 29844
rect 10008 29804 10232 29832
rect 10008 29792 10014 29804
rect 10226 29792 10232 29804
rect 10284 29792 10290 29844
rect 12526 29792 12532 29844
rect 12584 29832 12590 29844
rect 21450 29832 21456 29844
rect 12584 29804 21456 29832
rect 12584 29792 12590 29804
rect 21450 29792 21456 29804
rect 21508 29792 21514 29844
rect 22922 29792 22928 29844
rect 22980 29792 22986 29844
rect 23201 29835 23259 29841
rect 23201 29801 23213 29835
rect 23247 29832 23259 29835
rect 23566 29832 23572 29844
rect 23247 29804 23572 29832
rect 23247 29801 23259 29804
rect 23201 29795 23259 29801
rect 23566 29792 23572 29804
rect 23624 29792 23630 29844
rect 23658 29792 23664 29844
rect 23716 29792 23722 29844
rect 2682 29724 2688 29776
rect 2740 29764 2746 29776
rect 2740 29724 2774 29764
rect 4430 29724 4436 29776
rect 4488 29724 4494 29776
rect 5905 29767 5963 29773
rect 5905 29733 5917 29767
rect 5951 29733 5963 29767
rect 5905 29727 5963 29733
rect 1394 29656 1400 29708
rect 1452 29696 1458 29708
rect 1857 29699 1915 29705
rect 1857 29696 1869 29699
rect 1452 29668 1869 29696
rect 1452 29656 1458 29668
rect 1857 29665 1869 29668
rect 1903 29665 1915 29699
rect 2746 29696 2774 29724
rect 3789 29699 3847 29705
rect 3789 29696 3801 29699
rect 2746 29668 3801 29696
rect 1857 29659 1915 29665
rect 3789 29665 3801 29668
rect 3835 29665 3847 29699
rect 5920 29696 5948 29727
rect 11790 29724 11796 29776
rect 11848 29764 11854 29776
rect 14918 29764 14924 29776
rect 11848 29736 14924 29764
rect 11848 29724 11854 29736
rect 14918 29724 14924 29736
rect 14976 29764 14982 29776
rect 15746 29764 15752 29776
rect 14976 29736 15752 29764
rect 14976 29724 14982 29736
rect 15746 29724 15752 29736
rect 15804 29724 15810 29776
rect 16758 29724 16764 29776
rect 16816 29724 16822 29776
rect 19521 29767 19579 29773
rect 19521 29733 19533 29767
rect 19567 29764 19579 29767
rect 20714 29764 20720 29776
rect 19567 29736 20720 29764
rect 19567 29733 19579 29736
rect 19521 29727 19579 29733
rect 20714 29724 20720 29736
rect 20772 29724 20778 29776
rect 5920 29668 6302 29696
rect 3789 29659 3847 29665
rect 11054 29656 11060 29708
rect 11112 29656 11118 29708
rect 11606 29656 11612 29708
rect 11664 29696 11670 29708
rect 12526 29696 12532 29708
rect 11664 29668 12532 29696
rect 11664 29656 11670 29668
rect 12526 29656 12532 29668
rect 12584 29656 12590 29708
rect 16666 29656 16672 29708
rect 16724 29656 16730 29708
rect 22370 29696 22376 29708
rect 19306 29668 22376 29696
rect 750 29588 756 29640
rect 808 29628 814 29640
rect 1489 29631 1547 29637
rect 1489 29628 1501 29631
rect 808 29600 1501 29628
rect 808 29588 814 29600
rect 1489 29597 1501 29600
rect 1535 29597 1547 29631
rect 1489 29591 1547 29597
rect 2130 29588 2136 29640
rect 2188 29588 2194 29640
rect 3237 29631 3295 29637
rect 3237 29597 3249 29631
rect 3283 29597 3295 29631
rect 4065 29631 4123 29637
rect 4065 29628 4077 29631
rect 3237 29591 3295 29597
rect 3528 29600 4077 29628
rect 1302 29520 1308 29572
rect 1360 29560 1366 29572
rect 3252 29560 3280 29591
rect 3528 29560 3556 29600
rect 4065 29597 4077 29600
rect 4111 29597 4123 29631
rect 4065 29591 4123 29597
rect 4893 29631 4951 29637
rect 4893 29597 4905 29631
rect 4939 29597 4951 29631
rect 7193 29631 7251 29637
rect 7193 29628 7205 29631
rect 4893 29591 4951 29597
rect 5151 29601 5209 29607
rect 1360 29532 3280 29560
rect 3344 29532 3556 29560
rect 1360 29520 1366 29532
rect 1581 29495 1639 29501
rect 1581 29461 1593 29495
rect 1627 29492 1639 29495
rect 2406 29492 2412 29504
rect 1627 29464 2412 29492
rect 1627 29461 1639 29464
rect 1581 29455 1639 29461
rect 2406 29452 2412 29464
rect 2464 29452 2470 29504
rect 2498 29452 2504 29504
rect 2556 29492 2562 29504
rect 3344 29492 3372 29532
rect 3528 29504 3556 29532
rect 2556 29464 3372 29492
rect 2556 29452 2562 29464
rect 3418 29452 3424 29504
rect 3476 29452 3482 29504
rect 3510 29452 3516 29504
rect 3568 29452 3574 29504
rect 4908 29492 4936 29591
rect 5151 29567 5163 29601
rect 5197 29598 5209 29601
rect 5644 29600 7205 29628
rect 5197 29572 5212 29598
rect 5644 29572 5672 29600
rect 7193 29597 7205 29600
rect 7239 29597 7251 29631
rect 7193 29591 7251 29597
rect 7374 29588 7380 29640
rect 7432 29628 7438 29640
rect 8754 29628 8760 29640
rect 7432 29600 8760 29628
rect 7432 29588 7438 29600
rect 8754 29588 8760 29600
rect 8812 29628 8818 29640
rect 8941 29631 8999 29637
rect 8941 29628 8953 29631
rect 8812 29600 8953 29628
rect 8812 29588 8818 29600
rect 8941 29597 8953 29600
rect 8987 29597 8999 29631
rect 9214 29628 9220 29640
rect 9175 29600 9220 29628
rect 8941 29591 8999 29597
rect 9214 29588 9220 29600
rect 9272 29588 9278 29640
rect 10594 29588 10600 29640
rect 10652 29588 10658 29640
rect 10686 29588 10692 29640
rect 10744 29628 10750 29640
rect 10781 29631 10839 29637
rect 10781 29628 10793 29631
rect 10744 29600 10793 29628
rect 10744 29588 10750 29600
rect 10781 29597 10793 29600
rect 10827 29597 10839 29631
rect 10781 29591 10839 29597
rect 10873 29631 10931 29637
rect 10873 29597 10885 29631
rect 10919 29628 10931 29631
rect 11698 29628 11704 29640
rect 10919 29600 11704 29628
rect 10919 29597 10931 29600
rect 10873 29591 10931 29597
rect 11698 29588 11704 29600
rect 11756 29588 11762 29640
rect 12544 29628 12572 29656
rect 15654 29628 15660 29640
rect 12544 29600 15660 29628
rect 15654 29588 15660 29600
rect 15712 29628 15718 29640
rect 15749 29631 15807 29637
rect 15749 29628 15761 29631
rect 15712 29600 15761 29628
rect 15712 29588 15718 29600
rect 15749 29597 15761 29600
rect 15795 29597 15807 29631
rect 15749 29591 15807 29597
rect 16023 29631 16081 29637
rect 16023 29597 16035 29631
rect 16069 29624 16081 29631
rect 16684 29628 16712 29656
rect 17129 29631 17187 29637
rect 17129 29628 17141 29631
rect 16069 29597 16160 29624
rect 16684 29600 17141 29628
rect 16023 29596 16160 29597
rect 16023 29591 16081 29596
rect 5151 29561 5172 29567
rect 5166 29520 5172 29561
rect 5224 29520 5230 29572
rect 5626 29520 5632 29572
rect 5684 29520 5690 29572
rect 6086 29520 6092 29572
rect 6144 29520 6150 29572
rect 6270 29520 6276 29572
rect 6328 29560 6334 29572
rect 6457 29563 6515 29569
rect 6457 29560 6469 29563
rect 6328 29532 6469 29560
rect 6328 29520 6334 29532
rect 6457 29529 6469 29532
rect 6503 29529 6515 29563
rect 6457 29523 6515 29529
rect 6546 29520 6552 29572
rect 6604 29560 6610 29572
rect 6733 29563 6791 29569
rect 6733 29560 6745 29563
rect 6604 29532 6745 29560
rect 6604 29520 6610 29532
rect 6733 29529 6745 29532
rect 6779 29529 6791 29563
rect 6733 29523 6791 29529
rect 6822 29520 6828 29572
rect 6880 29520 6886 29572
rect 7282 29560 7288 29572
rect 6932 29532 7288 29560
rect 6104 29492 6132 29520
rect 4908 29464 6132 29492
rect 6362 29452 6368 29504
rect 6420 29492 6426 29504
rect 6932 29492 6960 29532
rect 7282 29520 7288 29532
rect 7340 29560 7346 29572
rect 7561 29563 7619 29569
rect 7561 29560 7573 29563
rect 7340 29532 7573 29560
rect 7340 29520 7346 29532
rect 7561 29529 7573 29532
rect 7607 29529 7619 29563
rect 10226 29560 10232 29572
rect 7561 29523 7619 29529
rect 7760 29532 10232 29560
rect 7760 29501 7788 29532
rect 10226 29520 10232 29532
rect 10284 29520 10290 29572
rect 10505 29563 10563 29569
rect 10505 29529 10517 29563
rect 10551 29529 10563 29563
rect 10612 29560 10640 29588
rect 11054 29560 11060 29572
rect 10612 29532 11060 29560
rect 10505 29523 10563 29529
rect 6420 29464 6960 29492
rect 7745 29495 7803 29501
rect 6420 29452 6426 29464
rect 7745 29461 7757 29495
rect 7791 29461 7803 29495
rect 7745 29455 7803 29461
rect 8938 29452 8944 29504
rect 8996 29492 9002 29504
rect 9953 29495 10011 29501
rect 9953 29492 9965 29495
rect 8996 29464 9965 29492
rect 8996 29452 9002 29464
rect 9953 29461 9965 29464
rect 9999 29461 10011 29495
rect 10520 29492 10548 29523
rect 11054 29520 11060 29532
rect 11112 29520 11118 29572
rect 11238 29520 11244 29572
rect 11296 29520 11302 29572
rect 13262 29560 13268 29572
rect 11440 29532 13268 29560
rect 11440 29492 11468 29532
rect 13262 29520 13268 29532
rect 13320 29520 13326 29572
rect 15562 29520 15568 29572
rect 15620 29520 15626 29572
rect 10520 29464 11468 29492
rect 9953 29455 10011 29461
rect 11514 29452 11520 29504
rect 11572 29492 11578 29504
rect 11609 29495 11667 29501
rect 11609 29492 11621 29495
rect 11572 29464 11621 29492
rect 11572 29452 11578 29464
rect 11609 29461 11621 29464
rect 11655 29461 11667 29495
rect 11609 29455 11667 29461
rect 11790 29452 11796 29504
rect 11848 29452 11854 29504
rect 12066 29452 12072 29504
rect 12124 29492 12130 29504
rect 15470 29492 15476 29504
rect 12124 29464 15476 29492
rect 12124 29452 12130 29464
rect 15470 29452 15476 29464
rect 15528 29452 15534 29504
rect 15580 29492 15608 29520
rect 16132 29492 16160 29596
rect 17129 29597 17141 29600
rect 17175 29597 17187 29631
rect 17402 29628 17408 29640
rect 17363 29600 17408 29628
rect 17129 29591 17187 29597
rect 17402 29588 17408 29600
rect 17460 29588 17466 29640
rect 18874 29628 18880 29640
rect 17604 29600 18880 29628
rect 16758 29520 16764 29572
rect 16816 29560 16822 29572
rect 17310 29560 17316 29572
rect 16816 29532 17316 29560
rect 16816 29520 16822 29532
rect 17310 29520 17316 29532
rect 17368 29520 17374 29572
rect 17604 29492 17632 29600
rect 18874 29588 18880 29600
rect 18932 29628 18938 29640
rect 19306 29628 19334 29668
rect 22370 29656 22376 29668
rect 22428 29656 22434 29708
rect 18932 29600 19334 29628
rect 19705 29631 19763 29637
rect 18932 29588 18938 29600
rect 19705 29597 19717 29631
rect 19751 29597 19763 29631
rect 19705 29591 19763 29597
rect 17678 29520 17684 29572
rect 17736 29560 17742 29572
rect 19242 29560 19248 29572
rect 17736 29532 19248 29560
rect 17736 29520 17742 29532
rect 19242 29520 19248 29532
rect 19300 29560 19306 29572
rect 19720 29560 19748 29591
rect 20346 29588 20352 29640
rect 20404 29628 20410 29640
rect 20625 29631 20683 29637
rect 20625 29628 20637 29631
rect 20404 29600 20637 29628
rect 20404 29588 20410 29600
rect 20625 29597 20637 29600
rect 20671 29597 20683 29631
rect 20625 29591 20683 29597
rect 19300 29532 19748 29560
rect 19300 29520 19306 29532
rect 20070 29520 20076 29572
rect 20128 29560 20134 29572
rect 21358 29560 21364 29572
rect 20128 29532 21364 29560
rect 20128 29520 20134 29532
rect 21358 29520 21364 29532
rect 21416 29520 21422 29572
rect 22940 29560 22968 29792
rect 23676 29696 23704 29792
rect 23676 29668 23980 29696
rect 23106 29588 23112 29640
rect 23164 29628 23170 29640
rect 23385 29631 23443 29637
rect 23385 29628 23397 29631
rect 23164 29600 23397 29628
rect 23164 29588 23170 29600
rect 23385 29597 23397 29600
rect 23431 29597 23443 29631
rect 23385 29591 23443 29597
rect 23474 29588 23480 29640
rect 23532 29628 23538 29640
rect 23952 29637 23980 29668
rect 23845 29631 23903 29637
rect 23845 29628 23857 29631
rect 23532 29600 23857 29628
rect 23532 29588 23538 29600
rect 23845 29597 23857 29600
rect 23891 29597 23903 29631
rect 23845 29591 23903 29597
rect 23937 29631 23995 29637
rect 23937 29597 23949 29631
rect 23983 29597 23995 29631
rect 23937 29591 23995 29597
rect 23750 29560 23756 29572
rect 22940 29532 23756 29560
rect 23750 29520 23756 29532
rect 23808 29520 23814 29572
rect 15580 29464 17632 29492
rect 17862 29452 17868 29504
rect 17920 29492 17926 29504
rect 18141 29495 18199 29501
rect 18141 29492 18153 29495
rect 17920 29464 18153 29492
rect 17920 29452 17926 29464
rect 18141 29461 18153 29464
rect 18187 29461 18199 29495
rect 18141 29455 18199 29461
rect 20441 29495 20499 29501
rect 20441 29461 20453 29495
rect 20487 29492 20499 29495
rect 21082 29492 21088 29504
rect 20487 29464 21088 29492
rect 20487 29461 20499 29464
rect 20441 29455 20499 29461
rect 21082 29452 21088 29464
rect 21140 29452 21146 29504
rect 23658 29452 23664 29504
rect 23716 29452 23722 29504
rect 24121 29495 24179 29501
rect 24121 29461 24133 29495
rect 24167 29492 24179 29495
rect 24854 29492 24860 29504
rect 24167 29464 24860 29492
rect 24167 29461 24179 29464
rect 24121 29455 24179 29461
rect 24854 29452 24860 29464
rect 24912 29452 24918 29504
rect 1104 29402 24723 29424
rect 1104 29350 6814 29402
rect 6866 29350 6878 29402
rect 6930 29350 6942 29402
rect 6994 29350 7006 29402
rect 7058 29350 7070 29402
rect 7122 29350 12679 29402
rect 12731 29350 12743 29402
rect 12795 29350 12807 29402
rect 12859 29350 12871 29402
rect 12923 29350 12935 29402
rect 12987 29350 18544 29402
rect 18596 29350 18608 29402
rect 18660 29350 18672 29402
rect 18724 29350 18736 29402
rect 18788 29350 18800 29402
rect 18852 29350 24409 29402
rect 24461 29350 24473 29402
rect 24525 29350 24537 29402
rect 24589 29350 24601 29402
rect 24653 29350 24665 29402
rect 24717 29350 24723 29402
rect 1104 29328 24723 29350
rect 1578 29248 1584 29300
rect 1636 29288 1642 29300
rect 3418 29288 3424 29300
rect 1636 29260 3424 29288
rect 1636 29248 1642 29260
rect 3418 29248 3424 29260
rect 3476 29288 3482 29300
rect 3476 29260 7236 29288
rect 3476 29248 3482 29260
rect 7208 29232 7236 29260
rect 7282 29248 7288 29300
rect 7340 29288 7346 29300
rect 7377 29291 7435 29297
rect 7377 29288 7389 29291
rect 7340 29260 7389 29288
rect 7340 29248 7346 29260
rect 7377 29257 7389 29260
rect 7423 29257 7435 29291
rect 7377 29251 7435 29257
rect 10137 29291 10195 29297
rect 10137 29257 10149 29291
rect 10183 29257 10195 29291
rect 10137 29251 10195 29257
rect 1302 29180 1308 29232
rect 1360 29220 1366 29232
rect 2682 29220 2688 29232
rect 1360 29192 2688 29220
rect 1360 29180 1366 29192
rect 2682 29180 2688 29192
rect 2740 29180 2746 29232
rect 4798 29220 4804 29232
rect 3068 29192 4804 29220
rect 2406 29112 2412 29164
rect 2464 29112 2470 29164
rect 1394 29044 1400 29096
rect 1452 29044 1458 29096
rect 1670 29044 1676 29096
rect 1728 29084 1734 29096
rect 3068 29084 3096 29192
rect 4798 29180 4804 29192
rect 4856 29180 4862 29232
rect 5258 29180 5264 29232
rect 5316 29220 5322 29232
rect 5316 29192 7144 29220
rect 5316 29180 5322 29192
rect 3142 29112 3148 29164
rect 3200 29152 3206 29164
rect 3421 29155 3479 29161
rect 3421 29152 3433 29155
rect 3200 29124 3433 29152
rect 3200 29112 3206 29124
rect 3421 29121 3433 29124
rect 3467 29121 3479 29155
rect 3421 29115 3479 29121
rect 3695 29155 3753 29161
rect 3695 29121 3707 29155
rect 3741 29152 3753 29155
rect 5276 29152 5304 29180
rect 3741 29124 5304 29152
rect 3741 29121 3753 29124
rect 3695 29115 3753 29121
rect 6086 29112 6092 29164
rect 6144 29112 6150 29164
rect 6178 29112 6184 29164
rect 6236 29152 6242 29164
rect 6607 29155 6665 29161
rect 6607 29152 6619 29155
rect 6236 29124 6619 29152
rect 6236 29112 6242 29124
rect 6607 29121 6619 29124
rect 6653 29121 6665 29155
rect 7116 29152 7144 29192
rect 7190 29180 7196 29232
rect 7248 29180 7254 29232
rect 10152 29220 10180 29251
rect 10226 29248 10232 29300
rect 10284 29288 10290 29300
rect 16666 29288 16672 29300
rect 10284 29260 16672 29288
rect 10284 29248 10290 29260
rect 16666 29248 16672 29260
rect 16724 29248 16730 29300
rect 17678 29288 17684 29300
rect 16776 29260 17684 29288
rect 14737 29223 14795 29229
rect 10152 29192 10640 29220
rect 8110 29152 8116 29164
rect 7116 29124 8116 29152
rect 6607 29115 6665 29121
rect 8110 29112 8116 29124
rect 8168 29112 8174 29164
rect 8662 29112 8668 29164
rect 8720 29112 8726 29164
rect 8938 29112 8944 29164
rect 8996 29112 9002 29164
rect 10612 29161 10640 29192
rect 14737 29189 14749 29223
rect 14783 29220 14795 29223
rect 15378 29220 15384 29232
rect 14783 29192 15384 29220
rect 14783 29189 14795 29192
rect 14737 29183 14795 29189
rect 15378 29180 15384 29192
rect 15436 29220 15442 29232
rect 16776 29220 16804 29260
rect 17678 29248 17684 29260
rect 17736 29248 17742 29300
rect 17954 29248 17960 29300
rect 18012 29288 18018 29300
rect 18012 29260 19012 29288
rect 18012 29248 18018 29260
rect 15436 29192 16804 29220
rect 15436 29180 15442 29192
rect 9585 29155 9643 29161
rect 9585 29121 9597 29155
rect 9631 29152 9643 29155
rect 10045 29155 10103 29161
rect 10045 29152 10057 29155
rect 9631 29124 10057 29152
rect 9631 29121 9643 29124
rect 9585 29115 9643 29121
rect 10045 29121 10057 29124
rect 10091 29121 10103 29155
rect 10045 29115 10103 29121
rect 10321 29155 10379 29161
rect 10321 29121 10333 29155
rect 10367 29121 10379 29155
rect 10321 29115 10379 29121
rect 10413 29155 10471 29161
rect 10413 29121 10425 29155
rect 10459 29121 10471 29155
rect 10413 29115 10471 29121
rect 10597 29155 10655 29161
rect 10597 29121 10609 29155
rect 10643 29121 10655 29155
rect 10597 29115 10655 29121
rect 10689 29155 10747 29161
rect 10689 29121 10701 29155
rect 10735 29121 10747 29155
rect 10689 29115 10747 29121
rect 1728 29056 3096 29084
rect 1728 29044 1734 29056
rect 4246 29044 4252 29096
rect 4304 29084 4310 29096
rect 4430 29084 4436 29096
rect 4304 29056 4436 29084
rect 4304 29044 4310 29056
rect 4430 29044 4436 29056
rect 4488 29044 4494 29096
rect 6104 29084 6132 29112
rect 6270 29084 6276 29096
rect 6104 29056 6276 29084
rect 6270 29044 6276 29056
rect 6328 29084 6334 29096
rect 6365 29087 6423 29093
rect 6365 29084 6377 29087
rect 6328 29056 6377 29084
rect 6328 29044 6334 29056
rect 6365 29053 6377 29056
rect 6411 29053 6423 29087
rect 6365 29047 6423 29053
rect 7466 29044 7472 29096
rect 7524 29084 7530 29096
rect 7745 29087 7803 29093
rect 7745 29084 7757 29087
rect 7524 29056 7757 29084
rect 7524 29044 7530 29056
rect 7745 29053 7757 29056
rect 7791 29053 7803 29087
rect 7745 29047 7803 29053
rect 7929 29087 7987 29093
rect 7929 29053 7941 29087
rect 7975 29084 7987 29087
rect 8018 29084 8024 29096
rect 7975 29056 8024 29084
rect 7975 29053 7987 29056
rect 7929 29047 7987 29053
rect 8018 29044 8024 29056
rect 8076 29044 8082 29096
rect 8386 29044 8392 29096
rect 8444 29044 8450 29096
rect 8782 29087 8840 29093
rect 8782 29084 8794 29087
rect 8496 29056 8794 29084
rect 2222 28976 2228 29028
rect 2280 29016 2286 29028
rect 2593 29019 2651 29025
rect 2593 29016 2605 29019
rect 2280 28988 2605 29016
rect 2280 28976 2286 28988
rect 2593 28985 2605 28988
rect 2639 29016 2651 29019
rect 2682 29016 2688 29028
rect 2639 28988 2688 29016
rect 2639 28985 2651 28988
rect 2593 28979 2651 28985
rect 2682 28976 2688 28988
rect 2740 28976 2746 29028
rect 7190 28976 7196 29028
rect 7248 29016 7254 29028
rect 8496 29016 8524 29056
rect 8782 29053 8794 29056
rect 8828 29053 8840 29087
rect 8782 29047 8840 29053
rect 10134 29044 10140 29096
rect 10192 29084 10198 29096
rect 10336 29084 10364 29115
rect 10192 29056 10364 29084
rect 10428 29084 10456 29115
rect 10502 29084 10508 29096
rect 10428 29056 10508 29084
rect 10192 29044 10198 29056
rect 10502 29044 10508 29056
rect 10560 29044 10566 29096
rect 7248 28988 8524 29016
rect 9861 29019 9919 29025
rect 7248 28976 7254 28988
rect 9861 28985 9873 29019
rect 9907 29016 9919 29019
rect 10704 29016 10732 29115
rect 10778 29112 10784 29164
rect 10836 29152 10842 29164
rect 12897 29155 12955 29161
rect 12897 29152 12909 29155
rect 10836 29124 12909 29152
rect 10836 29112 10842 29124
rect 12897 29121 12909 29124
rect 12943 29121 12955 29155
rect 12897 29115 12955 29121
rect 16485 29158 16543 29161
rect 16485 29155 16618 29158
rect 16485 29121 16497 29155
rect 16531 29152 16618 29155
rect 16531 29130 16804 29152
rect 16531 29121 16543 29130
rect 16590 29124 16804 29130
rect 16485 29115 16543 29121
rect 9907 28988 10732 29016
rect 12912 29016 12940 29115
rect 13078 29044 13084 29096
rect 13136 29044 13142 29096
rect 13814 29044 13820 29096
rect 13872 29044 13878 29096
rect 13906 29044 13912 29096
rect 13964 29093 13970 29096
rect 13964 29087 13992 29093
rect 13980 29053 13992 29087
rect 13964 29047 13992 29053
rect 13964 29044 13970 29047
rect 14090 29044 14096 29096
rect 14148 29044 14154 29096
rect 14274 29044 14280 29096
rect 14332 29084 14338 29096
rect 14332 29056 16066 29084
rect 14332 29044 14338 29056
rect 12912 28988 13492 29016
rect 9907 28985 9919 28988
rect 9861 28979 9919 28985
rect 3694 28908 3700 28960
rect 3752 28948 3758 28960
rect 4154 28948 4160 28960
rect 3752 28920 4160 28948
rect 3752 28908 3758 28920
rect 4154 28908 4160 28920
rect 4212 28908 4218 28960
rect 4430 28908 4436 28960
rect 4488 28908 4494 28960
rect 5258 28908 5264 28960
rect 5316 28948 5322 28960
rect 7834 28948 7840 28960
rect 5316 28920 7840 28948
rect 5316 28908 5322 28920
rect 7834 28908 7840 28920
rect 7892 28948 7898 28960
rect 8662 28948 8668 28960
rect 7892 28920 8668 28948
rect 7892 28908 7898 28920
rect 8662 28908 8668 28920
rect 8720 28908 8726 28960
rect 9490 28908 9496 28960
rect 9548 28948 9554 28960
rect 10042 28948 10048 28960
rect 9548 28920 10048 28948
rect 9548 28908 9554 28920
rect 10042 28908 10048 28920
rect 10100 28908 10106 28960
rect 10502 28908 10508 28960
rect 10560 28908 10566 28960
rect 10778 28908 10784 28960
rect 10836 28908 10842 28960
rect 11054 28908 11060 28960
rect 11112 28948 11118 28960
rect 11422 28948 11428 28960
rect 11112 28920 11428 28948
rect 11112 28908 11118 28920
rect 11422 28908 11428 28920
rect 11480 28908 11486 28960
rect 13464 28948 13492 28988
rect 13538 28976 13544 29028
rect 13596 28976 13602 29028
rect 15930 29016 15936 29028
rect 14476 28988 15936 29016
rect 14476 28948 14504 28988
rect 15930 28976 15936 28988
rect 15988 28976 15994 29028
rect 16038 29016 16066 29056
rect 16666 29044 16672 29096
rect 16724 29044 16730 29096
rect 16776 29016 16804 29124
rect 16850 29112 16856 29164
rect 16908 29112 16914 29164
rect 17678 29112 17684 29164
rect 17736 29161 17742 29164
rect 17736 29155 17764 29161
rect 17752 29121 17764 29155
rect 17736 29115 17764 29121
rect 17736 29112 17742 29115
rect 17862 29112 17868 29164
rect 17920 29112 17926 29164
rect 18984 29161 19012 29260
rect 20346 29248 20352 29300
rect 20404 29248 20410 29300
rect 20901 29291 20959 29297
rect 20901 29288 20913 29291
rect 20548 29260 20913 29288
rect 19242 29229 19248 29232
rect 19236 29220 19248 29229
rect 19203 29192 19248 29220
rect 19236 29183 19248 29192
rect 19242 29180 19248 29183
rect 19300 29180 19306 29232
rect 18969 29155 19027 29161
rect 18969 29121 18981 29155
rect 19015 29121 19027 29155
rect 18969 29115 19027 29121
rect 20346 29112 20352 29164
rect 20404 29152 20410 29164
rect 20441 29155 20499 29161
rect 20441 29152 20453 29155
rect 20404 29124 20453 29152
rect 20404 29112 20410 29124
rect 20441 29121 20453 29124
rect 20487 29121 20499 29155
rect 20441 29115 20499 29121
rect 17310 29044 17316 29096
rect 17368 29044 17374 29096
rect 20548 29093 20576 29260
rect 20901 29257 20913 29260
rect 20947 29257 20959 29291
rect 20901 29251 20959 29257
rect 21082 29248 21088 29300
rect 21140 29248 21146 29300
rect 22278 29248 22284 29300
rect 22336 29288 22342 29300
rect 22922 29288 22928 29300
rect 22336 29260 22928 29288
rect 22336 29248 22342 29260
rect 22922 29248 22928 29260
rect 22980 29288 22986 29300
rect 23106 29288 23112 29300
rect 22980 29260 23112 29288
rect 22980 29248 22986 29260
rect 23106 29248 23112 29260
rect 23164 29248 23170 29300
rect 23474 29248 23480 29300
rect 23532 29248 23538 29300
rect 23658 29248 23664 29300
rect 23716 29248 23722 29300
rect 20714 29180 20720 29232
rect 20772 29220 20778 29232
rect 21100 29220 21128 29248
rect 20772 29192 20852 29220
rect 21100 29192 21312 29220
rect 20772 29180 20778 29192
rect 20824 29159 20852 29192
rect 20809 29153 20867 29159
rect 20809 29119 20821 29153
rect 20855 29119 20867 29153
rect 20809 29113 20867 29119
rect 21082 29112 21088 29164
rect 21140 29112 21146 29164
rect 21284 29161 21312 29192
rect 21450 29180 21456 29232
rect 21508 29220 21514 29232
rect 23676 29220 23704 29248
rect 23845 29223 23903 29229
rect 23845 29220 23857 29223
rect 21508 29192 23520 29220
rect 23676 29192 23857 29220
rect 21508 29180 21514 29192
rect 21269 29155 21327 29161
rect 21269 29121 21281 29155
rect 21315 29121 21327 29155
rect 21269 29115 21327 29121
rect 21358 29112 21364 29164
rect 21416 29152 21422 29164
rect 23385 29155 23443 29161
rect 23385 29152 23397 29155
rect 21416 29124 23397 29152
rect 21416 29112 21422 29124
rect 23385 29121 23397 29124
rect 23431 29121 23443 29155
rect 23492 29152 23520 29192
rect 23845 29189 23857 29192
rect 23891 29189 23903 29223
rect 23845 29183 23903 29189
rect 23661 29155 23719 29161
rect 23661 29152 23673 29155
rect 23492 29124 23673 29152
rect 23385 29115 23443 29121
rect 23661 29121 23673 29124
rect 23707 29121 23719 29155
rect 23661 29115 23719 29121
rect 17589 29087 17647 29093
rect 17589 29084 17601 29087
rect 17418 29056 17601 29084
rect 17418 29016 17446 29056
rect 17589 29053 17601 29056
rect 17635 29053 17647 29087
rect 17589 29047 17647 29053
rect 20533 29087 20591 29093
rect 20533 29053 20545 29087
rect 20579 29053 20591 29087
rect 20533 29047 20591 29053
rect 20717 29087 20775 29093
rect 20717 29053 20729 29087
rect 20763 29053 20775 29087
rect 21177 29087 21235 29093
rect 21177 29084 21189 29087
rect 21008 29076 21189 29084
rect 20717 29047 20775 29053
rect 20916 29056 21189 29076
rect 20916 29048 21036 29056
rect 21177 29053 21189 29056
rect 21223 29053 21235 29087
rect 16038 28988 16436 29016
rect 16776 28988 17446 29016
rect 18509 29019 18567 29025
rect 13464 28920 14504 28948
rect 14550 28908 14556 28960
rect 14608 28948 14614 28960
rect 16206 28948 16212 28960
rect 14608 28920 16212 28948
rect 14608 28908 14614 28920
rect 16206 28908 16212 28920
rect 16264 28908 16270 28960
rect 16408 28948 16436 28988
rect 18509 28985 18521 29019
rect 18555 29016 18567 29019
rect 18966 29016 18972 29028
rect 18555 28988 18972 29016
rect 18555 28985 18567 28988
rect 18509 28979 18567 28985
rect 18966 28976 18972 28988
rect 19024 28976 19030 29028
rect 20732 29016 20760 29047
rect 20916 29016 20944 29048
rect 21177 29047 21235 29053
rect 21910 29016 21916 29028
rect 20732 28988 20944 29016
rect 21008 28988 21916 29016
rect 17034 28948 17040 28960
rect 16408 28920 17040 28948
rect 17034 28908 17040 28920
rect 17092 28908 17098 28960
rect 20625 28951 20683 28957
rect 20625 28917 20637 28951
rect 20671 28948 20683 28951
rect 21008 28948 21036 28988
rect 21910 28976 21916 28988
rect 21968 28976 21974 29028
rect 23198 28976 23204 29028
rect 23256 28976 23262 29028
rect 24118 28976 24124 29028
rect 24176 28976 24182 29028
rect 20671 28920 21036 28948
rect 20671 28917 20683 28920
rect 20625 28911 20683 28917
rect 1104 28858 24564 28880
rect 1104 28806 3882 28858
rect 3934 28806 3946 28858
rect 3998 28806 4010 28858
rect 4062 28806 4074 28858
rect 4126 28806 4138 28858
rect 4190 28806 9747 28858
rect 9799 28806 9811 28858
rect 9863 28806 9875 28858
rect 9927 28806 9939 28858
rect 9991 28806 10003 28858
rect 10055 28806 15612 28858
rect 15664 28806 15676 28858
rect 15728 28806 15740 28858
rect 15792 28806 15804 28858
rect 15856 28806 15868 28858
rect 15920 28806 21477 28858
rect 21529 28806 21541 28858
rect 21593 28806 21605 28858
rect 21657 28806 21669 28858
rect 21721 28806 21733 28858
rect 21785 28806 24564 28858
rect 1104 28784 24564 28806
rect 3142 28744 3148 28756
rect 2332 28716 3148 28744
rect 2332 28617 2360 28716
rect 3142 28704 3148 28716
rect 3200 28704 3206 28756
rect 8754 28704 8760 28756
rect 8812 28744 8818 28756
rect 10597 28747 10655 28753
rect 8812 28716 10548 28744
rect 8812 28704 8818 28716
rect 3329 28679 3387 28685
rect 3329 28645 3341 28679
rect 3375 28676 3387 28679
rect 3375 28648 3832 28676
rect 3375 28645 3387 28648
rect 3329 28639 3387 28645
rect 2317 28611 2375 28617
rect 2317 28577 2329 28611
rect 2363 28577 2375 28611
rect 3804 28594 3832 28648
rect 9490 28608 9496 28620
rect 2317 28571 2375 28577
rect 8864 28580 9496 28608
rect 1210 28500 1216 28552
rect 1268 28540 1274 28552
rect 2591 28543 2649 28549
rect 1268 28512 2452 28540
rect 1268 28500 1274 28512
rect 750 28432 756 28484
rect 808 28472 814 28484
rect 1489 28475 1547 28481
rect 1489 28472 1501 28475
rect 808 28444 1501 28472
rect 808 28432 814 28444
rect 1489 28441 1501 28444
rect 1535 28441 1547 28475
rect 1489 28435 1547 28441
rect 1673 28475 1731 28481
rect 1673 28441 1685 28475
rect 1719 28472 1731 28475
rect 2314 28472 2320 28484
rect 1719 28444 2320 28472
rect 1719 28441 1731 28444
rect 1673 28435 1731 28441
rect 2314 28432 2320 28444
rect 2372 28432 2378 28484
rect 2424 28472 2452 28512
rect 2591 28509 2603 28543
rect 2637 28540 2649 28543
rect 3694 28540 3700 28552
rect 2637 28512 3700 28540
rect 2637 28509 2649 28512
rect 2591 28503 2649 28509
rect 3694 28500 3700 28512
rect 3752 28500 3758 28552
rect 4341 28543 4399 28549
rect 4341 28509 4353 28543
rect 4387 28540 4399 28543
rect 4430 28540 4436 28552
rect 4387 28512 4436 28540
rect 4387 28509 4399 28512
rect 4341 28503 4399 28509
rect 4430 28500 4436 28512
rect 4488 28500 4494 28552
rect 4522 28500 4528 28552
rect 4580 28540 4586 28552
rect 4580 28512 4936 28540
rect 4580 28500 4586 28512
rect 3234 28472 3240 28484
rect 2424 28444 3240 28472
rect 3234 28432 3240 28444
rect 3292 28432 3298 28484
rect 3786 28432 3792 28484
rect 3844 28472 3850 28484
rect 4249 28475 4307 28481
rect 4249 28472 4261 28475
rect 3844 28444 4261 28472
rect 3844 28432 3850 28444
rect 4249 28441 4261 28444
rect 4295 28441 4307 28475
rect 4249 28435 4307 28441
rect 4706 28432 4712 28484
rect 4764 28432 4770 28484
rect 4908 28416 4936 28512
rect 5442 28500 5448 28552
rect 5500 28500 5506 28552
rect 5719 28543 5777 28549
rect 5719 28509 5731 28543
rect 5765 28540 5777 28543
rect 8864 28540 8892 28580
rect 9490 28568 9496 28580
rect 9548 28568 9554 28620
rect 9600 28617 9628 28716
rect 10520 28676 10548 28716
rect 10597 28713 10609 28747
rect 10643 28744 10655 28747
rect 10686 28744 10692 28756
rect 10643 28716 10692 28744
rect 10643 28713 10655 28716
rect 10597 28707 10655 28713
rect 10686 28704 10692 28716
rect 10744 28704 10750 28756
rect 11514 28704 11520 28756
rect 11572 28744 11578 28756
rect 13449 28747 13507 28753
rect 11572 28716 12480 28744
rect 11572 28704 11578 28716
rect 10520 28648 10640 28676
rect 9585 28611 9643 28617
rect 9585 28577 9597 28611
rect 9631 28577 9643 28611
rect 9585 28571 9643 28577
rect 10612 28552 10640 28648
rect 12066 28636 12072 28688
rect 12124 28636 12130 28688
rect 5765 28512 8892 28540
rect 5765 28509 5777 28512
rect 5719 28503 5777 28509
rect 8938 28500 8944 28552
rect 8996 28540 9002 28552
rect 9827 28543 9885 28549
rect 9827 28540 9839 28543
rect 8996 28512 9839 28540
rect 8996 28500 9002 28512
rect 9827 28509 9839 28512
rect 9873 28509 9885 28543
rect 9827 28503 9885 28509
rect 10594 28500 10600 28552
rect 10652 28540 10658 28552
rect 11057 28543 11115 28549
rect 11057 28540 11069 28543
rect 10652 28512 11069 28540
rect 10652 28500 10658 28512
rect 11057 28509 11069 28512
rect 11103 28540 11115 28543
rect 11238 28540 11244 28552
rect 11103 28512 11244 28540
rect 11103 28509 11115 28512
rect 11057 28503 11115 28509
rect 11238 28500 11244 28512
rect 11296 28500 11302 28552
rect 11331 28543 11389 28549
rect 11331 28509 11343 28543
rect 11377 28540 11389 28543
rect 11422 28540 11428 28552
rect 11377 28512 11428 28540
rect 11377 28509 11389 28512
rect 11331 28503 11389 28509
rect 11422 28500 11428 28512
rect 11480 28500 11486 28552
rect 12452 28549 12480 28716
rect 13449 28713 13461 28747
rect 13495 28744 13507 28747
rect 13538 28744 13544 28756
rect 13495 28716 13544 28744
rect 13495 28713 13507 28716
rect 13449 28707 13507 28713
rect 13538 28704 13544 28716
rect 13596 28704 13602 28756
rect 13814 28704 13820 28756
rect 13872 28744 13878 28756
rect 14277 28747 14335 28753
rect 14277 28744 14289 28747
rect 13872 28716 14289 28744
rect 13872 28704 13878 28716
rect 14277 28713 14289 28716
rect 14323 28713 14335 28747
rect 14277 28707 14335 28713
rect 15304 28716 20576 28744
rect 12437 28543 12495 28549
rect 12437 28509 12449 28543
rect 12483 28540 12495 28543
rect 12711 28543 12769 28549
rect 12483 28512 12664 28540
rect 12483 28509 12495 28512
rect 12437 28503 12495 28509
rect 6086 28432 6092 28484
rect 6144 28472 6150 28484
rect 12636 28472 12664 28512
rect 12711 28509 12723 28543
rect 12757 28540 12769 28543
rect 12757 28512 13584 28540
rect 12757 28509 12769 28512
rect 12711 28503 12769 28509
rect 13170 28472 13176 28484
rect 6144 28444 12597 28472
rect 12636 28444 13176 28472
rect 6144 28432 6150 28444
rect 3326 28364 3332 28416
rect 3384 28404 3390 28416
rect 3973 28407 4031 28413
rect 3973 28404 3985 28407
rect 3384 28376 3985 28404
rect 3384 28364 3390 28376
rect 3973 28373 3985 28376
rect 4019 28404 4031 28407
rect 4614 28404 4620 28416
rect 4019 28376 4620 28404
rect 4019 28373 4031 28376
rect 3973 28367 4031 28373
rect 4614 28364 4620 28376
rect 4672 28364 4678 28416
rect 4890 28364 4896 28416
rect 4948 28404 4954 28416
rect 5077 28407 5135 28413
rect 5077 28404 5089 28407
rect 4948 28376 5089 28404
rect 4948 28364 4954 28376
rect 5077 28373 5089 28376
rect 5123 28373 5135 28407
rect 5077 28367 5135 28373
rect 5258 28364 5264 28416
rect 5316 28364 5322 28416
rect 6178 28364 6184 28416
rect 6236 28404 6242 28416
rect 6457 28407 6515 28413
rect 6457 28404 6469 28407
rect 6236 28376 6469 28404
rect 6236 28364 6242 28376
rect 6457 28373 6469 28376
rect 6503 28373 6515 28407
rect 6457 28367 6515 28373
rect 7650 28364 7656 28416
rect 7708 28404 7714 28416
rect 11606 28404 11612 28416
rect 7708 28376 11612 28404
rect 7708 28364 7714 28376
rect 11606 28364 11612 28376
rect 11664 28364 11670 28416
rect 12569 28404 12597 28444
rect 13170 28432 13176 28444
rect 13228 28432 13234 28484
rect 13556 28472 13584 28512
rect 13630 28500 13636 28552
rect 13688 28540 13694 28552
rect 13906 28540 13912 28552
rect 13688 28512 13912 28540
rect 13688 28500 13694 28512
rect 13906 28500 13912 28512
rect 13964 28500 13970 28552
rect 14182 28500 14188 28552
rect 14240 28500 14246 28552
rect 14550 28500 14556 28552
rect 14608 28540 14614 28552
rect 14645 28543 14703 28549
rect 14645 28540 14657 28543
rect 14608 28512 14657 28540
rect 14608 28500 14614 28512
rect 14645 28509 14657 28512
rect 14691 28509 14703 28543
rect 14887 28543 14945 28549
rect 14887 28540 14899 28543
rect 14645 28503 14703 28509
rect 14869 28509 14899 28540
rect 14933 28509 14945 28543
rect 14869 28503 14945 28509
rect 13814 28472 13820 28484
rect 13556 28444 13820 28472
rect 13814 28432 13820 28444
rect 13872 28432 13878 28484
rect 14200 28472 14228 28500
rect 14366 28472 14372 28484
rect 14200 28444 14372 28472
rect 14366 28432 14372 28444
rect 14424 28472 14430 28484
rect 14869 28472 14897 28503
rect 14424 28444 14897 28472
rect 14424 28432 14430 28444
rect 15304 28404 15332 28716
rect 18693 28679 18751 28685
rect 18693 28645 18705 28679
rect 18739 28645 18751 28679
rect 20548 28676 20576 28716
rect 20622 28704 20628 28756
rect 20680 28704 20686 28756
rect 23124 28716 23704 28744
rect 20714 28676 20720 28688
rect 20548 28648 20720 28676
rect 18693 28639 18751 28645
rect 17313 28543 17371 28549
rect 17313 28509 17325 28543
rect 17359 28540 17371 28543
rect 17954 28540 17960 28552
rect 17359 28512 17960 28540
rect 17359 28509 17371 28512
rect 17313 28503 17371 28509
rect 17954 28500 17960 28512
rect 18012 28500 18018 28552
rect 18708 28540 18736 28639
rect 20714 28636 20720 28648
rect 20772 28636 20778 28688
rect 23124 28685 23152 28716
rect 23109 28679 23167 28685
rect 23109 28676 23121 28679
rect 21100 28648 23121 28676
rect 20990 28568 20996 28620
rect 21048 28568 21054 28620
rect 18969 28543 19027 28549
rect 18969 28540 18981 28543
rect 18708 28512 18981 28540
rect 18969 28509 18981 28512
rect 19015 28509 19027 28543
rect 18969 28503 19027 28509
rect 19613 28543 19671 28549
rect 19613 28509 19625 28543
rect 19659 28509 19671 28543
rect 19613 28503 19671 28509
rect 19887 28543 19945 28549
rect 19887 28509 19899 28543
rect 19933 28540 19945 28543
rect 19978 28540 19984 28552
rect 19933 28512 19984 28540
rect 19933 28509 19945 28512
rect 19887 28503 19945 28509
rect 17586 28481 17592 28484
rect 17580 28435 17592 28481
rect 17644 28472 17650 28484
rect 19628 28472 19656 28503
rect 19978 28500 19984 28512
rect 20036 28500 20042 28552
rect 20070 28472 20076 28484
rect 17644 28444 17680 28472
rect 18708 28444 19564 28472
rect 19628 28444 20076 28472
rect 17586 28432 17592 28435
rect 17644 28432 17650 28444
rect 12569 28376 15332 28404
rect 15378 28364 15384 28416
rect 15436 28404 15442 28416
rect 15657 28407 15715 28413
rect 15657 28404 15669 28407
rect 15436 28376 15669 28404
rect 15436 28364 15442 28376
rect 15657 28373 15669 28376
rect 15703 28373 15715 28407
rect 15657 28367 15715 28373
rect 16482 28364 16488 28416
rect 16540 28404 16546 28416
rect 18708 28404 18736 28444
rect 16540 28376 18736 28404
rect 18785 28407 18843 28413
rect 16540 28364 16546 28376
rect 18785 28373 18797 28407
rect 18831 28404 18843 28407
rect 18966 28404 18972 28416
rect 18831 28376 18972 28404
rect 18831 28373 18843 28376
rect 18785 28367 18843 28373
rect 18966 28364 18972 28376
rect 19024 28364 19030 28416
rect 19536 28404 19564 28444
rect 20070 28432 20076 28444
rect 20128 28472 20134 28484
rect 21008 28472 21036 28568
rect 20128 28444 21036 28472
rect 20128 28432 20134 28444
rect 21100 28404 21128 28648
rect 23109 28645 23121 28648
rect 23155 28645 23167 28679
rect 23109 28639 23167 28645
rect 23477 28679 23535 28685
rect 23477 28645 23489 28679
rect 23523 28645 23535 28679
rect 23477 28639 23535 28645
rect 22094 28500 22100 28552
rect 22152 28500 22158 28552
rect 22833 28543 22891 28549
rect 22833 28509 22845 28543
rect 22879 28540 22891 28543
rect 23492 28540 23520 28639
rect 23676 28549 23704 28716
rect 22879 28512 23520 28540
rect 23661 28543 23719 28549
rect 22879 28509 22891 28512
rect 22833 28503 22891 28509
rect 23661 28509 23673 28543
rect 23707 28509 23719 28543
rect 23661 28503 23719 28509
rect 23937 28543 23995 28549
rect 23937 28509 23949 28543
rect 23983 28509 23995 28543
rect 23937 28503 23995 28509
rect 23952 28472 23980 28503
rect 22664 28444 23980 28472
rect 19536 28376 21128 28404
rect 22186 28364 22192 28416
rect 22244 28364 22250 28416
rect 22664 28413 22692 28444
rect 22649 28407 22707 28413
rect 22649 28373 22661 28407
rect 22695 28373 22707 28407
rect 22649 28367 22707 28373
rect 24121 28407 24179 28413
rect 24121 28373 24133 28407
rect 24167 28404 24179 28407
rect 24854 28404 24860 28416
rect 24167 28376 24860 28404
rect 24167 28373 24179 28376
rect 24121 28367 24179 28373
rect 24854 28364 24860 28376
rect 24912 28364 24918 28416
rect 1104 28314 24723 28336
rect 1104 28262 6814 28314
rect 6866 28262 6878 28314
rect 6930 28262 6942 28314
rect 6994 28262 7006 28314
rect 7058 28262 7070 28314
rect 7122 28262 12679 28314
rect 12731 28262 12743 28314
rect 12795 28262 12807 28314
rect 12859 28262 12871 28314
rect 12923 28262 12935 28314
rect 12987 28262 18544 28314
rect 18596 28262 18608 28314
rect 18660 28262 18672 28314
rect 18724 28262 18736 28314
rect 18788 28262 18800 28314
rect 18852 28262 24409 28314
rect 24461 28262 24473 28314
rect 24525 28262 24537 28314
rect 24589 28262 24601 28314
rect 24653 28262 24665 28314
rect 24717 28262 24723 28314
rect 1104 28240 24723 28262
rect 2314 28160 2320 28212
rect 2372 28200 2378 28212
rect 2372 28172 3188 28200
rect 2372 28160 2378 28172
rect 3160 28132 3188 28172
rect 3234 28160 3240 28212
rect 3292 28160 3298 28212
rect 3881 28203 3939 28209
rect 3881 28169 3893 28203
rect 3927 28200 3939 28203
rect 3927 28172 6040 28200
rect 3927 28169 3939 28172
rect 3881 28163 3939 28169
rect 4522 28132 4528 28144
rect 3160 28104 4528 28132
rect 4522 28092 4528 28104
rect 4580 28092 4586 28144
rect 4798 28092 4804 28144
rect 4856 28092 4862 28144
rect 5169 28135 5227 28141
rect 5169 28101 5181 28135
rect 5215 28132 5227 28135
rect 5810 28132 5816 28144
rect 5215 28104 5816 28132
rect 5215 28101 5227 28104
rect 5169 28095 5227 28101
rect 5810 28092 5816 28104
rect 5868 28092 5874 28144
rect 5905 28135 5963 28141
rect 5905 28101 5917 28135
rect 5951 28101 5963 28135
rect 6012 28132 6040 28172
rect 6086 28160 6092 28212
rect 6144 28160 6150 28212
rect 9677 28203 9735 28209
rect 8036 28172 9536 28200
rect 8036 28132 8064 28172
rect 6012 28104 8064 28132
rect 9508 28132 9536 28172
rect 9677 28169 9689 28203
rect 9723 28200 9735 28203
rect 10134 28200 10140 28212
rect 9723 28172 10140 28200
rect 9723 28169 9735 28172
rect 9677 28163 9735 28169
rect 10134 28160 10140 28172
rect 10192 28160 10198 28212
rect 11054 28200 11060 28212
rect 10428 28172 11060 28200
rect 10428 28132 10456 28172
rect 11054 28160 11060 28172
rect 11112 28160 11118 28212
rect 11624 28172 13490 28200
rect 11624 28144 11652 28172
rect 9508 28104 10456 28132
rect 5905 28095 5963 28101
rect 2314 28024 2320 28076
rect 2372 28024 2378 28076
rect 2406 28024 2412 28076
rect 2464 28073 2470 28076
rect 2464 28067 2492 28073
rect 2480 28033 2492 28067
rect 2464 28027 2492 28033
rect 3421 28067 3479 28073
rect 3421 28033 3433 28067
rect 3467 28033 3479 28067
rect 3421 28027 3479 28033
rect 2464 28024 2470 28027
rect 1397 27999 1455 28005
rect 1397 27965 1409 27999
rect 1443 27965 1455 27999
rect 1397 27959 1455 27965
rect 1581 27999 1639 28005
rect 1581 27965 1593 27999
rect 1627 27996 1639 27999
rect 2130 27996 2136 28008
rect 1627 27968 2136 27996
rect 1627 27965 1639 27968
rect 1581 27959 1639 27965
rect 1412 27928 1440 27959
rect 2130 27956 2136 27968
rect 2188 27956 2194 28008
rect 2590 27956 2596 28008
rect 2648 27956 2654 28008
rect 1486 27928 1492 27940
rect 1412 27900 1492 27928
rect 1486 27888 1492 27900
rect 1544 27928 1550 27940
rect 1762 27928 1768 27940
rect 1544 27900 1768 27928
rect 1544 27888 1550 27900
rect 1762 27888 1768 27900
rect 1820 27888 1826 27940
rect 2038 27888 2044 27940
rect 2096 27888 2102 27940
rect 3436 27928 3464 28027
rect 3694 28024 3700 28076
rect 3752 28024 3758 28076
rect 5077 28067 5135 28073
rect 5077 28033 5089 28067
rect 5123 28064 5135 28067
rect 5258 28064 5264 28076
rect 5123 28036 5264 28064
rect 5123 28033 5135 28036
rect 5077 28027 5135 28033
rect 5258 28024 5264 28036
rect 5316 28024 5322 28076
rect 5537 28067 5595 28073
rect 5537 28033 5549 28067
rect 5583 28064 5595 28067
rect 5626 28064 5632 28076
rect 5583 28036 5632 28064
rect 5583 28033 5595 28036
rect 5537 28027 5595 28033
rect 5626 28024 5632 28036
rect 5684 28024 5690 28076
rect 5920 28064 5948 28095
rect 10502 28092 10508 28144
rect 10560 28132 10566 28144
rect 10965 28135 11023 28141
rect 10965 28132 10977 28135
rect 10560 28104 10977 28132
rect 10560 28092 10566 28104
rect 10965 28101 10977 28104
rect 11011 28101 11023 28135
rect 10965 28095 11023 28101
rect 11606 28092 11612 28144
rect 11664 28092 11670 28144
rect 11698 28092 11704 28144
rect 11756 28092 11762 28144
rect 12805 28135 12863 28141
rect 12805 28101 12817 28135
rect 12851 28132 12863 28135
rect 12894 28132 12900 28144
rect 12851 28104 12900 28132
rect 12851 28101 12863 28104
rect 12805 28095 12863 28101
rect 12894 28092 12900 28104
rect 12952 28092 12958 28144
rect 13462 28103 13490 28172
rect 14090 28160 14096 28212
rect 14148 28200 14154 28212
rect 14185 28203 14243 28209
rect 14185 28200 14197 28203
rect 14148 28172 14197 28200
rect 14148 28160 14154 28172
rect 14185 28169 14197 28172
rect 14231 28169 14243 28203
rect 15194 28200 15200 28212
rect 14185 28163 14243 28169
rect 14660 28172 15200 28200
rect 13431 28097 13490 28103
rect 6362 28064 6368 28076
rect 5920 28036 6368 28064
rect 6362 28024 6368 28036
rect 6420 28024 6426 28076
rect 6546 28024 6552 28076
rect 6604 28064 6610 28076
rect 8202 28064 8208 28076
rect 6604 28036 8208 28064
rect 6604 28024 6610 28036
rect 8202 28024 8208 28036
rect 8260 28024 8266 28076
rect 8754 28024 8760 28076
rect 8812 28024 8818 28076
rect 9030 28024 9036 28076
rect 9088 28024 9094 28076
rect 10597 28067 10655 28073
rect 10597 28033 10609 28067
rect 10643 28064 10655 28067
rect 10778 28064 10784 28076
rect 10643 28036 10784 28064
rect 10643 28033 10655 28036
rect 10597 28027 10655 28033
rect 10778 28024 10784 28036
rect 10836 28024 10842 28076
rect 10888 28062 11744 28064
rect 11790 28062 11796 28076
rect 10888 28036 11796 28062
rect 6178 27996 6184 28008
rect 5842 27968 6184 27996
rect 6178 27956 6184 27968
rect 6236 27956 6242 28008
rect 6638 27956 6644 28008
rect 6696 27996 6702 28008
rect 7650 27996 7656 28008
rect 6696 27968 7656 27996
rect 6696 27956 6702 27968
rect 7650 27956 7656 27968
rect 7708 27996 7714 28008
rect 7837 27999 7895 28005
rect 7837 27996 7849 27999
rect 7708 27968 7849 27996
rect 7708 27956 7714 27968
rect 7837 27965 7849 27968
rect 7883 27965 7895 27999
rect 7837 27959 7895 27965
rect 8021 27999 8079 28005
rect 8021 27965 8033 27999
rect 8067 27965 8079 27999
rect 8021 27959 8079 27965
rect 3068 27900 3464 27928
rect 1302 27820 1308 27872
rect 1360 27860 1366 27872
rect 3068 27860 3096 27900
rect 7742 27888 7748 27940
rect 7800 27928 7806 27940
rect 8036 27928 8064 27959
rect 8386 27956 8392 28008
rect 8444 27996 8450 28008
rect 8481 27999 8539 28005
rect 8481 27996 8493 27999
rect 8444 27968 8493 27996
rect 8444 27956 8450 27968
rect 8481 27965 8493 27968
rect 8527 27965 8539 27999
rect 8481 27959 8539 27965
rect 8570 27956 8576 28008
rect 8628 27996 8634 28008
rect 8874 27999 8932 28005
rect 8874 27996 8886 27999
rect 8628 27968 8886 27996
rect 8628 27956 8634 27968
rect 8874 27965 8886 27968
rect 8920 27996 8932 27999
rect 9214 27996 9220 28008
rect 8920 27968 9220 27996
rect 8920 27965 8932 27968
rect 8874 27959 8932 27965
rect 9214 27956 9220 27968
rect 9272 27996 9278 28008
rect 9398 27996 9404 28008
rect 9272 27968 9404 27996
rect 9272 27956 9278 27968
rect 9398 27956 9404 27968
rect 9456 27956 9462 28008
rect 10686 27956 10692 28008
rect 10744 27956 10750 28008
rect 10888 27928 10916 28036
rect 11716 28034 11796 28036
rect 11790 28024 11796 28034
rect 11848 28064 11854 28076
rect 11977 28067 12035 28073
rect 11977 28064 11989 28067
rect 11848 28036 11989 28064
rect 11848 28024 11854 28036
rect 11977 28033 11989 28036
rect 12023 28033 12035 28067
rect 11977 28027 12035 28033
rect 12066 28024 12072 28076
rect 12124 28024 12130 28076
rect 12434 28024 12440 28076
rect 12492 28024 12498 28076
rect 13170 28024 13176 28076
rect 13228 28024 13234 28076
rect 13431 28063 13443 28097
rect 13477 28064 13490 28097
rect 14660 28073 14688 28172
rect 15194 28160 15200 28172
rect 15252 28160 15258 28212
rect 16390 28160 16396 28212
rect 16448 28200 16454 28212
rect 16758 28200 16764 28212
rect 16448 28172 16764 28200
rect 16448 28160 16454 28172
rect 16758 28160 16764 28172
rect 16816 28160 16822 28212
rect 17681 28203 17739 28209
rect 17681 28169 17693 28203
rect 17727 28169 17739 28203
rect 17681 28163 17739 28169
rect 16485 28135 16543 28141
rect 16485 28101 16497 28135
rect 16531 28101 16543 28135
rect 17696 28132 17724 28163
rect 18966 28160 18972 28212
rect 19024 28160 19030 28212
rect 21453 28203 21511 28209
rect 21453 28169 21465 28203
rect 21499 28200 21511 28203
rect 22094 28200 22100 28212
rect 21499 28172 22100 28200
rect 21499 28169 21511 28172
rect 21453 28163 21511 28169
rect 22094 28160 22100 28172
rect 22152 28160 22158 28212
rect 22186 28160 22192 28212
rect 22244 28160 22250 28212
rect 17696 28104 18276 28132
rect 16485 28095 16543 28101
rect 15746 28073 15752 28076
rect 14645 28067 14703 28073
rect 13477 28063 13860 28064
rect 13431 28057 13860 28063
rect 13462 28036 13860 28057
rect 11606 27956 11612 28008
rect 11664 27956 11670 28008
rect 7800 27900 8064 27928
rect 10152 27900 10916 27928
rect 7800 27888 7806 27900
rect 10152 27872 10180 27900
rect 12986 27888 12992 27940
rect 13044 27888 13050 27940
rect 1360 27832 3096 27860
rect 1360 27820 1366 27832
rect 3326 27820 3332 27872
rect 3384 27860 3390 27872
rect 3513 27863 3571 27869
rect 3513 27860 3525 27863
rect 3384 27832 3525 27860
rect 3384 27820 3390 27832
rect 3513 27829 3525 27832
rect 3559 27829 3571 27863
rect 3513 27823 3571 27829
rect 6086 27820 6092 27872
rect 6144 27860 6150 27872
rect 8754 27860 8760 27872
rect 6144 27832 8760 27860
rect 6144 27820 6150 27832
rect 8754 27820 8760 27832
rect 8812 27860 8818 27872
rect 10134 27860 10140 27872
rect 8812 27832 10140 27860
rect 8812 27820 8818 27832
rect 10134 27820 10140 27832
rect 10192 27820 10198 27872
rect 10778 27820 10784 27872
rect 10836 27860 10842 27872
rect 10873 27863 10931 27869
rect 10873 27860 10885 27863
rect 10836 27832 10885 27860
rect 10836 27820 10842 27832
rect 10873 27829 10885 27832
rect 10919 27829 10931 27863
rect 13832 27860 13860 28036
rect 14645 28033 14657 28067
rect 14691 28033 14703 28067
rect 14645 28027 14703 28033
rect 15703 28067 15752 28073
rect 15703 28033 15715 28067
rect 15749 28033 15752 28067
rect 15703 28027 15752 28033
rect 15746 28024 15752 28027
rect 15804 28024 15810 28076
rect 16500 28064 16528 28095
rect 17586 28064 17592 28076
rect 16500 28036 17592 28064
rect 17586 28024 17592 28036
rect 17644 28064 17650 28076
rect 18248 28073 18276 28104
rect 17865 28067 17923 28073
rect 17865 28064 17877 28067
rect 17644 28036 17877 28064
rect 17644 28024 17650 28036
rect 17865 28033 17877 28036
rect 17911 28033 17923 28067
rect 17865 28027 17923 28033
rect 18233 28067 18291 28073
rect 18233 28033 18245 28067
rect 18279 28033 18291 28067
rect 18233 28027 18291 28033
rect 18509 28067 18567 28073
rect 18509 28033 18521 28067
rect 18555 28064 18567 28067
rect 18877 28067 18935 28073
rect 18877 28064 18889 28067
rect 18555 28036 18889 28064
rect 18555 28033 18567 28036
rect 18509 28027 18567 28033
rect 18616 28008 18644 28036
rect 18877 28033 18889 28036
rect 18923 28033 18935 28067
rect 18984 28064 19012 28160
rect 20714 28092 20720 28144
rect 20772 28132 20778 28144
rect 21082 28132 21088 28144
rect 20772 28104 21088 28132
rect 20772 28092 20778 28104
rect 21082 28092 21088 28104
rect 21140 28132 21146 28144
rect 22204 28132 22232 28160
rect 21140 28104 21680 28132
rect 22204 28104 23520 28132
rect 21140 28092 21146 28104
rect 19061 28067 19119 28073
rect 19061 28064 19073 28067
rect 18984 28036 19073 28064
rect 18877 28027 18935 28033
rect 19061 28033 19073 28036
rect 19107 28033 19119 28067
rect 19061 28027 19119 28033
rect 20990 28024 20996 28076
rect 21048 28024 21054 28076
rect 21652 28073 21680 28104
rect 21637 28067 21695 28073
rect 21637 28033 21649 28067
rect 21683 28033 21695 28067
rect 21637 28027 21695 28033
rect 22279 28067 22337 28073
rect 22279 28033 22291 28067
rect 22325 28064 22337 28067
rect 22646 28064 22652 28076
rect 22325 28036 22652 28064
rect 22325 28033 22337 28036
rect 22279 28027 22337 28033
rect 22646 28024 22652 28036
rect 22704 28024 22710 28076
rect 23492 28073 23520 28104
rect 23385 28067 23443 28073
rect 23385 28064 23397 28067
rect 23032 28036 23397 28064
rect 13906 27956 13912 28008
rect 13964 27996 13970 28008
rect 14826 27996 14832 28008
rect 13964 27968 14832 27996
rect 13964 27956 13970 27968
rect 14826 27956 14832 27968
rect 14884 27956 14890 28008
rect 15289 27999 15347 28005
rect 15289 27965 15301 27999
rect 15335 27996 15347 27999
rect 15378 27996 15384 28008
rect 15335 27968 15384 27996
rect 15335 27965 15347 27968
rect 15289 27959 15347 27965
rect 15378 27956 15384 27968
rect 15436 27956 15442 28008
rect 15562 27956 15568 28008
rect 15620 27956 15626 28008
rect 15841 27999 15899 28005
rect 15841 27965 15853 27999
rect 15887 27996 15899 27999
rect 16482 27996 16488 28008
rect 15887 27968 16488 27996
rect 15887 27965 15899 27968
rect 15841 27959 15899 27965
rect 16482 27956 16488 27968
rect 16540 27956 16546 28008
rect 18598 27956 18604 28008
rect 18656 27956 18662 28008
rect 18785 27999 18843 28005
rect 18785 27965 18797 27999
rect 18831 27996 18843 27999
rect 18969 27999 19027 28005
rect 18969 27996 18981 27999
rect 18831 27968 18981 27996
rect 18831 27965 18843 27968
rect 18785 27959 18843 27965
rect 18969 27965 18981 27968
rect 19015 27965 19027 27999
rect 21008 27996 21036 28024
rect 22005 27999 22063 28005
rect 22005 27996 22017 27999
rect 21008 27968 22017 27996
rect 18969 27959 19027 27965
rect 22005 27965 22017 27968
rect 22051 27965 22063 27999
rect 22005 27959 22063 27965
rect 18230 27888 18236 27940
rect 18288 27928 18294 27940
rect 19702 27928 19708 27940
rect 18288 27900 19708 27928
rect 18288 27888 18294 27900
rect 19702 27888 19708 27900
rect 19760 27888 19766 27940
rect 14826 27860 14832 27872
rect 13832 27832 14832 27860
rect 10873 27823 10931 27829
rect 14826 27820 14832 27832
rect 14884 27820 14890 27872
rect 15562 27820 15568 27872
rect 15620 27860 15626 27872
rect 16022 27860 16028 27872
rect 15620 27832 16028 27860
rect 15620 27820 15626 27832
rect 16022 27820 16028 27832
rect 16080 27860 16086 27872
rect 16390 27860 16396 27872
rect 16080 27832 16396 27860
rect 16080 27820 16086 27832
rect 16390 27820 16396 27832
rect 16448 27820 16454 27872
rect 16758 27820 16764 27872
rect 16816 27860 16822 27872
rect 17586 27860 17592 27872
rect 16816 27832 17592 27860
rect 16816 27820 16822 27832
rect 17586 27820 17592 27832
rect 17644 27820 17650 27872
rect 18325 27863 18383 27869
rect 18325 27829 18337 27863
rect 18371 27860 18383 27863
rect 18601 27863 18659 27869
rect 18601 27860 18613 27863
rect 18371 27832 18613 27860
rect 18371 27829 18383 27832
rect 18325 27823 18383 27829
rect 18601 27829 18613 27832
rect 18647 27829 18659 27863
rect 18601 27823 18659 27829
rect 18693 27863 18751 27869
rect 18693 27829 18705 27863
rect 18739 27860 18751 27863
rect 22002 27860 22008 27872
rect 18739 27832 22008 27860
rect 18739 27829 18751 27832
rect 18693 27823 18751 27829
rect 22002 27820 22008 27832
rect 22060 27820 22066 27872
rect 22738 27820 22744 27872
rect 22796 27860 22802 27872
rect 23032 27869 23060 28036
rect 23385 28033 23397 28036
rect 23431 28033 23443 28067
rect 23385 28027 23443 28033
rect 23477 28067 23535 28073
rect 23477 28033 23489 28067
rect 23523 28033 23535 28067
rect 23477 28027 23535 28033
rect 23934 28024 23940 28076
rect 23992 28024 23998 28076
rect 23106 27956 23112 28008
rect 23164 27996 23170 28008
rect 23661 27999 23719 28005
rect 23661 27996 23673 27999
rect 23164 27968 23673 27996
rect 23164 27956 23170 27968
rect 23661 27965 23673 27968
rect 23707 27965 23719 27999
rect 23661 27959 23719 27965
rect 23017 27863 23075 27869
rect 23017 27860 23029 27863
rect 22796 27832 23029 27860
rect 22796 27820 22802 27832
rect 23017 27829 23029 27832
rect 23063 27829 23075 27863
rect 23017 27823 23075 27829
rect 23566 27820 23572 27872
rect 23624 27820 23630 27872
rect 24118 27820 24124 27872
rect 24176 27820 24182 27872
rect 1104 27770 24564 27792
rect 1104 27718 3882 27770
rect 3934 27718 3946 27770
rect 3998 27718 4010 27770
rect 4062 27718 4074 27770
rect 4126 27718 4138 27770
rect 4190 27718 9747 27770
rect 9799 27718 9811 27770
rect 9863 27718 9875 27770
rect 9927 27718 9939 27770
rect 9991 27718 10003 27770
rect 10055 27718 15612 27770
rect 15664 27718 15676 27770
rect 15728 27718 15740 27770
rect 15792 27718 15804 27770
rect 15856 27718 15868 27770
rect 15920 27718 21477 27770
rect 21529 27718 21541 27770
rect 21593 27718 21605 27770
rect 21657 27718 21669 27770
rect 21721 27718 21733 27770
rect 21785 27718 24564 27770
rect 1104 27696 24564 27718
rect 1688 27628 2268 27656
rect 842 27548 848 27600
rect 900 27588 906 27600
rect 1688 27588 1716 27628
rect 900 27560 1716 27588
rect 900 27548 906 27560
rect 2240 27520 2268 27628
rect 2590 27616 2596 27668
rect 2648 27616 2654 27668
rect 5442 27656 5448 27668
rect 5092 27628 5448 27656
rect 3421 27591 3479 27597
rect 3421 27557 3433 27591
rect 3467 27588 3479 27591
rect 3467 27560 4108 27588
rect 3467 27557 3479 27560
rect 3421 27551 3479 27557
rect 2240 27492 3832 27520
rect 1394 27412 1400 27464
rect 1452 27452 1458 27464
rect 1581 27455 1639 27461
rect 1581 27452 1593 27455
rect 1452 27424 1593 27452
rect 1452 27412 1458 27424
rect 1581 27421 1593 27424
rect 1627 27421 1639 27455
rect 1855 27455 1913 27461
rect 1855 27452 1867 27455
rect 1581 27415 1639 27421
rect 1780 27424 1867 27452
rect 1780 27396 1808 27424
rect 1855 27421 1867 27424
rect 1901 27452 1913 27455
rect 2866 27452 2872 27464
rect 1901 27442 2176 27452
rect 2240 27442 2872 27452
rect 1901 27424 2872 27442
rect 1901 27421 1913 27424
rect 1855 27415 1913 27421
rect 2148 27414 2268 27424
rect 2866 27412 2872 27424
rect 2924 27412 2930 27464
rect 2958 27412 2964 27464
rect 3016 27412 3022 27464
rect 3804 27461 3832 27492
rect 4080 27464 4108 27560
rect 5092 27529 5120 27628
rect 5442 27616 5448 27628
rect 5500 27656 5506 27668
rect 5500 27628 5762 27656
rect 5500 27616 5506 27628
rect 5077 27523 5135 27529
rect 5077 27489 5089 27523
rect 5123 27489 5135 27523
rect 5734 27520 5762 27628
rect 5810 27616 5816 27668
rect 5868 27616 5874 27668
rect 6546 27616 6552 27668
rect 6604 27656 6610 27668
rect 15194 27656 15200 27668
rect 6604 27628 15200 27656
rect 6604 27616 6610 27628
rect 15194 27616 15200 27628
rect 15252 27616 15258 27668
rect 16482 27616 16488 27668
rect 16540 27616 16546 27668
rect 18598 27616 18604 27668
rect 18656 27616 18662 27668
rect 23106 27656 23112 27668
rect 22756 27628 23112 27656
rect 5828 27588 5856 27616
rect 6089 27591 6147 27597
rect 6089 27588 6101 27591
rect 5828 27560 6101 27588
rect 6089 27557 6101 27560
rect 6135 27557 6147 27591
rect 8570 27588 8576 27600
rect 6089 27551 6147 27557
rect 8036 27560 8576 27588
rect 7009 27523 7067 27529
rect 7009 27520 7021 27523
rect 5734 27492 7021 27520
rect 5077 27483 5135 27489
rect 7009 27489 7021 27492
rect 7055 27489 7067 27523
rect 7009 27483 7067 27489
rect 3237 27455 3295 27461
rect 3237 27421 3249 27455
rect 3283 27421 3295 27455
rect 3237 27415 3295 27421
rect 3789 27455 3847 27461
rect 3789 27421 3801 27455
rect 3835 27421 3847 27455
rect 3789 27415 3847 27421
rect 1762 27344 1768 27396
rect 1820 27344 1826 27396
rect 3252 27384 3280 27415
rect 4062 27412 4068 27464
rect 4120 27412 4126 27464
rect 4982 27412 4988 27464
rect 5040 27452 5046 27464
rect 5319 27455 5377 27461
rect 5319 27452 5331 27455
rect 5040 27424 5331 27452
rect 5040 27412 5046 27424
rect 5319 27421 5331 27424
rect 5365 27421 5377 27455
rect 7282 27452 7288 27464
rect 7243 27424 7288 27452
rect 5319 27415 5377 27421
rect 7282 27412 7288 27424
rect 7340 27412 7346 27464
rect 8036 27384 8064 27560
rect 8570 27548 8576 27560
rect 8628 27548 8634 27600
rect 11606 27548 11612 27600
rect 11664 27588 11670 27600
rect 22756 27597 22784 27628
rect 23106 27616 23112 27628
rect 23164 27616 23170 27668
rect 23934 27616 23940 27668
rect 23992 27616 23998 27668
rect 11793 27591 11851 27597
rect 11793 27588 11805 27591
rect 11664 27560 11805 27588
rect 11664 27548 11670 27560
rect 11793 27557 11805 27560
rect 11839 27557 11851 27591
rect 11793 27551 11851 27557
rect 22189 27591 22247 27597
rect 22189 27557 22201 27591
rect 22235 27557 22247 27591
rect 22189 27551 22247 27557
rect 22373 27591 22431 27597
rect 22373 27557 22385 27591
rect 22419 27557 22431 27591
rect 22373 27551 22431 27557
rect 22741 27591 22799 27597
rect 22741 27557 22753 27591
rect 22787 27557 22799 27591
rect 22741 27551 22799 27557
rect 22925 27591 22983 27597
rect 22925 27557 22937 27591
rect 22971 27588 22983 27591
rect 23952 27588 23980 27616
rect 22971 27560 23980 27588
rect 22971 27557 22983 27560
rect 22925 27551 22983 27557
rect 8110 27480 8116 27532
rect 8168 27520 8174 27532
rect 9398 27520 9404 27532
rect 8168 27492 9404 27520
rect 8168 27480 8174 27492
rect 9398 27480 9404 27492
rect 9456 27480 9462 27532
rect 10134 27480 10140 27532
rect 10192 27520 10198 27532
rect 10410 27520 10416 27532
rect 10192 27492 10416 27520
rect 10192 27480 10198 27492
rect 10410 27480 10416 27492
rect 10468 27480 10474 27532
rect 10502 27480 10508 27532
rect 10560 27520 10566 27532
rect 10781 27523 10839 27529
rect 10781 27520 10793 27523
rect 10560 27492 10793 27520
rect 10560 27480 10566 27492
rect 10781 27489 10793 27492
rect 10827 27489 10839 27523
rect 10781 27483 10839 27489
rect 17494 27480 17500 27532
rect 17552 27520 17558 27532
rect 17589 27523 17647 27529
rect 17589 27520 17601 27523
rect 17552 27492 17601 27520
rect 17552 27480 17558 27492
rect 17589 27489 17601 27492
rect 17635 27489 17647 27523
rect 17589 27483 17647 27489
rect 2746 27356 3280 27384
rect 3896 27356 8064 27384
rect 1302 27276 1308 27328
rect 1360 27316 1366 27328
rect 2746 27316 2774 27356
rect 1360 27288 2774 27316
rect 3145 27319 3203 27325
rect 1360 27276 1366 27288
rect 3145 27285 3157 27319
rect 3191 27316 3203 27319
rect 3896 27316 3924 27356
rect 8128 27328 8156 27480
rect 11055 27455 11113 27461
rect 11055 27421 11067 27455
rect 11101 27452 11113 27455
rect 11790 27452 11796 27464
rect 11101 27424 11796 27452
rect 11101 27421 11113 27424
rect 11055 27415 11113 27421
rect 11790 27412 11796 27424
rect 11848 27452 11854 27464
rect 11848 27424 13584 27452
rect 11848 27412 11854 27424
rect 10410 27344 10416 27396
rect 10468 27384 10474 27396
rect 13446 27384 13452 27396
rect 10468 27356 13452 27384
rect 10468 27344 10474 27356
rect 13446 27344 13452 27356
rect 13504 27344 13510 27396
rect 13556 27384 13584 27424
rect 14090 27412 14096 27464
rect 14148 27412 14154 27464
rect 15473 27455 15531 27461
rect 15473 27452 15485 27455
rect 14367 27445 14425 27451
rect 14367 27411 14379 27445
rect 14413 27442 14425 27445
rect 14413 27414 14504 27442
rect 14413 27411 14425 27414
rect 14367 27405 14425 27411
rect 14182 27384 14188 27396
rect 13556 27356 14188 27384
rect 14182 27344 14188 27356
rect 14240 27344 14246 27396
rect 3191 27288 3924 27316
rect 3191 27285 3203 27288
rect 3145 27279 3203 27285
rect 3970 27276 3976 27328
rect 4028 27276 4034 27328
rect 5074 27276 5080 27328
rect 5132 27316 5138 27328
rect 6362 27316 6368 27328
rect 5132 27288 6368 27316
rect 5132 27276 5138 27288
rect 6362 27276 6368 27288
rect 6420 27276 6426 27328
rect 6638 27276 6644 27328
rect 6696 27316 6702 27328
rect 7190 27316 7196 27328
rect 6696 27288 7196 27316
rect 6696 27276 6702 27288
rect 7190 27276 7196 27288
rect 7248 27276 7254 27328
rect 7282 27276 7288 27328
rect 7340 27316 7346 27328
rect 7742 27316 7748 27328
rect 7340 27288 7748 27316
rect 7340 27276 7346 27288
rect 7742 27276 7748 27288
rect 7800 27276 7806 27328
rect 8018 27276 8024 27328
rect 8076 27276 8082 27328
rect 8110 27276 8116 27328
rect 8168 27276 8174 27328
rect 8662 27276 8668 27328
rect 8720 27316 8726 27328
rect 9030 27316 9036 27328
rect 8720 27288 9036 27316
rect 8720 27276 8726 27288
rect 9030 27276 9036 27288
rect 9088 27316 9094 27328
rect 14090 27316 14096 27328
rect 9088 27288 14096 27316
rect 9088 27276 9094 27288
rect 14090 27276 14096 27288
rect 14148 27316 14154 27328
rect 14476 27316 14504 27414
rect 14568 27424 15485 27452
rect 14568 27328 14596 27424
rect 15473 27421 15485 27424
rect 15519 27421 15531 27455
rect 15473 27415 15531 27421
rect 15715 27455 15773 27461
rect 15715 27421 15727 27455
rect 15761 27421 15773 27455
rect 17831 27455 17889 27461
rect 17831 27452 17843 27455
rect 15715 27415 15773 27421
rect 17696 27424 17843 27452
rect 15286 27344 15292 27396
rect 15344 27384 15350 27396
rect 15718 27384 15746 27415
rect 16022 27384 16028 27396
rect 15344 27356 16028 27384
rect 15344 27344 15350 27356
rect 16022 27344 16028 27356
rect 16080 27344 16086 27396
rect 17218 27344 17224 27396
rect 17276 27384 17282 27396
rect 17696 27384 17724 27424
rect 17831 27421 17843 27424
rect 17877 27421 17889 27455
rect 17831 27415 17889 27421
rect 17954 27412 17960 27464
rect 18012 27452 18018 27464
rect 21082 27461 21088 27464
rect 20809 27455 20867 27461
rect 20809 27452 20821 27455
rect 18012 27424 20821 27452
rect 18012 27412 18018 27424
rect 20809 27421 20821 27424
rect 20855 27421 20867 27455
rect 21076 27452 21088 27461
rect 21043 27424 21088 27452
rect 20809 27415 20867 27421
rect 21076 27415 21088 27424
rect 21082 27412 21088 27415
rect 21140 27412 21146 27464
rect 22204 27452 22232 27551
rect 22388 27520 22416 27551
rect 22388 27492 22876 27520
rect 22557 27455 22615 27461
rect 22557 27452 22569 27455
rect 22204 27424 22569 27452
rect 22557 27421 22569 27424
rect 22603 27421 22615 27455
rect 22557 27415 22615 27421
rect 22649 27455 22707 27461
rect 22649 27421 22661 27455
rect 22695 27452 22707 27455
rect 22738 27452 22744 27464
rect 22695 27424 22744 27452
rect 22695 27421 22707 27424
rect 22649 27415 22707 27421
rect 22738 27412 22744 27424
rect 22796 27412 22802 27464
rect 22848 27461 22876 27492
rect 23198 27480 23204 27532
rect 23256 27480 23262 27532
rect 22833 27455 22891 27461
rect 22833 27421 22845 27455
rect 22879 27421 22891 27455
rect 22833 27415 22891 27421
rect 23109 27455 23167 27461
rect 23109 27421 23121 27455
rect 23155 27452 23167 27455
rect 23216 27452 23244 27480
rect 23155 27424 23244 27452
rect 23155 27421 23167 27424
rect 23109 27415 23167 27421
rect 23290 27412 23296 27464
rect 23348 27452 23354 27464
rect 23385 27455 23443 27461
rect 23385 27452 23397 27455
rect 23348 27424 23397 27452
rect 23348 27412 23354 27424
rect 23385 27421 23397 27424
rect 23431 27421 23443 27455
rect 23845 27455 23903 27461
rect 23845 27452 23857 27455
rect 23385 27415 23443 27421
rect 23584 27424 23857 27452
rect 23584 27384 23612 27424
rect 23845 27421 23857 27424
rect 23891 27421 23903 27455
rect 23845 27415 23903 27421
rect 23937 27455 23995 27461
rect 23937 27421 23949 27455
rect 23983 27421 23995 27455
rect 23937 27415 23995 27421
rect 23952 27384 23980 27415
rect 17276 27356 17724 27384
rect 23216 27356 23612 27384
rect 23676 27356 23980 27384
rect 17276 27344 17282 27356
rect 14148 27288 14504 27316
rect 14148 27276 14154 27288
rect 14550 27276 14556 27328
rect 14608 27276 14614 27328
rect 15102 27276 15108 27328
rect 15160 27276 15166 27328
rect 16206 27276 16212 27328
rect 16264 27316 16270 27328
rect 19334 27316 19340 27328
rect 16264 27288 19340 27316
rect 16264 27276 16270 27288
rect 19334 27276 19340 27288
rect 19392 27316 19398 27328
rect 20990 27316 20996 27328
rect 19392 27288 20996 27316
rect 19392 27276 19398 27288
rect 20990 27276 20996 27288
rect 21048 27276 21054 27328
rect 23216 27325 23244 27356
rect 23676 27325 23704 27356
rect 23201 27319 23259 27325
rect 23201 27285 23213 27319
rect 23247 27285 23259 27319
rect 23201 27279 23259 27285
rect 23661 27319 23719 27325
rect 23661 27285 23673 27319
rect 23707 27285 23719 27319
rect 23661 27279 23719 27285
rect 24121 27319 24179 27325
rect 24121 27285 24133 27319
rect 24167 27316 24179 27319
rect 24854 27316 24860 27328
rect 24167 27288 24860 27316
rect 24167 27285 24179 27288
rect 24121 27279 24179 27285
rect 24854 27276 24860 27288
rect 24912 27276 24918 27328
rect 1104 27226 24723 27248
rect 1104 27174 6814 27226
rect 6866 27174 6878 27226
rect 6930 27174 6942 27226
rect 6994 27174 7006 27226
rect 7058 27174 7070 27226
rect 7122 27174 12679 27226
rect 12731 27174 12743 27226
rect 12795 27174 12807 27226
rect 12859 27174 12871 27226
rect 12923 27174 12935 27226
rect 12987 27174 18544 27226
rect 18596 27174 18608 27226
rect 18660 27174 18672 27226
rect 18724 27174 18736 27226
rect 18788 27174 18800 27226
rect 18852 27174 24409 27226
rect 24461 27174 24473 27226
rect 24525 27174 24537 27226
rect 24589 27174 24601 27226
rect 24653 27174 24665 27226
rect 24717 27174 24723 27226
rect 1104 27152 24723 27174
rect 2038 27072 2044 27124
rect 2096 27112 2102 27124
rect 2409 27115 2467 27121
rect 2409 27112 2421 27115
rect 2096 27084 2421 27112
rect 2096 27072 2102 27084
rect 2409 27081 2421 27084
rect 2455 27081 2467 27115
rect 2958 27112 2964 27124
rect 2409 27075 2467 27081
rect 2746 27084 2964 27112
rect 1210 27004 1216 27056
rect 1268 27044 1274 27056
rect 2746 27044 2774 27084
rect 2958 27072 2964 27084
rect 3016 27072 3022 27124
rect 3237 27115 3295 27121
rect 3237 27081 3249 27115
rect 3283 27081 3295 27115
rect 3237 27075 3295 27081
rect 3513 27115 3571 27121
rect 3513 27081 3525 27115
rect 3559 27112 3571 27115
rect 6546 27112 6552 27124
rect 3559 27084 6552 27112
rect 3559 27081 3571 27084
rect 3513 27075 3571 27081
rect 1268 27016 2774 27044
rect 3252 27044 3280 27075
rect 6546 27072 6552 27084
rect 6604 27072 6610 27124
rect 6638 27072 6644 27124
rect 6696 27112 6702 27124
rect 7009 27115 7067 27121
rect 7009 27112 7021 27115
rect 6696 27084 7021 27112
rect 6696 27072 6702 27084
rect 7009 27081 7021 27084
rect 7055 27081 7067 27115
rect 7834 27112 7840 27124
rect 7009 27075 7067 27081
rect 7116 27084 7840 27112
rect 5626 27044 5632 27056
rect 3252 27016 5632 27044
rect 1268 27004 1274 27016
rect 5626 27004 5632 27016
rect 5684 27004 5690 27056
rect 6822 27004 6828 27056
rect 6880 27044 6886 27056
rect 7116 27044 7144 27084
rect 7834 27072 7840 27084
rect 7892 27112 7898 27124
rect 7892 27084 8156 27112
rect 7892 27072 7898 27084
rect 6880 27016 7144 27044
rect 6880 27004 6886 27016
rect 7282 27004 7288 27056
rect 7340 27004 7346 27056
rect 7377 27047 7435 27053
rect 7377 27013 7389 27047
rect 7423 27044 7435 27047
rect 8018 27044 8024 27056
rect 7423 27016 8024 27044
rect 7423 27013 7435 27016
rect 7377 27007 7435 27013
rect 8018 27004 8024 27016
rect 8076 27004 8082 27056
rect 8128 27053 8156 27084
rect 8386 27072 8392 27124
rect 8444 27072 8450 27124
rect 8754 27072 8760 27124
rect 8812 27112 8818 27124
rect 11330 27112 11336 27124
rect 8812 27084 11336 27112
rect 8812 27072 8818 27084
rect 11330 27072 11336 27084
rect 11388 27072 11394 27124
rect 14182 27072 14188 27124
rect 14240 27112 14246 27124
rect 14240 27084 23336 27112
rect 14240 27072 14246 27084
rect 8113 27047 8171 27053
rect 8113 27013 8125 27047
rect 8159 27013 8171 27047
rect 8113 27007 8171 27013
rect 1671 26979 1729 26985
rect 1671 26945 1683 26979
rect 1717 26976 1729 26979
rect 2682 26976 2688 26988
rect 1717 26948 2688 26976
rect 1717 26945 1729 26948
rect 1671 26939 1729 26945
rect 2682 26936 2688 26948
rect 2740 26936 2746 26988
rect 2774 26936 2780 26988
rect 2832 26936 2838 26988
rect 2866 26936 2872 26988
rect 2924 26976 2930 26988
rect 3053 26979 3111 26985
rect 3053 26976 3065 26979
rect 2924 26948 3065 26976
rect 2924 26936 2930 26948
rect 3053 26945 3065 26948
rect 3099 26945 3111 26979
rect 3053 26939 3111 26945
rect 3329 26979 3387 26985
rect 3329 26945 3341 26979
rect 3375 26945 3387 26979
rect 3329 26939 3387 26945
rect 1394 26868 1400 26920
rect 1452 26868 1458 26920
rect 3344 26840 3372 26939
rect 3602 26936 3608 26988
rect 3660 26936 3666 26988
rect 3878 26976 3884 26988
rect 3839 26948 3884 26976
rect 3878 26936 3884 26948
rect 3936 26936 3942 26988
rect 3970 26936 3976 26988
rect 4028 26976 4034 26988
rect 7466 26976 7472 26988
rect 4028 26948 7472 26976
rect 4028 26936 4034 26948
rect 7466 26936 7472 26948
rect 7524 26976 7530 26988
rect 7745 26979 7803 26985
rect 7745 26976 7757 26979
rect 7524 26948 7757 26976
rect 7524 26936 7530 26948
rect 7745 26945 7757 26948
rect 7791 26945 7803 26979
rect 7745 26939 7803 26945
rect 8404 26920 8432 27072
rect 8662 27004 8668 27056
rect 8720 27044 8726 27056
rect 8720 27016 9674 27044
rect 8720 27004 8726 27016
rect 8999 26979 9057 26985
rect 8999 26945 9011 26979
rect 9045 26976 9057 26979
rect 9398 26976 9404 26988
rect 9045 26948 9404 26976
rect 9045 26945 9057 26948
rect 8999 26939 9057 26945
rect 9398 26936 9404 26948
rect 9456 26936 9462 26988
rect 7190 26868 7196 26920
rect 7248 26868 7254 26920
rect 8386 26868 8392 26920
rect 8444 26868 8450 26920
rect 8662 26868 8668 26920
rect 8720 26908 8726 26920
rect 8757 26911 8815 26917
rect 8757 26908 8769 26911
rect 8720 26880 8769 26908
rect 8720 26868 8726 26880
rect 8757 26877 8769 26880
rect 8803 26877 8815 26911
rect 9646 26908 9674 27016
rect 13814 27004 13820 27056
rect 13872 27044 13878 27056
rect 15930 27044 15936 27056
rect 13872 27016 15936 27044
rect 13872 27004 13878 27016
rect 15930 27004 15936 27016
rect 15988 27004 15994 27056
rect 16206 27004 16212 27056
rect 16264 27004 16270 27056
rect 20438 27044 20444 27056
rect 17420 27016 20444 27044
rect 12527 26979 12585 26985
rect 12527 26976 12539 26979
rect 11716 26948 12539 26976
rect 9646 26880 11376 26908
rect 8757 26871 8815 26877
rect 5350 26840 5356 26852
rect 2746 26812 3372 26840
rect 4540 26812 5356 26840
rect 1302 26732 1308 26784
rect 1360 26772 1366 26784
rect 2746 26772 2774 26812
rect 1360 26744 2774 26772
rect 2961 26775 3019 26781
rect 1360 26732 1366 26744
rect 2961 26741 2973 26775
rect 3007 26772 3019 26775
rect 3510 26772 3516 26784
rect 3007 26744 3516 26772
rect 3007 26741 3019 26744
rect 2961 26735 3019 26741
rect 3510 26732 3516 26744
rect 3568 26732 3574 26784
rect 4062 26732 4068 26784
rect 4120 26772 4126 26784
rect 4540 26772 4568 26812
rect 5350 26800 5356 26812
rect 5408 26800 5414 26852
rect 11348 26840 11376 26880
rect 11422 26868 11428 26920
rect 11480 26908 11486 26920
rect 11716 26908 11744 26948
rect 12527 26945 12539 26948
rect 12573 26976 12585 26979
rect 16224 26976 16252 27004
rect 12573 26948 16252 26976
rect 12573 26945 12585 26948
rect 12527 26939 12585 26945
rect 11480 26880 11744 26908
rect 12253 26911 12311 26917
rect 11480 26868 11486 26880
rect 12253 26877 12265 26911
rect 12299 26877 12311 26911
rect 17420 26908 17448 27016
rect 20438 27004 20444 27016
rect 20496 27044 20502 27056
rect 20496 27016 20944 27044
rect 20496 27004 20502 27016
rect 17494 26936 17500 26988
rect 17552 26936 17558 26988
rect 18138 26936 18144 26988
rect 18196 26976 18202 26988
rect 19150 26976 19156 26988
rect 18196 26948 19156 26976
rect 18196 26936 18202 26948
rect 19150 26936 19156 26948
rect 19208 26976 19214 26988
rect 19243 26979 19301 26985
rect 19243 26976 19255 26979
rect 19208 26948 19255 26976
rect 19208 26936 19214 26948
rect 19243 26945 19255 26948
rect 19289 26945 19301 26979
rect 20349 26979 20407 26985
rect 20349 26976 20361 26979
rect 19243 26939 19301 26945
rect 19996 26948 20361 26976
rect 12253 26871 12311 26877
rect 13096 26880 17448 26908
rect 17512 26908 17540 26936
rect 18969 26911 19027 26917
rect 18969 26908 18981 26911
rect 17512 26880 18981 26908
rect 11606 26840 11612 26852
rect 9416 26812 10364 26840
rect 11348 26812 11612 26840
rect 4120 26744 4568 26772
rect 4617 26775 4675 26781
rect 4120 26732 4126 26744
rect 4617 26741 4629 26775
rect 4663 26772 4675 26775
rect 4982 26772 4988 26784
rect 4663 26744 4988 26772
rect 4663 26741 4675 26744
rect 4617 26735 4675 26741
rect 4982 26732 4988 26744
rect 5040 26732 5046 26784
rect 5166 26732 5172 26784
rect 5224 26772 5230 26784
rect 6362 26772 6368 26784
rect 5224 26744 6368 26772
rect 5224 26732 5230 26744
rect 6362 26732 6368 26744
rect 6420 26732 6426 26784
rect 8297 26775 8355 26781
rect 8297 26741 8309 26775
rect 8343 26772 8355 26775
rect 9416 26772 9444 26812
rect 8343 26744 9444 26772
rect 8343 26741 8355 26744
rect 8297 26735 8355 26741
rect 9490 26732 9496 26784
rect 9548 26772 9554 26784
rect 9769 26775 9827 26781
rect 9769 26772 9781 26775
rect 9548 26744 9781 26772
rect 9548 26732 9554 26744
rect 9769 26741 9781 26744
rect 9815 26741 9827 26775
rect 10336 26772 10364 26812
rect 11606 26800 11612 26812
rect 11664 26840 11670 26852
rect 12268 26840 12296 26871
rect 11664 26812 12296 26840
rect 11664 26800 11670 26812
rect 13096 26772 13124 26880
rect 18969 26877 18981 26880
rect 19015 26877 19027 26911
rect 18969 26871 19027 26877
rect 16482 26800 16488 26852
rect 16540 26840 16546 26852
rect 16850 26840 16856 26852
rect 16540 26812 16856 26840
rect 16540 26800 16546 26812
rect 16850 26800 16856 26812
rect 16908 26800 16914 26852
rect 10336 26744 13124 26772
rect 9769 26735 9827 26741
rect 13170 26732 13176 26784
rect 13228 26772 13234 26784
rect 13265 26775 13323 26781
rect 13265 26772 13277 26775
rect 13228 26744 13277 26772
rect 13228 26732 13234 26744
rect 13265 26741 13277 26744
rect 13311 26741 13323 26775
rect 13265 26735 13323 26741
rect 15010 26732 15016 26784
rect 15068 26772 15074 26784
rect 17402 26772 17408 26784
rect 15068 26744 17408 26772
rect 15068 26732 15074 26744
rect 17402 26732 17408 26744
rect 17460 26732 17466 26784
rect 19794 26732 19800 26784
rect 19852 26772 19858 26784
rect 19996 26781 20024 26948
rect 20349 26945 20361 26948
rect 20395 26945 20407 26979
rect 20349 26939 20407 26945
rect 20530 26936 20536 26988
rect 20588 26936 20594 26988
rect 20916 26985 20944 27016
rect 20990 27004 20996 27056
rect 21048 27044 21054 27056
rect 23198 27044 23204 27056
rect 21048 27016 23204 27044
rect 21048 27004 21054 27016
rect 23198 27004 23204 27016
rect 23256 27004 23262 27056
rect 23308 26985 23336 27084
rect 25130 27072 25136 27124
rect 25188 27072 25194 27124
rect 20901 26979 20959 26985
rect 20901 26945 20913 26979
rect 20947 26945 20959 26979
rect 20901 26939 20959 26945
rect 23293 26979 23351 26985
rect 23293 26945 23305 26979
rect 23339 26945 23351 26979
rect 23845 26979 23903 26985
rect 23845 26976 23857 26979
rect 23293 26939 23351 26945
rect 23492 26948 23857 26976
rect 23492 26908 23520 26948
rect 23845 26945 23857 26948
rect 23891 26945 23903 26979
rect 23845 26939 23903 26945
rect 23937 26979 23995 26985
rect 23937 26945 23949 26979
rect 23983 26945 23995 26979
rect 23937 26939 23995 26945
rect 23952 26908 23980 26939
rect 25148 26920 25176 27072
rect 23124 26880 23520 26908
rect 23676 26880 23980 26908
rect 23124 26849 23152 26880
rect 23676 26849 23704 26880
rect 25130 26868 25136 26920
rect 25188 26868 25194 26920
rect 23109 26843 23167 26849
rect 23109 26809 23121 26843
rect 23155 26809 23167 26843
rect 23109 26803 23167 26809
rect 23661 26843 23719 26849
rect 23661 26809 23673 26843
rect 23707 26809 23719 26843
rect 23661 26803 23719 26809
rect 19981 26775 20039 26781
rect 19981 26772 19993 26775
rect 19852 26744 19993 26772
rect 19852 26732 19858 26744
rect 19981 26741 19993 26744
rect 20027 26741 20039 26775
rect 19981 26735 20039 26741
rect 20162 26732 20168 26784
rect 20220 26772 20226 26784
rect 20441 26775 20499 26781
rect 20441 26772 20453 26775
rect 20220 26744 20453 26772
rect 20220 26732 20226 26744
rect 20441 26741 20453 26744
rect 20487 26741 20499 26775
rect 20441 26735 20499 26741
rect 20714 26732 20720 26784
rect 20772 26732 20778 26784
rect 24118 26732 24124 26784
rect 24176 26732 24182 26784
rect 24210 26732 24216 26784
rect 24268 26772 24274 26784
rect 25222 26772 25228 26784
rect 24268 26744 25228 26772
rect 24268 26732 24274 26744
rect 25222 26732 25228 26744
rect 25280 26732 25286 26784
rect 1104 26682 24564 26704
rect 1104 26630 3882 26682
rect 3934 26630 3946 26682
rect 3998 26630 4010 26682
rect 4062 26630 4074 26682
rect 4126 26630 4138 26682
rect 4190 26630 9747 26682
rect 9799 26630 9811 26682
rect 9863 26630 9875 26682
rect 9927 26630 9939 26682
rect 9991 26630 10003 26682
rect 10055 26630 15612 26682
rect 15664 26630 15676 26682
rect 15728 26630 15740 26682
rect 15792 26630 15804 26682
rect 15856 26630 15868 26682
rect 15920 26630 21477 26682
rect 21529 26630 21541 26682
rect 21593 26630 21605 26682
rect 21657 26630 21669 26682
rect 21721 26630 21733 26682
rect 21785 26630 24564 26682
rect 1104 26608 24564 26630
rect 1857 26571 1915 26577
rect 1857 26537 1869 26571
rect 1903 26568 1915 26571
rect 6822 26568 6828 26580
rect 1903 26540 6828 26568
rect 1903 26537 1915 26540
rect 1857 26531 1915 26537
rect 6822 26528 6828 26540
rect 6880 26528 6886 26580
rect 7101 26571 7159 26577
rect 7101 26537 7113 26571
rect 7147 26568 7159 26571
rect 7190 26568 7196 26580
rect 7147 26540 7196 26568
rect 7147 26537 7159 26540
rect 7101 26531 7159 26537
rect 7190 26528 7196 26540
rect 7248 26528 7254 26580
rect 10410 26528 10416 26580
rect 10468 26528 10474 26580
rect 13078 26568 13084 26580
rect 10520 26540 13084 26568
rect 1394 26460 1400 26512
rect 1452 26460 1458 26512
rect 1581 26503 1639 26509
rect 1581 26469 1593 26503
rect 1627 26500 1639 26503
rect 2038 26500 2044 26512
rect 1627 26472 2044 26500
rect 1627 26469 1639 26472
rect 1581 26463 1639 26469
rect 2038 26460 2044 26472
rect 2096 26460 2102 26512
rect 3145 26503 3203 26509
rect 3145 26500 3157 26503
rect 3068 26472 3157 26500
rect 1412 26432 1440 26460
rect 3068 26444 3096 26472
rect 3145 26469 3157 26472
rect 3191 26469 3203 26503
rect 3145 26463 3203 26469
rect 4430 26460 4436 26512
rect 4488 26460 4494 26512
rect 5442 26460 5448 26512
rect 5500 26500 5506 26512
rect 8481 26503 8539 26509
rect 5500 26472 6132 26500
rect 5500 26460 5506 26472
rect 2133 26435 2191 26441
rect 2133 26432 2145 26435
rect 1228 26404 2145 26432
rect 1228 26376 1256 26404
rect 2133 26401 2145 26404
rect 2179 26401 2191 26435
rect 2133 26395 2191 26401
rect 3050 26392 3056 26444
rect 3108 26392 3114 26444
rect 3786 26392 3792 26444
rect 3844 26392 3850 26444
rect 4338 26392 4344 26444
rect 4396 26432 4402 26444
rect 6104 26441 6132 26472
rect 8481 26469 8493 26503
rect 8527 26500 8539 26503
rect 10520 26500 10548 26540
rect 13078 26528 13084 26540
rect 13136 26528 13142 26580
rect 13446 26528 13452 26580
rect 13504 26568 13510 26580
rect 19886 26568 19892 26580
rect 13504 26540 19892 26568
rect 13504 26528 13510 26540
rect 19886 26528 19892 26540
rect 19944 26528 19950 26580
rect 8527 26472 8984 26500
rect 8527 26469 8539 26472
rect 8481 26463 8539 26469
rect 4709 26435 4767 26441
rect 4709 26432 4721 26435
rect 4396 26404 4721 26432
rect 4396 26392 4402 26404
rect 4709 26401 4721 26404
rect 4755 26401 4767 26435
rect 4709 26395 4767 26401
rect 4847 26435 4905 26441
rect 4847 26401 4859 26435
rect 4893 26432 4905 26435
rect 6089 26435 6147 26441
rect 4893 26404 5764 26432
rect 4893 26401 4905 26404
rect 4847 26395 4905 26401
rect 5736 26376 5764 26404
rect 6089 26401 6101 26435
rect 6135 26401 6147 26435
rect 7374 26432 7380 26444
rect 6089 26395 6147 26401
rect 7300 26404 7380 26432
rect 1210 26324 1216 26376
rect 1268 26324 1274 26376
rect 1394 26324 1400 26376
rect 1452 26324 1458 26376
rect 1670 26324 1676 26376
rect 1728 26324 1734 26376
rect 2407 26367 2465 26373
rect 2407 26333 2419 26367
rect 2453 26364 2465 26367
rect 2498 26364 2504 26376
rect 2453 26336 2504 26364
rect 2453 26333 2465 26336
rect 2407 26327 2465 26333
rect 2498 26324 2504 26336
rect 2556 26324 2562 26376
rect 3973 26367 4031 26373
rect 3973 26333 3985 26367
rect 4019 26333 4031 26367
rect 3973 26327 4031 26333
rect 1946 26188 1952 26240
rect 2004 26228 2010 26240
rect 3142 26228 3148 26240
rect 2004 26200 3148 26228
rect 2004 26188 2010 26200
rect 3142 26188 3148 26200
rect 3200 26188 3206 26240
rect 3988 26228 4016 26327
rect 4982 26324 4988 26376
rect 5040 26324 5046 26376
rect 5718 26324 5724 26376
rect 5776 26324 5782 26376
rect 5810 26324 5816 26376
rect 5868 26364 5874 26376
rect 6331 26367 6389 26373
rect 6331 26364 6343 26367
rect 5868 26336 6343 26364
rect 5868 26324 5874 26336
rect 6331 26333 6343 26336
rect 6377 26333 6389 26367
rect 6331 26327 6389 26333
rect 5626 26256 5632 26308
rect 5684 26256 5690 26308
rect 4706 26228 4712 26240
rect 3988 26200 4712 26228
rect 4706 26188 4712 26200
rect 4764 26228 4770 26240
rect 5994 26228 6000 26240
rect 4764 26200 6000 26228
rect 4764 26188 4770 26200
rect 5994 26188 6000 26200
rect 6052 26188 6058 26240
rect 6270 26188 6276 26240
rect 6328 26228 6334 26240
rect 6638 26228 6644 26240
rect 6328 26200 6644 26228
rect 6328 26188 6334 26200
rect 6638 26188 6644 26200
rect 6696 26228 6702 26240
rect 7300 26228 7328 26404
rect 7374 26392 7380 26404
rect 7432 26432 7438 26444
rect 7469 26435 7527 26441
rect 7469 26432 7481 26435
rect 7432 26404 7481 26432
rect 7432 26392 7438 26404
rect 7469 26401 7481 26404
rect 7515 26401 7527 26435
rect 8956 26418 8984 26472
rect 10244 26472 10548 26500
rect 10689 26503 10747 26509
rect 7469 26395 7527 26401
rect 7711 26367 7769 26373
rect 7711 26364 7723 26367
rect 7392 26336 7723 26364
rect 7392 26240 7420 26336
rect 7711 26333 7723 26336
rect 7757 26333 7769 26367
rect 7711 26327 7769 26333
rect 7834 26324 7840 26376
rect 7892 26364 7898 26376
rect 9861 26367 9919 26373
rect 9861 26364 9873 26367
rect 7892 26336 9873 26364
rect 7892 26324 7898 26336
rect 9861 26333 9873 26336
rect 9907 26333 9919 26367
rect 9861 26327 9919 26333
rect 8478 26256 8484 26308
rect 8536 26296 8542 26308
rect 9125 26299 9183 26305
rect 9125 26296 9137 26299
rect 8536 26268 9137 26296
rect 8536 26256 8542 26268
rect 9125 26265 9137 26268
rect 9171 26265 9183 26299
rect 9125 26259 9183 26265
rect 9214 26256 9220 26308
rect 9272 26296 9278 26308
rect 9401 26299 9459 26305
rect 9401 26296 9413 26299
rect 9272 26268 9413 26296
rect 9272 26256 9278 26268
rect 9401 26265 9413 26268
rect 9447 26265 9459 26299
rect 9401 26259 9459 26265
rect 9490 26256 9496 26308
rect 9548 26256 9554 26308
rect 10244 26305 10272 26472
rect 10689 26469 10701 26503
rect 10735 26500 10747 26503
rect 11057 26503 11115 26509
rect 11057 26500 11069 26503
rect 10735 26472 11069 26500
rect 10735 26469 10747 26472
rect 10689 26463 10747 26469
rect 11057 26469 11069 26472
rect 11103 26469 11115 26503
rect 21637 26503 21695 26509
rect 11057 26463 11115 26469
rect 17972 26472 20300 26500
rect 17972 26444 18000 26472
rect 10873 26435 10931 26441
rect 10873 26401 10885 26435
rect 10919 26432 10931 26435
rect 11333 26435 11391 26441
rect 11333 26432 11345 26435
rect 10919 26404 11345 26432
rect 10919 26401 10931 26404
rect 10873 26395 10931 26401
rect 11333 26401 11345 26404
rect 11379 26401 11391 26435
rect 14550 26432 14556 26444
rect 11333 26395 11391 26401
rect 14108 26404 14556 26432
rect 10597 26367 10655 26373
rect 10597 26333 10609 26367
rect 10643 26333 10655 26367
rect 10597 26327 10655 26333
rect 10229 26299 10287 26305
rect 10229 26296 10241 26299
rect 9692 26268 10241 26296
rect 6696 26200 7328 26228
rect 6696 26188 6702 26200
rect 7374 26188 7380 26240
rect 7432 26188 7438 26240
rect 7742 26188 7748 26240
rect 7800 26228 7806 26240
rect 8202 26228 8208 26240
rect 7800 26200 8208 26228
rect 7800 26188 7806 26200
rect 8202 26188 8208 26200
rect 8260 26228 8266 26240
rect 9692 26228 9720 26268
rect 10229 26265 10241 26268
rect 10275 26265 10287 26299
rect 10612 26296 10640 26327
rect 10962 26324 10968 26376
rect 11020 26324 11026 26376
rect 11241 26367 11299 26373
rect 11241 26333 11253 26367
rect 11287 26333 11299 26367
rect 11241 26327 11299 26333
rect 10686 26296 10692 26308
rect 10612 26268 10692 26296
rect 10229 26259 10287 26265
rect 10686 26256 10692 26268
rect 10744 26296 10750 26308
rect 11256 26296 11284 26327
rect 11422 26324 11428 26376
rect 11480 26324 11486 26376
rect 11885 26367 11943 26373
rect 11885 26333 11897 26367
rect 11931 26333 11943 26367
rect 11885 26327 11943 26333
rect 12159 26367 12217 26373
rect 12159 26333 12171 26367
rect 12205 26364 12217 26367
rect 12250 26364 12256 26376
rect 12205 26336 12256 26364
rect 12205 26333 12217 26336
rect 12159 26327 12217 26333
rect 10744 26268 11284 26296
rect 10744 26256 10750 26268
rect 11514 26256 11520 26308
rect 11572 26296 11578 26308
rect 11900 26296 11928 26327
rect 12250 26324 12256 26336
rect 12308 26324 12314 26376
rect 14108 26296 14136 26404
rect 14550 26392 14556 26404
rect 14608 26392 14614 26444
rect 16209 26435 16267 26441
rect 16209 26432 16221 26435
rect 15212 26404 16221 26432
rect 15212 26376 15240 26404
rect 16209 26401 16221 26404
rect 16255 26432 16267 26435
rect 16298 26432 16304 26444
rect 16255 26404 16304 26432
rect 16255 26401 16267 26404
rect 16209 26395 16267 26401
rect 16298 26392 16304 26404
rect 16356 26392 16362 26444
rect 16666 26392 16672 26444
rect 16724 26392 16730 26444
rect 17402 26432 17408 26444
rect 17144 26404 17408 26432
rect 17144 26398 17172 26404
rect 14182 26324 14188 26376
rect 14240 26364 14246 26376
rect 14240 26337 14872 26364
rect 14240 26336 14823 26337
rect 14240 26324 14246 26336
rect 14811 26303 14823 26336
rect 14857 26306 14872 26337
rect 15194 26324 15200 26376
rect 15252 26324 15258 26376
rect 15286 26324 15292 26376
rect 15344 26364 15350 26376
rect 16025 26367 16083 26373
rect 16025 26364 16037 26367
rect 15344 26336 16037 26364
rect 15344 26324 15350 26336
rect 16025 26333 16037 26336
rect 16071 26333 16083 26367
rect 16025 26327 16083 26333
rect 14857 26303 14869 26306
rect 14811 26297 14869 26303
rect 11572 26268 14136 26296
rect 11572 26256 11578 26268
rect 8260 26200 9720 26228
rect 8260 26188 8266 26200
rect 10870 26188 10876 26240
rect 10928 26188 10934 26240
rect 12897 26231 12955 26237
rect 12897 26197 12909 26231
rect 12943 26228 12955 26231
rect 13078 26228 13084 26240
rect 12943 26200 13084 26228
rect 12943 26197 12955 26200
rect 12897 26191 12955 26197
rect 13078 26188 13084 26200
rect 13136 26188 13142 26240
rect 13814 26188 13820 26240
rect 13872 26228 13878 26240
rect 14182 26228 14188 26240
rect 13872 26200 14188 26228
rect 13872 26188 13878 26200
rect 14182 26188 14188 26200
rect 14240 26188 14246 26240
rect 15470 26188 15476 26240
rect 15528 26228 15534 26240
rect 15565 26231 15623 26237
rect 15565 26228 15577 26231
rect 15528 26200 15577 26228
rect 15528 26188 15534 26200
rect 15565 26197 15577 26200
rect 15611 26197 15623 26231
rect 16040 26228 16068 26327
rect 16942 26324 16948 26376
rect 17000 26373 17006 26376
rect 17077 26373 17172 26398
rect 17402 26392 17408 26404
rect 17460 26392 17466 26444
rect 17954 26392 17960 26444
rect 18012 26392 18018 26444
rect 19521 26435 19579 26441
rect 19521 26401 19533 26435
rect 19567 26432 19579 26435
rect 19889 26435 19947 26441
rect 19889 26432 19901 26435
rect 19567 26404 19901 26432
rect 19567 26401 19579 26404
rect 19521 26395 19579 26401
rect 19889 26401 19901 26404
rect 19935 26401 19947 26435
rect 19889 26395 19947 26401
rect 20073 26435 20131 26441
rect 20073 26401 20085 26435
rect 20119 26432 20131 26435
rect 20162 26432 20168 26444
rect 20119 26404 20168 26432
rect 20119 26401 20131 26404
rect 20073 26395 20131 26401
rect 20162 26392 20168 26404
rect 20220 26392 20226 26444
rect 20272 26441 20300 26472
rect 21637 26469 21649 26503
rect 21683 26469 21695 26503
rect 21637 26463 21695 26469
rect 21729 26503 21787 26509
rect 21729 26469 21741 26503
rect 21775 26500 21787 26503
rect 22370 26500 22376 26512
rect 21775 26472 22376 26500
rect 21775 26469 21787 26472
rect 21729 26463 21787 26469
rect 20257 26435 20315 26441
rect 20257 26401 20269 26435
rect 20303 26401 20315 26435
rect 20257 26395 20315 26401
rect 17000 26367 17021 26373
rect 17009 26333 17021 26367
rect 17000 26327 17021 26333
rect 17062 26370 17172 26373
rect 17062 26367 17120 26370
rect 17062 26333 17074 26367
rect 17108 26333 17120 26367
rect 17062 26327 17120 26333
rect 17000 26324 17006 26327
rect 17218 26324 17224 26376
rect 17276 26324 17282 26376
rect 17865 26367 17923 26373
rect 17865 26333 17877 26367
rect 17911 26364 17923 26367
rect 18414 26364 18420 26376
rect 17911 26336 18420 26364
rect 17911 26333 17923 26336
rect 17865 26327 17923 26333
rect 18414 26324 18420 26336
rect 18472 26364 18478 26376
rect 18969 26367 19027 26373
rect 18969 26364 18981 26367
rect 18472 26336 18981 26364
rect 18472 26324 18478 26336
rect 18969 26333 18981 26336
rect 19015 26333 19027 26367
rect 18969 26327 19027 26333
rect 19429 26367 19487 26373
rect 19429 26333 19441 26367
rect 19475 26333 19487 26367
rect 19429 26327 19487 26333
rect 19444 26296 19472 26327
rect 19794 26324 19800 26376
rect 19852 26324 19858 26376
rect 20524 26367 20582 26373
rect 20524 26364 20536 26367
rect 20456 26336 20536 26364
rect 20456 26308 20484 26336
rect 20524 26333 20536 26336
rect 20570 26333 20582 26367
rect 21652 26364 21680 26463
rect 22370 26460 22376 26472
rect 22428 26460 22434 26512
rect 21913 26367 21971 26373
rect 21913 26364 21925 26367
rect 21652 26336 21925 26364
rect 20524 26327 20582 26333
rect 21913 26333 21925 26336
rect 21959 26333 21971 26367
rect 21913 26327 21971 26333
rect 22002 26324 22008 26376
rect 22060 26364 22066 26376
rect 23845 26367 23903 26373
rect 23845 26364 23857 26367
rect 22060 26336 23857 26364
rect 22060 26324 22066 26336
rect 23845 26333 23857 26336
rect 23891 26333 23903 26367
rect 23845 26327 23903 26333
rect 18800 26268 19472 26296
rect 20073 26299 20131 26305
rect 17678 26228 17684 26240
rect 16040 26200 17684 26228
rect 15565 26191 15623 26197
rect 17678 26188 17684 26200
rect 17736 26188 17742 26240
rect 18800 26237 18828 26268
rect 20073 26265 20085 26299
rect 20119 26296 20131 26299
rect 20119 26268 20392 26296
rect 20119 26265 20131 26268
rect 20073 26259 20131 26265
rect 18785 26231 18843 26237
rect 18785 26197 18797 26231
rect 18831 26197 18843 26231
rect 20364 26228 20392 26268
rect 20438 26256 20444 26308
rect 20496 26256 20502 26308
rect 24118 26296 24124 26308
rect 20640 26268 24124 26296
rect 20640 26228 20668 26268
rect 24118 26256 24124 26268
rect 24176 26256 24182 26308
rect 24213 26299 24271 26305
rect 24213 26265 24225 26299
rect 24259 26296 24271 26299
rect 24854 26296 24860 26308
rect 24259 26268 24860 26296
rect 24259 26265 24271 26268
rect 24213 26259 24271 26265
rect 24854 26256 24860 26268
rect 24912 26256 24918 26308
rect 20364 26200 20668 26228
rect 18785 26191 18843 26197
rect 1104 26138 24723 26160
rect 1104 26086 6814 26138
rect 6866 26086 6878 26138
rect 6930 26086 6942 26138
rect 6994 26086 7006 26138
rect 7058 26086 7070 26138
rect 7122 26086 12679 26138
rect 12731 26086 12743 26138
rect 12795 26086 12807 26138
rect 12859 26086 12871 26138
rect 12923 26086 12935 26138
rect 12987 26086 18544 26138
rect 18596 26086 18608 26138
rect 18660 26086 18672 26138
rect 18724 26086 18736 26138
rect 18788 26086 18800 26138
rect 18852 26086 24409 26138
rect 24461 26086 24473 26138
rect 24525 26086 24537 26138
rect 24589 26086 24601 26138
rect 24653 26086 24665 26138
rect 24717 26086 24723 26138
rect 1104 26064 24723 26086
rect 1854 25984 1860 26036
rect 1912 26024 1918 26036
rect 2498 26024 2504 26036
rect 1912 25996 2504 26024
rect 1912 25984 1918 25996
rect 2498 25984 2504 25996
rect 2556 25984 2562 26036
rect 2961 26027 3019 26033
rect 2961 25993 2973 26027
rect 3007 25993 3019 26027
rect 2961 25987 3019 25993
rect 4157 26027 4215 26033
rect 4157 25993 4169 26027
rect 4203 26024 4215 26027
rect 4430 26024 4436 26036
rect 4203 25996 4436 26024
rect 4203 25993 4215 25996
rect 4157 25987 4215 25993
rect 842 25916 848 25968
rect 900 25956 906 25968
rect 2976 25956 3004 25987
rect 4430 25984 4436 25996
rect 4488 25984 4494 26036
rect 4908 25996 6224 26024
rect 4908 25956 4936 25996
rect 900 25928 2820 25956
rect 2976 25928 4936 25956
rect 6196 25956 6224 25996
rect 6270 25984 6276 26036
rect 6328 26024 6334 26036
rect 9030 26024 9036 26036
rect 6328 25996 9036 26024
rect 6328 25984 6334 25996
rect 9030 25984 9036 25996
rect 9088 25984 9094 26036
rect 9674 25984 9680 26036
rect 9732 26024 9738 26036
rect 10318 26024 10324 26036
rect 9732 25996 10324 26024
rect 9732 25984 9738 25996
rect 10318 25984 10324 25996
rect 10376 25984 10382 26036
rect 10686 25984 10692 26036
rect 10744 25984 10750 26036
rect 11057 26027 11115 26033
rect 11057 25993 11069 26027
rect 11103 26024 11115 26027
rect 11422 26024 11428 26036
rect 11103 25996 11428 26024
rect 11103 25993 11115 25996
rect 11057 25987 11115 25993
rect 11422 25984 11428 25996
rect 11480 25984 11486 26036
rect 11606 25984 11612 26036
rect 11664 26024 11670 26036
rect 13814 26024 13820 26036
rect 11664 25996 13820 26024
rect 11664 25984 11670 25996
rect 13814 25984 13820 25996
rect 13872 25984 13878 26036
rect 15194 26024 15200 26036
rect 14108 25996 15200 26024
rect 14108 25956 14136 25996
rect 15194 25984 15200 25996
rect 15252 25984 15258 26036
rect 16482 25984 16488 26036
rect 16540 26024 16546 26036
rect 16666 26024 16672 26036
rect 16540 25996 16672 26024
rect 16540 25984 16546 25996
rect 16666 25984 16672 25996
rect 16724 25984 16730 26036
rect 17218 25984 17224 26036
rect 17276 26024 17282 26036
rect 17681 26027 17739 26033
rect 17681 26024 17693 26027
rect 17276 25996 17693 26024
rect 17276 25984 17282 25996
rect 17681 25993 17693 25996
rect 17727 25993 17739 26027
rect 17681 25987 17739 25993
rect 19705 26027 19763 26033
rect 19705 25993 19717 26027
rect 19751 25993 19763 26027
rect 19705 25987 19763 25993
rect 19889 26027 19947 26033
rect 19889 25993 19901 26027
rect 19935 26024 19947 26027
rect 20530 26024 20536 26036
rect 19935 25996 20536 26024
rect 19935 25993 19947 25996
rect 19889 25987 19947 25993
rect 14458 25956 14464 25968
rect 6196 25928 14136 25956
rect 14200 25928 14464 25956
rect 900 25916 906 25928
rect 1671 25891 1729 25897
rect 1671 25857 1683 25891
rect 1717 25888 1729 25891
rect 2406 25888 2412 25900
rect 1717 25860 2412 25888
rect 1717 25857 1729 25860
rect 1671 25851 1729 25857
rect 2406 25848 2412 25860
rect 2464 25848 2470 25900
rect 2792 25897 2820 25928
rect 5151 25921 5209 25927
rect 2777 25891 2835 25897
rect 2777 25857 2789 25891
rect 2823 25857 2835 25891
rect 3387 25891 3445 25897
rect 3387 25888 3399 25891
rect 2777 25851 2835 25857
rect 3068 25860 3399 25888
rect 1210 25780 1216 25832
rect 1268 25820 1274 25832
rect 1397 25823 1455 25829
rect 1397 25820 1409 25823
rect 1268 25792 1409 25820
rect 1268 25780 1274 25792
rect 1397 25789 1409 25792
rect 1443 25789 1455 25823
rect 3068 25820 3096 25860
rect 3387 25857 3399 25860
rect 3433 25888 3445 25891
rect 4154 25888 4160 25900
rect 3433 25860 4160 25888
rect 3433 25857 3445 25860
rect 3387 25851 3445 25857
rect 4154 25848 4160 25860
rect 4212 25848 4218 25900
rect 5151 25887 5163 25921
rect 5197 25918 5209 25921
rect 5197 25900 5212 25918
rect 5151 25881 5172 25887
rect 5166 25848 5172 25881
rect 5224 25848 5230 25900
rect 7374 25848 7380 25900
rect 7432 25888 7438 25900
rect 8938 25888 8944 25900
rect 7432 25860 8944 25888
rect 7432 25848 7438 25860
rect 8938 25848 8944 25860
rect 8996 25848 9002 25900
rect 9858 25848 9864 25900
rect 9916 25888 9922 25900
rect 9951 25891 10009 25897
rect 9951 25888 9963 25891
rect 9916 25860 9963 25888
rect 9916 25848 9922 25860
rect 9951 25857 9963 25860
rect 9997 25888 10009 25891
rect 10318 25888 10324 25900
rect 9997 25860 10324 25888
rect 9997 25857 10009 25860
rect 9951 25851 10009 25857
rect 10318 25848 10324 25860
rect 10376 25848 10382 25900
rect 10870 25848 10876 25900
rect 10928 25888 10934 25900
rect 11241 25891 11299 25897
rect 11241 25888 11253 25891
rect 10928 25860 11253 25888
rect 10928 25848 10934 25860
rect 11241 25857 11253 25860
rect 11287 25857 11299 25891
rect 11241 25851 11299 25857
rect 11514 25848 11520 25900
rect 11572 25848 11578 25900
rect 11698 25848 11704 25900
rect 11756 25888 11762 25900
rect 11791 25891 11849 25897
rect 11791 25888 11803 25891
rect 11756 25860 11803 25888
rect 11756 25848 11762 25860
rect 11791 25857 11803 25860
rect 11837 25888 11849 25891
rect 12342 25888 12348 25900
rect 11837 25860 12348 25888
rect 11837 25857 11849 25860
rect 11791 25851 11849 25857
rect 12342 25848 12348 25860
rect 12400 25848 12406 25900
rect 13814 25848 13820 25900
rect 13872 25888 13878 25900
rect 14200 25897 14228 25928
rect 14458 25916 14464 25928
rect 14516 25956 14522 25968
rect 14734 25956 14740 25968
rect 14516 25928 14740 25956
rect 14516 25916 14522 25928
rect 14734 25916 14740 25928
rect 14792 25916 14798 25968
rect 14826 25916 14832 25968
rect 14884 25956 14890 25968
rect 14884 25928 16618 25956
rect 14884 25916 14890 25928
rect 13909 25891 13967 25897
rect 13909 25888 13921 25891
rect 13872 25860 13921 25888
rect 13872 25848 13878 25860
rect 13909 25857 13921 25860
rect 13955 25857 13967 25891
rect 13909 25851 13967 25857
rect 14183 25891 14241 25897
rect 14183 25857 14195 25891
rect 14229 25857 14241 25891
rect 14183 25851 14241 25857
rect 14550 25848 14556 25900
rect 14608 25888 14614 25900
rect 16590 25888 16618 25928
rect 18414 25916 18420 25968
rect 18472 25956 18478 25968
rect 18570 25959 18628 25965
rect 18570 25956 18582 25959
rect 18472 25928 18582 25956
rect 18472 25916 18478 25928
rect 18570 25925 18582 25928
rect 18616 25925 18628 25959
rect 18570 25919 18628 25925
rect 16911 25891 16969 25897
rect 16911 25888 16923 25891
rect 14608 25860 16528 25888
rect 16590 25860 16923 25888
rect 14608 25848 14614 25860
rect 16500 25832 16528 25860
rect 16911 25857 16923 25860
rect 16957 25888 16969 25891
rect 17218 25888 17224 25910
rect 16957 25860 17224 25888
rect 16957 25857 16969 25860
rect 17218 25858 17224 25860
rect 17276 25858 17282 25910
rect 16911 25851 16969 25857
rect 17954 25848 17960 25900
rect 18012 25888 18018 25900
rect 18325 25891 18383 25897
rect 18325 25888 18337 25891
rect 18012 25860 18337 25888
rect 18012 25848 18018 25860
rect 18325 25857 18337 25860
rect 18371 25857 18383 25891
rect 19720 25888 19748 25987
rect 20530 25984 20536 25996
rect 20588 25984 20594 26036
rect 21818 25984 21824 26036
rect 21876 25984 21882 26036
rect 21836 25956 21864 25984
rect 24026 25956 24032 25968
rect 21836 25928 22876 25956
rect 20073 25891 20131 25897
rect 20073 25888 20085 25891
rect 18325 25851 18383 25857
rect 18423 25860 19656 25888
rect 19720 25860 20085 25888
rect 1397 25783 1455 25789
rect 2792 25792 3096 25820
rect 3145 25823 3203 25829
rect 2792 25696 2820 25792
rect 3145 25789 3157 25823
rect 3191 25789 3203 25823
rect 3145 25783 3203 25789
rect 2406 25644 2412 25696
rect 2464 25644 2470 25696
rect 2774 25644 2780 25696
rect 2832 25644 2838 25696
rect 3160 25684 3188 25783
rect 4890 25780 4896 25832
rect 4948 25780 4954 25832
rect 9306 25780 9312 25832
rect 9364 25820 9370 25832
rect 9490 25820 9496 25832
rect 9364 25792 9496 25820
rect 9364 25780 9370 25792
rect 9490 25780 9496 25792
rect 9548 25780 9554 25832
rect 9582 25780 9588 25832
rect 9640 25820 9646 25832
rect 9677 25823 9735 25829
rect 9677 25820 9689 25823
rect 9640 25792 9689 25820
rect 9640 25780 9646 25792
rect 9677 25789 9689 25792
rect 9723 25789 9735 25823
rect 9677 25783 9735 25789
rect 16482 25780 16488 25832
rect 16540 25820 16546 25832
rect 16669 25823 16727 25829
rect 16669 25820 16681 25823
rect 16540 25792 16681 25820
rect 16540 25780 16546 25792
rect 16669 25789 16681 25792
rect 16715 25789 16727 25823
rect 18423 25820 18451 25860
rect 16669 25783 16727 25789
rect 17604 25792 18451 25820
rect 19628 25820 19656 25860
rect 20073 25857 20085 25860
rect 20119 25857 20131 25891
rect 20591 25891 20649 25897
rect 20591 25888 20603 25891
rect 20073 25851 20131 25857
rect 20180 25860 20603 25888
rect 20180 25820 20208 25860
rect 20591 25857 20603 25860
rect 20637 25857 20649 25891
rect 21821 25891 21879 25897
rect 21821 25888 21833 25891
rect 20591 25851 20649 25857
rect 21376 25860 21833 25888
rect 19628 25792 20208 25820
rect 20349 25823 20407 25829
rect 17604 25764 17632 25792
rect 20349 25789 20361 25823
rect 20395 25789 20407 25823
rect 20349 25783 20407 25789
rect 5552 25724 6040 25752
rect 3510 25684 3516 25696
rect 3160 25656 3516 25684
rect 3510 25644 3516 25656
rect 3568 25644 3574 25696
rect 3602 25644 3608 25696
rect 3660 25684 3666 25696
rect 5552 25684 5580 25724
rect 3660 25656 5580 25684
rect 3660 25644 3666 25656
rect 5902 25644 5908 25696
rect 5960 25644 5966 25696
rect 6012 25684 6040 25724
rect 6086 25712 6092 25764
rect 6144 25752 6150 25764
rect 6822 25752 6828 25764
rect 6144 25724 6828 25752
rect 6144 25712 6150 25724
rect 6822 25712 6828 25724
rect 6880 25712 6886 25764
rect 13814 25752 13820 25764
rect 12452 25724 13820 25752
rect 12452 25684 12480 25724
rect 13814 25712 13820 25724
rect 13872 25712 13878 25764
rect 14642 25712 14648 25764
rect 14700 25752 14706 25764
rect 14700 25724 15056 25752
rect 14700 25712 14706 25724
rect 6012 25656 12480 25684
rect 12526 25644 12532 25696
rect 12584 25644 12590 25696
rect 14826 25644 14832 25696
rect 14884 25684 14890 25696
rect 14921 25687 14979 25693
rect 14921 25684 14933 25687
rect 14884 25656 14933 25684
rect 14884 25644 14890 25656
rect 14921 25653 14933 25656
rect 14967 25653 14979 25687
rect 15028 25684 15056 25724
rect 17586 25712 17592 25764
rect 17644 25712 17650 25764
rect 19334 25712 19340 25764
rect 19392 25752 19398 25764
rect 20070 25752 20076 25764
rect 19392 25724 20076 25752
rect 19392 25712 19398 25724
rect 20070 25712 20076 25724
rect 20128 25752 20134 25764
rect 20364 25752 20392 25783
rect 21376 25761 21404 25860
rect 21821 25857 21833 25860
rect 21867 25888 21879 25891
rect 22189 25891 22247 25897
rect 22189 25888 22201 25891
rect 21867 25860 22201 25888
rect 21867 25857 21879 25860
rect 21821 25851 21879 25857
rect 22189 25857 22201 25860
rect 22235 25857 22247 25891
rect 22189 25851 22247 25857
rect 22370 25848 22376 25900
rect 22428 25848 22434 25900
rect 22848 25897 22876 25928
rect 23492 25928 24032 25956
rect 23492 25897 23520 25928
rect 24026 25916 24032 25928
rect 24084 25916 24090 25968
rect 22833 25891 22891 25897
rect 22833 25857 22845 25891
rect 22879 25857 22891 25891
rect 22833 25851 22891 25857
rect 23293 25891 23351 25897
rect 23293 25857 23305 25891
rect 23339 25857 23351 25891
rect 23293 25851 23351 25857
rect 23477 25891 23535 25897
rect 23477 25857 23489 25891
rect 23523 25857 23535 25891
rect 23477 25851 23535 25857
rect 22097 25823 22155 25829
rect 22097 25789 22109 25823
rect 22143 25820 22155 25823
rect 22281 25823 22339 25829
rect 22281 25820 22293 25823
rect 22143 25792 22293 25820
rect 22143 25789 22155 25792
rect 22097 25783 22155 25789
rect 22281 25789 22293 25792
rect 22327 25789 22339 25823
rect 23308 25820 23336 25851
rect 23566 25848 23572 25900
rect 23624 25848 23630 25900
rect 23750 25848 23756 25900
rect 23808 25888 23814 25900
rect 23937 25891 23995 25897
rect 23937 25888 23949 25891
rect 23808 25860 23949 25888
rect 23808 25848 23814 25860
rect 23937 25857 23949 25860
rect 23983 25857 23995 25891
rect 23937 25851 23995 25857
rect 23658 25820 23664 25832
rect 23308 25792 23664 25820
rect 22281 25783 22339 25789
rect 23658 25780 23664 25792
rect 23716 25780 23722 25832
rect 20128 25724 20392 25752
rect 21361 25755 21419 25761
rect 20128 25712 20134 25724
rect 21361 25721 21373 25755
rect 21407 25721 21419 25755
rect 21361 25715 21419 25721
rect 22005 25755 22063 25761
rect 22005 25721 22017 25755
rect 22051 25752 22063 25755
rect 23934 25752 23940 25764
rect 22051 25724 23940 25752
rect 22051 25721 22063 25724
rect 22005 25715 22063 25721
rect 23934 25712 23940 25724
rect 23992 25712 23998 25764
rect 21818 25684 21824 25696
rect 15028 25656 21824 25684
rect 14921 25647 14979 25653
rect 21818 25644 21824 25656
rect 21876 25644 21882 25696
rect 21910 25644 21916 25696
rect 21968 25644 21974 25696
rect 22646 25644 22652 25696
rect 22704 25644 22710 25696
rect 23382 25644 23388 25696
rect 23440 25644 23446 25696
rect 23750 25644 23756 25696
rect 23808 25644 23814 25696
rect 24121 25687 24179 25693
rect 24121 25653 24133 25687
rect 24167 25684 24179 25687
rect 24854 25684 24860 25696
rect 24167 25656 24860 25684
rect 24167 25653 24179 25656
rect 24121 25647 24179 25653
rect 24854 25644 24860 25656
rect 24912 25644 24918 25696
rect 1104 25594 24564 25616
rect 1104 25542 3882 25594
rect 3934 25542 3946 25594
rect 3998 25542 4010 25594
rect 4062 25542 4074 25594
rect 4126 25542 4138 25594
rect 4190 25542 9747 25594
rect 9799 25542 9811 25594
rect 9863 25542 9875 25594
rect 9927 25542 9939 25594
rect 9991 25542 10003 25594
rect 10055 25542 15612 25594
rect 15664 25542 15676 25594
rect 15728 25542 15740 25594
rect 15792 25542 15804 25594
rect 15856 25542 15868 25594
rect 15920 25542 21477 25594
rect 21529 25542 21541 25594
rect 21593 25542 21605 25594
rect 21657 25542 21669 25594
rect 21721 25542 21733 25594
rect 21785 25542 24564 25594
rect 1104 25520 24564 25542
rect 3326 25440 3332 25492
rect 3384 25480 3390 25492
rect 10781 25483 10839 25489
rect 3384 25452 10732 25480
rect 3384 25440 3390 25452
rect 6546 25372 6552 25424
rect 6604 25372 6610 25424
rect 10704 25412 10732 25452
rect 10781 25449 10793 25483
rect 10827 25480 10839 25483
rect 10962 25480 10968 25492
rect 10827 25452 10968 25480
rect 10827 25449 10839 25452
rect 10781 25443 10839 25449
rect 10962 25440 10968 25452
rect 11020 25440 11026 25492
rect 12526 25480 12532 25492
rect 12176 25452 12532 25480
rect 12066 25412 12072 25424
rect 10704 25384 12072 25412
rect 12066 25372 12072 25384
rect 12124 25372 12130 25424
rect 12176 25421 12204 25452
rect 12526 25440 12532 25452
rect 12584 25440 12590 25492
rect 13357 25483 13415 25489
rect 13357 25449 13369 25483
rect 13403 25480 13415 25483
rect 14642 25480 14648 25492
rect 13403 25452 14648 25480
rect 13403 25449 13415 25452
rect 13357 25443 13415 25449
rect 14642 25440 14648 25452
rect 14700 25440 14706 25492
rect 15102 25480 15108 25492
rect 14752 25452 15108 25480
rect 14752 25421 14780 25452
rect 15102 25440 15108 25452
rect 15160 25440 15166 25492
rect 16482 25480 16488 25492
rect 16040 25452 16488 25480
rect 12161 25415 12219 25421
rect 12161 25381 12173 25415
rect 12207 25381 12219 25415
rect 12161 25375 12219 25381
rect 14737 25415 14795 25421
rect 14737 25381 14749 25415
rect 14783 25381 14795 25415
rect 14737 25375 14795 25381
rect 2406 25304 2412 25356
rect 2464 25304 2470 25356
rect 6564 25344 6592 25372
rect 6288 25316 6592 25344
rect 1302 25236 1308 25288
rect 1360 25276 1366 25288
rect 3053 25279 3111 25285
rect 3053 25276 3065 25279
rect 1360 25248 3065 25276
rect 1360 25236 1366 25248
rect 3053 25245 3065 25248
rect 3099 25245 3111 25279
rect 3053 25239 3111 25245
rect 4890 25236 4896 25288
rect 4948 25276 4954 25288
rect 5442 25276 5448 25288
rect 4948 25248 5448 25276
rect 4948 25236 4954 25248
rect 5442 25236 5448 25248
rect 5500 25276 5506 25288
rect 5629 25279 5687 25285
rect 5629 25276 5641 25279
rect 5500 25248 5641 25276
rect 5500 25236 5506 25248
rect 5629 25245 5641 25248
rect 5675 25245 5687 25279
rect 5629 25239 5687 25245
rect 5903 25279 5961 25285
rect 5903 25245 5915 25279
rect 5949 25276 5961 25279
rect 6288 25276 6316 25316
rect 6822 25304 6828 25356
rect 6880 25344 6886 25356
rect 8938 25344 8944 25356
rect 6880 25316 8944 25344
rect 6880 25304 6886 25316
rect 8938 25304 8944 25316
rect 8996 25304 9002 25356
rect 9950 25304 9956 25356
rect 10008 25344 10014 25356
rect 11330 25344 11336 25356
rect 10008 25316 11336 25344
rect 10008 25304 10014 25316
rect 11330 25304 11336 25316
rect 11388 25304 11394 25356
rect 11514 25344 11520 25356
rect 11440 25316 11520 25344
rect 5949 25248 6316 25276
rect 5949 25245 5961 25248
rect 5903 25239 5961 25245
rect 6362 25236 6368 25288
rect 6420 25276 6426 25288
rect 7374 25276 7380 25288
rect 6420 25248 7380 25276
rect 6420 25236 6426 25248
rect 7374 25236 7380 25248
rect 7432 25236 7438 25288
rect 8294 25236 8300 25288
rect 8352 25276 8358 25288
rect 10686 25276 10692 25288
rect 8352 25248 10692 25276
rect 8352 25236 8358 25248
rect 10686 25236 10692 25248
rect 10744 25236 10750 25288
rect 10962 25236 10968 25288
rect 11020 25236 11026 25288
rect 11440 25276 11468 25316
rect 11514 25304 11520 25316
rect 11572 25304 11578 25356
rect 12250 25304 12256 25356
rect 12308 25344 12314 25356
rect 12437 25347 12495 25353
rect 12437 25344 12449 25347
rect 12308 25316 12449 25344
rect 12308 25304 12314 25316
rect 12437 25313 12449 25316
rect 12483 25313 12495 25347
rect 12437 25307 12495 25313
rect 12526 25304 12532 25356
rect 12584 25353 12590 25356
rect 12584 25347 12612 25353
rect 12600 25313 12612 25347
rect 12584 25307 12612 25313
rect 12713 25347 12771 25353
rect 12713 25313 12725 25347
rect 12759 25344 12771 25347
rect 13078 25344 13084 25356
rect 12759 25316 13084 25344
rect 12759 25313 12771 25316
rect 12713 25307 12771 25313
rect 12584 25304 12590 25307
rect 13078 25304 13084 25316
rect 13136 25304 13142 25356
rect 14277 25347 14335 25353
rect 14277 25344 14289 25347
rect 13832 25316 14289 25344
rect 13832 25288 13860 25316
rect 14277 25313 14289 25316
rect 14323 25313 14335 25347
rect 14277 25307 14335 25313
rect 15289 25347 15347 25353
rect 15289 25313 15301 25347
rect 15335 25344 15347 25347
rect 15470 25344 15476 25356
rect 15335 25316 15476 25344
rect 15335 25313 15347 25316
rect 15289 25307 15347 25313
rect 15470 25304 15476 25316
rect 15528 25304 15534 25356
rect 15838 25304 15844 25356
rect 15896 25344 15902 25356
rect 16040 25353 16068 25452
rect 16482 25440 16488 25452
rect 16540 25440 16546 25492
rect 16758 25440 16764 25492
rect 16816 25480 16822 25492
rect 17037 25483 17095 25489
rect 17037 25480 17049 25483
rect 16816 25452 17049 25480
rect 16816 25440 16822 25452
rect 17037 25449 17049 25452
rect 17083 25449 17095 25483
rect 17037 25443 17095 25449
rect 21361 25483 21419 25489
rect 21361 25449 21373 25483
rect 21407 25480 21419 25483
rect 21910 25480 21916 25492
rect 21407 25452 21916 25480
rect 21407 25449 21419 25452
rect 21361 25443 21419 25449
rect 21910 25440 21916 25452
rect 21968 25440 21974 25492
rect 23382 25440 23388 25492
rect 23440 25440 23446 25492
rect 16942 25372 16948 25424
rect 17000 25412 17006 25424
rect 17402 25412 17408 25424
rect 17000 25384 17408 25412
rect 17000 25372 17006 25384
rect 17402 25372 17408 25384
rect 17460 25372 17466 25424
rect 16025 25347 16083 25353
rect 16025 25344 16037 25347
rect 15896 25316 16037 25344
rect 15896 25304 15902 25316
rect 16025 25313 16037 25316
rect 16071 25313 16083 25347
rect 23400 25344 23428 25440
rect 23753 25415 23811 25421
rect 23753 25381 23765 25415
rect 23799 25412 23811 25415
rect 24121 25415 24179 25421
rect 24121 25412 24133 25415
rect 23799 25384 24133 25412
rect 23799 25381 23811 25384
rect 23753 25375 23811 25381
rect 24121 25381 24133 25384
rect 24167 25381 24179 25415
rect 24121 25375 24179 25381
rect 23937 25347 23995 25353
rect 23937 25344 23949 25347
rect 23400 25316 23949 25344
rect 16025 25307 16083 25313
rect 23937 25313 23949 25316
rect 23983 25313 23995 25347
rect 23937 25307 23995 25313
rect 11070 25248 11468 25276
rect 1578 25168 1584 25220
rect 1636 25168 1642 25220
rect 1854 25168 1860 25220
rect 1912 25168 1918 25220
rect 1946 25168 1952 25220
rect 2004 25168 2010 25220
rect 2314 25168 2320 25220
rect 2372 25168 2378 25220
rect 2685 25211 2743 25217
rect 2685 25177 2697 25211
rect 2731 25208 2743 25211
rect 2958 25208 2964 25220
rect 2731 25180 2964 25208
rect 2731 25177 2743 25180
rect 2685 25171 2743 25177
rect 2958 25168 2964 25180
rect 3016 25168 3022 25220
rect 11070 25208 11098 25248
rect 11698 25236 11704 25288
rect 11756 25236 11762 25288
rect 13814 25236 13820 25288
rect 13872 25236 13878 25288
rect 14093 25279 14151 25285
rect 14093 25276 14105 25279
rect 13924 25248 14105 25276
rect 3252 25180 11098 25208
rect 2866 25100 2872 25152
rect 2924 25100 2930 25152
rect 3252 25149 3280 25180
rect 3237 25143 3295 25149
rect 3237 25109 3249 25143
rect 3283 25109 3295 25143
rect 3237 25103 3295 25109
rect 4246 25100 4252 25152
rect 4304 25140 4310 25152
rect 5166 25140 5172 25152
rect 4304 25112 5172 25140
rect 4304 25100 4310 25112
rect 5166 25100 5172 25112
rect 5224 25100 5230 25152
rect 6641 25143 6699 25149
rect 6641 25109 6653 25143
rect 6687 25140 6699 25143
rect 7190 25140 7196 25152
rect 6687 25112 7196 25140
rect 6687 25109 6699 25112
rect 6641 25103 6699 25109
rect 7190 25100 7196 25112
rect 7248 25100 7254 25152
rect 8570 25100 8576 25152
rect 8628 25140 8634 25152
rect 13924 25140 13952 25248
rect 14093 25245 14105 25248
rect 14139 25245 14151 25279
rect 14093 25239 14151 25245
rect 15010 25236 15016 25288
rect 15068 25236 15074 25288
rect 15102 25236 15108 25288
rect 15160 25285 15166 25288
rect 15160 25279 15188 25285
rect 15176 25245 15188 25279
rect 15160 25239 15188 25245
rect 15160 25236 15166 25239
rect 15930 25236 15936 25288
rect 15988 25276 15994 25288
rect 16267 25279 16325 25285
rect 16267 25276 16279 25279
rect 15988 25248 16279 25276
rect 15988 25236 15994 25248
rect 16267 25245 16279 25248
rect 16313 25245 16325 25279
rect 16267 25239 16325 25245
rect 20714 25236 20720 25288
rect 20772 25276 20778 25288
rect 21269 25279 21327 25285
rect 21269 25276 21281 25279
rect 20772 25248 21281 25276
rect 20772 25236 20778 25248
rect 21269 25245 21281 25248
rect 21315 25245 21327 25279
rect 21269 25239 21327 25245
rect 21818 25236 21824 25288
rect 21876 25236 21882 25288
rect 22094 25236 22100 25288
rect 22152 25236 22158 25288
rect 22646 25236 22652 25288
rect 22704 25236 22710 25288
rect 23658 25236 23664 25288
rect 23716 25236 23722 25288
rect 24029 25279 24087 25285
rect 24029 25245 24041 25279
rect 24075 25245 24087 25279
rect 24029 25239 24087 25245
rect 15948 25208 15976 25236
rect 15746 25180 15976 25208
rect 21836 25208 21864 25236
rect 22342 25211 22400 25217
rect 22342 25208 22354 25211
rect 21836 25180 22354 25208
rect 13998 25140 14004 25152
rect 8628 25112 14004 25140
rect 8628 25100 8634 25112
rect 13998 25100 14004 25112
rect 14056 25140 14062 25152
rect 14642 25140 14648 25152
rect 14056 25112 14648 25140
rect 14056 25100 14062 25112
rect 14642 25100 14648 25112
rect 14700 25100 14706 25152
rect 15378 25100 15384 25152
rect 15436 25140 15442 25152
rect 15746 25140 15774 25180
rect 22342 25177 22354 25180
rect 22388 25177 22400 25211
rect 22664 25208 22692 25236
rect 24044 25208 24072 25239
rect 22664 25180 24072 25208
rect 22342 25171 22400 25177
rect 15436 25112 15774 25140
rect 15933 25143 15991 25149
rect 15436 25100 15442 25112
rect 15933 25109 15945 25143
rect 15979 25140 15991 25143
rect 17770 25140 17776 25152
rect 15979 25112 17776 25140
rect 15979 25109 15991 25112
rect 15933 25103 15991 25109
rect 17770 25100 17776 25112
rect 17828 25100 17834 25152
rect 20254 25100 20260 25152
rect 20312 25140 20318 25152
rect 20714 25140 20720 25152
rect 20312 25112 20720 25140
rect 20312 25100 20318 25112
rect 20714 25100 20720 25112
rect 20772 25100 20778 25152
rect 23474 25100 23480 25152
rect 23532 25100 23538 25152
rect 23658 25100 23664 25152
rect 23716 25140 23722 25152
rect 23937 25143 23995 25149
rect 23937 25140 23949 25143
rect 23716 25112 23949 25140
rect 23716 25100 23722 25112
rect 23937 25109 23949 25112
rect 23983 25109 23995 25143
rect 23937 25103 23995 25109
rect 1104 25050 24723 25072
rect 1104 24998 6814 25050
rect 6866 24998 6878 25050
rect 6930 24998 6942 25050
rect 6994 24998 7006 25050
rect 7058 24998 7070 25050
rect 7122 24998 12679 25050
rect 12731 24998 12743 25050
rect 12795 24998 12807 25050
rect 12859 24998 12871 25050
rect 12923 24998 12935 25050
rect 12987 24998 18544 25050
rect 18596 24998 18608 25050
rect 18660 24998 18672 25050
rect 18724 24998 18736 25050
rect 18788 24998 18800 25050
rect 18852 24998 24409 25050
rect 24461 24998 24473 25050
rect 24525 24998 24537 25050
rect 24589 24998 24601 25050
rect 24653 24998 24665 25050
rect 24717 24998 24723 25050
rect 1104 24976 24723 24998
rect 1946 24896 1952 24948
rect 2004 24936 2010 24948
rect 2685 24939 2743 24945
rect 2685 24936 2697 24939
rect 2004 24908 2697 24936
rect 2004 24896 2010 24908
rect 2685 24905 2697 24908
rect 2731 24905 2743 24939
rect 2685 24899 2743 24905
rect 3418 24896 3424 24948
rect 3476 24936 3482 24948
rect 6178 24936 6184 24948
rect 3476 24908 5304 24936
rect 3476 24896 3482 24908
rect 2774 24828 2780 24880
rect 2832 24868 2838 24880
rect 5074 24868 5080 24880
rect 2832 24840 5080 24868
rect 2832 24828 2838 24840
rect 5074 24828 5080 24840
rect 5132 24828 5138 24880
rect 842 24760 848 24812
rect 900 24800 906 24812
rect 1397 24803 1455 24809
rect 1397 24800 1409 24803
rect 900 24772 1409 24800
rect 900 24760 906 24772
rect 1397 24769 1409 24772
rect 1443 24769 1455 24803
rect 1397 24763 1455 24769
rect 1578 24760 1584 24812
rect 1636 24800 1642 24812
rect 1915 24803 1973 24809
rect 1915 24800 1927 24803
rect 1636 24772 1927 24800
rect 1636 24760 1642 24772
rect 1915 24769 1927 24772
rect 1961 24769 1973 24803
rect 1915 24763 1973 24769
rect 4063 24803 4121 24809
rect 4063 24769 4075 24803
rect 4109 24800 4121 24803
rect 5276 24800 5304 24908
rect 5368 24908 6184 24936
rect 5368 24880 5396 24908
rect 6178 24896 6184 24908
rect 6236 24936 6242 24948
rect 7098 24936 7104 24948
rect 6236 24908 7104 24936
rect 6236 24896 6242 24908
rect 7098 24896 7104 24908
rect 7156 24936 7162 24948
rect 7156 24908 7328 24936
rect 7156 24896 7162 24908
rect 5350 24828 5356 24880
rect 5408 24828 5414 24880
rect 6546 24828 6552 24880
rect 6604 24828 6610 24880
rect 7190 24828 7196 24880
rect 7248 24828 7254 24880
rect 7300 24877 7328 24908
rect 7466 24896 7472 24948
rect 7524 24936 7530 24948
rect 7650 24936 7656 24948
rect 7524 24908 7656 24936
rect 7524 24896 7530 24908
rect 7650 24896 7656 24908
rect 7708 24896 7714 24948
rect 8662 24896 8668 24948
rect 8720 24896 8726 24948
rect 14274 24936 14280 24948
rect 13556 24908 14280 24936
rect 7285 24871 7343 24877
rect 7285 24837 7297 24871
rect 7331 24837 7343 24871
rect 8680 24868 8708 24896
rect 7285 24831 7343 24837
rect 8036 24840 8708 24868
rect 6564 24800 6592 24828
rect 4109 24772 4476 24800
rect 5276 24772 6592 24800
rect 4109 24769 4121 24772
rect 4063 24763 4121 24769
rect 1210 24692 1216 24744
rect 1268 24732 1274 24744
rect 1673 24735 1731 24741
rect 1673 24732 1685 24735
rect 1268 24704 1685 24732
rect 1268 24692 1274 24704
rect 1673 24701 1685 24704
rect 1719 24701 1731 24735
rect 1673 24695 1731 24701
rect 1578 24624 1584 24676
rect 1636 24624 1642 24676
rect 1688 24596 1716 24695
rect 3786 24692 3792 24744
rect 3844 24692 3850 24744
rect 4448 24732 4476 24772
rect 6730 24760 6736 24812
rect 6788 24800 6794 24812
rect 6825 24803 6883 24809
rect 6825 24800 6837 24803
rect 6788 24772 6837 24800
rect 6788 24760 6794 24772
rect 6825 24769 6837 24772
rect 6871 24769 6883 24803
rect 6825 24763 6883 24769
rect 6917 24803 6975 24809
rect 6917 24769 6929 24803
rect 6963 24800 6975 24803
rect 7208 24800 7236 24828
rect 8036 24809 8064 24840
rect 9122 24828 9128 24880
rect 9180 24828 9186 24880
rect 9582 24828 9588 24880
rect 9640 24868 9646 24880
rect 11422 24868 11428 24880
rect 9640 24840 11428 24868
rect 9640 24828 9646 24840
rect 11422 24828 11428 24840
rect 11480 24868 11486 24880
rect 11882 24868 11888 24880
rect 11480 24840 11888 24868
rect 11480 24828 11486 24840
rect 11882 24828 11888 24840
rect 11940 24828 11946 24880
rect 12250 24828 12256 24880
rect 12308 24868 12314 24880
rect 13446 24868 13452 24880
rect 12308 24840 13452 24868
rect 12308 24828 12314 24840
rect 13446 24828 13452 24840
rect 13504 24828 13510 24880
rect 6963 24772 7236 24800
rect 8021 24803 8079 24809
rect 6963 24769 6975 24772
rect 6917 24763 6975 24769
rect 8021 24769 8033 24803
rect 8067 24769 8079 24803
rect 8021 24763 8079 24769
rect 8295 24803 8353 24809
rect 8295 24769 8307 24803
rect 8341 24800 8353 24803
rect 8662 24800 8668 24812
rect 8341 24772 8668 24800
rect 8341 24769 8353 24772
rect 8295 24763 8353 24769
rect 8662 24760 8668 24772
rect 8720 24800 8726 24812
rect 9140 24800 9168 24828
rect 8720 24772 9168 24800
rect 8720 24760 8726 24772
rect 4448 24704 5856 24732
rect 2038 24596 2044 24608
rect 1688 24568 2044 24596
rect 2038 24556 2044 24568
rect 2096 24596 2102 24608
rect 3804 24596 3832 24692
rect 5828 24664 5856 24704
rect 5902 24692 5908 24744
rect 5960 24732 5966 24744
rect 5960 24704 6394 24732
rect 5960 24692 5966 24704
rect 8754 24692 8760 24744
rect 8812 24732 8818 24744
rect 9600 24741 9628 24828
rect 9859 24803 9917 24809
rect 9859 24769 9871 24803
rect 9905 24800 9917 24803
rect 9950 24800 9956 24812
rect 9905 24772 9956 24800
rect 9905 24769 9917 24772
rect 9859 24763 9917 24769
rect 9950 24760 9956 24772
rect 10008 24760 10014 24812
rect 12527 24803 12585 24809
rect 12527 24800 12539 24803
rect 12084 24772 12539 24800
rect 9585 24735 9643 24741
rect 9585 24732 9597 24735
rect 8812 24704 9597 24732
rect 8812 24692 8818 24704
rect 9585 24701 9597 24704
rect 9631 24701 9643 24735
rect 9585 24695 9643 24701
rect 11606 24692 11612 24744
rect 11664 24692 11670 24744
rect 11974 24692 11980 24744
rect 12032 24732 12038 24744
rect 12084 24732 12112 24772
rect 12527 24769 12539 24772
rect 12573 24800 12585 24803
rect 13556 24800 13584 24908
rect 14274 24896 14280 24908
rect 14332 24896 14338 24948
rect 23474 24896 23480 24948
rect 23532 24896 23538 24948
rect 23566 24896 23572 24948
rect 23624 24936 23630 24948
rect 23661 24939 23719 24945
rect 23661 24936 23673 24939
rect 23624 24908 23673 24936
rect 23624 24896 23630 24908
rect 23661 24905 23673 24908
rect 23707 24905 23719 24939
rect 23661 24899 23719 24905
rect 24026 24896 24032 24948
rect 24084 24896 24090 24948
rect 13814 24828 13820 24880
rect 13872 24828 13878 24880
rect 17236 24840 17540 24868
rect 12573 24772 13584 24800
rect 13633 24803 13691 24809
rect 12573 24769 12585 24772
rect 12527 24763 12585 24769
rect 13633 24769 13645 24803
rect 13679 24800 13691 24803
rect 13832 24800 13860 24828
rect 13679 24772 13860 24800
rect 13679 24769 13691 24772
rect 13633 24763 13691 24769
rect 14642 24760 14648 24812
rect 14700 24809 14706 24812
rect 14700 24803 14728 24809
rect 14716 24769 14728 24803
rect 14700 24763 14728 24769
rect 14700 24760 14706 24763
rect 14826 24760 14832 24812
rect 14884 24760 14890 24812
rect 17129 24803 17187 24809
rect 17129 24769 17141 24803
rect 17175 24800 17187 24803
rect 17236 24800 17264 24840
rect 17402 24809 17408 24812
rect 17396 24800 17408 24809
rect 17175 24772 17264 24800
rect 17363 24772 17408 24800
rect 17175 24769 17187 24772
rect 17129 24763 17187 24769
rect 17396 24763 17408 24772
rect 17402 24760 17408 24763
rect 17460 24760 17466 24812
rect 17512 24800 17540 24840
rect 18248 24840 19472 24868
rect 17954 24800 17960 24812
rect 17512 24772 17960 24800
rect 17954 24760 17960 24772
rect 18012 24760 18018 24812
rect 12032 24704 12112 24732
rect 12253 24735 12311 24741
rect 12032 24692 12038 24704
rect 12253 24701 12265 24735
rect 12299 24701 12311 24735
rect 12253 24695 12311 24701
rect 13817 24735 13875 24741
rect 13817 24701 13829 24735
rect 13863 24732 13875 24735
rect 13906 24732 13912 24744
rect 13863 24704 13912 24732
rect 13863 24701 13875 24704
rect 13817 24695 13875 24701
rect 6270 24664 6276 24676
rect 5828 24636 6276 24664
rect 6270 24624 6276 24636
rect 6328 24624 6334 24676
rect 7834 24624 7840 24676
rect 7892 24624 7898 24676
rect 11624 24664 11652 24692
rect 12268 24664 12296 24695
rect 13906 24692 13912 24704
rect 13964 24692 13970 24744
rect 14550 24692 14556 24744
rect 14608 24732 14614 24744
rect 15010 24732 15016 24744
rect 14608 24704 15016 24732
rect 14608 24692 14614 24704
rect 15010 24692 15016 24704
rect 15068 24692 15074 24744
rect 10244 24636 10732 24664
rect 11624 24636 12296 24664
rect 13265 24667 13323 24673
rect 2096 24568 3832 24596
rect 2096 24556 2102 24568
rect 4798 24556 4804 24608
rect 4856 24556 4862 24608
rect 9030 24556 9036 24608
rect 9088 24556 9094 24608
rect 9306 24556 9312 24608
rect 9364 24596 9370 24608
rect 10244 24596 10272 24636
rect 9364 24568 10272 24596
rect 9364 24556 9370 24568
rect 10502 24556 10508 24608
rect 10560 24596 10566 24608
rect 10597 24599 10655 24605
rect 10597 24596 10609 24599
rect 10560 24568 10609 24596
rect 10560 24556 10566 24568
rect 10597 24565 10609 24568
rect 10643 24565 10655 24599
rect 10704 24596 10732 24636
rect 13265 24633 13277 24667
rect 13311 24664 13323 24667
rect 14277 24667 14335 24673
rect 14277 24664 14289 24667
rect 13311 24636 14289 24664
rect 13311 24633 13323 24636
rect 13265 24627 13323 24633
rect 14277 24633 14289 24636
rect 14323 24633 14335 24667
rect 14277 24627 14335 24633
rect 14182 24596 14188 24608
rect 10704 24568 14188 24596
rect 10597 24559 10655 24565
rect 14182 24556 14188 24568
rect 14240 24596 14246 24608
rect 14918 24596 14924 24608
rect 14240 24568 14924 24596
rect 14240 24556 14246 24568
rect 14918 24556 14924 24568
rect 14976 24556 14982 24608
rect 15473 24599 15531 24605
rect 15473 24565 15485 24599
rect 15519 24596 15531 24599
rect 18248 24596 18276 24840
rect 18601 24803 18659 24809
rect 18601 24769 18613 24803
rect 18647 24769 18659 24803
rect 19061 24803 19119 24809
rect 19061 24800 19073 24803
rect 18601 24763 18659 24769
rect 18800 24772 19073 24800
rect 18322 24692 18328 24744
rect 18380 24732 18386 24744
rect 18616 24732 18644 24763
rect 18380 24704 18644 24732
rect 18380 24692 18386 24704
rect 18509 24667 18567 24673
rect 18509 24633 18521 24667
rect 18555 24664 18567 24667
rect 18800 24664 18828 24772
rect 19061 24769 19073 24772
rect 19107 24769 19119 24803
rect 19061 24763 19119 24769
rect 19150 24760 19156 24812
rect 19208 24760 19214 24812
rect 19337 24803 19395 24809
rect 19337 24800 19349 24803
rect 19260 24772 19349 24800
rect 19260 24664 19288 24772
rect 19337 24769 19349 24772
rect 19383 24769 19395 24803
rect 19444 24800 19472 24840
rect 19518 24800 19524 24812
rect 19444 24772 19524 24800
rect 19337 24763 19395 24769
rect 19518 24760 19524 24772
rect 19576 24800 19582 24812
rect 19613 24803 19671 24809
rect 19613 24800 19625 24803
rect 19576 24772 19625 24800
rect 19576 24760 19582 24772
rect 19613 24769 19625 24772
rect 19659 24769 19671 24803
rect 19613 24763 19671 24769
rect 20073 24803 20131 24809
rect 20073 24769 20085 24803
rect 20119 24769 20131 24803
rect 20073 24763 20131 24769
rect 20088 24732 20116 24763
rect 21174 24760 21180 24812
rect 21232 24800 21238 24812
rect 22923 24803 22981 24809
rect 22923 24800 22935 24803
rect 21232 24772 22935 24800
rect 21232 24760 21238 24772
rect 22923 24769 22935 24772
rect 22969 24800 22981 24803
rect 23492 24800 23520 24896
rect 24213 24803 24271 24809
rect 24213 24800 24225 24803
rect 22969 24772 23336 24800
rect 23492 24772 24225 24800
rect 22969 24769 22981 24772
rect 22923 24763 22981 24769
rect 19444 24704 20116 24732
rect 19444 24673 19472 24704
rect 22646 24692 22652 24744
rect 22704 24692 22710 24744
rect 23308 24732 23336 24772
rect 24213 24769 24225 24772
rect 24259 24769 24271 24803
rect 24213 24763 24271 24769
rect 23308 24704 24256 24732
rect 24228 24676 24256 24704
rect 18555 24636 18828 24664
rect 18892 24636 19288 24664
rect 19429 24667 19487 24673
rect 18555 24633 18567 24636
rect 18509 24627 18567 24633
rect 15519 24568 18276 24596
rect 18693 24599 18751 24605
rect 15519 24565 15531 24568
rect 15473 24559 15531 24565
rect 18693 24565 18705 24599
rect 18739 24596 18751 24599
rect 18782 24596 18788 24608
rect 18739 24568 18788 24596
rect 18739 24565 18751 24568
rect 18693 24559 18751 24565
rect 18782 24556 18788 24568
rect 18840 24556 18846 24608
rect 18892 24605 18920 24636
rect 19429 24633 19441 24667
rect 19475 24633 19487 24667
rect 19429 24627 19487 24633
rect 24210 24624 24216 24676
rect 24268 24624 24274 24676
rect 18877 24599 18935 24605
rect 18877 24565 18889 24599
rect 18923 24565 18935 24599
rect 18877 24559 18935 24565
rect 19242 24556 19248 24608
rect 19300 24556 19306 24608
rect 20162 24556 20168 24608
rect 20220 24556 20226 24608
rect 1104 24506 24564 24528
rect 1104 24454 3882 24506
rect 3934 24454 3946 24506
rect 3998 24454 4010 24506
rect 4062 24454 4074 24506
rect 4126 24454 4138 24506
rect 4190 24454 9747 24506
rect 9799 24454 9811 24506
rect 9863 24454 9875 24506
rect 9927 24454 9939 24506
rect 9991 24454 10003 24506
rect 10055 24454 15612 24506
rect 15664 24454 15676 24506
rect 15728 24454 15740 24506
rect 15792 24454 15804 24506
rect 15856 24454 15868 24506
rect 15920 24454 21477 24506
rect 21529 24454 21541 24506
rect 21593 24454 21605 24506
rect 21657 24454 21669 24506
rect 21721 24454 21733 24506
rect 21785 24454 24564 24506
rect 1104 24432 24564 24454
rect 3602 24392 3608 24404
rect 1688 24364 3608 24392
rect 750 24216 756 24268
rect 808 24256 814 24268
rect 1688 24265 1716 24364
rect 3602 24352 3608 24364
rect 3660 24352 3666 24404
rect 5166 24392 5172 24404
rect 5000 24364 5172 24392
rect 2774 24284 2780 24336
rect 2832 24284 2838 24336
rect 4614 24324 4620 24336
rect 4264 24296 4620 24324
rect 1397 24259 1455 24265
rect 1397 24256 1409 24259
rect 808 24228 1409 24256
rect 808 24216 814 24228
rect 1397 24225 1409 24228
rect 1443 24225 1455 24259
rect 1397 24219 1455 24225
rect 1673 24259 1731 24265
rect 1673 24225 1685 24259
rect 1719 24225 1731 24259
rect 1673 24219 1731 24225
rect 2130 24216 2136 24268
rect 2188 24256 2194 24268
rect 4264 24265 4292 24296
rect 4614 24284 4620 24296
rect 4672 24284 4678 24336
rect 4798 24284 4804 24336
rect 4856 24324 4862 24336
rect 4893 24327 4951 24333
rect 4893 24324 4905 24327
rect 4856 24296 4905 24324
rect 4856 24284 4862 24296
rect 4893 24293 4905 24296
rect 4939 24293 4951 24327
rect 4893 24287 4951 24293
rect 4249 24259 4307 24265
rect 4249 24256 4261 24259
rect 2188 24228 4261 24256
rect 2188 24216 2194 24228
rect 4249 24225 4261 24228
rect 4295 24225 4307 24259
rect 5000 24256 5028 24364
rect 5166 24352 5172 24364
rect 5224 24352 5230 24404
rect 6086 24352 6092 24404
rect 6144 24352 6150 24404
rect 9030 24352 9036 24404
rect 9088 24352 9094 24404
rect 10870 24352 10876 24404
rect 10928 24392 10934 24404
rect 10965 24395 11023 24401
rect 10965 24392 10977 24395
rect 10928 24364 10977 24392
rect 10928 24352 10934 24364
rect 10965 24361 10977 24364
rect 11011 24361 11023 24395
rect 10965 24355 11023 24361
rect 12342 24352 12348 24404
rect 12400 24392 12406 24404
rect 17313 24395 17371 24401
rect 12400 24364 13584 24392
rect 12400 24352 12406 24364
rect 5307 24259 5365 24265
rect 5307 24256 5319 24259
rect 5000 24228 5319 24256
rect 4249 24219 4307 24225
rect 5307 24225 5319 24228
rect 5353 24225 5365 24259
rect 5307 24219 5365 24225
rect 7374 24216 7380 24268
rect 7432 24216 7438 24268
rect 1210 24148 1216 24200
rect 1268 24188 1274 24200
rect 2317 24191 2375 24197
rect 2317 24188 2329 24191
rect 1268 24160 2329 24188
rect 1268 24148 1274 24160
rect 2317 24157 2329 24160
rect 2363 24157 2375 24191
rect 2317 24151 2375 24157
rect 2593 24191 2651 24197
rect 2593 24157 2605 24191
rect 2639 24157 2651 24191
rect 2593 24151 2651 24157
rect 1302 24080 1308 24132
rect 1360 24120 1366 24132
rect 2608 24120 2636 24151
rect 4062 24148 4068 24200
rect 4120 24188 4126 24200
rect 4433 24191 4491 24197
rect 4433 24188 4445 24191
rect 4120 24160 4445 24188
rect 4120 24148 4126 24160
rect 4433 24157 4445 24160
rect 4479 24157 4491 24191
rect 4433 24151 4491 24157
rect 5166 24148 5172 24200
rect 5224 24148 5230 24200
rect 5442 24148 5448 24200
rect 5500 24148 5506 24200
rect 7561 24191 7619 24197
rect 7561 24157 7573 24191
rect 7607 24188 7619 24191
rect 9048 24188 9076 24352
rect 9582 24284 9588 24336
rect 9640 24324 9646 24336
rect 9640 24296 9904 24324
rect 9640 24284 9674 24296
rect 9646 24268 9674 24284
rect 9306 24216 9312 24268
rect 9364 24216 9370 24268
rect 9646 24228 9680 24268
rect 9674 24216 9680 24228
rect 9732 24216 9738 24268
rect 9766 24216 9772 24268
rect 9824 24216 9830 24268
rect 9876 24256 9904 24296
rect 12360 24296 12597 24324
rect 12360 24268 12388 24296
rect 10226 24265 10232 24268
rect 10045 24259 10103 24265
rect 10045 24256 10057 24259
rect 9876 24228 10057 24256
rect 10045 24225 10057 24228
rect 10091 24225 10103 24259
rect 10045 24219 10103 24225
rect 10183 24259 10232 24265
rect 10183 24225 10195 24259
rect 10229 24225 10232 24259
rect 10183 24219 10232 24225
rect 10226 24216 10232 24219
rect 10284 24216 10290 24268
rect 10502 24256 10508 24268
rect 10336 24228 10508 24256
rect 7607 24160 9076 24188
rect 7607 24157 7619 24160
rect 7561 24151 7619 24157
rect 9122 24148 9128 24200
rect 9180 24148 9186 24200
rect 10336 24197 10364 24228
rect 10502 24216 10508 24228
rect 10560 24256 10566 24268
rect 10870 24256 10876 24268
rect 10560 24228 10876 24256
rect 10560 24216 10566 24228
rect 10870 24216 10876 24228
rect 10928 24216 10934 24268
rect 11514 24216 11520 24268
rect 11572 24256 11578 24268
rect 11793 24259 11851 24265
rect 11793 24256 11805 24259
rect 11572 24228 11805 24256
rect 11572 24216 11578 24228
rect 11793 24225 11805 24228
rect 11839 24225 11851 24259
rect 11793 24219 11851 24225
rect 12342 24216 12348 24268
rect 12400 24216 12406 24268
rect 12434 24216 12440 24268
rect 12492 24216 12498 24268
rect 12569 24256 12597 24296
rect 12830 24259 12888 24265
rect 12830 24256 12842 24259
rect 12569 24228 12842 24256
rect 12830 24225 12842 24228
rect 12876 24225 12888 24259
rect 12830 24219 12888 24225
rect 12989 24259 13047 24265
rect 12989 24225 13001 24259
rect 13035 24256 13047 24259
rect 13170 24256 13176 24268
rect 13035 24228 13176 24256
rect 13035 24225 13047 24228
rect 12989 24219 13047 24225
rect 13170 24216 13176 24228
rect 13228 24216 13234 24268
rect 10321 24191 10379 24197
rect 10321 24157 10333 24191
rect 10367 24157 10379 24191
rect 10321 24151 10379 24157
rect 11054 24148 11060 24200
rect 11112 24188 11118 24200
rect 11698 24188 11704 24200
rect 11112 24160 11704 24188
rect 11112 24148 11118 24160
rect 11698 24148 11704 24160
rect 11756 24188 11762 24200
rect 11977 24191 12035 24197
rect 11977 24188 11989 24191
rect 11756 24160 11989 24188
rect 11756 24148 11762 24160
rect 11977 24157 11989 24160
rect 12023 24157 12035 24191
rect 11977 24151 12035 24157
rect 12710 24148 12716 24200
rect 12768 24148 12774 24200
rect 1360 24092 2636 24120
rect 6012 24092 7328 24120
rect 1360 24080 1366 24092
rect 2501 24055 2559 24061
rect 2501 24021 2513 24055
rect 2547 24052 2559 24055
rect 6012 24052 6040 24092
rect 2547 24024 6040 24052
rect 2547 24021 2559 24024
rect 2501 24015 2559 24021
rect 6270 24012 6276 24064
rect 6328 24052 6334 24064
rect 6638 24052 6644 24064
rect 6328 24024 6644 24052
rect 6328 24012 6334 24024
rect 6638 24012 6644 24024
rect 6696 24012 6702 24064
rect 7098 24012 7104 24064
rect 7156 24052 7162 24064
rect 7193 24055 7251 24061
rect 7193 24052 7205 24055
rect 7156 24024 7205 24052
rect 7156 24012 7162 24024
rect 7193 24021 7205 24024
rect 7239 24021 7251 24055
rect 7300 24052 7328 24092
rect 7466 24080 7472 24132
rect 7524 24080 7530 24132
rect 7650 24080 7656 24132
rect 7708 24120 7714 24132
rect 7929 24123 7987 24129
rect 7929 24120 7941 24123
rect 7708 24092 7941 24120
rect 7708 24080 7714 24092
rect 7929 24089 7941 24092
rect 7975 24089 7987 24123
rect 13556 24120 13584 24364
rect 17313 24361 17325 24395
rect 17359 24392 17371 24395
rect 18322 24392 18328 24404
rect 17359 24364 18328 24392
rect 17359 24361 17371 24364
rect 17313 24355 17371 24361
rect 18322 24352 18328 24364
rect 18380 24352 18386 24404
rect 18601 24395 18659 24401
rect 18601 24361 18613 24395
rect 18647 24392 18659 24395
rect 19150 24392 19156 24404
rect 18647 24364 19156 24392
rect 18647 24361 18659 24364
rect 18601 24355 18659 24361
rect 19150 24352 19156 24364
rect 19208 24352 19214 24404
rect 20162 24352 20168 24404
rect 20220 24392 20226 24404
rect 20809 24395 20867 24401
rect 20809 24392 20821 24395
rect 20220 24364 20821 24392
rect 20220 24352 20226 24364
rect 20809 24361 20821 24364
rect 20855 24361 20867 24395
rect 20809 24355 20867 24361
rect 21174 24352 21180 24404
rect 21232 24352 21238 24404
rect 23753 24395 23811 24401
rect 23753 24361 23765 24395
rect 23799 24392 23811 24395
rect 23842 24392 23848 24404
rect 23799 24364 23848 24392
rect 23799 24361 23811 24364
rect 23753 24355 23811 24361
rect 23842 24352 23848 24364
rect 23900 24352 23906 24404
rect 17494 24284 17500 24336
rect 17552 24284 17558 24336
rect 21192 24324 21220 24352
rect 20272 24296 21220 24324
rect 21361 24327 21419 24333
rect 14274 24216 14280 24268
rect 14332 24256 14338 24268
rect 14458 24256 14464 24268
rect 14332 24228 14464 24256
rect 14332 24216 14338 24228
rect 14458 24216 14464 24228
rect 14516 24216 14522 24268
rect 17512 24256 17540 24284
rect 17589 24259 17647 24265
rect 17589 24256 17601 24259
rect 17512 24228 17601 24256
rect 17589 24225 17601 24228
rect 17635 24225 17647 24259
rect 17589 24219 17647 24225
rect 13633 24191 13691 24197
rect 13633 24157 13645 24191
rect 13679 24188 13691 24191
rect 17402 24188 17408 24200
rect 13679 24160 17408 24188
rect 13679 24157 13691 24160
rect 13633 24151 13691 24157
rect 17402 24148 17408 24160
rect 17460 24188 17466 24200
rect 17497 24191 17555 24197
rect 17497 24188 17509 24191
rect 17460 24160 17509 24188
rect 17460 24148 17466 24160
rect 17497 24157 17509 24160
rect 17543 24157 17555 24191
rect 17847 24161 17905 24167
rect 17847 24158 17859 24161
rect 17497 24151 17555 24157
rect 14274 24120 14280 24132
rect 7929 24083 7987 24089
rect 8036 24092 8616 24120
rect 13556 24092 14280 24120
rect 8036 24052 8064 24092
rect 7300 24024 8064 24052
rect 8297 24055 8355 24061
rect 7193 24015 7251 24021
rect 8297 24021 8309 24055
rect 8343 24052 8355 24055
rect 8386 24052 8392 24064
rect 8343 24024 8392 24052
rect 8343 24021 8355 24024
rect 8297 24015 8355 24021
rect 8386 24012 8392 24024
rect 8444 24012 8450 24064
rect 8478 24012 8484 24064
rect 8536 24012 8542 24064
rect 8588 24052 8616 24092
rect 14274 24080 14280 24092
rect 14332 24120 14338 24132
rect 17846 24127 17859 24158
rect 17893 24127 17905 24161
rect 17954 24148 17960 24200
rect 18012 24188 18018 24200
rect 19518 24197 19524 24200
rect 19245 24191 19303 24197
rect 19245 24188 19257 24191
rect 18012 24160 19257 24188
rect 18012 24148 18018 24160
rect 19245 24157 19257 24160
rect 19291 24157 19303 24191
rect 19512 24188 19524 24197
rect 19479 24160 19524 24188
rect 19245 24151 19303 24157
rect 19512 24151 19524 24160
rect 19518 24148 19524 24151
rect 19576 24148 19582 24200
rect 17846 24121 17905 24127
rect 17846 24120 17874 24121
rect 14332 24092 17874 24120
rect 14332 24080 14338 24092
rect 13814 24052 13820 24064
rect 8588 24024 13820 24052
rect 13814 24012 13820 24024
rect 13872 24012 13878 24064
rect 14458 24012 14464 24064
rect 14516 24052 14522 24064
rect 20272 24052 20300 24296
rect 21361 24293 21373 24327
rect 21407 24293 21419 24327
rect 21361 24287 21419 24293
rect 20993 24259 21051 24265
rect 20993 24225 21005 24259
rect 21039 24256 21051 24259
rect 21177 24259 21235 24265
rect 21177 24256 21189 24259
rect 21039 24228 21189 24256
rect 21039 24225 21051 24228
rect 20993 24219 21051 24225
rect 21177 24225 21189 24228
rect 21223 24225 21235 24259
rect 21177 24219 21235 24225
rect 20717 24191 20775 24197
rect 20717 24188 20729 24191
rect 20456 24160 20729 24188
rect 20456 24064 20484 24160
rect 20717 24157 20729 24160
rect 20763 24188 20775 24191
rect 21085 24191 21143 24197
rect 21085 24188 21097 24191
rect 20763 24160 21097 24188
rect 20763 24157 20775 24160
rect 20717 24151 20775 24157
rect 21085 24157 21097 24160
rect 21131 24157 21143 24191
rect 21085 24151 21143 24157
rect 21269 24191 21327 24197
rect 21269 24157 21281 24191
rect 21315 24188 21327 24191
rect 21376 24188 21404 24287
rect 21315 24160 21404 24188
rect 21545 24191 21603 24197
rect 21315 24157 21327 24160
rect 21269 24151 21327 24157
rect 21545 24157 21557 24191
rect 21591 24157 21603 24191
rect 21545 24151 21603 24157
rect 22741 24191 22799 24197
rect 22741 24157 22753 24191
rect 22787 24157 22799 24191
rect 22741 24151 22799 24157
rect 23477 24191 23535 24197
rect 23477 24157 23489 24191
rect 23523 24188 23535 24191
rect 23658 24188 23664 24200
rect 23523 24160 23664 24188
rect 23523 24157 23535 24160
rect 23477 24151 23535 24157
rect 21560 24120 21588 24151
rect 20640 24092 21588 24120
rect 14516 24024 20300 24052
rect 14516 24012 14522 24024
rect 20438 24012 20444 24064
rect 20496 24012 20502 24064
rect 20640 24061 20668 24092
rect 22370 24080 22376 24132
rect 22428 24120 22434 24132
rect 22756 24120 22784 24151
rect 23658 24148 23664 24160
rect 23716 24148 23722 24200
rect 23937 24191 23995 24197
rect 23937 24157 23949 24191
rect 23983 24188 23995 24191
rect 24118 24188 24124 24200
rect 23983 24160 24124 24188
rect 23983 24157 23995 24160
rect 23937 24151 23995 24157
rect 24118 24148 24124 24160
rect 24176 24148 24182 24200
rect 22428 24092 22784 24120
rect 22428 24080 22434 24092
rect 20625 24055 20683 24061
rect 20625 24021 20637 24055
rect 20671 24021 20683 24055
rect 20625 24015 20683 24021
rect 20993 24055 21051 24061
rect 20993 24021 21005 24055
rect 21039 24052 21051 24055
rect 21818 24052 21824 24064
rect 21039 24024 21824 24052
rect 21039 24021 21051 24024
rect 20993 24015 21051 24021
rect 21818 24012 21824 24024
rect 21876 24012 21882 24064
rect 22557 24055 22615 24061
rect 22557 24021 22569 24055
rect 22603 24052 22615 24055
rect 23198 24052 23204 24064
rect 22603 24024 23204 24052
rect 22603 24021 22615 24024
rect 22557 24015 22615 24021
rect 23198 24012 23204 24024
rect 23256 24012 23262 24064
rect 24121 24055 24179 24061
rect 24121 24021 24133 24055
rect 24167 24052 24179 24055
rect 24854 24052 24860 24064
rect 24167 24024 24860 24052
rect 24167 24021 24179 24024
rect 24121 24015 24179 24021
rect 24854 24012 24860 24024
rect 24912 24012 24918 24064
rect 1104 23962 24723 23984
rect 1104 23910 6814 23962
rect 6866 23910 6878 23962
rect 6930 23910 6942 23962
rect 6994 23910 7006 23962
rect 7058 23910 7070 23962
rect 7122 23910 12679 23962
rect 12731 23910 12743 23962
rect 12795 23910 12807 23962
rect 12859 23910 12871 23962
rect 12923 23910 12935 23962
rect 12987 23910 18544 23962
rect 18596 23910 18608 23962
rect 18660 23910 18672 23962
rect 18724 23910 18736 23962
rect 18788 23910 18800 23962
rect 18852 23910 24409 23962
rect 24461 23910 24473 23962
rect 24525 23910 24537 23962
rect 24589 23910 24601 23962
rect 24653 23910 24665 23962
rect 24717 23910 24723 23962
rect 1104 23888 24723 23910
rect 1581 23851 1639 23857
rect 1581 23817 1593 23851
rect 1627 23817 1639 23851
rect 1581 23811 1639 23817
rect 1857 23851 1915 23857
rect 1857 23817 1869 23851
rect 1903 23848 1915 23851
rect 1903 23820 3096 23848
rect 1903 23817 1915 23820
rect 1857 23811 1915 23817
rect 1596 23780 1624 23811
rect 2498 23780 2504 23792
rect 1596 23752 2504 23780
rect 2498 23740 2504 23752
rect 2556 23740 2562 23792
rect 2590 23740 2596 23792
rect 2648 23740 2654 23792
rect 3068 23780 3096 23820
rect 3142 23808 3148 23860
rect 3200 23848 3206 23860
rect 3200 23820 7144 23848
rect 3200 23808 3206 23820
rect 3068 23752 3372 23780
rect 750 23672 756 23724
rect 808 23712 814 23724
rect 1397 23715 1455 23721
rect 1397 23712 1409 23715
rect 808 23684 1409 23712
rect 808 23672 814 23684
rect 1397 23681 1409 23684
rect 1443 23681 1455 23715
rect 1397 23675 1455 23681
rect 1670 23672 1676 23724
rect 1728 23672 1734 23724
rect 1946 23672 1952 23724
rect 2004 23672 2010 23724
rect 2130 23672 2136 23724
rect 2188 23672 2194 23724
rect 2774 23672 2780 23724
rect 2832 23712 2838 23724
rect 2869 23715 2927 23721
rect 2869 23712 2881 23715
rect 2832 23684 2881 23712
rect 2832 23672 2838 23684
rect 2869 23681 2881 23684
rect 2915 23681 2927 23715
rect 2869 23675 2927 23681
rect 2961 23715 3019 23721
rect 2961 23681 2973 23715
rect 3007 23712 3019 23715
rect 3142 23712 3148 23724
rect 3007 23684 3148 23712
rect 3007 23681 3019 23684
rect 2961 23675 3019 23681
rect 3142 23672 3148 23684
rect 3200 23672 3206 23724
rect 3344 23721 3372 23752
rect 3694 23740 3700 23792
rect 3752 23740 3758 23792
rect 4062 23740 4068 23792
rect 4120 23780 4126 23792
rect 4798 23780 4804 23792
rect 4120 23752 4804 23780
rect 4120 23740 4126 23752
rect 4798 23740 4804 23752
rect 4856 23740 4862 23792
rect 7116 23780 7144 23820
rect 7190 23808 7196 23860
rect 7248 23848 7254 23860
rect 8386 23848 8392 23860
rect 7248 23820 8392 23848
rect 7248 23808 7254 23820
rect 8386 23808 8392 23820
rect 8444 23808 8450 23860
rect 9122 23808 9128 23860
rect 9180 23848 9186 23860
rect 9180 23820 10916 23848
rect 9180 23808 9186 23820
rect 7116 23752 7972 23780
rect 3329 23715 3387 23721
rect 3329 23681 3341 23715
rect 3375 23712 3387 23715
rect 3786 23712 3792 23724
rect 3375 23684 3792 23712
rect 3375 23681 3387 23684
rect 3329 23675 3387 23681
rect 3786 23672 3792 23684
rect 3844 23672 3850 23724
rect 4154 23672 4160 23724
rect 4212 23712 4218 23724
rect 4675 23715 4733 23721
rect 4675 23712 4687 23715
rect 4212 23684 4687 23712
rect 4212 23672 4218 23684
rect 4675 23681 4687 23684
rect 4721 23681 4733 23715
rect 4675 23675 4733 23681
rect 5074 23672 5080 23724
rect 5132 23712 5138 23724
rect 6607 23715 6665 23721
rect 6607 23712 6619 23715
rect 5132 23684 6619 23712
rect 5132 23672 5138 23684
rect 6607 23681 6619 23684
rect 6653 23712 6665 23715
rect 7558 23712 7564 23724
rect 6653 23684 7564 23712
rect 6653 23681 6665 23684
rect 6607 23675 6665 23681
rect 7558 23672 7564 23684
rect 7616 23672 7622 23724
rect 7650 23672 7656 23724
rect 7708 23712 7714 23724
rect 7745 23715 7803 23721
rect 7745 23712 7757 23715
rect 7708 23684 7757 23712
rect 7708 23672 7714 23684
rect 7745 23681 7757 23684
rect 7791 23681 7803 23715
rect 7944 23712 7972 23752
rect 8202 23740 8208 23792
rect 8260 23780 8266 23792
rect 10888 23780 10916 23820
rect 10962 23808 10968 23860
rect 11020 23808 11026 23860
rect 11238 23808 11244 23860
rect 11296 23848 11302 23860
rect 11698 23848 11704 23860
rect 11296 23820 11704 23848
rect 11296 23808 11302 23820
rect 11698 23808 11704 23820
rect 11756 23808 11762 23860
rect 12434 23808 12440 23860
rect 12492 23848 12498 23860
rect 12621 23851 12679 23857
rect 12621 23848 12633 23851
rect 12492 23820 12633 23848
rect 12492 23808 12498 23820
rect 12621 23817 12633 23820
rect 12667 23817 12679 23851
rect 12621 23811 12679 23817
rect 13078 23808 13084 23860
rect 13136 23808 13142 23860
rect 20438 23808 20444 23860
rect 20496 23808 20502 23860
rect 13096 23780 13124 23808
rect 8260 23752 9168 23780
rect 10888 23752 13124 23780
rect 18432 23752 19334 23780
rect 8260 23740 8266 23752
rect 8003 23715 8061 23721
rect 8003 23712 8015 23715
rect 7944 23684 8015 23712
rect 7745 23675 7803 23681
rect 8003 23681 8015 23684
rect 8049 23712 8061 23715
rect 8386 23712 8392 23724
rect 8049 23684 8392 23712
rect 8049 23681 8061 23684
rect 8003 23675 8061 23681
rect 8386 23672 8392 23684
rect 8444 23672 8450 23724
rect 9140 23721 9168 23752
rect 9125 23715 9183 23721
rect 9125 23681 9137 23715
rect 9171 23712 9183 23715
rect 9171 23684 9444 23712
rect 9171 23681 9183 23684
rect 9125 23675 9183 23681
rect 2148 23585 2176 23672
rect 3050 23604 3056 23656
rect 3108 23604 3114 23656
rect 3878 23604 3884 23656
rect 3936 23644 3942 23656
rect 4433 23647 4491 23653
rect 4433 23644 4445 23647
rect 3936 23616 4445 23644
rect 3936 23604 3942 23616
rect 4433 23613 4445 23616
rect 4479 23613 4491 23647
rect 4433 23607 4491 23613
rect 2133 23579 2191 23585
rect 2133 23545 2145 23579
rect 2179 23545 2191 23579
rect 4448 23576 4476 23607
rect 6270 23604 6276 23656
rect 6328 23644 6334 23656
rect 6365 23647 6423 23653
rect 6365 23644 6377 23647
rect 6328 23616 6377 23644
rect 6328 23604 6334 23616
rect 6365 23613 6377 23616
rect 6411 23613 6423 23647
rect 6365 23607 6423 23613
rect 9306 23604 9312 23656
rect 9364 23604 9370 23656
rect 9416 23644 9444 23684
rect 11606 23672 11612 23724
rect 11664 23672 11670 23724
rect 11882 23712 11888 23724
rect 11843 23684 11888 23712
rect 11882 23672 11888 23684
rect 11940 23672 11946 23724
rect 15471 23715 15529 23721
rect 15471 23681 15483 23715
rect 15517 23712 15529 23715
rect 15517 23684 16160 23712
rect 15517 23681 15529 23684
rect 15471 23675 15529 23681
rect 9858 23655 9864 23656
rect 9842 23644 9864 23655
rect 9416 23616 9864 23644
rect 9858 23604 9864 23616
rect 9916 23604 9922 23656
rect 10042 23604 10048 23656
rect 10100 23604 10106 23656
rect 10226 23653 10232 23656
rect 10183 23647 10232 23653
rect 10183 23613 10195 23647
rect 10229 23613 10232 23647
rect 10183 23607 10232 23613
rect 10226 23604 10232 23607
rect 10284 23604 10290 23656
rect 10321 23647 10379 23653
rect 10321 23613 10333 23647
rect 10367 23636 10379 23647
rect 10520 23644 10640 23655
rect 10870 23644 10876 23656
rect 10520 23636 10876 23644
rect 10367 23627 10876 23636
rect 10367 23613 10548 23627
rect 10612 23616 10876 23627
rect 10321 23608 10548 23613
rect 10321 23607 10379 23608
rect 10870 23604 10876 23616
rect 10928 23604 10934 23656
rect 4448 23548 4568 23576
rect 2133 23539 2191 23545
rect 3881 23511 3939 23517
rect 3881 23477 3893 23511
rect 3927 23508 3939 23511
rect 4430 23508 4436 23520
rect 3927 23480 4436 23508
rect 3927 23477 3939 23480
rect 3881 23471 3939 23477
rect 4430 23468 4436 23480
rect 4488 23468 4494 23520
rect 4540 23508 4568 23548
rect 5092 23548 5580 23576
rect 5092 23508 5120 23548
rect 4540 23480 5120 23508
rect 5442 23468 5448 23520
rect 5500 23468 5506 23520
rect 5552 23508 5580 23548
rect 7098 23536 7104 23588
rect 7156 23576 7162 23588
rect 7282 23576 7288 23588
rect 7156 23548 7288 23576
rect 7156 23536 7162 23548
rect 7282 23536 7288 23548
rect 7340 23536 7346 23588
rect 7374 23536 7380 23588
rect 7432 23536 7438 23588
rect 9766 23585 9772 23588
rect 8757 23579 8815 23585
rect 8757 23545 8769 23579
rect 8803 23576 8815 23579
rect 9749 23579 9772 23585
rect 9749 23576 9761 23579
rect 8803 23548 9761 23576
rect 8803 23545 8815 23548
rect 8757 23539 8815 23545
rect 9749 23545 9761 23548
rect 9749 23539 9772 23545
rect 9766 23536 9772 23539
rect 9824 23536 9830 23588
rect 9582 23508 9588 23520
rect 5552 23480 9588 23508
rect 9582 23468 9588 23480
rect 9640 23468 9646 23520
rect 9858 23468 9864 23520
rect 9916 23508 9922 23520
rect 11054 23508 11060 23520
rect 9916 23480 11060 23508
rect 9916 23468 9922 23480
rect 11054 23468 11060 23480
rect 11112 23468 11118 23520
rect 11624 23508 11652 23672
rect 15197 23647 15255 23653
rect 15197 23613 15209 23647
rect 15243 23613 15255 23647
rect 15197 23607 15255 23613
rect 15212 23520 15240 23607
rect 14642 23508 14648 23520
rect 11624 23480 14648 23508
rect 14642 23468 14648 23480
rect 14700 23508 14706 23520
rect 15194 23508 15200 23520
rect 14700 23480 15200 23508
rect 14700 23468 14706 23480
rect 15194 23468 15200 23480
rect 15252 23468 15258 23520
rect 16132 23508 16160 23684
rect 16298 23672 16304 23724
rect 16356 23712 16362 23724
rect 16669 23715 16727 23721
rect 16669 23712 16681 23715
rect 16356 23684 16681 23712
rect 16356 23672 16362 23684
rect 16669 23681 16681 23684
rect 16715 23681 16727 23715
rect 16669 23675 16727 23681
rect 16758 23672 16764 23724
rect 16816 23712 16822 23724
rect 16853 23715 16911 23721
rect 16853 23712 16865 23715
rect 16816 23684 16865 23712
rect 16816 23672 16822 23684
rect 16853 23681 16865 23684
rect 16899 23681 16911 23715
rect 16853 23675 16911 23681
rect 17678 23672 17684 23724
rect 17736 23721 17742 23724
rect 17736 23715 17764 23721
rect 17752 23681 17764 23715
rect 17736 23675 17764 23681
rect 17736 23672 17742 23675
rect 18432 23656 18460 23752
rect 18601 23715 18659 23721
rect 18601 23681 18613 23715
rect 18647 23681 18659 23715
rect 18601 23675 18659 23681
rect 18693 23715 18751 23721
rect 18693 23681 18705 23715
rect 18739 23712 18751 23715
rect 18782 23712 18788 23724
rect 18739 23684 18788 23712
rect 18739 23681 18751 23684
rect 18693 23675 18751 23681
rect 17034 23604 17040 23656
rect 17092 23644 17098 23656
rect 17402 23644 17408 23656
rect 17092 23616 17408 23644
rect 17092 23604 17098 23616
rect 17402 23604 17408 23616
rect 17460 23644 17466 23656
rect 17589 23647 17647 23653
rect 17589 23644 17601 23647
rect 17460 23616 17601 23644
rect 17460 23604 17466 23616
rect 17589 23613 17601 23616
rect 17635 23613 17647 23647
rect 17589 23607 17647 23613
rect 17862 23604 17868 23656
rect 17920 23604 17926 23656
rect 18414 23604 18420 23656
rect 18472 23604 18478 23656
rect 16209 23579 16267 23585
rect 16209 23545 16221 23579
rect 16255 23576 16267 23579
rect 17313 23579 17371 23585
rect 17313 23576 17325 23579
rect 16255 23548 17325 23576
rect 16255 23545 16267 23548
rect 16209 23539 16267 23545
rect 17313 23545 17325 23548
rect 17359 23545 17371 23579
rect 18616 23576 18644 23675
rect 18782 23672 18788 23684
rect 18840 23672 18846 23724
rect 19306 23712 19334 23752
rect 21082 23740 21088 23792
rect 21140 23780 21146 23792
rect 22250 23783 22308 23789
rect 22250 23780 22262 23783
rect 21140 23752 22262 23780
rect 21140 23740 21146 23752
rect 22250 23749 22262 23752
rect 22296 23780 22308 23783
rect 22370 23780 22376 23792
rect 22296 23752 22376 23780
rect 22296 23749 22308 23752
rect 22250 23743 22308 23749
rect 22370 23740 22376 23752
rect 22428 23740 22434 23792
rect 23845 23783 23903 23789
rect 23845 23749 23857 23783
rect 23891 23780 23903 23783
rect 23934 23780 23940 23792
rect 23891 23752 23940 23780
rect 23891 23749 23903 23752
rect 23845 23743 23903 23749
rect 23934 23740 23940 23752
rect 23992 23740 23998 23792
rect 19671 23715 19729 23721
rect 19671 23712 19683 23715
rect 19306 23684 19683 23712
rect 19671 23681 19683 23684
rect 19717 23681 19729 23715
rect 19671 23675 19729 23681
rect 21358 23672 21364 23724
rect 21416 23672 21422 23724
rect 22005 23715 22063 23721
rect 22005 23681 22017 23715
rect 22051 23712 22063 23715
rect 22094 23712 22100 23724
rect 22051 23684 22100 23712
rect 22051 23681 22063 23684
rect 22005 23675 22063 23681
rect 18877 23647 18935 23653
rect 18877 23613 18889 23647
rect 18923 23644 18935 23647
rect 19242 23644 19248 23656
rect 18923 23616 19248 23644
rect 18923 23613 18935 23616
rect 18877 23607 18935 23613
rect 19242 23604 19248 23616
rect 19300 23604 19306 23656
rect 19334 23604 19340 23656
rect 19392 23644 19398 23656
rect 19429 23647 19487 23653
rect 19429 23644 19441 23647
rect 19392 23616 19441 23644
rect 19392 23604 19398 23616
rect 19429 23613 19441 23616
rect 19475 23613 19487 23647
rect 19429 23607 19487 23613
rect 20254 23604 20260 23656
rect 20312 23644 20318 23656
rect 22020 23644 22048 23675
rect 22094 23672 22100 23684
rect 22152 23672 22158 23724
rect 23661 23715 23719 23721
rect 23661 23712 23673 23715
rect 23400 23684 23673 23712
rect 20312 23616 22048 23644
rect 20312 23604 20318 23616
rect 19150 23576 19156 23588
rect 18616 23548 19156 23576
rect 17313 23539 17371 23545
rect 19150 23536 19156 23548
rect 19208 23536 19214 23588
rect 23400 23585 23428 23684
rect 23661 23681 23673 23684
rect 23707 23681 23719 23715
rect 23661 23675 23719 23681
rect 23385 23579 23443 23585
rect 23385 23545 23397 23579
rect 23431 23545 23443 23579
rect 23385 23539 23443 23545
rect 16758 23508 16764 23520
rect 16132 23480 16764 23508
rect 16758 23468 16764 23480
rect 16816 23508 16822 23520
rect 17586 23508 17592 23520
rect 16816 23480 17592 23508
rect 16816 23468 16822 23480
rect 17586 23468 17592 23480
rect 17644 23468 17650 23520
rect 18414 23468 18420 23520
rect 18472 23508 18478 23520
rect 18509 23511 18567 23517
rect 18509 23508 18521 23511
rect 18472 23480 18521 23508
rect 18472 23468 18478 23480
rect 18509 23477 18521 23480
rect 18555 23477 18567 23511
rect 18509 23471 18567 23477
rect 18785 23511 18843 23517
rect 18785 23477 18797 23511
rect 18831 23508 18843 23511
rect 20530 23508 20536 23520
rect 18831 23480 20536 23508
rect 18831 23477 18843 23480
rect 18785 23471 18843 23477
rect 20530 23468 20536 23480
rect 20588 23468 20594 23520
rect 21453 23511 21511 23517
rect 21453 23477 21465 23511
rect 21499 23508 21511 23511
rect 21910 23508 21916 23520
rect 21499 23480 21916 23508
rect 21499 23477 21511 23480
rect 21453 23471 21511 23477
rect 21910 23468 21916 23480
rect 21968 23468 21974 23520
rect 23290 23468 23296 23520
rect 23348 23508 23354 23520
rect 23477 23511 23535 23517
rect 23477 23508 23489 23511
rect 23348 23480 23489 23508
rect 23348 23468 23354 23480
rect 23477 23477 23489 23480
rect 23523 23477 23535 23511
rect 23477 23471 23535 23477
rect 24118 23468 24124 23520
rect 24176 23468 24182 23520
rect 1104 23418 24564 23440
rect 1104 23366 3882 23418
rect 3934 23366 3946 23418
rect 3998 23366 4010 23418
rect 4062 23366 4074 23418
rect 4126 23366 4138 23418
rect 4190 23366 9747 23418
rect 9799 23366 9811 23418
rect 9863 23366 9875 23418
rect 9927 23366 9939 23418
rect 9991 23366 10003 23418
rect 10055 23366 15612 23418
rect 15664 23366 15676 23418
rect 15728 23366 15740 23418
rect 15792 23366 15804 23418
rect 15856 23366 15868 23418
rect 15920 23366 21477 23418
rect 21529 23366 21541 23418
rect 21593 23366 21605 23418
rect 21657 23366 21669 23418
rect 21721 23366 21733 23418
rect 21785 23366 24564 23418
rect 1104 23344 24564 23366
rect 1949 23307 2007 23313
rect 1949 23273 1961 23307
rect 1995 23304 2007 23307
rect 2590 23304 2596 23316
rect 1995 23276 2596 23304
rect 1995 23273 2007 23276
rect 1949 23267 2007 23273
rect 2590 23264 2596 23276
rect 2648 23304 2654 23316
rect 2648 23276 3096 23304
rect 2648 23264 2654 23276
rect 3068 23236 3096 23276
rect 3142 23264 3148 23316
rect 3200 23304 3206 23316
rect 3329 23307 3387 23313
rect 3329 23304 3341 23307
rect 3200 23276 3341 23304
rect 3200 23264 3206 23276
rect 3329 23273 3341 23276
rect 3375 23273 3387 23307
rect 3329 23267 3387 23273
rect 5626 23264 5632 23316
rect 5684 23304 5690 23316
rect 5810 23304 5816 23316
rect 5684 23276 5816 23304
rect 5684 23264 5690 23276
rect 5810 23264 5816 23276
rect 5868 23264 5874 23316
rect 7098 23264 7104 23316
rect 7156 23304 7162 23316
rect 7374 23304 7380 23316
rect 7156 23276 7380 23304
rect 7156 23264 7162 23276
rect 7374 23264 7380 23276
rect 7432 23264 7438 23316
rect 8386 23264 8392 23316
rect 8444 23264 8450 23316
rect 10686 23264 10692 23316
rect 10744 23304 10750 23316
rect 10962 23304 10968 23316
rect 10744 23276 10968 23304
rect 10744 23264 10750 23276
rect 10962 23264 10968 23276
rect 11020 23264 11026 23316
rect 11514 23264 11520 23316
rect 11572 23304 11578 23316
rect 14458 23304 14464 23316
rect 11572 23276 14464 23304
rect 11572 23264 11578 23276
rect 14458 23264 14464 23276
rect 14516 23264 14522 23316
rect 17129 23307 17187 23313
rect 17129 23273 17141 23307
rect 17175 23304 17187 23307
rect 17862 23304 17868 23316
rect 17175 23276 17868 23304
rect 17175 23273 17187 23276
rect 17129 23267 17187 23273
rect 17862 23264 17868 23276
rect 17920 23264 17926 23316
rect 20717 23307 20775 23313
rect 20717 23273 20729 23307
rect 20763 23304 20775 23307
rect 21358 23304 21364 23316
rect 20763 23276 21364 23304
rect 20763 23273 20775 23276
rect 20717 23267 20775 23273
rect 21358 23264 21364 23276
rect 21416 23264 21422 23316
rect 22646 23264 22652 23316
rect 22704 23264 22710 23316
rect 8404 23236 8432 23264
rect 3068 23208 8432 23236
rect 8662 23196 8668 23248
rect 8720 23196 8726 23248
rect 8938 23196 8944 23248
rect 8996 23236 9002 23248
rect 10226 23236 10232 23248
rect 8996 23208 10232 23236
rect 8996 23196 9002 23208
rect 10226 23196 10232 23208
rect 10284 23236 10290 23248
rect 12342 23236 12348 23248
rect 10284 23208 12348 23236
rect 10284 23196 10290 23208
rect 12342 23196 12348 23208
rect 12400 23196 12406 23248
rect 17770 23196 17776 23248
rect 17828 23196 17834 23248
rect 22664 23236 22692 23264
rect 22572 23208 22692 23236
rect 2038 23128 2044 23180
rect 2096 23168 2102 23180
rect 2317 23171 2375 23177
rect 2317 23168 2329 23171
rect 2096 23140 2329 23168
rect 2096 23128 2102 23140
rect 2317 23137 2329 23140
rect 2363 23137 2375 23171
rect 2317 23131 2375 23137
rect 2332 23100 2360 23131
rect 6454 23128 6460 23180
rect 6512 23168 6518 23180
rect 8680 23168 8708 23196
rect 6512 23140 8708 23168
rect 6512 23128 6518 23140
rect 9490 23128 9496 23180
rect 9548 23168 9554 23180
rect 10686 23168 10692 23180
rect 9548 23140 10692 23168
rect 9548 23128 9554 23140
rect 10686 23128 10692 23140
rect 10744 23128 10750 23180
rect 15194 23128 15200 23180
rect 15252 23168 15258 23180
rect 16117 23171 16175 23177
rect 16117 23168 16129 23171
rect 15252 23140 16129 23168
rect 15252 23128 15258 23140
rect 2498 23100 2504 23112
rect 1688 23072 2176 23100
rect 2332 23072 2504 23100
rect 750 22992 756 23044
rect 808 23032 814 23044
rect 1688 23041 1716 23072
rect 1489 23035 1547 23041
rect 1489 23032 1501 23035
rect 808 23004 1501 23032
rect 808 22992 814 23004
rect 1489 23001 1501 23004
rect 1535 23001 1547 23035
rect 1489 22995 1547 23001
rect 1673 23035 1731 23041
rect 1673 23001 1685 23035
rect 1719 23001 1731 23035
rect 1673 22995 1731 23001
rect 1857 23035 1915 23041
rect 1857 23001 1869 23035
rect 1903 23001 1915 23035
rect 1857 22995 1915 23001
rect 842 22924 848 22976
rect 900 22964 906 22976
rect 1872 22964 1900 22995
rect 900 22936 1900 22964
rect 2148 22964 2176 23072
rect 2498 23060 2504 23072
rect 2556 23060 2562 23112
rect 2591 23103 2649 23109
rect 2591 23069 2603 23103
rect 2637 23100 2649 23103
rect 2682 23100 2688 23112
rect 2637 23072 2688 23100
rect 2637 23069 2649 23072
rect 2591 23063 2649 23069
rect 2682 23060 2688 23072
rect 2740 23060 2746 23112
rect 3786 23060 3792 23112
rect 3844 23100 3850 23112
rect 12526 23100 12532 23112
rect 3844 23072 12532 23100
rect 3844 23060 3850 23072
rect 12526 23060 12532 23072
rect 12584 23060 12590 23112
rect 13814 23060 13820 23112
rect 13872 23100 13878 23112
rect 13998 23100 14004 23112
rect 13872 23072 14004 23100
rect 13872 23060 13878 23072
rect 13998 23060 14004 23072
rect 14056 23060 14062 23112
rect 14461 23103 14519 23109
rect 14461 23069 14473 23103
rect 14507 23069 14519 23103
rect 14461 23063 14519 23069
rect 14735 23103 14793 23109
rect 14735 23069 14747 23103
rect 14781 23100 14793 23103
rect 14826 23100 14832 23112
rect 14781 23072 14832 23100
rect 14781 23069 14793 23072
rect 14735 23063 14793 23069
rect 2774 22992 2780 23044
rect 2832 23032 2838 23044
rect 7926 23032 7932 23044
rect 2832 23004 7932 23032
rect 2832 22992 2838 23004
rect 7926 22992 7932 23004
rect 7984 22992 7990 23044
rect 9398 22992 9404 23044
rect 9456 23032 9462 23044
rect 10226 23032 10232 23044
rect 9456 23004 10232 23032
rect 9456 22992 9462 23004
rect 10226 22992 10232 23004
rect 10284 22992 10290 23044
rect 11606 23032 11612 23044
rect 10520 23004 11612 23032
rect 3602 22964 3608 22976
rect 2148 22936 3608 22964
rect 900 22924 906 22936
rect 3602 22924 3608 22936
rect 3660 22964 3666 22976
rect 6270 22964 6276 22976
rect 3660 22936 6276 22964
rect 3660 22924 3666 22936
rect 6270 22924 6276 22936
rect 6328 22924 6334 22976
rect 6546 22924 6552 22976
rect 6604 22964 6610 22976
rect 7558 22964 7564 22976
rect 6604 22936 7564 22964
rect 6604 22924 6610 22936
rect 7558 22924 7564 22936
rect 7616 22924 7622 22976
rect 7742 22924 7748 22976
rect 7800 22964 7806 22976
rect 10520 22964 10548 23004
rect 11606 22992 11612 23004
rect 11664 22992 11670 23044
rect 14476 23032 14504 23063
rect 14826 23060 14832 23072
rect 14884 23060 14890 23112
rect 14016 23004 14504 23032
rect 14016 22976 14044 23004
rect 7800 22936 10548 22964
rect 7800 22924 7806 22936
rect 10594 22924 10600 22976
rect 10652 22964 10658 22976
rect 12250 22964 12256 22976
rect 10652 22936 12256 22964
rect 10652 22924 10658 22936
rect 12250 22924 12256 22936
rect 12308 22924 12314 22976
rect 12434 22924 12440 22976
rect 12492 22964 12498 22976
rect 13998 22964 14004 22976
rect 12492 22936 14004 22964
rect 12492 22924 12498 22936
rect 13998 22924 14004 22936
rect 14056 22924 14062 22976
rect 15194 22924 15200 22976
rect 15252 22964 15258 22976
rect 15473 22967 15531 22973
rect 15473 22964 15485 22967
rect 15252 22936 15485 22964
rect 15252 22924 15258 22936
rect 15473 22933 15485 22936
rect 15519 22933 15531 22967
rect 16040 22964 16068 23140
rect 16117 23137 16129 23140
rect 16163 23137 16175 23171
rect 16117 23131 16175 23137
rect 16391 23103 16449 23109
rect 16391 23069 16403 23103
rect 16437 23100 16449 23103
rect 17788 23100 17816 23196
rect 19334 23128 19340 23180
rect 19392 23168 19398 23180
rect 22572 23177 22600 23208
rect 20993 23171 21051 23177
rect 20993 23168 21005 23171
rect 19392 23140 21005 23168
rect 19392 23128 19398 23140
rect 20993 23137 21005 23140
rect 21039 23137 21051 23171
rect 22557 23171 22615 23177
rect 22557 23168 22569 23171
rect 20993 23131 21051 23137
rect 22066 23140 22569 23168
rect 20438 23100 20444 23112
rect 16437 23072 17749 23100
rect 17788 23072 20444 23100
rect 16437 23069 16449 23072
rect 16391 23063 16449 23069
rect 16114 22992 16120 23044
rect 16172 23032 16178 23044
rect 16298 23032 16304 23044
rect 16172 23004 16304 23032
rect 16172 22992 16178 23004
rect 16298 22992 16304 23004
rect 16356 22992 16362 23044
rect 17721 23032 17749 23072
rect 20438 23060 20444 23072
rect 20496 23100 20502 23112
rect 20901 23103 20959 23109
rect 20901 23100 20913 23103
rect 20496 23072 20913 23100
rect 20496 23060 20502 23072
rect 20901 23069 20913 23072
rect 20947 23069 20959 23103
rect 20901 23063 20959 23069
rect 18138 23032 18144 23044
rect 17721 23004 18144 23032
rect 18138 22992 18144 23004
rect 18196 22992 18202 23044
rect 21008 23032 21036 23131
rect 21266 23060 21272 23112
rect 21324 23060 21330 23112
rect 22066 23032 22094 23140
rect 22557 23137 22569 23140
rect 22603 23137 22615 23171
rect 24213 23171 24271 23177
rect 24213 23168 24225 23171
rect 22557 23131 22615 23137
rect 23216 23140 24225 23168
rect 22830 23109 22836 23112
rect 22799 23103 22836 23109
rect 22799 23069 22811 23103
rect 22799 23063 22836 23069
rect 22830 23060 22836 23063
rect 22888 23060 22894 23112
rect 21008 23004 22094 23032
rect 23106 22992 23112 23044
rect 23164 23032 23170 23044
rect 23216 23032 23244 23140
rect 24213 23137 24225 23140
rect 24259 23137 24271 23171
rect 24213 23131 24271 23137
rect 23937 23103 23995 23109
rect 23937 23100 23949 23103
rect 23164 23004 23244 23032
rect 23584 23072 23949 23100
rect 23164 22992 23170 23004
rect 16482 22964 16488 22976
rect 16040 22936 16488 22964
rect 15473 22927 15531 22933
rect 16482 22924 16488 22936
rect 16540 22924 16546 22976
rect 22002 22924 22008 22976
rect 22060 22924 22066 22976
rect 23474 22924 23480 22976
rect 23532 22964 23538 22976
rect 23584 22973 23612 23072
rect 23937 23069 23949 23072
rect 23983 23069 23995 23103
rect 23937 23063 23995 23069
rect 24026 23060 24032 23112
rect 24084 23060 24090 23112
rect 23569 22967 23627 22973
rect 23569 22964 23581 22967
rect 23532 22936 23581 22964
rect 23532 22924 23538 22936
rect 23569 22933 23581 22936
rect 23615 22933 23627 22967
rect 23569 22927 23627 22933
rect 24213 22967 24271 22973
rect 24213 22933 24225 22967
rect 24259 22964 24271 22967
rect 24259 22936 24808 22964
rect 24259 22933 24271 22936
rect 24213 22927 24271 22933
rect 1104 22874 24723 22896
rect 1104 22822 6814 22874
rect 6866 22822 6878 22874
rect 6930 22822 6942 22874
rect 6994 22822 7006 22874
rect 7058 22822 7070 22874
rect 7122 22822 12679 22874
rect 12731 22822 12743 22874
rect 12795 22822 12807 22874
rect 12859 22822 12871 22874
rect 12923 22822 12935 22874
rect 12987 22822 18544 22874
rect 18596 22822 18608 22874
rect 18660 22822 18672 22874
rect 18724 22822 18736 22874
rect 18788 22822 18800 22874
rect 18852 22822 24409 22874
rect 24461 22822 24473 22874
rect 24525 22822 24537 22874
rect 24589 22822 24601 22874
rect 24653 22822 24665 22874
rect 24717 22822 24723 22874
rect 1104 22800 24723 22822
rect 2961 22763 3019 22769
rect 2961 22729 2973 22763
rect 3007 22760 3019 22763
rect 3234 22760 3240 22772
rect 3007 22732 3240 22760
rect 3007 22729 3019 22732
rect 2961 22723 3019 22729
rect 3234 22720 3240 22732
rect 3292 22720 3298 22772
rect 3510 22720 3516 22772
rect 3568 22720 3574 22772
rect 5810 22720 5816 22772
rect 5868 22760 5874 22772
rect 5905 22763 5963 22769
rect 5905 22760 5917 22763
rect 5868 22732 5917 22760
rect 5868 22720 5874 22732
rect 5905 22729 5917 22732
rect 5951 22729 5963 22763
rect 7190 22760 7196 22772
rect 5905 22723 5963 22729
rect 6748 22732 7196 22760
rect 1302 22652 1308 22704
rect 1360 22692 1366 22704
rect 2869 22695 2927 22701
rect 2869 22692 2881 22695
rect 1360 22664 2881 22692
rect 1360 22652 1366 22664
rect 2869 22661 2881 22664
rect 2915 22661 2927 22695
rect 3528 22692 3556 22720
rect 6362 22692 6368 22704
rect 2869 22655 2927 22661
rect 3344 22664 3556 22692
rect 5166 22664 6368 22692
rect 1671 22627 1729 22633
rect 1671 22593 1683 22627
rect 1717 22624 1729 22627
rect 1762 22624 1768 22636
rect 1717 22596 1768 22624
rect 1717 22593 1729 22596
rect 1671 22587 1729 22593
rect 1762 22584 1768 22596
rect 1820 22624 1826 22636
rect 3344 22633 3372 22664
rect 3602 22633 3608 22636
rect 3329 22627 3387 22633
rect 1820 22596 2912 22624
rect 1820 22584 1826 22596
rect 1394 22516 1400 22568
rect 1452 22516 1458 22568
rect 2884 22432 2912 22596
rect 3329 22593 3341 22627
rect 3375 22593 3387 22627
rect 3329 22587 3387 22593
rect 3571 22627 3608 22633
rect 3571 22593 3583 22627
rect 3571 22587 3608 22593
rect 3602 22584 3608 22587
rect 3660 22584 3666 22636
rect 4706 22584 4712 22636
rect 4764 22624 4770 22636
rect 5166 22633 5194 22664
rect 6362 22652 6368 22664
rect 6420 22652 6426 22704
rect 6748 22636 6776 22732
rect 7190 22720 7196 22732
rect 7248 22720 7254 22772
rect 8478 22720 8484 22772
rect 8536 22760 8542 22772
rect 14734 22760 14740 22772
rect 8536 22732 13768 22760
rect 8536 22720 8542 22732
rect 10502 22652 10508 22704
rect 10560 22692 10566 22704
rect 10778 22692 10784 22704
rect 10560 22664 10784 22692
rect 10560 22652 10566 22664
rect 10778 22652 10784 22664
rect 10836 22652 10842 22704
rect 11514 22652 11520 22704
rect 11572 22652 11578 22704
rect 12710 22663 12716 22704
rect 12695 22657 12716 22663
rect 5151 22627 5209 22633
rect 5151 22624 5163 22627
rect 4764 22596 5163 22624
rect 4764 22584 4770 22596
rect 5151 22593 5163 22596
rect 5197 22593 5209 22627
rect 5151 22587 5209 22593
rect 5718 22584 5724 22636
rect 5776 22624 5782 22636
rect 5994 22624 6000 22636
rect 5776 22596 6000 22624
rect 5776 22584 5782 22596
rect 5994 22584 6000 22596
rect 6052 22584 6058 22636
rect 6178 22584 6184 22636
rect 6236 22624 6242 22636
rect 6549 22627 6607 22633
rect 6549 22624 6561 22627
rect 6236 22596 6561 22624
rect 6236 22584 6242 22596
rect 6549 22593 6561 22596
rect 6595 22593 6607 22627
rect 6549 22587 6607 22593
rect 6730 22584 6736 22636
rect 6788 22584 6794 22636
rect 7558 22584 7564 22636
rect 7616 22633 7622 22636
rect 7616 22627 7644 22633
rect 7632 22593 7644 22627
rect 7616 22587 7644 22593
rect 8389 22627 8447 22633
rect 8389 22593 8401 22627
rect 8435 22624 8447 22627
rect 8849 22627 8907 22633
rect 8849 22624 8861 22627
rect 8435 22596 8861 22624
rect 8435 22593 8447 22596
rect 8389 22587 8447 22593
rect 8849 22593 8861 22596
rect 8895 22593 8907 22627
rect 10043 22627 10101 22633
rect 10043 22624 10055 22627
rect 8849 22587 8907 22593
rect 8956 22596 10055 22624
rect 7616 22584 7622 22587
rect 4890 22516 4896 22568
rect 4948 22516 4954 22568
rect 5902 22516 5908 22568
rect 5960 22556 5966 22568
rect 6638 22556 6644 22568
rect 5960 22528 6644 22556
rect 5960 22516 5966 22528
rect 6638 22516 6644 22528
rect 6696 22516 6702 22568
rect 7469 22559 7527 22565
rect 7469 22556 7481 22559
rect 6932 22528 7481 22556
rect 4264 22460 5028 22488
rect 2409 22423 2467 22429
rect 2409 22389 2421 22423
rect 2455 22420 2467 22423
rect 2682 22420 2688 22432
rect 2455 22392 2688 22420
rect 2455 22389 2467 22392
rect 2409 22383 2467 22389
rect 2682 22380 2688 22392
rect 2740 22380 2746 22432
rect 2866 22380 2872 22432
rect 2924 22380 2930 22432
rect 3234 22380 3240 22432
rect 3292 22420 3298 22432
rect 4264 22420 4292 22460
rect 3292 22392 4292 22420
rect 3292 22380 3298 22392
rect 4338 22380 4344 22432
rect 4396 22380 4402 22432
rect 5000 22420 5028 22460
rect 5626 22448 5632 22500
rect 5684 22488 5690 22500
rect 6932 22488 6960 22528
rect 7469 22525 7481 22528
rect 7515 22525 7527 22559
rect 7469 22519 7527 22525
rect 7745 22559 7803 22565
rect 7745 22525 7757 22559
rect 7791 22556 7803 22559
rect 7926 22556 7932 22568
rect 7791 22528 7932 22556
rect 7791 22525 7803 22528
rect 7745 22519 7803 22525
rect 7926 22516 7932 22528
rect 7984 22516 7990 22568
rect 5684 22460 6960 22488
rect 5684 22448 5690 22460
rect 7190 22448 7196 22500
rect 7248 22448 7254 22500
rect 8202 22448 8208 22500
rect 8260 22488 8266 22500
rect 8956 22488 8984 22596
rect 10043 22593 10055 22596
rect 10089 22624 10101 22627
rect 11532 22624 11560 22652
rect 10089 22596 11560 22624
rect 10089 22593 10101 22596
rect 10043 22587 10101 22593
rect 11790 22584 11796 22636
rect 11848 22624 11854 22636
rect 12342 22624 12348 22636
rect 11848 22596 12348 22624
rect 11848 22584 11854 22596
rect 12342 22584 12348 22596
rect 12400 22584 12406 22636
rect 12434 22584 12440 22636
rect 12492 22584 12498 22636
rect 12695 22623 12707 22657
rect 12768 22652 12774 22704
rect 13740 22692 13768 22732
rect 14016 22732 14740 22760
rect 14016 22692 14044 22732
rect 14734 22720 14740 22732
rect 14792 22720 14798 22772
rect 14826 22720 14832 22772
rect 14884 22760 14890 22772
rect 15102 22760 15108 22772
rect 14884 22732 15108 22760
rect 14884 22720 14890 22732
rect 15102 22720 15108 22732
rect 15160 22720 15166 22772
rect 16850 22720 16856 22772
rect 16908 22760 16914 22772
rect 17402 22760 17408 22772
rect 16908 22732 17408 22760
rect 16908 22720 16914 22732
rect 17402 22720 17408 22732
rect 17460 22720 17466 22772
rect 20438 22720 20444 22772
rect 20496 22720 20502 22772
rect 22002 22720 22008 22772
rect 22060 22720 22066 22772
rect 23106 22720 23112 22772
rect 23164 22720 23170 22772
rect 23290 22720 23296 22772
rect 23348 22720 23354 22772
rect 24026 22720 24032 22772
rect 24084 22720 24090 22772
rect 19242 22692 19248 22704
rect 13740 22664 14044 22692
rect 18156 22664 19248 22692
rect 12741 22626 12756 22652
rect 12741 22623 12753 22626
rect 12695 22617 12753 22623
rect 13446 22584 13452 22636
rect 13504 22624 13510 22636
rect 13504 22596 14136 22624
rect 13504 22584 13510 22596
rect 9582 22516 9588 22568
rect 9640 22556 9646 22568
rect 9769 22559 9827 22565
rect 9769 22556 9781 22559
rect 9640 22528 9781 22556
rect 9640 22516 9646 22528
rect 9769 22525 9781 22528
rect 9815 22525 9827 22559
rect 9769 22519 9827 22525
rect 13814 22516 13820 22568
rect 13872 22516 13878 22568
rect 13906 22516 13912 22568
rect 13964 22556 13970 22568
rect 14001 22559 14059 22565
rect 14001 22556 14013 22559
rect 13964 22528 14013 22556
rect 13964 22516 13970 22528
rect 14001 22525 14013 22528
rect 14047 22525 14059 22559
rect 14108 22556 14136 22596
rect 14826 22584 14832 22636
rect 14884 22633 14890 22636
rect 14884 22627 14912 22633
rect 14900 22593 14912 22627
rect 14884 22587 14912 22593
rect 15657 22627 15715 22633
rect 15657 22593 15669 22627
rect 15703 22624 15715 22627
rect 16853 22627 16911 22633
rect 16853 22624 16865 22627
rect 15703 22596 16865 22624
rect 15703 22593 15715 22596
rect 15657 22587 15715 22593
rect 16853 22593 16865 22596
rect 16899 22593 16911 22627
rect 16853 22587 16911 22593
rect 14884 22584 14890 22587
rect 17954 22584 17960 22636
rect 18012 22624 18018 22636
rect 18156 22633 18184 22664
rect 19242 22652 19248 22664
rect 19300 22692 19306 22704
rect 19300 22664 20266 22692
rect 19300 22652 19306 22664
rect 20238 22636 20266 22664
rect 18414 22633 18420 22636
rect 18141 22627 18199 22633
rect 18141 22624 18153 22627
rect 18012 22596 18153 22624
rect 18012 22584 18018 22596
rect 18141 22593 18153 22596
rect 18187 22593 18199 22627
rect 18408 22624 18420 22633
rect 18375 22596 18420 22624
rect 18141 22587 18199 22593
rect 18408 22587 18420 22596
rect 18414 22584 18420 22587
rect 18472 22584 18478 22636
rect 19797 22627 19855 22633
rect 19797 22624 19809 22627
rect 19536 22596 19809 22624
rect 14737 22559 14795 22565
rect 14737 22556 14749 22559
rect 14108 22528 14749 22556
rect 14001 22519 14059 22525
rect 14737 22525 14749 22528
rect 14783 22525 14795 22559
rect 14737 22519 14795 22525
rect 15013 22559 15071 22565
rect 15013 22525 15025 22559
rect 15059 22556 15071 22559
rect 15194 22556 15200 22568
rect 15059 22528 15200 22556
rect 15059 22525 15071 22528
rect 15013 22519 15071 22525
rect 15194 22516 15200 22528
rect 15252 22516 15258 22568
rect 8260 22460 8984 22488
rect 8260 22448 8266 22460
rect 10594 22448 10600 22500
rect 10652 22448 10658 22500
rect 11514 22448 11520 22500
rect 11572 22488 11578 22500
rect 12158 22488 12164 22500
rect 11572 22460 12164 22488
rect 11572 22448 11578 22460
rect 12158 22448 12164 22460
rect 12216 22448 12222 22500
rect 13449 22491 13507 22497
rect 13449 22457 13461 22491
rect 13495 22488 13507 22491
rect 14458 22488 14464 22500
rect 13495 22460 14464 22488
rect 13495 22457 13507 22460
rect 13449 22451 13507 22457
rect 14458 22448 14464 22460
rect 14516 22448 14522 22500
rect 19536 22497 19564 22596
rect 19797 22593 19809 22596
rect 19843 22593 19855 22627
rect 20238 22596 20260 22636
rect 20312 22633 20318 22636
rect 19797 22587 19855 22593
rect 20254 22584 20260 22596
rect 20312 22624 20322 22633
rect 20456 22624 20484 22720
rect 22020 22692 22048 22720
rect 23308 22692 23336 22720
rect 24044 22692 24072 22720
rect 21836 22664 22508 22692
rect 21836 22633 21864 22664
rect 20513 22627 20571 22633
rect 20513 22624 20525 22627
rect 20312 22596 20357 22624
rect 20456 22596 20525 22624
rect 20312 22587 20322 22596
rect 20513 22593 20525 22596
rect 20559 22593 20571 22627
rect 20513 22587 20571 22593
rect 21821 22627 21879 22633
rect 21821 22593 21833 22627
rect 21867 22593 21879 22627
rect 21821 22587 21879 22593
rect 20312 22584 20318 22587
rect 21910 22584 21916 22636
rect 21968 22584 21974 22636
rect 22480 22633 22508 22664
rect 23124 22664 23336 22692
rect 23492 22664 24072 22692
rect 23124 22633 23152 22664
rect 22373 22627 22431 22633
rect 22373 22624 22385 22627
rect 22020 22596 22385 22624
rect 22020 22556 22048 22596
rect 22373 22593 22385 22596
rect 22419 22593 22431 22627
rect 22373 22587 22431 22593
rect 22465 22627 22523 22633
rect 22465 22593 22477 22627
rect 22511 22593 22523 22627
rect 22465 22587 22523 22593
rect 22649 22627 22707 22633
rect 22649 22593 22661 22627
rect 22695 22593 22707 22627
rect 22649 22587 22707 22593
rect 22925 22627 22983 22633
rect 22925 22593 22937 22627
rect 22971 22593 22983 22627
rect 22925 22587 22983 22593
rect 23109 22627 23167 22633
rect 23109 22593 23121 22627
rect 23155 22593 23167 22627
rect 23109 22587 23167 22593
rect 21652 22528 22048 22556
rect 22097 22559 22155 22565
rect 21652 22497 21680 22528
rect 22097 22525 22109 22559
rect 22143 22556 22155 22559
rect 22557 22559 22615 22565
rect 22557 22556 22569 22559
rect 22143 22528 22569 22556
rect 22143 22525 22155 22528
rect 22097 22519 22155 22525
rect 22557 22525 22569 22528
rect 22603 22525 22615 22559
rect 22557 22519 22615 22525
rect 19521 22491 19579 22497
rect 19521 22457 19533 22491
rect 19567 22457 19579 22491
rect 19521 22451 19579 22457
rect 21637 22491 21695 22497
rect 21637 22457 21649 22491
rect 21683 22457 21695 22491
rect 21637 22451 21695 22457
rect 22189 22491 22247 22497
rect 22189 22457 22201 22491
rect 22235 22488 22247 22491
rect 22664 22488 22692 22587
rect 22940 22556 22968 22587
rect 23198 22584 23204 22636
rect 23256 22584 23262 22636
rect 23293 22627 23351 22633
rect 23293 22593 23305 22627
rect 23339 22624 23351 22627
rect 23492 22624 23520 22664
rect 23339 22596 23520 22624
rect 23569 22627 23627 22633
rect 23339 22593 23351 22596
rect 23293 22587 23351 22593
rect 23569 22593 23581 22627
rect 23615 22593 23627 22627
rect 23569 22587 23627 22593
rect 23937 22627 23995 22633
rect 23937 22593 23949 22627
rect 23983 22624 23995 22627
rect 24780 22624 24808 22936
rect 23983 22596 24808 22624
rect 23983 22593 23995 22596
rect 23937 22587 23995 22593
rect 23474 22556 23480 22568
rect 22940 22528 23480 22556
rect 23474 22516 23480 22528
rect 23532 22516 23538 22568
rect 22235 22460 22692 22488
rect 22235 22457 22247 22460
rect 22189 22451 22247 22457
rect 22922 22448 22928 22500
rect 22980 22488 22986 22500
rect 23382 22488 23388 22500
rect 22980 22460 23388 22488
rect 22980 22448 22986 22460
rect 23382 22448 23388 22460
rect 23440 22448 23446 22500
rect 8570 22420 8576 22432
rect 5000 22392 8576 22420
rect 8570 22380 8576 22392
rect 8628 22380 8634 22432
rect 8662 22380 8668 22432
rect 8720 22380 8726 22432
rect 9030 22380 9036 22432
rect 9088 22420 9094 22432
rect 10612 22420 10640 22448
rect 9088 22392 10640 22420
rect 9088 22380 9094 22392
rect 10778 22380 10784 22432
rect 10836 22380 10842 22432
rect 10962 22380 10968 22432
rect 11020 22420 11026 22432
rect 14826 22420 14832 22432
rect 11020 22392 14832 22420
rect 11020 22380 11026 22392
rect 14826 22380 14832 22392
rect 14884 22380 14890 22432
rect 16669 22423 16727 22429
rect 16669 22389 16681 22423
rect 16715 22420 16727 22423
rect 17310 22420 17316 22432
rect 16715 22392 17316 22420
rect 16715 22389 16727 22392
rect 16669 22383 16727 22389
rect 17310 22380 17316 22392
rect 17368 22380 17374 22432
rect 19613 22423 19671 22429
rect 19613 22389 19625 22423
rect 19659 22420 19671 22423
rect 20898 22420 20904 22432
rect 19659 22392 20904 22420
rect 19659 22389 19671 22392
rect 19613 22383 19671 22389
rect 20898 22380 20904 22392
rect 20956 22380 20962 22432
rect 22005 22423 22063 22429
rect 22005 22389 22017 22423
rect 22051 22420 22063 22423
rect 23584 22420 23612 22587
rect 22051 22392 23612 22420
rect 22051 22389 22063 22392
rect 22005 22383 22063 22389
rect 23750 22380 23756 22432
rect 23808 22380 23814 22432
rect 24121 22423 24179 22429
rect 24121 22389 24133 22423
rect 24167 22420 24179 22423
rect 24854 22420 24860 22432
rect 24167 22392 24860 22420
rect 24167 22389 24179 22392
rect 24121 22383 24179 22389
rect 24854 22380 24860 22392
rect 24912 22380 24918 22432
rect 1104 22330 24564 22352
rect 1104 22278 3882 22330
rect 3934 22278 3946 22330
rect 3998 22278 4010 22330
rect 4062 22278 4074 22330
rect 4126 22278 4138 22330
rect 4190 22278 9747 22330
rect 9799 22278 9811 22330
rect 9863 22278 9875 22330
rect 9927 22278 9939 22330
rect 9991 22278 10003 22330
rect 10055 22278 15612 22330
rect 15664 22278 15676 22330
rect 15728 22278 15740 22330
rect 15792 22278 15804 22330
rect 15856 22278 15868 22330
rect 15920 22278 21477 22330
rect 21529 22278 21541 22330
rect 21593 22278 21605 22330
rect 21657 22278 21669 22330
rect 21721 22278 21733 22330
rect 21785 22278 24564 22330
rect 1104 22256 24564 22278
rect 24854 22244 24860 22296
rect 24912 22284 24918 22296
rect 25130 22284 25136 22296
rect 24912 22256 25136 22284
rect 24912 22244 24918 22256
rect 25130 22244 25136 22256
rect 25188 22244 25194 22296
rect 2240 22188 3372 22216
rect 2240 22148 2268 22188
rect 1872 22120 2268 22148
rect 3344 22148 3372 22188
rect 3418 22176 3424 22228
rect 3476 22216 3482 22228
rect 3602 22216 3608 22228
rect 3476 22188 3608 22216
rect 3476 22176 3482 22188
rect 3602 22176 3608 22188
rect 3660 22176 3666 22228
rect 4080 22188 4844 22216
rect 4080 22148 4108 22188
rect 3344 22120 4108 22148
rect 4816 22148 4844 22188
rect 4890 22176 4896 22228
rect 4948 22216 4954 22228
rect 5350 22216 5356 22228
rect 4948 22188 5356 22216
rect 4948 22176 4954 22188
rect 5350 22176 5356 22188
rect 5408 22176 5414 22228
rect 7742 22216 7748 22228
rect 5552 22188 7748 22216
rect 5552 22148 5580 22188
rect 7742 22176 7748 22188
rect 7800 22216 7806 22228
rect 7800 22188 8432 22216
rect 7800 22176 7806 22188
rect 4816 22120 5580 22148
rect 1872 22092 1900 22120
rect 1854 22040 1860 22092
rect 1912 22040 1918 22092
rect 2130 22040 2136 22092
rect 2188 22040 2194 22092
rect 2240 22080 2268 22120
rect 6270 22108 6276 22160
rect 6328 22148 6334 22160
rect 7282 22148 7288 22160
rect 6328 22120 7288 22148
rect 6328 22108 6334 22120
rect 7282 22108 7288 22120
rect 7340 22148 7346 22160
rect 8404 22148 8432 22188
rect 11514 22176 11520 22228
rect 11572 22176 11578 22228
rect 14826 22176 14832 22228
rect 14884 22216 14890 22228
rect 21450 22216 21456 22228
rect 14884 22188 21456 22216
rect 14884 22176 14890 22188
rect 21450 22176 21456 22188
rect 21508 22176 21514 22228
rect 8754 22148 8760 22160
rect 7340 22120 7604 22148
rect 8404 22120 8760 22148
rect 7340 22108 7346 22120
rect 2590 22089 2596 22092
rect 2409 22083 2467 22089
rect 2409 22080 2421 22083
rect 2240 22052 2421 22080
rect 2409 22049 2421 22052
rect 2455 22049 2467 22083
rect 2409 22043 2467 22049
rect 2547 22083 2596 22089
rect 2547 22049 2559 22083
rect 2593 22049 2596 22083
rect 2547 22043 2596 22049
rect 2590 22040 2596 22043
rect 2648 22040 2654 22092
rect 2682 22040 2688 22092
rect 2740 22040 2746 22092
rect 7190 22080 7196 22092
rect 6288 22052 7196 22080
rect 1489 22015 1547 22021
rect 1489 21981 1501 22015
rect 1535 21981 1547 22015
rect 1489 21975 1547 21981
rect 1673 22015 1731 22021
rect 1673 21981 1685 22015
rect 1719 21981 1731 22015
rect 1673 21975 1731 21981
rect 290 21904 296 21956
rect 348 21944 354 21956
rect 934 21944 940 21956
rect 348 21916 940 21944
rect 348 21904 354 21916
rect 934 21904 940 21916
rect 992 21904 998 21956
rect 1504 21888 1532 21975
rect 1486 21836 1492 21888
rect 1544 21836 1550 21888
rect 1688 21876 1716 21975
rect 3602 21972 3608 22024
rect 3660 22012 3666 22024
rect 3973 22015 4031 22021
rect 3973 22012 3985 22015
rect 3660 21984 3985 22012
rect 3660 21972 3666 21984
rect 3973 21981 3985 21984
rect 4019 21981 4031 22015
rect 4982 22012 4988 22024
rect 3973 21975 4031 21981
rect 4231 21985 4289 21991
rect 4231 21951 4243 21985
rect 4277 21982 4289 21985
rect 4690 21984 4988 22012
rect 4277 21951 4290 21982
rect 4231 21945 4290 21951
rect 4262 21944 4290 21945
rect 4430 21944 4436 21956
rect 4262 21916 4436 21944
rect 4430 21904 4436 21916
rect 4488 21904 4494 21956
rect 1946 21876 1952 21888
rect 1688 21848 1952 21876
rect 1946 21836 1952 21848
rect 2004 21836 2010 21888
rect 3326 21836 3332 21888
rect 3384 21836 3390 21888
rect 4154 21836 4160 21888
rect 4212 21876 4218 21888
rect 4690 21876 4718 21984
rect 4982 21972 4988 21984
rect 5040 21972 5046 22024
rect 5445 22015 5503 22021
rect 5445 21981 5457 22015
rect 5491 21981 5503 22015
rect 5445 21975 5503 21981
rect 5719 22015 5777 22021
rect 5719 21981 5731 22015
rect 5765 22012 5777 22015
rect 6178 22012 6184 22024
rect 5765 21984 6184 22012
rect 5765 21981 5777 21984
rect 5719 21975 5777 21981
rect 4890 21904 4896 21956
rect 4948 21944 4954 21956
rect 5460 21944 5488 21975
rect 6178 21972 6184 21984
rect 6236 21972 6242 22024
rect 4948 21916 6040 21944
rect 4948 21904 4954 21916
rect 6012 21888 6040 21916
rect 4212 21848 4718 21876
rect 4212 21836 4218 21848
rect 4982 21836 4988 21888
rect 5040 21836 5046 21888
rect 5994 21836 6000 21888
rect 6052 21836 6058 21888
rect 6288 21876 6316 22052
rect 7190 22040 7196 22052
rect 7248 22080 7254 22092
rect 7469 22083 7527 22089
rect 7469 22080 7481 22083
rect 7248 22052 7481 22080
rect 7248 22040 7254 22052
rect 7469 22049 7481 22052
rect 7515 22049 7527 22083
rect 7576 22080 7604 22120
rect 8754 22108 8760 22120
rect 8812 22108 8818 22160
rect 13262 22108 13268 22160
rect 13320 22108 13326 22160
rect 14458 22108 14464 22160
rect 14516 22148 14522 22160
rect 14737 22151 14795 22157
rect 14737 22148 14749 22151
rect 14516 22120 14749 22148
rect 14516 22108 14522 22120
rect 14737 22117 14749 22120
rect 14783 22117 14795 22151
rect 14737 22111 14795 22117
rect 19150 22108 19156 22160
rect 19208 22148 19214 22160
rect 19208 22120 19288 22148
rect 19208 22108 19214 22120
rect 7576 22052 7926 22080
rect 7469 22043 7527 22049
rect 6546 21972 6552 22024
rect 6604 21972 6610 22024
rect 6638 21972 6644 22024
rect 6696 22012 6702 22024
rect 6825 22015 6883 22021
rect 6825 22012 6837 22015
rect 6696 21984 6837 22012
rect 6696 21972 6702 21984
rect 6825 21981 6837 21984
rect 6871 21981 6883 22015
rect 6825 21975 6883 21981
rect 7009 22015 7067 22021
rect 7009 21981 7021 22015
rect 7055 21981 7067 22015
rect 7009 21975 7067 21981
rect 6564 21944 6592 21972
rect 7024 21944 7052 21975
rect 7742 21972 7748 22024
rect 7800 21972 7806 22024
rect 7898 22021 7926 22052
rect 9306 22040 9312 22092
rect 9364 22080 9370 22092
rect 9364 22052 9996 22080
rect 9364 22040 9370 22052
rect 7883 22015 7941 22021
rect 7883 21981 7895 22015
rect 7929 21981 7941 22015
rect 7883 21975 7941 21981
rect 8018 21972 8024 22024
rect 8076 21972 8082 22024
rect 8665 22015 8723 22021
rect 8665 21981 8677 22015
rect 8711 22012 8723 22015
rect 9217 22015 9275 22021
rect 9217 22012 9229 22015
rect 8711 21984 9229 22012
rect 8711 21981 8723 21984
rect 8665 21975 8723 21981
rect 9217 21981 9229 21984
rect 9263 21981 9275 22015
rect 9217 21975 9275 21981
rect 9398 21972 9404 22024
rect 9456 21972 9462 22024
rect 9585 22015 9643 22021
rect 9585 21981 9597 22015
rect 9631 21981 9643 22015
rect 9968 22012 9996 22052
rect 10778 22040 10784 22092
rect 10836 22040 10842 22092
rect 12434 22040 12440 22092
rect 12492 22040 12498 22092
rect 13078 22040 13084 22092
rect 13136 22080 13142 22092
rect 13446 22080 13452 22092
rect 13136 22052 13452 22080
rect 13136 22040 13142 22052
rect 13446 22040 13452 22052
rect 13504 22080 13510 22092
rect 14093 22083 14151 22089
rect 14093 22080 14105 22083
rect 13504 22052 14105 22080
rect 13504 22040 13510 22052
rect 14093 22049 14105 22052
rect 14139 22049 14151 22083
rect 14093 22043 14151 22049
rect 14182 22040 14188 22092
rect 14240 22080 14246 22092
rect 14277 22083 14335 22089
rect 14277 22080 14289 22083
rect 14240 22052 14289 22080
rect 14240 22040 14246 22052
rect 14277 22049 14289 22052
rect 14323 22049 14335 22083
rect 14826 22080 14832 22092
rect 14277 22043 14335 22049
rect 14366 22052 14832 22080
rect 9968 21984 10732 22012
rect 9585 21975 9643 21981
rect 9600 21944 9628 21975
rect 6564 21916 7052 21944
rect 9048 21916 9628 21944
rect 9048 21885 9076 21916
rect 10318 21904 10324 21956
rect 10376 21944 10382 21956
rect 10505 21947 10563 21953
rect 10505 21944 10517 21947
rect 10376 21916 10517 21944
rect 10376 21904 10382 21916
rect 10505 21913 10517 21916
rect 10551 21913 10563 21947
rect 10505 21907 10563 21913
rect 10594 21904 10600 21956
rect 10652 21904 10658 21956
rect 10704 21944 10732 21984
rect 10962 21972 10968 22024
rect 11020 21972 11026 22024
rect 12250 21972 12256 22024
rect 12308 22012 12314 22024
rect 14366 22012 14394 22052
rect 14826 22040 14832 22052
rect 14884 22040 14890 22092
rect 15102 22040 15108 22092
rect 15160 22089 15166 22092
rect 15160 22083 15188 22089
rect 15176 22049 15188 22083
rect 15160 22043 15188 22049
rect 15160 22040 15166 22043
rect 15286 22040 15292 22092
rect 15344 22040 15350 22092
rect 19260 22089 19288 22120
rect 15933 22083 15991 22089
rect 15933 22049 15945 22083
rect 15979 22080 15991 22083
rect 19245 22083 19303 22089
rect 15979 22052 18000 22080
rect 15979 22049 15991 22052
rect 15933 22043 15991 22049
rect 12308 21984 14394 22012
rect 12308 21972 12314 21984
rect 15010 21972 15016 22024
rect 15068 21972 15074 22024
rect 17034 21972 17040 22024
rect 17092 22012 17098 22024
rect 17221 22015 17279 22021
rect 17221 22012 17233 22015
rect 17092 21984 17233 22012
rect 17092 21972 17098 21984
rect 17221 21981 17233 21984
rect 17267 21981 17279 22015
rect 17221 21975 17279 21981
rect 17310 21972 17316 22024
rect 17368 22012 17374 22024
rect 17497 22015 17555 22021
rect 17497 22012 17509 22015
rect 17368 21984 17509 22012
rect 17368 21972 17374 21984
rect 17497 21981 17509 21984
rect 17543 21981 17555 22015
rect 17497 21975 17555 21981
rect 17589 22015 17647 22021
rect 17589 21981 17601 22015
rect 17635 22012 17647 22015
rect 17862 22012 17868 22024
rect 17635 21984 17868 22012
rect 17635 21981 17647 21984
rect 17589 21975 17647 21981
rect 17862 21972 17868 21984
rect 17920 21972 17926 22024
rect 17972 22021 18000 22052
rect 18156 22052 19196 22080
rect 18156 22021 18184 22052
rect 17957 22015 18015 22021
rect 17957 21981 17969 22015
rect 18003 21981 18015 22015
rect 17957 21975 18015 21981
rect 18141 22015 18199 22021
rect 18141 21981 18153 22015
rect 18187 21981 18199 22015
rect 18141 21975 18199 21981
rect 18325 22015 18383 22021
rect 18325 21981 18337 22015
rect 18371 21981 18383 22015
rect 18325 21975 18383 21981
rect 11333 21947 11391 21953
rect 11333 21944 11345 21947
rect 10704 21916 11345 21944
rect 11333 21913 11345 21916
rect 11379 21944 11391 21947
rect 11379 21916 12112 21944
rect 11379 21913 11391 21916
rect 11333 21907 11391 21913
rect 12084 21888 12112 21916
rect 12342 21904 12348 21956
rect 12400 21904 12406 21956
rect 12526 21904 12532 21956
rect 12584 21944 12590 21956
rect 12713 21947 12771 21953
rect 12713 21944 12725 21947
rect 12584 21916 12725 21944
rect 12584 21904 12590 21916
rect 12713 21913 12725 21916
rect 12759 21913 12771 21947
rect 14182 21944 14188 21956
rect 12713 21907 12771 21913
rect 13096 21916 14188 21944
rect 6457 21879 6515 21885
rect 6457 21876 6469 21879
rect 6288 21848 6469 21876
rect 6457 21845 6469 21848
rect 6503 21845 6515 21879
rect 6457 21839 6515 21845
rect 9033 21879 9091 21885
rect 9033 21845 9045 21879
rect 9079 21845 9091 21879
rect 9033 21839 9091 21845
rect 9582 21836 9588 21888
rect 9640 21836 9646 21888
rect 10229 21879 10287 21885
rect 10229 21845 10241 21879
rect 10275 21876 10287 21879
rect 10410 21876 10416 21888
rect 10275 21848 10416 21876
rect 10275 21845 10287 21848
rect 10229 21839 10287 21845
rect 10410 21836 10416 21848
rect 10468 21876 10474 21888
rect 10686 21876 10692 21888
rect 10468 21848 10692 21876
rect 10468 21836 10474 21848
rect 10686 21836 10692 21848
rect 10744 21836 10750 21888
rect 11422 21836 11428 21888
rect 11480 21876 11486 21888
rect 11790 21876 11796 21888
rect 11480 21848 11796 21876
rect 11480 21836 11486 21848
rect 11790 21836 11796 21848
rect 11848 21876 11854 21888
rect 11977 21879 12035 21885
rect 11977 21876 11989 21879
rect 11848 21848 11989 21876
rect 11848 21836 11854 21848
rect 11977 21845 11989 21848
rect 12023 21845 12035 21879
rect 11977 21839 12035 21845
rect 12066 21836 12072 21888
rect 12124 21836 12130 21888
rect 13096 21885 13124 21916
rect 14182 21904 14188 21916
rect 14240 21904 14246 21956
rect 18340 21944 18368 21975
rect 18506 21972 18512 22024
rect 18564 22012 18570 22024
rect 18785 22015 18843 22021
rect 18785 22012 18797 22015
rect 18564 21984 18797 22012
rect 18564 21972 18570 21984
rect 18785 21981 18797 21984
rect 18831 21981 18843 22015
rect 18785 21975 18843 21981
rect 18877 22015 18935 22021
rect 18877 21981 18889 22015
rect 18923 21981 18935 22015
rect 18877 21975 18935 21981
rect 17788 21916 18368 21944
rect 13081 21879 13139 21885
rect 13081 21845 13093 21879
rect 13127 21845 13139 21879
rect 13081 21839 13139 21845
rect 13170 21836 13176 21888
rect 13228 21876 13234 21888
rect 15010 21876 15016 21888
rect 13228 21848 15016 21876
rect 13228 21836 13234 21848
rect 15010 21836 15016 21848
rect 15068 21836 15074 21888
rect 17788 21885 17816 21916
rect 17773 21879 17831 21885
rect 17773 21845 17785 21879
rect 17819 21845 17831 21879
rect 17773 21839 17831 21845
rect 18322 21836 18328 21888
rect 18380 21836 18386 21888
rect 18601 21879 18659 21885
rect 18601 21845 18613 21879
rect 18647 21876 18659 21879
rect 18892 21876 18920 21975
rect 19168 21888 19196 22052
rect 19245 22049 19257 22083
rect 19291 22049 19303 22083
rect 25498 22080 25504 22092
rect 19245 22043 19303 22049
rect 23952 22052 25504 22080
rect 20625 22015 20683 22021
rect 20625 22012 20637 22015
rect 19503 21985 19561 21991
rect 19503 21982 19515 21985
rect 19502 21951 19515 21982
rect 19549 21951 19561 21985
rect 19502 21945 19561 21951
rect 20272 21984 20637 22012
rect 19502 21944 19530 21945
rect 19352 21916 19530 21944
rect 19352 21888 19380 21916
rect 18647 21848 18920 21876
rect 18647 21845 18659 21848
rect 18601 21839 18659 21845
rect 18966 21836 18972 21888
rect 19024 21836 19030 21888
rect 19150 21836 19156 21888
rect 19208 21836 19214 21888
rect 19334 21836 19340 21888
rect 19392 21836 19398 21888
rect 19610 21836 19616 21888
rect 19668 21876 19674 21888
rect 20272 21885 20300 21984
rect 20625 21981 20637 21984
rect 20671 21981 20683 22015
rect 20625 21975 20683 21981
rect 20806 21972 20812 22024
rect 20864 21972 20870 22024
rect 21174 21972 21180 22024
rect 21232 21972 21238 22024
rect 23952 22021 23980 22052
rect 25498 22040 25504 22052
rect 25556 22040 25562 22092
rect 23937 22015 23995 22021
rect 23937 21981 23949 22015
rect 23983 21981 23995 22015
rect 23937 21975 23995 21981
rect 24854 21972 24860 22024
rect 24912 21972 24918 22024
rect 25130 21972 25136 22024
rect 25188 22012 25194 22024
rect 25590 22012 25596 22024
rect 25188 21984 25596 22012
rect 25188 21972 25194 21984
rect 25590 21972 25596 21984
rect 25648 21972 25654 22024
rect 24872 21944 24900 21972
rect 24872 21916 25636 21944
rect 25608 21888 25636 21916
rect 20257 21879 20315 21885
rect 20257 21876 20269 21879
rect 19668 21848 20269 21876
rect 19668 21836 19674 21848
rect 20257 21845 20269 21848
rect 20303 21845 20315 21879
rect 20257 21839 20315 21845
rect 20714 21836 20720 21888
rect 20772 21836 20778 21888
rect 21358 21836 21364 21888
rect 21416 21836 21422 21888
rect 24121 21879 24179 21885
rect 24121 21845 24133 21879
rect 24167 21876 24179 21879
rect 24854 21876 24860 21888
rect 24167 21848 24860 21876
rect 24167 21845 24179 21848
rect 24121 21839 24179 21845
rect 24854 21836 24860 21848
rect 24912 21836 24918 21888
rect 25590 21836 25596 21888
rect 25648 21836 25654 21888
rect 1104 21786 24723 21808
rect 1104 21734 6814 21786
rect 6866 21734 6878 21786
rect 6930 21734 6942 21786
rect 6994 21734 7006 21786
rect 7058 21734 7070 21786
rect 7122 21734 12679 21786
rect 12731 21734 12743 21786
rect 12795 21734 12807 21786
rect 12859 21734 12871 21786
rect 12923 21734 12935 21786
rect 12987 21734 18544 21786
rect 18596 21734 18608 21786
rect 18660 21734 18672 21786
rect 18724 21734 18736 21786
rect 18788 21734 18800 21786
rect 18852 21734 24409 21786
rect 24461 21734 24473 21786
rect 24525 21734 24537 21786
rect 24589 21734 24601 21786
rect 24653 21734 24665 21786
rect 24717 21734 24723 21786
rect 1104 21712 24723 21734
rect 2130 21632 2136 21684
rect 2188 21672 2194 21684
rect 2409 21675 2467 21681
rect 2409 21672 2421 21675
rect 2188 21644 2421 21672
rect 2188 21632 2194 21644
rect 2409 21641 2421 21644
rect 2455 21641 2467 21675
rect 2409 21635 2467 21641
rect 3786 21632 3792 21684
rect 3844 21672 3850 21684
rect 3844 21644 5672 21672
rect 3844 21632 3850 21644
rect 1118 21564 1124 21616
rect 1176 21604 1182 21616
rect 1176 21576 2820 21604
rect 1176 21564 1182 21576
rect 1671 21539 1729 21545
rect 1671 21505 1683 21539
rect 1717 21536 1729 21539
rect 2038 21536 2044 21548
rect 1717 21508 2044 21536
rect 1717 21505 1729 21508
rect 1671 21499 1729 21505
rect 2038 21496 2044 21508
rect 2096 21536 2102 21548
rect 2406 21536 2412 21548
rect 2096 21508 2412 21536
rect 2096 21496 2102 21508
rect 2406 21496 2412 21508
rect 2464 21496 2470 21548
rect 2792 21545 2820 21576
rect 5534 21564 5540 21616
rect 5592 21564 5598 21616
rect 5644 21613 5672 21644
rect 7926 21632 7932 21684
rect 7984 21672 7990 21684
rect 8021 21675 8079 21681
rect 8021 21672 8033 21675
rect 7984 21644 8033 21672
rect 7984 21632 7990 21644
rect 8021 21641 8033 21644
rect 8067 21641 8079 21675
rect 10410 21672 10416 21684
rect 8021 21635 8079 21641
rect 8128 21644 10416 21672
rect 5629 21607 5687 21613
rect 5629 21573 5641 21607
rect 5675 21573 5687 21607
rect 8128 21604 8156 21644
rect 10410 21632 10416 21644
rect 10468 21632 10474 21684
rect 10594 21632 10600 21684
rect 10652 21672 10658 21684
rect 11057 21675 11115 21681
rect 11057 21672 11069 21675
rect 10652 21644 11069 21672
rect 10652 21632 10658 21644
rect 11057 21641 11069 21644
rect 11103 21641 11115 21675
rect 11057 21635 11115 21641
rect 12066 21632 12072 21684
rect 12124 21672 12130 21684
rect 12124 21644 12296 21672
rect 12124 21632 12130 21644
rect 5629 21567 5687 21573
rect 6104 21576 8156 21604
rect 2777 21539 2835 21545
rect 2777 21505 2789 21539
rect 2823 21505 2835 21539
rect 2777 21499 2835 21505
rect 3053 21539 3111 21545
rect 3053 21505 3065 21539
rect 3099 21505 3111 21539
rect 3053 21499 3111 21505
rect 1394 21428 1400 21480
rect 1452 21428 1458 21480
rect 3068 21468 3096 21499
rect 4982 21496 4988 21548
rect 5040 21496 5046 21548
rect 2056 21440 3096 21468
rect 1302 21292 1308 21344
rect 1360 21332 1366 21344
rect 2056 21332 2084 21440
rect 3234 21428 3240 21480
rect 3292 21468 3298 21480
rect 3789 21471 3847 21477
rect 3789 21468 3801 21471
rect 3292 21440 3801 21468
rect 3292 21428 3298 21440
rect 3789 21437 3801 21440
rect 3835 21437 3847 21471
rect 3789 21431 3847 21437
rect 3970 21428 3976 21480
rect 4028 21428 4034 21480
rect 4709 21471 4767 21477
rect 4709 21468 4721 21471
rect 4540 21440 4721 21468
rect 2130 21360 2136 21412
rect 2188 21400 2194 21412
rect 3988 21400 4016 21428
rect 2188 21372 4016 21400
rect 2188 21360 2194 21372
rect 4430 21360 4436 21412
rect 4488 21360 4494 21412
rect 1360 21304 2084 21332
rect 1360 21292 1366 21304
rect 2958 21292 2964 21344
rect 3016 21292 3022 21344
rect 3237 21335 3295 21341
rect 3237 21301 3249 21335
rect 3283 21332 3295 21335
rect 3694 21332 3700 21344
rect 3283 21304 3700 21332
rect 3283 21301 3295 21304
rect 3237 21295 3295 21301
rect 3694 21292 3700 21304
rect 3752 21292 3758 21344
rect 4154 21292 4160 21344
rect 4212 21332 4218 21344
rect 4540 21332 4568 21440
rect 4709 21437 4721 21440
rect 4755 21437 4767 21471
rect 4709 21431 4767 21437
rect 4847 21471 4905 21477
rect 4847 21437 4859 21471
rect 4893 21468 4905 21471
rect 5552 21468 5580 21564
rect 6104 21536 6132 21576
rect 11698 21564 11704 21616
rect 11756 21604 11762 21616
rect 12268 21604 12296 21644
rect 12342 21632 12348 21684
rect 12400 21672 12406 21684
rect 13081 21675 13139 21681
rect 13081 21672 13093 21675
rect 12400 21644 13093 21672
rect 12400 21632 12406 21644
rect 13081 21641 13093 21644
rect 13127 21641 13139 21675
rect 13081 21635 13139 21641
rect 13906 21632 13912 21684
rect 13964 21632 13970 21684
rect 15378 21632 15384 21684
rect 15436 21672 15442 21684
rect 15436 21644 15608 21672
rect 15436 21632 15442 21644
rect 13924 21604 13952 21632
rect 11756 21576 12202 21604
rect 12268 21576 13952 21604
rect 11756 21564 11762 21576
rect 4893 21440 5580 21468
rect 5920 21508 6132 21536
rect 4893 21437 4905 21440
rect 4847 21431 4905 21437
rect 5442 21360 5448 21412
rect 5500 21400 5506 21412
rect 5920 21400 5948 21508
rect 6178 21496 6184 21548
rect 6236 21536 6242 21548
rect 6546 21536 6552 21548
rect 6236 21508 6552 21536
rect 6236 21496 6242 21508
rect 6546 21496 6552 21508
rect 6604 21496 6610 21548
rect 7283 21539 7341 21545
rect 7283 21505 7295 21539
rect 7329 21536 7341 21539
rect 8018 21536 8024 21548
rect 7329 21508 8024 21536
rect 7329 21505 7341 21508
rect 7283 21499 7341 21505
rect 8018 21496 8024 21508
rect 8076 21496 8082 21548
rect 8939 21539 8997 21545
rect 8939 21505 8951 21539
rect 8985 21536 8997 21539
rect 10319 21539 10377 21545
rect 10319 21536 10331 21539
rect 8985 21508 10331 21536
rect 8985 21505 8997 21508
rect 8939 21499 8997 21505
rect 10319 21505 10331 21508
rect 10365 21536 10377 21539
rect 10962 21536 10968 21548
rect 10365 21508 10968 21536
rect 10365 21505 10377 21508
rect 10319 21499 10377 21505
rect 10962 21496 10968 21508
rect 11020 21496 11026 21548
rect 11514 21496 11520 21548
rect 11572 21536 11578 21548
rect 12066 21536 12072 21548
rect 11572 21508 12072 21536
rect 11572 21496 11578 21508
rect 12066 21496 12072 21508
rect 12124 21496 12130 21548
rect 12174 21536 12202 21576
rect 12343 21539 12401 21545
rect 12343 21536 12355 21539
rect 12174 21508 12355 21536
rect 12343 21505 12355 21508
rect 12389 21536 12401 21539
rect 12389 21508 12756 21536
rect 12389 21505 12401 21508
rect 12343 21499 12401 21505
rect 5994 21428 6000 21480
rect 6052 21468 6058 21480
rect 7009 21471 7067 21477
rect 7009 21468 7021 21471
rect 6052 21440 7021 21468
rect 6052 21428 6058 21440
rect 7009 21437 7021 21440
rect 7055 21437 7067 21471
rect 7009 21431 7067 21437
rect 8665 21471 8723 21477
rect 8665 21437 8677 21471
rect 8711 21437 8723 21471
rect 8665 21431 8723 21437
rect 5500 21372 5948 21400
rect 5500 21360 5506 21372
rect 6270 21360 6276 21412
rect 6328 21400 6334 21412
rect 6730 21400 6736 21412
rect 6328 21372 6736 21400
rect 6328 21360 6334 21372
rect 6730 21360 6736 21372
rect 6788 21360 6794 21412
rect 4212 21304 4568 21332
rect 4212 21292 4218 21304
rect 5166 21292 5172 21344
rect 5224 21332 5230 21344
rect 6546 21332 6552 21344
rect 5224 21304 6552 21332
rect 5224 21292 5230 21304
rect 6546 21292 6552 21304
rect 6604 21292 6610 21344
rect 7024 21332 7052 21431
rect 8680 21332 8708 21431
rect 9674 21428 9680 21480
rect 9732 21468 9738 21480
rect 10045 21471 10103 21477
rect 10045 21468 10057 21471
rect 9732 21440 10057 21468
rect 9732 21428 9738 21440
rect 10045 21437 10057 21440
rect 10091 21437 10103 21471
rect 10045 21431 10103 21437
rect 7024 21304 8708 21332
rect 9398 21292 9404 21344
rect 9456 21332 9462 21344
rect 9677 21335 9735 21341
rect 9677 21332 9689 21335
rect 9456 21304 9689 21332
rect 9456 21292 9462 21304
rect 9677 21301 9689 21304
rect 9723 21301 9735 21335
rect 10060 21332 10088 21431
rect 12158 21332 12164 21344
rect 10060 21304 12164 21332
rect 9677 21295 9735 21301
rect 12158 21292 12164 21304
rect 12216 21292 12222 21344
rect 12728 21332 12756 21508
rect 14458 21496 14464 21548
rect 14516 21536 14522 21548
rect 14642 21536 14648 21548
rect 14516 21508 14648 21536
rect 14516 21496 14522 21508
rect 14642 21496 14648 21508
rect 14700 21536 14706 21548
rect 15197 21539 15255 21545
rect 15197 21536 15209 21539
rect 14700 21508 15209 21536
rect 14700 21496 14706 21508
rect 15197 21505 15209 21508
rect 15243 21505 15255 21539
rect 15197 21499 15255 21505
rect 15471 21539 15529 21545
rect 15471 21505 15483 21539
rect 15517 21536 15529 21539
rect 15580 21536 15608 21644
rect 16850 21632 16856 21684
rect 16908 21672 16914 21684
rect 17678 21672 17684 21684
rect 16908 21644 17684 21672
rect 16908 21632 16914 21644
rect 17678 21632 17684 21644
rect 17736 21632 17742 21684
rect 17954 21632 17960 21684
rect 18012 21672 18018 21684
rect 18414 21672 18420 21684
rect 18012 21644 18420 21672
rect 18012 21632 18018 21644
rect 18414 21632 18420 21644
rect 18472 21632 18478 21684
rect 18966 21632 18972 21684
rect 19024 21632 19030 21684
rect 19061 21675 19119 21681
rect 19061 21641 19073 21675
rect 19107 21672 19119 21675
rect 19150 21672 19156 21684
rect 19107 21644 19156 21672
rect 19107 21641 19119 21644
rect 19061 21635 19119 21641
rect 19150 21632 19156 21644
rect 19208 21632 19214 21684
rect 20714 21632 20720 21684
rect 20772 21632 20778 21684
rect 22741 21675 22799 21681
rect 22741 21641 22753 21675
rect 22787 21641 22799 21675
rect 22741 21635 22799 21641
rect 16022 21564 16028 21616
rect 16080 21604 16086 21616
rect 18984 21604 19012 21632
rect 16080 21576 18828 21604
rect 18984 21576 19748 21604
rect 16080 21564 16086 21576
rect 15517 21508 15608 21536
rect 16669 21539 16727 21545
rect 15517 21505 15529 21508
rect 15471 21499 15529 21505
rect 16669 21505 16681 21539
rect 16715 21505 16727 21539
rect 16669 21502 16727 21505
rect 16592 21499 16727 21502
rect 16911 21539 16969 21545
rect 16911 21505 16923 21539
rect 16957 21536 16969 21539
rect 17310 21536 17316 21548
rect 16957 21508 17316 21536
rect 16957 21505 16969 21508
rect 16911 21499 16969 21505
rect 16482 21428 16488 21480
rect 16540 21468 16546 21480
rect 16592 21474 16712 21499
rect 17310 21496 17316 21508
rect 17368 21496 17374 21548
rect 18323 21539 18381 21545
rect 18323 21505 18335 21539
rect 18369 21536 18381 21539
rect 18800 21536 18828 21576
rect 19334 21536 19340 21548
rect 18369 21508 18736 21536
rect 18800 21508 19340 21536
rect 18369 21505 18381 21508
rect 18323 21499 18381 21505
rect 16592 21468 16620 21474
rect 16540 21440 16620 21468
rect 16540 21428 16546 21440
rect 18046 21428 18052 21480
rect 18104 21428 18110 21480
rect 12894 21360 12900 21412
rect 12952 21400 12958 21412
rect 17954 21400 17960 21412
rect 12952 21372 15332 21400
rect 12952 21360 12958 21372
rect 15194 21332 15200 21344
rect 12728 21304 15200 21332
rect 15194 21292 15200 21304
rect 15252 21292 15258 21344
rect 15304 21332 15332 21372
rect 16132 21372 16804 21400
rect 16132 21332 16160 21372
rect 15304 21304 16160 21332
rect 16206 21292 16212 21344
rect 16264 21292 16270 21344
rect 16776 21332 16804 21372
rect 17604 21372 17960 21400
rect 17604 21332 17632 21372
rect 17954 21360 17960 21372
rect 18012 21360 18018 21412
rect 16776 21304 17632 21332
rect 17678 21292 17684 21344
rect 17736 21292 17742 21344
rect 18064 21332 18092 21428
rect 18708 21400 18736 21508
rect 19334 21496 19340 21508
rect 19392 21496 19398 21548
rect 19610 21496 19616 21548
rect 19668 21496 19674 21548
rect 19720 21545 19748 21576
rect 19705 21539 19763 21545
rect 19705 21505 19717 21539
rect 19751 21505 19763 21539
rect 19705 21499 19763 21505
rect 19889 21471 19947 21477
rect 19889 21437 19901 21471
rect 19935 21468 19947 21471
rect 20732 21468 20760 21632
rect 22756 21604 22784 21635
rect 22756 21576 23428 21604
rect 21450 21496 21456 21548
rect 21508 21536 21514 21548
rect 22002 21536 22008 21548
rect 21508 21508 22008 21536
rect 21508 21496 21514 21508
rect 22002 21496 22008 21508
rect 22060 21536 22066 21548
rect 23400 21545 23428 21576
rect 22925 21539 22983 21545
rect 22925 21536 22937 21539
rect 22060 21508 22937 21536
rect 22060 21496 22066 21508
rect 22925 21505 22937 21508
rect 22971 21505 22983 21539
rect 22925 21499 22983 21505
rect 23385 21539 23443 21545
rect 23385 21505 23397 21539
rect 23431 21505 23443 21539
rect 23385 21499 23443 21505
rect 23842 21496 23848 21548
rect 23900 21496 23906 21548
rect 23937 21539 23995 21545
rect 23937 21505 23949 21539
rect 23983 21505 23995 21539
rect 23937 21499 23995 21505
rect 19935 21440 20760 21468
rect 19935 21437 19947 21440
rect 19889 21431 19947 21437
rect 21910 21428 21916 21480
rect 21968 21468 21974 21480
rect 23952 21468 23980 21499
rect 21968 21440 23980 21468
rect 21968 21428 21974 21440
rect 18874 21400 18880 21412
rect 18708 21372 18880 21400
rect 18874 21360 18880 21372
rect 18932 21400 18938 21412
rect 23198 21400 23204 21412
rect 18932 21372 23204 21400
rect 18932 21360 18938 21372
rect 23198 21360 23204 21372
rect 23256 21360 23262 21412
rect 23382 21360 23388 21412
rect 23440 21400 23446 21412
rect 23661 21403 23719 21409
rect 23661 21400 23673 21403
rect 23440 21372 23673 21400
rect 23440 21360 23446 21372
rect 23661 21369 23673 21372
rect 23707 21369 23719 21403
rect 23661 21363 23719 21369
rect 18414 21332 18420 21344
rect 18064 21304 18420 21332
rect 18414 21292 18420 21304
rect 18472 21292 18478 21344
rect 18506 21292 18512 21344
rect 18564 21332 18570 21344
rect 19518 21332 19524 21344
rect 18564 21304 19524 21332
rect 18564 21292 18570 21304
rect 19518 21292 19524 21304
rect 19576 21292 19582 21344
rect 19797 21335 19855 21341
rect 19797 21301 19809 21335
rect 19843 21332 19855 21335
rect 22738 21332 22744 21344
rect 19843 21304 22744 21332
rect 19843 21301 19855 21304
rect 19797 21295 19855 21301
rect 22738 21292 22744 21304
rect 22796 21292 22802 21344
rect 23477 21335 23535 21341
rect 23477 21301 23489 21335
rect 23523 21332 23535 21335
rect 24026 21332 24032 21344
rect 23523 21304 24032 21332
rect 23523 21301 23535 21304
rect 23477 21295 23535 21301
rect 24026 21292 24032 21304
rect 24084 21292 24090 21344
rect 24118 21292 24124 21344
rect 24176 21292 24182 21344
rect 1104 21242 24564 21264
rect 1104 21190 3882 21242
rect 3934 21190 3946 21242
rect 3998 21190 4010 21242
rect 4062 21190 4074 21242
rect 4126 21190 4138 21242
rect 4190 21190 9747 21242
rect 9799 21190 9811 21242
rect 9863 21190 9875 21242
rect 9927 21190 9939 21242
rect 9991 21190 10003 21242
rect 10055 21190 15612 21242
rect 15664 21190 15676 21242
rect 15728 21190 15740 21242
rect 15792 21190 15804 21242
rect 15856 21190 15868 21242
rect 15920 21190 21477 21242
rect 21529 21190 21541 21242
rect 21593 21190 21605 21242
rect 21657 21190 21669 21242
rect 21721 21190 21733 21242
rect 21785 21190 24564 21242
rect 1104 21168 24564 21190
rect 3513 21131 3571 21137
rect 3513 21097 3525 21131
rect 3559 21128 3571 21131
rect 4246 21128 4252 21140
rect 3559 21100 4252 21128
rect 3559 21097 3571 21100
rect 3513 21091 3571 21097
rect 4246 21088 4252 21100
rect 4304 21088 4310 21140
rect 5442 21128 5448 21140
rect 4356 21100 5448 21128
rect 3694 21020 3700 21072
rect 3752 21060 3758 21072
rect 4356 21060 4384 21100
rect 5442 21088 5448 21100
rect 5500 21088 5506 21140
rect 5534 21088 5540 21140
rect 5592 21088 5598 21140
rect 5810 21088 5816 21140
rect 5868 21128 5874 21140
rect 8021 21131 8079 21137
rect 8021 21128 8033 21131
rect 5868 21100 6960 21128
rect 5868 21088 5874 21100
rect 5552 21060 5580 21088
rect 3752 21032 4384 21060
rect 5368 21032 5580 21060
rect 3752 21020 3758 21032
rect 934 20952 940 21004
rect 992 20992 998 21004
rect 992 20964 1808 20992
rect 992 20952 998 20964
rect 750 20884 756 20936
rect 808 20924 814 20936
rect 1780 20933 1808 20964
rect 2682 20952 2688 21004
rect 2740 20952 2746 21004
rect 4338 20952 4344 21004
rect 4396 20992 4402 21004
rect 5261 20995 5319 21001
rect 5261 20992 5273 20995
rect 4396 20964 5273 20992
rect 4396 20952 4402 20964
rect 5261 20961 5273 20964
rect 5307 20961 5319 20995
rect 5261 20955 5319 20961
rect 1489 20927 1547 20933
rect 1489 20924 1501 20927
rect 808 20896 1501 20924
rect 808 20884 814 20896
rect 1489 20893 1501 20896
rect 1535 20893 1547 20927
rect 1489 20887 1547 20893
rect 1765 20927 1823 20933
rect 1765 20893 1777 20927
rect 1811 20893 1823 20927
rect 1765 20887 1823 20893
rect 2130 20884 2136 20936
rect 2188 20924 2194 20936
rect 2314 20924 2320 20936
rect 2188 20896 2320 20924
rect 2188 20884 2194 20896
rect 2314 20884 2320 20896
rect 2372 20884 2378 20936
rect 2958 20884 2964 20936
rect 3016 20924 3022 20936
rect 5077 20927 5135 20933
rect 3016 20896 5028 20924
rect 3016 20884 3022 20896
rect 934 20816 940 20868
rect 992 20856 998 20868
rect 2501 20859 2559 20865
rect 2501 20856 2513 20859
rect 992 20828 2513 20856
rect 992 20816 998 20828
rect 2501 20825 2513 20828
rect 2547 20825 2559 20859
rect 2501 20819 2559 20825
rect 2590 20816 2596 20868
rect 2648 20816 2654 20868
rect 3326 20816 3332 20868
rect 3384 20816 3390 20868
rect 5000 20856 5028 20896
rect 5077 20893 5089 20927
rect 5123 20924 5135 20927
rect 5368 20924 5396 21032
rect 5718 21020 5724 21072
rect 5776 21020 5782 21072
rect 6932 21069 6960 21100
rect 7024 21100 8033 21128
rect 6917 21063 6975 21069
rect 6917 21029 6929 21063
rect 6963 21029 6975 21063
rect 6917 21023 6975 21029
rect 5442 20952 5448 21004
rect 5500 20992 5506 21004
rect 5997 20995 6055 21001
rect 5997 20992 6009 20995
rect 5500 20964 6009 20992
rect 5500 20952 5506 20964
rect 5997 20961 6009 20964
rect 6043 20961 6055 20995
rect 5997 20955 6055 20961
rect 6273 20995 6331 21001
rect 6273 20961 6285 20995
rect 6319 20992 6331 20995
rect 7024 20992 7052 21100
rect 8021 21097 8033 21100
rect 8067 21097 8079 21131
rect 8021 21091 8079 21097
rect 9582 21088 9588 21140
rect 9640 21088 9646 21140
rect 10134 21088 10140 21140
rect 10192 21128 10198 21140
rect 10778 21128 10784 21140
rect 10192 21100 10784 21128
rect 10192 21088 10198 21100
rect 10778 21088 10784 21100
rect 10836 21088 10842 21140
rect 11514 21088 11520 21140
rect 11572 21088 11578 21140
rect 12434 21088 12440 21140
rect 12492 21088 12498 21140
rect 16206 21088 16212 21140
rect 16264 21088 16270 21140
rect 17678 21088 17684 21140
rect 17736 21088 17742 21140
rect 17862 21088 17868 21140
rect 17920 21128 17926 21140
rect 18141 21131 18199 21137
rect 18141 21128 18153 21131
rect 17920 21100 18153 21128
rect 17920 21088 17926 21100
rect 18141 21097 18153 21100
rect 18187 21097 18199 21131
rect 18141 21091 18199 21097
rect 18322 21088 18328 21140
rect 18380 21088 18386 21140
rect 19150 21088 19156 21140
rect 19208 21088 19214 21140
rect 23569 21131 23627 21137
rect 23569 21097 23581 21131
rect 23615 21128 23627 21131
rect 23842 21128 23848 21140
rect 23615 21100 23848 21128
rect 23615 21097 23627 21100
rect 23569 21091 23627 21097
rect 23842 21088 23848 21100
rect 23900 21088 23906 21140
rect 9600 21060 9628 21088
rect 11532 21060 11560 21088
rect 9600 21032 9996 21060
rect 6319 20964 7052 20992
rect 9217 20995 9275 21001
rect 6319 20961 6331 20964
rect 6273 20955 6331 20961
rect 9217 20961 9229 20995
rect 9263 20992 9275 20995
rect 9263 20964 9628 20992
rect 9263 20961 9275 20964
rect 9217 20955 9275 20961
rect 6178 20933 6184 20936
rect 5123 20896 5396 20924
rect 6135 20927 6184 20933
rect 5123 20893 5135 20896
rect 5077 20887 5135 20893
rect 6135 20893 6147 20927
rect 6181 20893 6184 20927
rect 6135 20887 6184 20893
rect 6178 20884 6184 20887
rect 6236 20884 6242 20936
rect 6914 20884 6920 20936
rect 6972 20924 6978 20936
rect 7009 20927 7067 20933
rect 7009 20924 7021 20927
rect 6972 20896 7021 20924
rect 6972 20884 6978 20896
rect 7009 20893 7021 20896
rect 7055 20893 7067 20927
rect 7009 20887 7067 20893
rect 7283 20927 7341 20933
rect 7283 20893 7295 20927
rect 7329 20924 7341 20927
rect 7834 20924 7840 20936
rect 7329 20896 7840 20924
rect 7329 20893 7341 20896
rect 7283 20887 7341 20893
rect 7834 20884 7840 20896
rect 7892 20924 7898 20936
rect 8202 20924 8208 20936
rect 7892 20896 8208 20924
rect 7892 20884 7898 20896
rect 8202 20884 8208 20896
rect 8260 20884 8266 20936
rect 8662 20884 8668 20936
rect 8720 20924 8726 20936
rect 9125 20927 9183 20933
rect 9125 20924 9137 20927
rect 8720 20896 9137 20924
rect 8720 20884 8726 20896
rect 9125 20893 9137 20896
rect 9171 20893 9183 20927
rect 9125 20887 9183 20893
rect 9398 20884 9404 20936
rect 9456 20884 9462 20936
rect 9600 20933 9628 20964
rect 9968 20933 9996 21032
rect 11440 21032 11560 21060
rect 11440 21001 11468 21032
rect 12158 21020 12164 21072
rect 12216 21060 12222 21072
rect 12894 21060 12900 21072
rect 12216 21032 12900 21060
rect 12216 21020 12222 21032
rect 12894 21020 12900 21032
rect 12952 21020 12958 21072
rect 16224 21060 16252 21088
rect 16761 21063 16819 21069
rect 16761 21060 16773 21063
rect 16224 21032 16773 21060
rect 16761 21029 16773 21032
rect 16807 21029 16819 21063
rect 16761 21023 16819 21029
rect 11425 20995 11483 21001
rect 11425 20961 11437 20995
rect 11471 20961 11483 20995
rect 11425 20955 11483 20961
rect 14182 20952 14188 21004
rect 14240 20992 14246 21004
rect 16301 20995 16359 21001
rect 16301 20992 16313 20995
rect 14240 20964 16313 20992
rect 14240 20952 14246 20964
rect 16301 20961 16313 20964
rect 16347 20961 16359 20995
rect 16301 20955 16359 20961
rect 17034 20952 17040 21004
rect 17092 20952 17098 21004
rect 17313 20995 17371 21001
rect 17313 20961 17325 20995
rect 17359 20992 17371 20995
rect 17696 20992 17724 21088
rect 18340 21001 18368 21088
rect 17359 20964 17724 20992
rect 18325 20995 18383 21001
rect 17359 20961 17371 20964
rect 17313 20955 17371 20961
rect 18325 20961 18337 20995
rect 18371 20961 18383 20995
rect 18325 20955 18383 20961
rect 9585 20927 9643 20933
rect 9585 20893 9597 20927
rect 9631 20893 9643 20927
rect 9585 20887 9643 20893
rect 9953 20927 10011 20933
rect 9953 20893 9965 20927
rect 9999 20893 10011 20927
rect 9953 20887 10011 20893
rect 11238 20884 11244 20936
rect 11296 20924 11302 20936
rect 11667 20927 11725 20933
rect 11667 20924 11679 20927
rect 11296 20896 11679 20924
rect 11296 20884 11302 20896
rect 11667 20893 11679 20896
rect 11713 20893 11725 20927
rect 11667 20887 11725 20893
rect 12526 20884 12532 20936
rect 12584 20924 12590 20936
rect 17218 20933 17224 20936
rect 16117 20927 16175 20933
rect 16117 20924 16129 20927
rect 12584 20896 16129 20924
rect 12584 20884 12590 20896
rect 16117 20893 16129 20896
rect 16163 20893 16175 20927
rect 16117 20887 16175 20893
rect 17175 20927 17224 20933
rect 17175 20893 17187 20927
rect 17221 20893 17224 20927
rect 17175 20887 17224 20893
rect 17218 20884 17224 20887
rect 17276 20884 17282 20936
rect 18049 20927 18107 20933
rect 18049 20893 18061 20927
rect 18095 20924 18107 20927
rect 19168 20924 19196 21088
rect 18095 20896 19196 20924
rect 18095 20893 18107 20896
rect 18049 20887 18107 20893
rect 19334 20884 19340 20936
rect 19392 20924 19398 20936
rect 20073 20927 20131 20933
rect 20073 20924 20085 20927
rect 19392 20896 20085 20924
rect 19392 20884 19398 20896
rect 20073 20893 20085 20896
rect 20119 20893 20131 20927
rect 20073 20887 20131 20893
rect 22186 20884 22192 20936
rect 22244 20884 22250 20936
rect 23845 20927 23903 20933
rect 23845 20893 23857 20927
rect 23891 20924 23903 20927
rect 25130 20924 25136 20936
rect 23891 20896 25136 20924
rect 23891 20893 23903 20896
rect 23845 20887 23903 20893
rect 25130 20884 25136 20896
rect 25188 20884 25194 20936
rect 9861 20859 9919 20865
rect 5000 20828 5304 20856
rect 1578 20748 1584 20800
rect 1636 20788 1642 20800
rect 1854 20788 1860 20800
rect 1636 20760 1860 20788
rect 1636 20748 1642 20760
rect 1854 20748 1860 20760
rect 1912 20748 1918 20800
rect 1949 20791 2007 20797
rect 1949 20757 1961 20791
rect 1995 20788 2007 20791
rect 2130 20788 2136 20800
rect 1995 20760 2136 20788
rect 1995 20757 2007 20760
rect 1949 20751 2007 20757
rect 2130 20748 2136 20760
rect 2188 20748 2194 20800
rect 2225 20791 2283 20797
rect 2225 20757 2237 20791
rect 2271 20788 2283 20791
rect 3418 20788 3424 20800
rect 2271 20760 3424 20788
rect 2271 20757 2283 20760
rect 2225 20751 2283 20757
rect 3418 20748 3424 20760
rect 3476 20748 3482 20800
rect 5276 20788 5304 20828
rect 9861 20825 9873 20859
rect 9907 20856 9919 20859
rect 10962 20856 10968 20868
rect 9907 20828 10968 20856
rect 9907 20825 9919 20828
rect 9861 20819 9919 20825
rect 10962 20816 10968 20828
rect 11020 20816 11026 20868
rect 12434 20856 12440 20868
rect 11072 20828 12440 20856
rect 6086 20788 6092 20800
rect 5276 20760 6092 20788
rect 6086 20748 6092 20760
rect 6144 20748 6150 20800
rect 6546 20748 6552 20800
rect 6604 20788 6610 20800
rect 11072 20788 11100 20828
rect 12434 20816 12440 20828
rect 12492 20856 12498 20868
rect 13170 20856 13176 20868
rect 12492 20828 13176 20856
rect 12492 20816 12498 20828
rect 13170 20816 13176 20828
rect 13228 20816 13234 20868
rect 16022 20816 16028 20868
rect 16080 20856 16086 20868
rect 16206 20856 16212 20868
rect 16080 20828 16212 20856
rect 16080 20816 16086 20828
rect 16206 20816 16212 20828
rect 16264 20816 16270 20868
rect 17788 20828 19656 20856
rect 6604 20760 11100 20788
rect 6604 20748 6610 20760
rect 17310 20748 17316 20800
rect 17368 20788 17374 20800
rect 17788 20788 17816 20828
rect 19628 20800 19656 20828
rect 19886 20816 19892 20868
rect 19944 20856 19950 20868
rect 20346 20865 20352 20868
rect 20318 20859 20352 20865
rect 20318 20856 20330 20859
rect 19944 20828 20330 20856
rect 19944 20816 19950 20828
rect 20318 20825 20330 20828
rect 20318 20819 20352 20825
rect 20346 20816 20352 20819
rect 20404 20816 20410 20868
rect 20714 20816 20720 20868
rect 20772 20856 20778 20868
rect 21910 20856 21916 20868
rect 20772 20828 21916 20856
rect 20772 20816 20778 20828
rect 21910 20816 21916 20828
rect 21968 20816 21974 20868
rect 22002 20816 22008 20868
rect 22060 20856 22066 20868
rect 22434 20859 22492 20865
rect 22434 20856 22446 20859
rect 22060 20828 22446 20856
rect 22060 20816 22066 20828
rect 22434 20825 22446 20828
rect 22480 20825 22492 20859
rect 22434 20819 22492 20825
rect 24213 20859 24271 20865
rect 24213 20825 24225 20859
rect 24259 20856 24271 20859
rect 24854 20856 24860 20868
rect 24259 20828 24860 20856
rect 24259 20825 24271 20828
rect 24213 20819 24271 20825
rect 24854 20816 24860 20828
rect 24912 20816 24918 20868
rect 17368 20760 17816 20788
rect 17368 20748 17374 20760
rect 17954 20748 17960 20800
rect 18012 20748 18018 20800
rect 18325 20791 18383 20797
rect 18325 20757 18337 20791
rect 18371 20788 18383 20791
rect 18874 20788 18880 20800
rect 18371 20760 18880 20788
rect 18371 20757 18383 20760
rect 18325 20751 18383 20757
rect 18874 20748 18880 20760
rect 18932 20748 18938 20800
rect 19610 20748 19616 20800
rect 19668 20748 19674 20800
rect 21450 20748 21456 20800
rect 21508 20748 21514 20800
rect 1104 20698 24723 20720
rect 1104 20646 6814 20698
rect 6866 20646 6878 20698
rect 6930 20646 6942 20698
rect 6994 20646 7006 20698
rect 7058 20646 7070 20698
rect 7122 20646 12679 20698
rect 12731 20646 12743 20698
rect 12795 20646 12807 20698
rect 12859 20646 12871 20698
rect 12923 20646 12935 20698
rect 12987 20646 18544 20698
rect 18596 20646 18608 20698
rect 18660 20646 18672 20698
rect 18724 20646 18736 20698
rect 18788 20646 18800 20698
rect 18852 20646 24409 20698
rect 24461 20646 24473 20698
rect 24525 20646 24537 20698
rect 24589 20646 24601 20698
rect 24653 20646 24665 20698
rect 24717 20646 24723 20698
rect 1104 20624 24723 20646
rect 658 20544 664 20596
rect 716 20584 722 20596
rect 1578 20584 1584 20596
rect 716 20556 1584 20584
rect 716 20544 722 20556
rect 1578 20544 1584 20556
rect 1636 20544 1642 20596
rect 1949 20587 2007 20593
rect 1949 20553 1961 20587
rect 1995 20584 2007 20587
rect 2038 20584 2044 20596
rect 1995 20556 2044 20584
rect 1995 20553 2007 20556
rect 1949 20547 2007 20553
rect 2038 20544 2044 20556
rect 2096 20544 2102 20596
rect 2222 20544 2228 20596
rect 2280 20584 2286 20596
rect 2317 20587 2375 20593
rect 2317 20584 2329 20587
rect 2280 20556 2329 20584
rect 2280 20544 2286 20556
rect 2317 20553 2329 20556
rect 2363 20553 2375 20587
rect 2317 20547 2375 20553
rect 2590 20544 2596 20596
rect 2648 20584 2654 20596
rect 3697 20587 3755 20593
rect 3697 20584 3709 20587
rect 2648 20556 3709 20584
rect 2648 20544 2654 20556
rect 3697 20553 3709 20556
rect 3743 20553 3755 20587
rect 5810 20584 5816 20596
rect 3697 20547 3755 20553
rect 3804 20556 5816 20584
rect 934 20476 940 20528
rect 992 20516 998 20528
rect 3510 20516 3516 20528
rect 992 20488 1900 20516
rect 992 20476 998 20488
rect 1486 20408 1492 20460
rect 1544 20408 1550 20460
rect 1872 20457 1900 20488
rect 2976 20488 3516 20516
rect 2976 20487 3004 20488
rect 2943 20481 3004 20487
rect 1857 20451 1915 20457
rect 1857 20417 1869 20451
rect 1903 20417 1915 20451
rect 1857 20411 1915 20417
rect 2225 20451 2283 20457
rect 2225 20417 2237 20451
rect 2271 20417 2283 20451
rect 2225 20411 2283 20417
rect 1118 20340 1124 20392
rect 1176 20380 1182 20392
rect 2240 20380 2268 20411
rect 2498 20408 2504 20460
rect 2556 20448 2562 20460
rect 2685 20451 2743 20457
rect 2685 20448 2697 20451
rect 2556 20420 2697 20448
rect 2556 20408 2562 20420
rect 2685 20417 2697 20420
rect 2731 20417 2743 20451
rect 2943 20447 2955 20481
rect 2989 20450 3004 20481
rect 3510 20476 3516 20488
rect 3568 20476 3574 20528
rect 2989 20447 3001 20450
rect 2943 20441 3001 20447
rect 2685 20411 2743 20417
rect 3694 20408 3700 20460
rect 3752 20448 3758 20460
rect 3804 20448 3832 20556
rect 5810 20544 5816 20556
rect 5868 20544 5874 20596
rect 6362 20544 6368 20596
rect 6420 20584 6426 20596
rect 6730 20584 6736 20596
rect 6420 20556 6736 20584
rect 6420 20544 6426 20556
rect 6730 20544 6736 20556
rect 6788 20544 6794 20596
rect 8294 20584 8300 20596
rect 7484 20556 8300 20584
rect 4798 20476 4804 20528
rect 4856 20516 4862 20528
rect 7484 20516 7512 20556
rect 8294 20544 8300 20556
rect 8352 20544 8358 20596
rect 14366 20544 14372 20596
rect 14424 20544 14430 20596
rect 20346 20544 20352 20596
rect 20404 20544 20410 20596
rect 20625 20587 20683 20593
rect 20625 20553 20637 20587
rect 20671 20553 20683 20587
rect 20625 20547 20683 20553
rect 8662 20516 8668 20528
rect 4856 20488 7512 20516
rect 7576 20488 8668 20516
rect 4856 20476 4862 20488
rect 3752 20420 3832 20448
rect 3752 20408 3758 20420
rect 4338 20408 4344 20460
rect 4396 20408 4402 20460
rect 5534 20408 5540 20460
rect 5592 20448 5598 20460
rect 6638 20448 6644 20460
rect 5592 20420 6644 20448
rect 5592 20408 5598 20420
rect 6638 20408 6644 20420
rect 6696 20408 6702 20460
rect 1176 20352 2268 20380
rect 4065 20383 4123 20389
rect 1176 20340 1182 20352
rect 4065 20349 4077 20383
rect 4111 20349 4123 20383
rect 4065 20343 4123 20349
rect 1302 20204 1308 20256
rect 1360 20244 1366 20256
rect 4078 20244 4106 20343
rect 7190 20340 7196 20392
rect 7248 20380 7254 20392
rect 7576 20389 7604 20488
rect 8662 20476 8668 20488
rect 8720 20516 8726 20528
rect 10226 20516 10232 20528
rect 8720 20488 10232 20516
rect 8720 20476 8726 20488
rect 10226 20476 10232 20488
rect 10284 20476 10290 20528
rect 11146 20476 11152 20528
rect 11204 20516 11210 20528
rect 12250 20516 12256 20528
rect 11204 20488 12256 20516
rect 11204 20476 11210 20488
rect 12250 20476 12256 20488
rect 12308 20516 12314 20528
rect 12989 20519 13047 20525
rect 12989 20516 13001 20519
rect 12308 20488 13001 20516
rect 12308 20476 12314 20488
rect 12989 20485 13001 20488
rect 13035 20485 13047 20519
rect 12989 20479 13047 20485
rect 13906 20476 13912 20528
rect 13964 20516 13970 20528
rect 14093 20519 14151 20525
rect 14093 20516 14105 20519
rect 13964 20488 14105 20516
rect 13964 20476 13970 20488
rect 14093 20485 14105 20488
rect 14139 20485 14151 20519
rect 14384 20516 14412 20544
rect 20364 20516 20392 20544
rect 20640 20516 20668 20547
rect 21450 20544 21456 20596
rect 21508 20544 21514 20596
rect 21821 20587 21879 20593
rect 21821 20553 21833 20587
rect 21867 20584 21879 20587
rect 21867 20556 22324 20584
rect 21867 20553 21879 20556
rect 21821 20547 21879 20553
rect 14384 20488 14688 20516
rect 20364 20488 20484 20516
rect 20640 20488 21220 20516
rect 14093 20479 14151 20485
rect 14660 20472 14688 20488
rect 14660 20467 14713 20472
rect 14660 20461 14761 20467
rect 7742 20408 7748 20460
rect 7800 20448 7806 20460
rect 7835 20451 7893 20457
rect 7835 20448 7847 20451
rect 7800 20420 7847 20448
rect 7800 20408 7806 20420
rect 7835 20417 7847 20420
rect 7881 20417 7893 20451
rect 7835 20411 7893 20417
rect 12342 20408 12348 20460
rect 12400 20408 12406 20460
rect 13170 20408 13176 20460
rect 13228 20448 13234 20460
rect 13265 20451 13323 20457
rect 13265 20448 13277 20451
rect 13228 20420 13277 20448
rect 13228 20408 13234 20420
rect 13265 20417 13277 20420
rect 13311 20417 13323 20451
rect 13265 20411 13323 20417
rect 13354 20408 13360 20460
rect 13412 20408 13418 20460
rect 13725 20451 13783 20457
rect 13725 20417 13737 20451
rect 13771 20448 13783 20451
rect 13814 20448 13820 20460
rect 13771 20420 13820 20448
rect 13771 20417 13783 20420
rect 13725 20411 13783 20417
rect 13814 20408 13820 20420
rect 13872 20408 13878 20460
rect 14458 20408 14464 20460
rect 14516 20408 14522 20460
rect 14660 20444 14715 20461
rect 14685 20430 14715 20444
rect 14703 20427 14715 20430
rect 14749 20458 14761 20461
rect 14749 20448 14778 20458
rect 15102 20448 15108 20460
rect 14749 20427 15108 20448
rect 14703 20421 15108 20427
rect 14750 20420 15108 20421
rect 15102 20408 15108 20420
rect 15160 20408 15166 20460
rect 18874 20408 18880 20460
rect 18932 20448 18938 20460
rect 19705 20451 19763 20457
rect 19705 20448 19717 20451
rect 18932 20420 19717 20448
rect 18932 20408 18938 20420
rect 19705 20417 19717 20420
rect 19751 20417 19763 20451
rect 19705 20411 19763 20417
rect 20346 20408 20352 20460
rect 20404 20408 20410 20460
rect 20456 20448 20484 20488
rect 21192 20457 21220 20488
rect 20809 20451 20867 20457
rect 20809 20448 20821 20451
rect 20456 20420 20821 20448
rect 20809 20417 20821 20420
rect 20855 20417 20867 20451
rect 20809 20411 20867 20417
rect 21177 20451 21235 20457
rect 21177 20417 21189 20451
rect 21223 20417 21235 20451
rect 21468 20448 21496 20544
rect 22005 20451 22063 20457
rect 22005 20448 22017 20451
rect 21468 20420 22017 20448
rect 21177 20411 21235 20417
rect 22005 20417 22017 20420
rect 22051 20417 22063 20451
rect 22005 20411 22063 20417
rect 22094 20408 22100 20460
rect 22152 20408 22158 20460
rect 22296 20457 22324 20556
rect 22281 20451 22339 20457
rect 22281 20417 22293 20451
rect 22327 20417 22339 20451
rect 23075 20451 23133 20457
rect 23075 20448 23087 20451
rect 22281 20411 22339 20417
rect 22572 20420 23087 20448
rect 7561 20383 7619 20389
rect 7561 20380 7573 20383
rect 7248 20352 7573 20380
rect 7248 20340 7254 20352
rect 7561 20349 7573 20352
rect 7607 20349 7619 20383
rect 7561 20343 7619 20349
rect 8294 20340 8300 20392
rect 8352 20380 8358 20392
rect 11514 20380 11520 20392
rect 8352 20352 11520 20380
rect 8352 20340 8358 20352
rect 11514 20340 11520 20352
rect 11572 20340 11578 20392
rect 13446 20340 13452 20392
rect 13504 20340 13510 20392
rect 14274 20340 14280 20392
rect 14332 20340 14338 20392
rect 14292 20312 14320 20340
rect 14458 20312 14464 20324
rect 14292 20284 14464 20312
rect 14458 20272 14464 20284
rect 14516 20272 14522 20324
rect 15120 20312 15148 20408
rect 15194 20340 15200 20392
rect 15252 20380 15258 20392
rect 22572 20380 22600 20420
rect 23075 20417 23087 20420
rect 23121 20417 23133 20451
rect 23075 20411 23133 20417
rect 15252 20352 22600 20380
rect 22833 20383 22891 20389
rect 15252 20340 15258 20352
rect 22833 20349 22845 20383
rect 22879 20349 22891 20383
rect 22833 20343 22891 20349
rect 20254 20312 20260 20324
rect 15120 20284 20260 20312
rect 20254 20272 20260 20284
rect 20312 20272 20318 20324
rect 20714 20272 20720 20324
rect 20772 20312 20778 20324
rect 22370 20312 22376 20324
rect 20772 20284 22376 20312
rect 20772 20272 20778 20284
rect 22370 20272 22376 20284
rect 22428 20312 22434 20324
rect 22554 20312 22560 20324
rect 22428 20284 22560 20312
rect 22428 20272 22434 20284
rect 22554 20272 22560 20284
rect 22612 20312 22618 20324
rect 22848 20312 22876 20343
rect 22612 20284 22876 20312
rect 22612 20272 22618 20284
rect 8294 20244 8300 20256
rect 1360 20216 8300 20244
rect 1360 20204 1366 20216
rect 8294 20204 8300 20216
rect 8352 20204 8358 20256
rect 8570 20204 8576 20256
rect 8628 20204 8634 20256
rect 11146 20204 11152 20256
rect 11204 20244 11210 20256
rect 11885 20247 11943 20253
rect 11885 20244 11897 20247
rect 11204 20216 11897 20244
rect 11204 20204 11210 20216
rect 11885 20213 11897 20216
rect 11931 20213 11943 20247
rect 11885 20207 11943 20213
rect 12526 20204 12532 20256
rect 12584 20204 12590 20256
rect 14274 20204 14280 20256
rect 14332 20204 14338 20256
rect 15378 20204 15384 20256
rect 15436 20244 15442 20256
rect 15473 20247 15531 20253
rect 15473 20244 15485 20247
rect 15436 20216 15485 20244
rect 15436 20204 15442 20216
rect 15473 20213 15485 20216
rect 15519 20213 15531 20247
rect 15473 20207 15531 20213
rect 16022 20204 16028 20256
rect 16080 20204 16086 20256
rect 19794 20204 19800 20256
rect 19852 20204 19858 20256
rect 20162 20204 20168 20256
rect 20220 20204 20226 20256
rect 21269 20247 21327 20253
rect 21269 20213 21281 20247
rect 21315 20244 21327 20247
rect 21358 20244 21364 20256
rect 21315 20216 21364 20244
rect 21315 20213 21327 20216
rect 21269 20207 21327 20213
rect 21358 20204 21364 20216
rect 21416 20204 21422 20256
rect 22189 20247 22247 20253
rect 22189 20213 22201 20247
rect 22235 20244 22247 20247
rect 22278 20244 22284 20256
rect 22235 20216 22284 20244
rect 22235 20213 22247 20216
rect 22189 20207 22247 20213
rect 22278 20204 22284 20216
rect 22336 20204 22342 20256
rect 23842 20204 23848 20256
rect 23900 20204 23906 20256
rect 1104 20154 24564 20176
rect 1104 20102 3882 20154
rect 3934 20102 3946 20154
rect 3998 20102 4010 20154
rect 4062 20102 4074 20154
rect 4126 20102 4138 20154
rect 4190 20102 9747 20154
rect 9799 20102 9811 20154
rect 9863 20102 9875 20154
rect 9927 20102 9939 20154
rect 9991 20102 10003 20154
rect 10055 20102 15612 20154
rect 15664 20102 15676 20154
rect 15728 20102 15740 20154
rect 15792 20102 15804 20154
rect 15856 20102 15868 20154
rect 15920 20102 21477 20154
rect 21529 20102 21541 20154
rect 21593 20102 21605 20154
rect 21657 20102 21669 20154
rect 21721 20102 21733 20154
rect 21785 20102 24564 20154
rect 1104 20080 24564 20102
rect 1210 20000 1216 20052
rect 1268 20000 1274 20052
rect 2406 20040 2412 20052
rect 1964 20012 2412 20040
rect 1228 19904 1256 20000
rect 1670 19932 1676 19984
rect 1728 19932 1734 19984
rect 1964 19913 1992 20012
rect 2406 20000 2412 20012
rect 2464 20000 2470 20052
rect 2682 20000 2688 20052
rect 2740 20040 2746 20052
rect 2961 20043 3019 20049
rect 2961 20040 2973 20043
rect 2740 20012 2973 20040
rect 2740 20000 2746 20012
rect 2961 20009 2973 20012
rect 3007 20009 3019 20043
rect 2961 20003 3019 20009
rect 3050 20000 3056 20052
rect 3108 20040 3114 20052
rect 3513 20043 3571 20049
rect 3513 20040 3525 20043
rect 3108 20012 3525 20040
rect 3108 20000 3114 20012
rect 3513 20009 3525 20012
rect 3559 20040 3571 20043
rect 4062 20040 4068 20052
rect 3559 20012 4068 20040
rect 3559 20009 3571 20012
rect 3513 20003 3571 20009
rect 4062 20000 4068 20012
rect 4120 20000 4126 20052
rect 4172 20012 6500 20040
rect 3234 19932 3240 19984
rect 3292 19972 3298 19984
rect 4172 19972 4200 20012
rect 3292 19944 4200 19972
rect 3292 19932 3298 19944
rect 1949 19907 2007 19913
rect 1228 19876 1900 19904
rect 750 19796 756 19848
rect 808 19836 814 19848
rect 1489 19839 1547 19845
rect 1489 19836 1501 19839
rect 808 19808 1501 19836
rect 808 19796 814 19808
rect 1489 19805 1501 19808
rect 1535 19805 1547 19839
rect 1872 19836 1900 19876
rect 1949 19873 1961 19907
rect 1995 19873 2007 19907
rect 1949 19867 2007 19873
rect 2682 19864 2688 19916
rect 2740 19904 2746 19916
rect 2740 19876 3464 19904
rect 2740 19864 2746 19876
rect 2130 19836 2136 19848
rect 1872 19808 2136 19836
rect 1489 19799 1547 19805
rect 2130 19796 2136 19808
rect 2188 19845 2194 19848
rect 2188 19839 2249 19845
rect 2188 19805 2203 19839
rect 2237 19805 2249 19839
rect 3329 19839 3387 19845
rect 3329 19836 3341 19839
rect 2188 19799 2249 19805
rect 2746 19808 3341 19836
rect 2188 19796 2194 19799
rect 1302 19728 1308 19780
rect 1360 19768 1366 19780
rect 2746 19768 2774 19808
rect 3329 19805 3341 19808
rect 3375 19805 3387 19839
rect 3436 19836 3464 19876
rect 4890 19864 4896 19916
rect 4948 19904 4954 19916
rect 5350 19904 5356 19916
rect 4948 19876 5356 19904
rect 4948 19864 4954 19876
rect 5350 19864 5356 19876
rect 5408 19904 5414 19916
rect 5408 19876 5856 19904
rect 5408 19864 5414 19876
rect 5828 19845 5856 19876
rect 5813 19839 5871 19845
rect 3436 19808 5488 19836
rect 3329 19799 3387 19805
rect 5350 19768 5356 19780
rect 1360 19740 2774 19768
rect 3436 19740 5356 19768
rect 1360 19728 1366 19740
rect 2222 19660 2228 19712
rect 2280 19700 2286 19712
rect 3436 19700 3464 19740
rect 5350 19728 5356 19740
rect 5408 19728 5414 19780
rect 2280 19672 3464 19700
rect 5460 19700 5488 19808
rect 5813 19805 5825 19839
rect 5859 19836 5871 19839
rect 6472 19836 6500 20012
rect 8570 20000 8576 20052
rect 8628 20000 8634 20052
rect 8665 20043 8723 20049
rect 8665 20009 8677 20043
rect 8711 20040 8723 20043
rect 8754 20040 8760 20052
rect 8711 20012 8760 20040
rect 8711 20009 8723 20012
rect 8665 20003 8723 20009
rect 8754 20000 8760 20012
rect 8812 20040 8818 20052
rect 8938 20040 8944 20052
rect 8812 20012 8944 20040
rect 8812 20000 8818 20012
rect 8938 20000 8944 20012
rect 8996 20000 9002 20052
rect 12250 20000 12256 20052
rect 12308 20040 12314 20052
rect 12308 20012 13308 20040
rect 12308 20000 12314 20012
rect 7926 19864 7932 19916
rect 7984 19864 7990 19916
rect 5859 19808 5948 19836
rect 5859 19805 5871 19808
rect 5813 19799 5871 19805
rect 5920 19780 5948 19808
rect 6071 19809 6129 19815
rect 5902 19728 5908 19780
rect 5960 19728 5966 19780
rect 6071 19775 6083 19809
rect 6117 19806 6129 19809
rect 6472 19808 7512 19836
rect 6117 19775 6130 19806
rect 6071 19769 6130 19775
rect 6102 19768 6130 19769
rect 6454 19768 6460 19780
rect 6102 19740 6460 19768
rect 6454 19728 6460 19740
rect 6512 19728 6518 19780
rect 6564 19740 6960 19768
rect 6564 19700 6592 19740
rect 5460 19672 6592 19700
rect 2280 19660 2286 19672
rect 6822 19660 6828 19712
rect 6880 19660 6886 19712
rect 6932 19700 6960 19740
rect 7374 19728 7380 19780
rect 7432 19728 7438 19780
rect 7484 19768 7512 19808
rect 7650 19796 7656 19848
rect 7708 19796 7714 19848
rect 7745 19839 7803 19845
rect 7745 19805 7757 19839
rect 7791 19836 7803 19839
rect 8588 19836 8616 20000
rect 10321 19975 10379 19981
rect 10321 19941 10333 19975
rect 10367 19972 10379 19975
rect 13280 19972 13308 20012
rect 13354 20000 13360 20052
rect 13412 20040 13418 20052
rect 13633 20043 13691 20049
rect 13633 20040 13645 20043
rect 13412 20012 13645 20040
rect 13412 20000 13418 20012
rect 13633 20009 13645 20012
rect 13679 20009 13691 20043
rect 13633 20003 13691 20009
rect 13814 20000 13820 20052
rect 13872 20040 13878 20052
rect 13872 20012 14872 20040
rect 13872 20000 13878 20012
rect 10367 19944 10732 19972
rect 13280 19944 14688 19972
rect 10367 19941 10379 19944
rect 10321 19935 10379 19941
rect 10704 19890 10732 19944
rect 12066 19864 12072 19916
rect 12124 19904 12130 19916
rect 14660 19913 14688 19944
rect 14844 19913 14872 20012
rect 18874 20000 18880 20052
rect 18932 20000 18938 20052
rect 19978 20040 19984 20052
rect 19260 20012 19984 20040
rect 15289 19975 15347 19981
rect 15289 19941 15301 19975
rect 15335 19972 15347 19975
rect 15378 19972 15384 19984
rect 15335 19944 15384 19972
rect 15335 19941 15347 19944
rect 15289 19935 15347 19941
rect 15378 19932 15384 19944
rect 15436 19932 15442 19984
rect 19260 19972 19288 20012
rect 19978 20000 19984 20012
rect 20036 20000 20042 20052
rect 20254 20000 20260 20052
rect 20312 20000 20318 20052
rect 20346 20000 20352 20052
rect 20404 20040 20410 20052
rect 20625 20043 20683 20049
rect 20625 20040 20637 20043
rect 20404 20012 20637 20040
rect 20404 20000 20410 20012
rect 20625 20009 20637 20012
rect 20671 20009 20683 20043
rect 22094 20040 22100 20052
rect 20625 20003 20683 20009
rect 22066 20000 22100 20040
rect 22152 20000 22158 20052
rect 22278 20000 22284 20052
rect 22336 20000 22342 20052
rect 23750 20000 23756 20052
rect 23808 20000 23814 20052
rect 24026 20000 24032 20052
rect 24084 20000 24090 20052
rect 16408 19944 19288 19972
rect 12621 19907 12679 19913
rect 12621 19904 12633 19907
rect 12124 19876 12633 19904
rect 12124 19864 12130 19876
rect 12621 19873 12633 19876
rect 12667 19873 12679 19907
rect 12621 19867 12679 19873
rect 14645 19907 14703 19913
rect 14645 19873 14657 19907
rect 14691 19873 14703 19907
rect 14645 19867 14703 19873
rect 14829 19907 14887 19913
rect 14829 19873 14841 19907
rect 14875 19873 14887 19907
rect 14829 19867 14887 19873
rect 15565 19907 15623 19913
rect 15565 19873 15577 19907
rect 15611 19904 15623 19907
rect 16022 19904 16028 19916
rect 15611 19876 16028 19904
rect 15611 19873 15623 19876
rect 15565 19867 15623 19873
rect 16022 19864 16028 19876
rect 16080 19864 16086 19916
rect 7791 19808 8616 19836
rect 7791 19805 7803 19808
rect 7745 19799 7803 19805
rect 9306 19796 9312 19848
rect 9364 19796 9370 19848
rect 9582 19845 9588 19848
rect 9567 19839 9588 19845
rect 9567 19805 9579 19839
rect 9567 19799 9588 19805
rect 9582 19796 9588 19799
rect 9640 19796 9646 19848
rect 11146 19796 11152 19848
rect 11204 19796 11210 19848
rect 11606 19796 11612 19848
rect 11664 19796 11670 19848
rect 12863 19839 12921 19845
rect 12863 19836 12875 19839
rect 12728 19808 12875 19836
rect 7834 19768 7840 19780
rect 7484 19740 7840 19768
rect 7834 19728 7840 19740
rect 7892 19728 7898 19780
rect 8110 19728 8116 19780
rect 8168 19728 8174 19780
rect 8294 19728 8300 19780
rect 8352 19768 8358 19780
rect 8481 19771 8539 19777
rect 8481 19768 8493 19771
rect 8352 19740 8493 19768
rect 8352 19728 8358 19740
rect 8481 19737 8493 19740
rect 8527 19737 8539 19771
rect 8481 19731 8539 19737
rect 10134 19728 10140 19780
rect 10192 19768 10198 19780
rect 10192 19740 11008 19768
rect 10192 19728 10198 19740
rect 9582 19700 9588 19712
rect 6932 19672 9588 19700
rect 9582 19660 9588 19672
rect 9640 19660 9646 19712
rect 10502 19660 10508 19712
rect 10560 19700 10566 19712
rect 10873 19703 10931 19709
rect 10873 19700 10885 19703
rect 10560 19672 10885 19700
rect 10560 19660 10566 19672
rect 10873 19669 10885 19672
rect 10919 19669 10931 19703
rect 10980 19700 11008 19740
rect 11238 19728 11244 19780
rect 11296 19728 11302 19780
rect 11977 19771 12035 19777
rect 11977 19737 11989 19771
rect 12023 19737 12035 19771
rect 11977 19731 12035 19737
rect 11992 19700 12020 19731
rect 12250 19728 12256 19780
rect 12308 19768 12314 19780
rect 12728 19768 12756 19808
rect 12863 19805 12875 19808
rect 12909 19805 12921 19839
rect 12863 19799 12921 19805
rect 15654 19796 15660 19848
rect 15712 19845 15718 19848
rect 15712 19839 15740 19845
rect 15728 19805 15740 19839
rect 15712 19799 15740 19805
rect 15712 19796 15718 19799
rect 15838 19796 15844 19848
rect 15896 19796 15902 19848
rect 12308 19740 12756 19768
rect 12308 19728 12314 19740
rect 10980 19672 12020 19700
rect 12161 19703 12219 19709
rect 10873 19663 10931 19669
rect 12161 19669 12173 19703
rect 12207 19700 12219 19703
rect 16408 19700 16436 19944
rect 19242 19904 19248 19916
rect 18892 19876 19248 19904
rect 18892 19848 18920 19876
rect 19242 19864 19248 19876
rect 19300 19864 19306 19916
rect 18874 19796 18880 19848
rect 18932 19796 18938 19848
rect 19058 19796 19064 19848
rect 19116 19836 19122 19848
rect 19501 19839 19559 19845
rect 19501 19836 19513 19839
rect 19116 19808 19513 19836
rect 19116 19796 19122 19808
rect 19501 19805 19513 19808
rect 19547 19805 19559 19839
rect 20272 19836 20300 20000
rect 21729 19975 21787 19981
rect 21729 19941 21741 19975
rect 21775 19972 21787 19975
rect 22066 19972 22094 20000
rect 21775 19944 22094 19972
rect 21775 19941 21787 19944
rect 21729 19935 21787 19941
rect 20622 19864 20628 19916
rect 20680 19904 20686 19916
rect 20717 19907 20775 19913
rect 20717 19904 20729 19907
rect 20680 19876 20729 19904
rect 20680 19864 20686 19876
rect 20717 19873 20729 19876
rect 20763 19873 20775 19907
rect 22066 19904 22094 19944
rect 22296 19904 22324 20000
rect 23201 19975 23259 19981
rect 23201 19941 23213 19975
rect 23247 19972 23259 19975
rect 23247 19944 24256 19972
rect 23247 19941 23259 19944
rect 23201 19935 23259 19941
rect 22373 19907 22431 19913
rect 22373 19904 22385 19907
rect 22066 19876 22140 19904
rect 22296 19876 22385 19904
rect 20717 19867 20775 19873
rect 20959 19839 21017 19845
rect 20959 19836 20971 19839
rect 20272 19808 20971 19836
rect 19501 19799 19559 19805
rect 20959 19805 20971 19808
rect 21005 19805 21017 19839
rect 20959 19799 21017 19805
rect 21358 19796 21364 19848
rect 21416 19796 21422 19848
rect 22112 19845 22140 19876
rect 22373 19873 22385 19876
rect 22419 19873 22431 19907
rect 23842 19904 23848 19916
rect 22373 19867 22431 19873
rect 23124 19876 23848 19904
rect 23124 19845 23152 19876
rect 23842 19864 23848 19876
rect 23900 19904 23906 19916
rect 24228 19913 24256 19944
rect 24213 19907 24271 19913
rect 23900 19876 23980 19904
rect 23900 19864 23906 19876
rect 22097 19839 22155 19845
rect 22097 19805 22109 19839
rect 22143 19805 22155 19839
rect 22097 19799 22155 19805
rect 22189 19839 22247 19845
rect 22189 19805 22201 19839
rect 22235 19805 22247 19839
rect 22189 19799 22247 19805
rect 23109 19839 23167 19845
rect 23109 19805 23121 19839
rect 23155 19805 23167 19839
rect 23109 19799 23167 19805
rect 23293 19839 23351 19845
rect 23293 19805 23305 19839
rect 23339 19836 23351 19839
rect 23382 19836 23388 19848
rect 23339 19808 23388 19836
rect 23339 19805 23351 19808
rect 23293 19799 23351 19805
rect 21376 19768 21404 19796
rect 22204 19768 22232 19799
rect 23382 19796 23388 19808
rect 23440 19796 23446 19848
rect 23952 19845 23980 19876
rect 24213 19873 24225 19907
rect 24259 19873 24271 19907
rect 24213 19867 24271 19873
rect 23477 19839 23535 19845
rect 23477 19805 23489 19839
rect 23523 19836 23535 19839
rect 23937 19839 23995 19845
rect 23523 19808 23704 19836
rect 23523 19805 23535 19808
rect 23477 19799 23535 19805
rect 16500 19740 19288 19768
rect 21376 19740 22232 19768
rect 22373 19771 22431 19777
rect 16500 19709 16528 19740
rect 12207 19672 16436 19700
rect 16485 19703 16543 19709
rect 12207 19669 12219 19672
rect 12161 19663 12219 19669
rect 16485 19669 16497 19703
rect 16531 19669 16543 19703
rect 19260 19700 19288 19740
rect 22373 19737 22385 19771
rect 22419 19768 22431 19771
rect 23566 19768 23572 19780
rect 22419 19740 23572 19768
rect 22419 19737 22431 19740
rect 22373 19731 22431 19737
rect 23566 19728 23572 19740
rect 23624 19728 23630 19780
rect 22094 19700 22100 19712
rect 19260 19672 22100 19700
rect 16485 19663 16543 19669
rect 22094 19660 22100 19672
rect 22152 19660 22158 19712
rect 22646 19660 22652 19712
rect 22704 19700 22710 19712
rect 23676 19700 23704 19808
rect 23937 19805 23949 19839
rect 23983 19805 23995 19839
rect 23937 19799 23995 19805
rect 22704 19672 23704 19700
rect 22704 19660 22710 19672
rect 24210 19660 24216 19712
rect 24268 19660 24274 19712
rect 1104 19610 24723 19632
rect 1104 19558 6814 19610
rect 6866 19558 6878 19610
rect 6930 19558 6942 19610
rect 6994 19558 7006 19610
rect 7058 19558 7070 19610
rect 7122 19558 12679 19610
rect 12731 19558 12743 19610
rect 12795 19558 12807 19610
rect 12859 19558 12871 19610
rect 12923 19558 12935 19610
rect 12987 19558 18544 19610
rect 18596 19558 18608 19610
rect 18660 19558 18672 19610
rect 18724 19558 18736 19610
rect 18788 19558 18800 19610
rect 18852 19558 24409 19610
rect 24461 19558 24473 19610
rect 24525 19558 24537 19610
rect 24589 19558 24601 19610
rect 24653 19558 24665 19610
rect 24717 19558 24723 19610
rect 1104 19536 24723 19558
rect 658 19456 664 19508
rect 716 19496 722 19508
rect 7650 19496 7656 19508
rect 716 19468 3614 19496
rect 716 19456 722 19468
rect 1854 19388 1860 19440
rect 1912 19428 1918 19440
rect 2130 19428 2136 19440
rect 1912 19400 2136 19428
rect 1912 19388 1918 19400
rect 2130 19388 2136 19400
rect 2188 19388 2194 19440
rect 2222 19388 2228 19440
rect 2280 19388 2286 19440
rect 3234 19428 3240 19440
rect 2976 19400 3240 19428
rect 1671 19363 1729 19369
rect 1671 19329 1683 19363
rect 1717 19360 1729 19363
rect 2240 19360 2268 19388
rect 1717 19332 2268 19360
rect 1717 19329 1729 19332
rect 1671 19323 1729 19329
rect 2774 19320 2780 19372
rect 2832 19320 2838 19372
rect 1397 19295 1455 19301
rect 1397 19261 1409 19295
rect 1443 19261 1455 19295
rect 1397 19255 1455 19261
rect 1412 19224 1440 19255
rect 2976 19233 3004 19400
rect 3234 19388 3240 19400
rect 3292 19388 3298 19440
rect 3586 19428 3614 19468
rect 7484 19468 7656 19496
rect 7484 19440 7512 19468
rect 7650 19456 7656 19468
rect 7708 19456 7714 19508
rect 7834 19456 7840 19508
rect 7892 19456 7898 19508
rect 7926 19456 7932 19508
rect 7984 19456 7990 19508
rect 8018 19468 13400 19496
rect 4522 19428 4528 19440
rect 3586 19400 4528 19428
rect 3586 19370 3614 19400
rect 4522 19388 4528 19400
rect 4580 19428 4586 19440
rect 4580 19400 4844 19428
rect 4580 19388 4586 19400
rect 3526 19369 3614 19370
rect 3511 19363 3614 19369
rect 3511 19329 3523 19363
rect 3557 19342 3614 19363
rect 3557 19329 3569 19342
rect 3511 19323 3569 19329
rect 3050 19252 3056 19304
rect 3108 19292 3114 19304
rect 3237 19295 3295 19301
rect 3237 19292 3249 19295
rect 3108 19264 3249 19292
rect 3108 19252 3114 19264
rect 3237 19261 3249 19264
rect 3283 19261 3295 19295
rect 3237 19255 3295 19261
rect 2961 19227 3019 19233
rect 1412 19196 1532 19224
rect 1504 19168 1532 19196
rect 2961 19193 2973 19227
rect 3007 19193 3019 19227
rect 2961 19187 3019 19193
rect 1486 19116 1492 19168
rect 1544 19116 1550 19168
rect 2406 19116 2412 19168
rect 2464 19116 2470 19168
rect 4246 19116 4252 19168
rect 4304 19116 4310 19168
rect 4816 19156 4844 19400
rect 5552 19400 7310 19428
rect 4890 19320 4896 19372
rect 4948 19320 4954 19372
rect 5074 19320 5080 19372
rect 5132 19360 5138 19372
rect 5167 19363 5225 19369
rect 5167 19360 5179 19363
rect 5132 19332 5179 19360
rect 5132 19320 5138 19332
rect 5167 19329 5179 19332
rect 5213 19329 5225 19363
rect 5167 19323 5225 19329
rect 5552 19156 5580 19400
rect 5626 19320 5632 19372
rect 5684 19360 5690 19372
rect 6638 19360 6644 19372
rect 5684 19332 6644 19360
rect 5684 19320 5690 19332
rect 6638 19320 6644 19332
rect 6696 19320 6702 19372
rect 6914 19320 6920 19372
rect 6972 19320 6978 19372
rect 7159 19363 7217 19369
rect 7159 19329 7171 19363
rect 7205 19360 7217 19363
rect 7282 19360 7310 19400
rect 7466 19388 7472 19440
rect 7524 19388 7530 19440
rect 7852 19428 7880 19456
rect 8018 19428 8046 19468
rect 9306 19428 9312 19440
rect 7852 19400 8046 19428
rect 8680 19400 9312 19428
rect 8680 19369 8708 19400
rect 9306 19388 9312 19400
rect 9364 19388 9370 19440
rect 9490 19388 9496 19440
rect 9548 19388 9554 19440
rect 9582 19388 9588 19440
rect 9640 19428 9646 19440
rect 9640 19400 12664 19428
rect 9640 19388 9646 19400
rect 8665 19363 8723 19369
rect 7205 19332 7972 19360
rect 7205 19329 7217 19332
rect 7159 19323 7217 19329
rect 7944 19236 7972 19332
rect 8665 19329 8677 19363
rect 8711 19329 8723 19363
rect 8665 19323 8723 19329
rect 8939 19363 8997 19369
rect 8939 19329 8951 19363
rect 8985 19360 8997 19363
rect 9508 19360 9536 19388
rect 8985 19332 9536 19360
rect 8985 19329 8997 19332
rect 8939 19323 8997 19329
rect 12066 19320 12072 19372
rect 12124 19360 12130 19372
rect 12437 19363 12495 19369
rect 12437 19360 12449 19363
rect 12124 19332 12449 19360
rect 12124 19320 12130 19332
rect 12437 19329 12449 19332
rect 12483 19329 12495 19363
rect 12636 19360 12664 19400
rect 12695 19393 12753 19399
rect 12695 19360 12707 19393
rect 12636 19359 12707 19360
rect 12741 19360 12753 19393
rect 13170 19388 13176 19440
rect 13228 19388 13234 19440
rect 13372 19428 13400 19468
rect 13446 19456 13452 19508
rect 13504 19456 13510 19508
rect 15838 19456 15844 19508
rect 15896 19496 15902 19508
rect 15933 19499 15991 19505
rect 15933 19496 15945 19499
rect 15896 19468 15945 19496
rect 15896 19456 15902 19468
rect 15933 19465 15945 19468
rect 15979 19465 15991 19499
rect 15933 19459 15991 19465
rect 16666 19456 16672 19508
rect 16724 19456 16730 19508
rect 16850 19456 16856 19508
rect 16908 19456 16914 19508
rect 18138 19456 18144 19508
rect 18196 19496 18202 19508
rect 18196 19468 18451 19496
rect 18196 19456 18202 19468
rect 16684 19428 16712 19456
rect 13372 19400 16712 19428
rect 13188 19360 13216 19388
rect 13464 19372 13492 19400
rect 12741 19359 13216 19360
rect 12636 19332 13216 19359
rect 12437 19323 12495 19329
rect 13446 19320 13452 19372
rect 13504 19320 13510 19372
rect 14921 19363 14979 19369
rect 14921 19360 14933 19363
rect 14292 19332 14933 19360
rect 9398 19252 9404 19304
rect 9456 19292 9462 19304
rect 10229 19295 10287 19301
rect 10229 19292 10241 19295
rect 9456 19264 10241 19292
rect 9456 19252 9462 19264
rect 10229 19261 10241 19264
rect 10275 19261 10287 19295
rect 10229 19255 10287 19261
rect 14292 19236 14320 19332
rect 14921 19329 14933 19332
rect 14967 19329 14979 19363
rect 14921 19323 14979 19329
rect 15195 19363 15253 19369
rect 15195 19329 15207 19363
rect 15241 19360 15253 19363
rect 15241 19332 15608 19360
rect 15241 19329 15253 19332
rect 15195 19323 15253 19329
rect 15580 19292 15608 19332
rect 15654 19320 15660 19372
rect 15712 19360 15718 19372
rect 16390 19360 16396 19372
rect 15712 19332 16396 19360
rect 15712 19320 15718 19332
rect 16390 19320 16396 19332
rect 16448 19320 16454 19372
rect 16206 19292 16212 19304
rect 15580 19264 16212 19292
rect 16206 19252 16212 19264
rect 16264 19252 16270 19304
rect 16592 19292 16620 19400
rect 16669 19363 16727 19369
rect 16669 19329 16681 19363
rect 16715 19360 16727 19363
rect 16868 19360 16896 19456
rect 16715 19332 16896 19360
rect 17589 19363 17647 19369
rect 16715 19329 16727 19332
rect 16669 19323 16727 19329
rect 17589 19329 17601 19363
rect 17635 19329 17647 19363
rect 18423 19360 18451 19468
rect 18874 19456 18880 19508
rect 18932 19456 18938 19508
rect 20622 19456 20628 19508
rect 20680 19496 20686 19508
rect 22646 19496 22652 19508
rect 20680 19468 22652 19496
rect 20680 19456 20686 19468
rect 22646 19456 22652 19468
rect 22704 19456 22710 19508
rect 23201 19499 23259 19505
rect 23201 19465 23213 19499
rect 23247 19465 23259 19499
rect 23201 19459 23259 19465
rect 18892 19428 18920 19456
rect 22186 19428 22192 19440
rect 18892 19400 22192 19428
rect 18843 19363 18901 19369
rect 18843 19360 18855 19363
rect 18423 19332 18855 19360
rect 17589 19323 17647 19329
rect 18843 19329 18855 19332
rect 18889 19329 18901 19363
rect 18843 19323 18901 19329
rect 16853 19295 16911 19301
rect 16853 19292 16865 19295
rect 16592 19264 16865 19292
rect 16853 19261 16865 19264
rect 16899 19261 16911 19295
rect 17034 19292 17040 19304
rect 16853 19255 16911 19261
rect 16942 19264 17040 19292
rect 5626 19184 5632 19236
rect 5684 19224 5690 19236
rect 6362 19224 6368 19236
rect 5684 19196 6368 19224
rect 5684 19184 5690 19196
rect 6362 19184 6368 19196
rect 6420 19184 6426 19236
rect 6546 19184 6552 19236
rect 6604 19224 6610 19236
rect 6730 19224 6736 19236
rect 6604 19196 6736 19224
rect 6604 19184 6610 19196
rect 6730 19184 6736 19196
rect 6788 19184 6794 19236
rect 7926 19184 7932 19236
rect 7984 19184 7990 19236
rect 9324 19196 12572 19224
rect 4816 19128 5580 19156
rect 5902 19116 5908 19168
rect 5960 19116 5966 19168
rect 6086 19116 6092 19168
rect 6144 19156 6150 19168
rect 9324 19156 9352 19196
rect 6144 19128 9352 19156
rect 6144 19116 6150 19128
rect 9674 19116 9680 19168
rect 9732 19116 9738 19168
rect 10962 19116 10968 19168
rect 11020 19156 11026 19168
rect 12434 19156 12440 19168
rect 11020 19128 12440 19156
rect 11020 19116 11026 19128
rect 12434 19116 12440 19128
rect 12492 19116 12498 19168
rect 12544 19156 12572 19196
rect 14274 19184 14280 19236
rect 14332 19184 14338 19236
rect 16482 19184 16488 19236
rect 16540 19224 16546 19236
rect 16942 19224 16970 19264
rect 17034 19252 17040 19264
rect 17092 19292 17098 19304
rect 17604 19292 17632 19323
rect 19518 19320 19524 19372
rect 19576 19360 19582 19372
rect 19576 19332 19840 19360
rect 19576 19320 19582 19332
rect 17092 19264 17632 19292
rect 17092 19252 17098 19264
rect 17678 19252 17684 19304
rect 17736 19301 17742 19304
rect 17736 19295 17764 19301
rect 17752 19261 17764 19295
rect 17736 19255 17764 19261
rect 17736 19252 17742 19255
rect 17862 19252 17868 19304
rect 17920 19252 17926 19304
rect 18598 19252 18604 19304
rect 18656 19252 18662 19304
rect 19812 19292 19840 19332
rect 19886 19320 19892 19372
rect 19944 19360 19950 19372
rect 20223 19363 20281 19369
rect 20223 19360 20235 19363
rect 19944 19332 20235 19360
rect 19944 19320 19950 19332
rect 20223 19329 20235 19332
rect 20269 19329 20281 19363
rect 20223 19323 20281 19329
rect 20346 19320 20352 19372
rect 20404 19360 20410 19372
rect 21266 19360 21272 19372
rect 20404 19332 21272 19360
rect 20404 19320 20410 19332
rect 21266 19320 21272 19332
rect 21324 19320 21330 19372
rect 21836 19369 21864 19400
rect 22186 19388 22192 19400
rect 22244 19388 22250 19440
rect 22094 19369 22100 19372
rect 21821 19363 21879 19369
rect 21821 19329 21833 19363
rect 21867 19329 21879 19363
rect 21821 19323 21879 19329
rect 22088 19323 22100 19369
rect 22152 19360 22158 19372
rect 22370 19360 22376 19372
rect 22152 19332 22376 19360
rect 22094 19320 22100 19323
rect 22152 19320 22158 19332
rect 22370 19320 22376 19332
rect 22428 19320 22434 19372
rect 23216 19360 23244 19459
rect 23566 19456 23572 19508
rect 23624 19456 23630 19508
rect 23584 19428 23612 19456
rect 23661 19431 23719 19437
rect 23661 19428 23673 19431
rect 23584 19400 23673 19428
rect 23661 19397 23673 19400
rect 23707 19397 23719 19431
rect 23661 19391 23719 19397
rect 23477 19363 23535 19369
rect 23477 19360 23489 19363
rect 23216 19332 23489 19360
rect 23477 19329 23489 19332
rect 23523 19329 23535 19363
rect 23477 19323 23535 19329
rect 19981 19295 20039 19301
rect 19981 19292 19993 19295
rect 19812 19264 19993 19292
rect 19981 19261 19993 19264
rect 20027 19261 20039 19295
rect 19981 19255 20039 19261
rect 16540 19196 16970 19224
rect 16540 19184 16546 19196
rect 17310 19184 17316 19236
rect 17368 19184 17374 19236
rect 14366 19156 14372 19168
rect 12544 19128 14372 19156
rect 14366 19116 14372 19128
rect 14424 19116 14430 19168
rect 18506 19116 18512 19168
rect 18564 19116 18570 19168
rect 19518 19116 19524 19168
rect 19576 19156 19582 19168
rect 19613 19159 19671 19165
rect 19613 19156 19625 19159
rect 19576 19128 19625 19156
rect 19576 19116 19582 19128
rect 19613 19125 19625 19128
rect 19659 19125 19671 19159
rect 19996 19156 20024 19255
rect 22830 19252 22836 19304
rect 22888 19292 22894 19304
rect 23106 19292 23112 19304
rect 22888 19264 23112 19292
rect 22888 19252 22894 19264
rect 23106 19252 23112 19264
rect 23164 19252 23170 19304
rect 20070 19156 20076 19168
rect 19996 19128 20076 19156
rect 19613 19119 19671 19125
rect 20070 19116 20076 19128
rect 20128 19116 20134 19168
rect 20990 19116 20996 19168
rect 21048 19116 21054 19168
rect 22830 19116 22836 19168
rect 22888 19156 22894 19168
rect 23293 19159 23351 19165
rect 23293 19156 23305 19159
rect 22888 19128 23305 19156
rect 22888 19116 22894 19128
rect 23293 19125 23305 19128
rect 23339 19125 23351 19159
rect 23293 19119 23351 19125
rect 23934 19116 23940 19168
rect 23992 19116 23998 19168
rect 1104 19066 24564 19088
rect 1104 19014 3882 19066
rect 3934 19014 3946 19066
rect 3998 19014 4010 19066
rect 4062 19014 4074 19066
rect 4126 19014 4138 19066
rect 4190 19014 9747 19066
rect 9799 19014 9811 19066
rect 9863 19014 9875 19066
rect 9927 19014 9939 19066
rect 9991 19014 10003 19066
rect 10055 19014 15612 19066
rect 15664 19014 15676 19066
rect 15728 19014 15740 19066
rect 15792 19014 15804 19066
rect 15856 19014 15868 19066
rect 15920 19014 21477 19066
rect 21529 19014 21541 19066
rect 21593 19014 21605 19066
rect 21657 19014 21669 19066
rect 21721 19014 21733 19066
rect 21785 19014 24564 19066
rect 1104 18992 24564 19014
rect 1581 18955 1639 18961
rect 1581 18921 1593 18955
rect 1627 18952 1639 18955
rect 4798 18952 4804 18964
rect 1627 18924 4804 18952
rect 1627 18921 1639 18924
rect 1581 18915 1639 18921
rect 4798 18912 4804 18924
rect 4856 18912 4862 18964
rect 6362 18912 6368 18964
rect 6420 18952 6426 18964
rect 7282 18952 7288 18964
rect 6420 18924 7288 18952
rect 6420 18912 6426 18924
rect 7282 18912 7288 18924
rect 7340 18912 7346 18964
rect 8754 18912 8760 18964
rect 8812 18912 8818 18964
rect 11238 18912 11244 18964
rect 11296 18952 11302 18964
rect 11885 18955 11943 18961
rect 11885 18952 11897 18955
rect 11296 18924 11897 18952
rect 11296 18912 11302 18924
rect 11885 18921 11897 18924
rect 11931 18921 11943 18955
rect 11885 18915 11943 18921
rect 12434 18912 12440 18964
rect 12492 18952 12498 18964
rect 18417 18955 18475 18961
rect 12492 18924 18092 18952
rect 12492 18912 12498 18924
rect 2317 18887 2375 18893
rect 2317 18853 2329 18887
rect 2363 18884 2375 18887
rect 2406 18884 2412 18896
rect 2363 18856 2412 18884
rect 2363 18853 2375 18856
rect 2317 18847 2375 18853
rect 2406 18844 2412 18856
rect 2464 18844 2470 18896
rect 5902 18844 5908 18896
rect 5960 18884 5966 18896
rect 5997 18887 6055 18893
rect 5997 18884 6009 18887
rect 5960 18856 6009 18884
rect 5960 18844 5966 18856
rect 5997 18853 6009 18856
rect 6043 18853 6055 18887
rect 5997 18847 6055 18853
rect 474 18776 480 18828
rect 532 18816 538 18828
rect 2710 18819 2768 18825
rect 2710 18816 2722 18819
rect 532 18788 2722 18816
rect 532 18776 538 18788
rect 2710 18785 2722 18788
rect 2756 18785 2768 18819
rect 2710 18779 2768 18785
rect 3050 18776 3056 18828
rect 3108 18816 3114 18828
rect 3602 18816 3608 18828
rect 3108 18788 3608 18816
rect 3108 18776 3114 18788
rect 3602 18776 3608 18788
rect 3660 18816 3666 18828
rect 3789 18819 3847 18825
rect 3789 18816 3801 18819
rect 3660 18788 3801 18816
rect 3660 18776 3666 18788
rect 3789 18785 3801 18788
rect 3835 18785 3847 18819
rect 3789 18779 3847 18785
rect 5258 18776 5264 18828
rect 5316 18816 5322 18828
rect 5353 18819 5411 18825
rect 5353 18816 5365 18819
rect 5316 18788 5365 18816
rect 5316 18776 5322 18788
rect 5353 18785 5365 18788
rect 5399 18785 5411 18819
rect 5353 18779 5411 18785
rect 6086 18776 6092 18828
rect 6144 18816 6150 18828
rect 6144 18788 6316 18816
rect 6144 18776 6150 18788
rect 1394 18708 1400 18760
rect 1452 18708 1458 18760
rect 1578 18708 1584 18760
rect 1636 18748 1642 18760
rect 1673 18751 1731 18757
rect 1673 18748 1685 18751
rect 1636 18720 1685 18748
rect 1636 18708 1642 18720
rect 1673 18717 1685 18720
rect 1719 18717 1731 18751
rect 1857 18751 1915 18757
rect 1857 18748 1869 18751
rect 1673 18711 1731 18717
rect 1780 18720 1869 18748
rect 1780 18612 1808 18720
rect 1857 18717 1869 18720
rect 1903 18717 1915 18751
rect 1857 18711 1915 18717
rect 2590 18708 2596 18760
rect 2648 18708 2654 18760
rect 2866 18708 2872 18760
rect 2924 18708 2930 18760
rect 4063 18751 4121 18757
rect 4063 18717 4075 18751
rect 4109 18748 4121 18751
rect 4522 18748 4528 18760
rect 4109 18720 4528 18748
rect 4109 18717 4121 18720
rect 4063 18711 4121 18717
rect 4522 18708 4528 18720
rect 4580 18708 4586 18760
rect 5442 18708 5448 18760
rect 5500 18748 5506 18760
rect 6288 18757 6316 18788
rect 6362 18776 6368 18828
rect 6420 18825 6426 18828
rect 6420 18819 6448 18825
rect 6436 18785 6448 18819
rect 6420 18779 6448 18785
rect 6420 18776 6426 18779
rect 6546 18776 6552 18828
rect 6604 18776 6610 18828
rect 5537 18751 5595 18757
rect 5537 18748 5549 18751
rect 5500 18720 5549 18748
rect 5500 18708 5506 18720
rect 5537 18717 5549 18720
rect 5583 18717 5595 18751
rect 5537 18711 5595 18717
rect 6273 18751 6331 18757
rect 6273 18717 6285 18751
rect 6319 18717 6331 18751
rect 6273 18711 6331 18717
rect 7558 18708 7564 18760
rect 7616 18748 7622 18760
rect 8570 18748 8576 18760
rect 7616 18720 8576 18748
rect 7616 18708 7622 18720
rect 8570 18708 8576 18720
rect 8628 18708 8634 18760
rect 3602 18640 3608 18692
rect 3660 18680 3666 18692
rect 8772 18680 8800 18912
rect 12452 18856 16896 18884
rect 9674 18776 9680 18828
rect 9732 18776 9738 18828
rect 9398 18708 9404 18760
rect 9456 18708 9462 18760
rect 9490 18708 9496 18760
rect 9548 18708 9554 18760
rect 9950 18757 9956 18760
rect 9907 18751 9956 18757
rect 9907 18717 9919 18751
rect 9953 18717 9956 18751
rect 9907 18711 9956 18717
rect 9950 18708 9956 18711
rect 10008 18708 10014 18760
rect 10502 18708 10508 18760
rect 10560 18748 10566 18760
rect 10873 18751 10931 18757
rect 10873 18748 10885 18751
rect 10560 18720 10885 18748
rect 10560 18708 10566 18720
rect 10873 18717 10885 18720
rect 10919 18717 10931 18751
rect 10873 18711 10931 18717
rect 11147 18751 11205 18757
rect 11147 18717 11159 18751
rect 11193 18748 11205 18751
rect 11238 18748 11244 18760
rect 11193 18720 11244 18748
rect 11193 18717 11205 18720
rect 11147 18711 11205 18717
rect 11238 18708 11244 18720
rect 11296 18748 11302 18760
rect 12250 18748 12256 18760
rect 11296 18720 12256 18748
rect 11296 18708 11302 18720
rect 12250 18708 12256 18720
rect 12308 18748 12314 18760
rect 12452 18748 12480 18856
rect 12308 18720 12480 18748
rect 12912 18788 16804 18816
rect 12308 18708 12314 18720
rect 3660 18652 5396 18680
rect 3660 18640 3666 18652
rect 5368 18624 5396 18652
rect 7300 18652 8800 18680
rect 7300 18624 7328 18652
rect 10226 18640 10232 18692
rect 10284 18640 10290 18692
rect 12912 18680 12940 18788
rect 10428 18652 12940 18680
rect 3418 18612 3424 18624
rect 952 18584 3424 18612
rect 952 18488 980 18584
rect 3418 18572 3424 18584
rect 3476 18572 3482 18624
rect 3510 18572 3516 18624
rect 3568 18572 3574 18624
rect 4798 18572 4804 18624
rect 4856 18572 4862 18624
rect 5350 18572 5356 18624
rect 5408 18572 5414 18624
rect 5534 18572 5540 18624
rect 5592 18612 5598 18624
rect 7193 18615 7251 18621
rect 7193 18612 7205 18615
rect 5592 18584 7205 18612
rect 5592 18572 5598 18584
rect 7193 18581 7205 18584
rect 7239 18581 7251 18615
rect 7193 18575 7251 18581
rect 7282 18572 7288 18624
rect 7340 18572 7346 18624
rect 8294 18572 8300 18624
rect 8352 18612 8358 18624
rect 10428 18621 10456 18652
rect 13354 18640 13360 18692
rect 13412 18680 13418 18692
rect 16776 18680 16804 18788
rect 16868 18748 16896 18856
rect 16942 18844 16948 18896
rect 17000 18884 17006 18896
rect 17678 18884 17684 18896
rect 17000 18856 17684 18884
rect 17000 18844 17006 18856
rect 17678 18844 17684 18856
rect 17736 18844 17742 18896
rect 18064 18828 18092 18924
rect 18417 18921 18429 18955
rect 18463 18952 18475 18955
rect 18463 18924 19656 18952
rect 18463 18921 18475 18924
rect 18417 18915 18475 18921
rect 18141 18887 18199 18893
rect 18141 18853 18153 18887
rect 18187 18884 18199 18887
rect 18785 18887 18843 18893
rect 18187 18856 18736 18884
rect 18187 18853 18199 18856
rect 18141 18847 18199 18853
rect 18046 18776 18052 18828
rect 18104 18776 18110 18828
rect 18506 18816 18512 18828
rect 18340 18788 18512 18816
rect 18138 18748 18144 18760
rect 16868 18720 18144 18748
rect 18138 18708 18144 18720
rect 18196 18708 18202 18760
rect 18340 18757 18368 18788
rect 18506 18776 18512 18788
rect 18564 18776 18570 18828
rect 18708 18816 18736 18856
rect 18785 18853 18797 18887
rect 18831 18884 18843 18887
rect 19337 18887 19395 18893
rect 19337 18884 19349 18887
rect 18831 18856 19349 18884
rect 18831 18853 18843 18856
rect 18785 18847 18843 18853
rect 19337 18853 19349 18856
rect 19383 18853 19395 18887
rect 19628 18884 19656 18924
rect 19794 18912 19800 18964
rect 19852 18952 19858 18964
rect 20257 18955 20315 18961
rect 20257 18952 20269 18955
rect 19852 18924 20269 18952
rect 19852 18912 19858 18924
rect 20257 18921 20269 18924
rect 20303 18921 20315 18955
rect 20257 18915 20315 18921
rect 22738 18912 22744 18964
rect 22796 18952 22802 18964
rect 23382 18952 23388 18964
rect 22796 18924 23388 18952
rect 22796 18912 22802 18924
rect 23382 18912 23388 18924
rect 23440 18912 23446 18964
rect 19628 18856 19748 18884
rect 19337 18847 19395 18853
rect 18969 18819 19027 18825
rect 18708 18788 18828 18816
rect 18325 18751 18383 18757
rect 18325 18717 18337 18751
rect 18371 18717 18383 18751
rect 18325 18711 18383 18717
rect 18414 18708 18420 18760
rect 18472 18748 18478 18760
rect 18601 18751 18659 18757
rect 18601 18748 18613 18751
rect 18472 18720 18613 18748
rect 18472 18708 18478 18720
rect 18601 18717 18613 18720
rect 18647 18717 18659 18751
rect 18601 18711 18659 18717
rect 18693 18751 18751 18757
rect 18693 18717 18705 18751
rect 18739 18717 18751 18751
rect 18800 18748 18828 18788
rect 18969 18785 18981 18819
rect 19015 18816 19027 18819
rect 19613 18819 19671 18825
rect 19613 18816 19625 18819
rect 19015 18788 19625 18816
rect 19015 18785 19027 18788
rect 18969 18779 19027 18785
rect 19613 18785 19625 18788
rect 19659 18785 19671 18819
rect 19613 18779 19671 18785
rect 19245 18751 19303 18757
rect 19245 18748 19257 18751
rect 18800 18720 19257 18748
rect 18693 18711 18751 18717
rect 19245 18717 19257 18720
rect 19291 18717 19303 18751
rect 19245 18711 19303 18717
rect 17678 18680 17684 18692
rect 13412 18652 15332 18680
rect 16776 18652 17684 18680
rect 13412 18640 13418 18652
rect 9125 18615 9183 18621
rect 9125 18612 9137 18615
rect 8352 18584 9137 18612
rect 8352 18572 8358 18584
rect 9125 18581 9137 18584
rect 9171 18581 9183 18615
rect 9125 18575 9183 18581
rect 10413 18615 10471 18621
rect 10413 18581 10425 18615
rect 10459 18581 10471 18615
rect 10413 18575 10471 18581
rect 11974 18572 11980 18624
rect 12032 18612 12038 18624
rect 13814 18612 13820 18624
rect 12032 18584 13820 18612
rect 12032 18572 12038 18584
rect 13814 18572 13820 18584
rect 13872 18572 13878 18624
rect 13906 18572 13912 18624
rect 13964 18612 13970 18624
rect 15194 18612 15200 18624
rect 13964 18584 15200 18612
rect 13964 18572 13970 18584
rect 15194 18572 15200 18584
rect 15252 18572 15258 18624
rect 15304 18612 15332 18652
rect 17678 18640 17684 18652
rect 17736 18640 17742 18692
rect 18708 18680 18736 18711
rect 19518 18708 19524 18760
rect 19576 18708 19582 18760
rect 19720 18757 19748 18856
rect 20162 18844 20168 18896
rect 20220 18884 20226 18896
rect 20220 18856 20760 18884
rect 20220 18844 20226 18856
rect 20441 18819 20499 18825
rect 20441 18785 20453 18819
rect 20487 18816 20499 18819
rect 20625 18819 20683 18825
rect 20625 18816 20637 18819
rect 20487 18788 20637 18816
rect 20487 18785 20499 18788
rect 20441 18779 20499 18785
rect 20625 18785 20637 18788
rect 20671 18785 20683 18819
rect 20625 18779 20683 18785
rect 20732 18757 20760 18856
rect 22465 18819 22523 18825
rect 22465 18816 22477 18819
rect 22296 18788 22477 18816
rect 22296 18760 22324 18788
rect 22465 18785 22477 18788
rect 22511 18785 22523 18819
rect 24121 18819 24179 18825
rect 24121 18816 24133 18819
rect 22465 18779 22523 18785
rect 23124 18788 24133 18816
rect 19705 18751 19763 18757
rect 19705 18717 19717 18751
rect 19751 18717 19763 18751
rect 19705 18711 19763 18717
rect 20165 18751 20223 18757
rect 20165 18717 20177 18751
rect 20211 18717 20223 18751
rect 20165 18711 20223 18717
rect 20533 18751 20591 18757
rect 20533 18717 20545 18751
rect 20579 18717 20591 18751
rect 20533 18711 20591 18717
rect 20717 18751 20775 18757
rect 20717 18717 20729 18751
rect 20763 18717 20775 18751
rect 20717 18711 20775 18717
rect 19536 18680 19564 18708
rect 18708 18652 19564 18680
rect 20180 18680 20208 18711
rect 20548 18680 20576 18711
rect 22278 18708 22284 18760
rect 22336 18708 22342 18760
rect 22370 18708 22376 18760
rect 22428 18708 22434 18760
rect 22738 18757 22744 18760
rect 22707 18751 22744 18757
rect 22707 18717 22719 18751
rect 22707 18711 22744 18717
rect 22738 18708 22744 18711
rect 22796 18708 22802 18760
rect 20990 18680 20996 18692
rect 20180 18652 20996 18680
rect 20990 18640 20996 18652
rect 21048 18640 21054 18692
rect 22554 18640 22560 18692
rect 22612 18680 22618 18692
rect 23124 18680 23152 18788
rect 24121 18785 24133 18788
rect 24167 18785 24179 18819
rect 24121 18779 24179 18785
rect 23845 18751 23903 18757
rect 23845 18748 23857 18751
rect 22612 18652 23152 18680
rect 23492 18720 23857 18748
rect 22612 18640 22618 18652
rect 18322 18612 18328 18624
rect 15304 18584 18328 18612
rect 18322 18572 18328 18584
rect 18380 18572 18386 18624
rect 18969 18615 19027 18621
rect 18969 18581 18981 18615
rect 19015 18612 19027 18615
rect 19242 18612 19248 18624
rect 19015 18584 19248 18612
rect 19015 18581 19027 18584
rect 18969 18575 19027 18581
rect 19242 18572 19248 18584
rect 19300 18572 19306 18624
rect 20438 18572 20444 18624
rect 20496 18572 20502 18624
rect 22186 18572 22192 18624
rect 22244 18572 22250 18624
rect 22646 18572 22652 18624
rect 22704 18612 22710 18624
rect 23492 18621 23520 18720
rect 23845 18717 23857 18720
rect 23891 18717 23903 18751
rect 23845 18711 23903 18717
rect 23934 18708 23940 18760
rect 23992 18708 23998 18760
rect 23477 18615 23535 18621
rect 23477 18612 23489 18615
rect 22704 18584 23489 18612
rect 22704 18572 22710 18584
rect 23477 18581 23489 18584
rect 23523 18581 23535 18615
rect 23477 18575 23535 18581
rect 23842 18572 23848 18624
rect 23900 18612 23906 18624
rect 24121 18615 24179 18621
rect 24121 18612 24133 18615
rect 23900 18584 24133 18612
rect 23900 18572 23906 18584
rect 24121 18581 24133 18584
rect 24167 18581 24179 18615
rect 24121 18575 24179 18581
rect 1104 18522 24723 18544
rect 934 18436 940 18488
rect 992 18436 998 18488
rect 1104 18470 6814 18522
rect 6866 18470 6878 18522
rect 6930 18470 6942 18522
rect 6994 18470 7006 18522
rect 7058 18470 7070 18522
rect 7122 18470 12679 18522
rect 12731 18470 12743 18522
rect 12795 18470 12807 18522
rect 12859 18470 12871 18522
rect 12923 18470 12935 18522
rect 12987 18470 18544 18522
rect 18596 18470 18608 18522
rect 18660 18470 18672 18522
rect 18724 18470 18736 18522
rect 18788 18470 18800 18522
rect 18852 18470 24409 18522
rect 24461 18470 24473 18522
rect 24525 18470 24537 18522
rect 24589 18470 24601 18522
rect 24653 18470 24665 18522
rect 24717 18470 24723 18522
rect 1104 18448 24723 18470
rect 2685 18411 2743 18417
rect 2685 18377 2697 18411
rect 2731 18408 2743 18411
rect 2866 18408 2872 18420
rect 2731 18380 2872 18408
rect 2731 18377 2743 18380
rect 2685 18371 2743 18377
rect 2866 18368 2872 18380
rect 2924 18368 2930 18420
rect 3418 18368 3424 18420
rect 3476 18408 3482 18420
rect 5442 18408 5448 18420
rect 3476 18380 5448 18408
rect 3476 18368 3482 18380
rect 1596 18312 3648 18340
rect 1596 18284 1624 18312
rect 750 18232 756 18284
rect 808 18272 814 18284
rect 1397 18275 1455 18281
rect 1397 18272 1409 18275
rect 808 18244 1409 18272
rect 808 18232 814 18244
rect 1397 18241 1409 18244
rect 1443 18241 1455 18275
rect 1397 18235 1455 18241
rect 1578 18232 1584 18284
rect 1636 18232 1642 18284
rect 1854 18232 1860 18284
rect 1912 18272 1918 18284
rect 3620 18281 3648 18312
rect 3804 18281 3832 18380
rect 5442 18368 5448 18380
rect 5500 18368 5506 18420
rect 6086 18368 6092 18420
rect 6144 18408 6150 18420
rect 6546 18408 6552 18420
rect 6144 18380 6552 18408
rect 6144 18368 6150 18380
rect 6546 18368 6552 18380
rect 6604 18368 6610 18420
rect 7558 18368 7564 18420
rect 7616 18408 7622 18420
rect 9030 18408 9036 18420
rect 7616 18380 9036 18408
rect 7616 18368 7622 18380
rect 9030 18368 9036 18380
rect 9088 18368 9094 18420
rect 9674 18368 9680 18420
rect 9732 18408 9738 18420
rect 10413 18411 10471 18417
rect 10413 18408 10425 18411
rect 9732 18380 10425 18408
rect 9732 18368 9738 18380
rect 10413 18377 10425 18380
rect 10459 18377 10471 18411
rect 10413 18371 10471 18377
rect 10962 18368 10968 18420
rect 11020 18408 11026 18420
rect 16114 18408 16120 18420
rect 11020 18380 16120 18408
rect 11020 18368 11026 18380
rect 16114 18368 16120 18380
rect 16172 18368 16178 18420
rect 17402 18408 17408 18420
rect 16776 18380 17408 18408
rect 5350 18300 5356 18352
rect 5408 18340 5414 18352
rect 11698 18340 11704 18352
rect 5408 18312 7880 18340
rect 5408 18300 5414 18312
rect 1947 18275 2005 18281
rect 1947 18272 1959 18275
rect 1912 18244 1959 18272
rect 1912 18232 1918 18244
rect 1947 18241 1959 18244
rect 1993 18241 2005 18275
rect 1947 18235 2005 18241
rect 3145 18275 3203 18281
rect 3145 18241 3157 18275
rect 3191 18272 3203 18275
rect 3605 18275 3663 18281
rect 3191 18244 3556 18272
rect 3191 18241 3203 18244
rect 3145 18235 3203 18241
rect 1486 18204 1492 18216
rect 1412 18176 1492 18204
rect 1412 18080 1440 18176
rect 1486 18164 1492 18176
rect 1544 18204 1550 18216
rect 1673 18207 1731 18213
rect 1673 18204 1685 18207
rect 1544 18176 1685 18204
rect 1544 18164 1550 18176
rect 1673 18173 1685 18176
rect 1719 18173 1731 18207
rect 1673 18167 1731 18173
rect 3326 18136 3332 18148
rect 2608 18108 3332 18136
rect 1394 18028 1400 18080
rect 1452 18028 1458 18080
rect 1581 18071 1639 18077
rect 1581 18037 1593 18071
rect 1627 18068 1639 18071
rect 2608 18068 2636 18108
rect 3326 18096 3332 18108
rect 3384 18096 3390 18148
rect 3528 18136 3556 18244
rect 3605 18241 3617 18275
rect 3651 18241 3663 18275
rect 3605 18235 3663 18241
rect 3789 18275 3847 18281
rect 3789 18241 3801 18275
rect 3835 18241 3847 18275
rect 3789 18235 3847 18241
rect 4798 18232 4804 18284
rect 4856 18232 4862 18284
rect 5718 18232 5724 18284
rect 5776 18272 5782 18284
rect 6362 18272 6368 18284
rect 5776 18244 6368 18272
rect 5776 18232 5782 18244
rect 6362 18232 6368 18244
rect 6420 18232 6426 18284
rect 6454 18232 6460 18284
rect 6512 18272 6518 18284
rect 7190 18272 7196 18284
rect 6512 18244 7196 18272
rect 6512 18232 6518 18244
rect 7190 18232 7196 18244
rect 7248 18232 7254 18284
rect 4246 18164 4252 18216
rect 4304 18164 4310 18216
rect 4338 18164 4344 18216
rect 4396 18204 4402 18216
rect 4525 18207 4583 18213
rect 4525 18204 4537 18207
rect 4396 18176 4537 18204
rect 4396 18164 4402 18176
rect 4525 18173 4537 18176
rect 4571 18173 4583 18207
rect 4525 18167 4583 18173
rect 4663 18207 4721 18213
rect 4663 18173 4675 18207
rect 4709 18204 4721 18207
rect 4709 18176 5304 18204
rect 4709 18173 4721 18176
rect 4663 18167 4721 18173
rect 5276 18148 5304 18176
rect 3528 18108 4384 18136
rect 1627 18040 2636 18068
rect 1627 18037 1639 18040
rect 1581 18031 1639 18037
rect 3234 18028 3240 18080
rect 3292 18028 3298 18080
rect 3602 18028 3608 18080
rect 3660 18068 3666 18080
rect 4246 18068 4252 18080
rect 3660 18040 4252 18068
rect 3660 18028 3666 18040
rect 4246 18028 4252 18040
rect 4304 18028 4310 18080
rect 4356 18068 4384 18108
rect 5258 18096 5264 18148
rect 5316 18096 5322 18148
rect 7742 18136 7748 18148
rect 5368 18108 7748 18136
rect 5368 18068 5396 18108
rect 7742 18096 7748 18108
rect 7800 18096 7806 18148
rect 4356 18040 5396 18068
rect 5442 18028 5448 18080
rect 5500 18028 5506 18080
rect 5626 18028 5632 18080
rect 5684 18068 5690 18080
rect 5902 18068 5908 18080
rect 5684 18040 5908 18068
rect 5684 18028 5690 18040
rect 5902 18028 5908 18040
rect 5960 18028 5966 18080
rect 7852 18068 7880 18312
rect 9784 18312 11704 18340
rect 7926 18232 7932 18284
rect 7984 18272 7990 18284
rect 9582 18272 9588 18284
rect 7984 18244 9588 18272
rect 7984 18232 7990 18244
rect 9582 18232 9588 18244
rect 9640 18232 9646 18284
rect 9784 18282 9812 18312
rect 11698 18300 11704 18312
rect 11756 18300 11762 18352
rect 11900 18312 12278 18340
rect 9692 18281 9812 18282
rect 9675 18275 9812 18281
rect 9675 18241 9687 18275
rect 9721 18254 9812 18275
rect 9721 18241 9733 18254
rect 9675 18235 9733 18241
rect 10594 18232 10600 18284
rect 10652 18272 10658 18284
rect 11514 18272 11520 18284
rect 10652 18244 11520 18272
rect 10652 18232 10658 18244
rect 11514 18232 11520 18244
rect 11572 18272 11578 18284
rect 11900 18272 11928 18312
rect 12250 18291 12278 18312
rect 13446 18300 13452 18352
rect 13504 18340 13510 18352
rect 13504 18312 13584 18340
rect 13504 18300 13510 18312
rect 12250 18285 12309 18291
rect 11572 18244 11928 18272
rect 11572 18232 11578 18244
rect 11974 18232 11980 18284
rect 12032 18232 12038 18284
rect 12250 18254 12263 18285
rect 12251 18251 12263 18254
rect 12297 18251 12309 18285
rect 13556 18281 13584 18312
rect 16574 18300 16580 18352
rect 16632 18340 16638 18352
rect 16776 18340 16804 18380
rect 17402 18368 17408 18380
rect 17460 18368 17466 18420
rect 17678 18368 17684 18420
rect 17736 18408 17742 18420
rect 17736 18380 18368 18408
rect 17736 18368 17742 18380
rect 16632 18312 16804 18340
rect 18340 18340 18368 18380
rect 18414 18368 18420 18420
rect 18472 18408 18478 18420
rect 18509 18411 18567 18417
rect 18509 18408 18521 18411
rect 18472 18380 18521 18408
rect 18472 18368 18478 18380
rect 18509 18377 18521 18380
rect 18555 18377 18567 18411
rect 18509 18371 18567 18377
rect 22186 18368 22192 18420
rect 22244 18368 22250 18420
rect 22554 18368 22560 18420
rect 22612 18408 22618 18420
rect 22741 18411 22799 18417
rect 22741 18408 22753 18411
rect 22612 18380 22753 18408
rect 22612 18368 22618 18380
rect 22741 18377 22753 18380
rect 22787 18377 22799 18411
rect 22741 18371 22799 18377
rect 23017 18411 23075 18417
rect 23017 18377 23029 18411
rect 23063 18408 23075 18411
rect 23934 18408 23940 18420
rect 23063 18380 23940 18408
rect 23063 18377 23075 18380
rect 23017 18371 23075 18377
rect 23934 18368 23940 18380
rect 23992 18368 23998 18420
rect 24121 18411 24179 18417
rect 24121 18377 24133 18411
rect 24167 18408 24179 18411
rect 25130 18408 25136 18420
rect 24167 18380 25136 18408
rect 24167 18377 24179 18380
rect 24121 18371 24179 18377
rect 25130 18368 25136 18380
rect 25188 18368 25194 18420
rect 20806 18340 20812 18352
rect 18340 18312 20812 18340
rect 16632 18300 16638 18312
rect 12251 18245 12309 18251
rect 13541 18275 13599 18281
rect 13541 18241 13553 18275
rect 13587 18241 13599 18275
rect 13541 18235 13599 18241
rect 14366 18232 14372 18284
rect 14424 18281 14430 18284
rect 14424 18275 14452 18281
rect 14440 18241 14452 18275
rect 14424 18235 14452 18241
rect 14424 18232 14430 18235
rect 14550 18232 14556 18284
rect 14608 18232 14614 18284
rect 16114 18232 16120 18284
rect 16172 18272 16178 18284
rect 16298 18272 16304 18284
rect 16172 18244 16304 18272
rect 16172 18232 16178 18244
rect 16298 18232 16304 18244
rect 16356 18272 16362 18284
rect 16669 18275 16727 18281
rect 16669 18272 16681 18275
rect 16356 18244 16681 18272
rect 16356 18232 16362 18244
rect 16669 18241 16681 18244
rect 16715 18241 16727 18275
rect 16776 18272 16804 18312
rect 20806 18300 20812 18312
rect 20864 18300 20870 18352
rect 22204 18340 22232 18368
rect 22204 18312 22968 18340
rect 16853 18275 16911 18281
rect 16853 18272 16865 18275
rect 16776 18244 16865 18272
rect 16669 18235 16727 18241
rect 16853 18241 16865 18244
rect 16899 18241 16911 18275
rect 16853 18235 16911 18241
rect 17862 18232 17868 18284
rect 17920 18232 17926 18284
rect 20901 18275 20959 18281
rect 20901 18272 20913 18275
rect 20732 18244 20913 18272
rect 20732 18216 20760 18244
rect 20901 18241 20913 18244
rect 20947 18241 20959 18275
rect 20901 18235 20959 18241
rect 22646 18232 22652 18284
rect 22704 18232 22710 18284
rect 22830 18232 22836 18284
rect 22888 18232 22894 18284
rect 22940 18281 22968 18312
rect 22925 18275 22983 18281
rect 22925 18241 22937 18275
rect 22971 18241 22983 18275
rect 22925 18235 22983 18241
rect 23293 18275 23351 18281
rect 23293 18241 23305 18275
rect 23339 18241 23351 18275
rect 23293 18235 23351 18241
rect 9306 18164 9312 18216
rect 9364 18204 9370 18216
rect 9401 18207 9459 18213
rect 9401 18204 9413 18207
rect 9364 18176 9413 18204
rect 9364 18164 9370 18176
rect 9401 18173 9413 18176
rect 9447 18173 9459 18207
rect 9401 18167 9459 18173
rect 11698 18164 11704 18216
rect 11756 18204 11762 18216
rect 11882 18204 11888 18216
rect 11756 18176 11888 18204
rect 11756 18164 11762 18176
rect 11882 18164 11888 18176
rect 11940 18164 11946 18216
rect 13357 18207 13415 18213
rect 13357 18204 13369 18207
rect 12912 18176 13369 18204
rect 10060 18108 12020 18136
rect 10060 18068 10088 18108
rect 7852 18040 10088 18068
rect 11882 18028 11888 18080
rect 11940 18028 11946 18080
rect 11992 18068 12020 18108
rect 12912 18068 12940 18176
rect 13357 18173 13369 18176
rect 13403 18204 13415 18207
rect 13446 18204 13452 18216
rect 13403 18176 13452 18204
rect 13403 18173 13415 18176
rect 13357 18167 13415 18173
rect 13446 18164 13452 18176
rect 13504 18164 13510 18216
rect 14277 18207 14335 18213
rect 14277 18173 14289 18207
rect 14323 18204 14335 18207
rect 14323 18176 16528 18204
rect 14323 18173 14335 18176
rect 14277 18167 14335 18173
rect 12989 18139 13047 18145
rect 12989 18105 13001 18139
rect 13035 18136 13047 18139
rect 14001 18139 14059 18145
rect 14001 18136 14013 18139
rect 13035 18108 14013 18136
rect 13035 18105 13047 18108
rect 12989 18099 13047 18105
rect 14001 18105 14013 18108
rect 14047 18105 14059 18139
rect 16500 18136 16528 18176
rect 17310 18164 17316 18216
rect 17368 18164 17374 18216
rect 17402 18164 17408 18216
rect 17460 18204 17466 18216
rect 17589 18207 17647 18213
rect 17589 18204 17601 18207
rect 17460 18176 17601 18204
rect 17460 18164 17466 18176
rect 17589 18173 17601 18176
rect 17635 18173 17647 18207
rect 17589 18167 17647 18173
rect 17678 18164 17684 18216
rect 17736 18213 17742 18216
rect 17736 18207 17764 18213
rect 17752 18173 17764 18207
rect 17736 18167 17764 18173
rect 17736 18164 17742 18167
rect 20714 18164 20720 18216
rect 20772 18164 20778 18216
rect 17218 18136 17224 18148
rect 16500 18108 17224 18136
rect 14001 18099 14059 18105
rect 17218 18096 17224 18108
rect 17276 18136 17282 18148
rect 17420 18136 17448 18164
rect 17276 18108 17448 18136
rect 17276 18096 17282 18108
rect 21818 18096 21824 18148
rect 21876 18136 21882 18148
rect 23308 18136 23336 18235
rect 23382 18232 23388 18284
rect 23440 18272 23446 18284
rect 23845 18275 23903 18281
rect 23845 18272 23857 18275
rect 23440 18244 23857 18272
rect 23440 18232 23446 18244
rect 23845 18241 23857 18244
rect 23891 18241 23903 18275
rect 23845 18235 23903 18241
rect 21876 18108 23336 18136
rect 21876 18096 21882 18108
rect 11992 18040 12940 18068
rect 15194 18028 15200 18080
rect 15252 18028 15258 18080
rect 18046 18028 18052 18080
rect 18104 18068 18110 18080
rect 20162 18068 20168 18080
rect 18104 18040 20168 18068
rect 18104 18028 18110 18040
rect 20162 18028 20168 18040
rect 20220 18028 20226 18080
rect 20717 18071 20775 18077
rect 20717 18037 20729 18071
rect 20763 18068 20775 18071
rect 22094 18068 22100 18080
rect 20763 18040 22100 18068
rect 20763 18037 20775 18040
rect 20717 18031 20775 18037
rect 22094 18028 22100 18040
rect 22152 18028 22158 18080
rect 23566 18028 23572 18080
rect 23624 18028 23630 18080
rect 24854 18028 24860 18080
rect 24912 18028 24918 18080
rect 750 17960 756 18012
rect 808 18000 814 18012
rect 934 18000 940 18012
rect 808 17972 940 18000
rect 808 17960 814 17972
rect 934 17960 940 17972
rect 992 17960 998 18012
rect 1104 17978 24564 18000
rect 1104 17926 3882 17978
rect 3934 17926 3946 17978
rect 3998 17926 4010 17978
rect 4062 17926 4074 17978
rect 4126 17926 4138 17978
rect 4190 17926 9747 17978
rect 9799 17926 9811 17978
rect 9863 17926 9875 17978
rect 9927 17926 9939 17978
rect 9991 17926 10003 17978
rect 10055 17926 15612 17978
rect 15664 17926 15676 17978
rect 15728 17926 15740 17978
rect 15792 17926 15804 17978
rect 15856 17926 15868 17978
rect 15920 17926 21477 17978
rect 21529 17926 21541 17978
rect 21593 17926 21605 17978
rect 21657 17926 21669 17978
rect 21721 17926 21733 17978
rect 21785 17926 24564 17978
rect 1104 17904 24564 17926
rect 2130 17824 2136 17876
rect 2188 17864 2194 17876
rect 5442 17864 5448 17876
rect 2188 17836 5448 17864
rect 2188 17824 2194 17836
rect 5442 17824 5448 17836
rect 5500 17824 5506 17876
rect 6270 17824 6276 17876
rect 6328 17824 6334 17876
rect 7190 17824 7196 17876
rect 7248 17864 7254 17876
rect 7248 17836 10548 17864
rect 7248 17824 7254 17836
rect 2961 17799 3019 17805
rect 2961 17765 2973 17799
rect 3007 17796 3019 17799
rect 6288 17796 6316 17824
rect 3007 17768 6316 17796
rect 3007 17765 3019 17768
rect 2961 17759 3019 17765
rect 8202 17756 8208 17808
rect 8260 17796 8266 17808
rect 9674 17796 9680 17808
rect 8260 17768 9680 17796
rect 8260 17756 8266 17768
rect 9674 17756 9680 17768
rect 9732 17756 9738 17808
rect 9858 17756 9864 17808
rect 9916 17756 9922 17808
rect 2700 17700 4752 17728
rect 1394 17620 1400 17672
rect 1452 17620 1458 17672
rect 1671 17663 1729 17669
rect 1671 17629 1683 17663
rect 1717 17660 1729 17663
rect 2700 17660 2728 17700
rect 4724 17672 4752 17700
rect 5460 17700 7144 17728
rect 1717 17632 2728 17660
rect 1717 17629 1729 17632
rect 1671 17623 1729 17629
rect 2774 17620 2780 17672
rect 2832 17620 2838 17672
rect 3237 17663 3295 17669
rect 3237 17629 3249 17663
rect 3283 17660 3295 17663
rect 3694 17660 3700 17672
rect 3283 17632 3700 17660
rect 3283 17629 3295 17632
rect 3237 17623 3295 17629
rect 3694 17620 3700 17632
rect 3752 17620 3758 17672
rect 4246 17620 4252 17672
rect 4304 17660 4310 17672
rect 4617 17663 4675 17669
rect 4617 17660 4629 17663
rect 4304 17632 4629 17660
rect 4304 17620 4310 17632
rect 4617 17629 4629 17632
rect 4663 17629 4675 17663
rect 4617 17623 4675 17629
rect 4706 17620 4712 17672
rect 4764 17620 4770 17672
rect 4801 17663 4859 17669
rect 4801 17629 4813 17663
rect 4847 17660 4859 17663
rect 5460 17660 5488 17700
rect 4847 17632 5488 17660
rect 4847 17629 4859 17632
rect 4801 17623 4859 17629
rect 5534 17620 5540 17672
rect 5592 17620 5598 17672
rect 1302 17552 1308 17604
rect 1360 17592 1366 17604
rect 4065 17595 4123 17601
rect 1360 17564 3096 17592
rect 1360 17552 1366 17564
rect 1854 17484 1860 17536
rect 1912 17524 1918 17536
rect 2409 17527 2467 17533
rect 2409 17524 2421 17527
rect 1912 17496 2421 17524
rect 1912 17484 1918 17496
rect 2409 17493 2421 17496
rect 2455 17493 2467 17527
rect 3068 17524 3096 17564
rect 4065 17561 4077 17595
rect 4111 17592 4123 17595
rect 5552 17592 5580 17620
rect 4111 17564 5580 17592
rect 4111 17561 4123 17564
rect 4065 17555 4123 17561
rect 3329 17527 3387 17533
rect 3329 17524 3341 17527
rect 3068 17496 3341 17524
rect 2409 17487 2467 17493
rect 3329 17493 3341 17496
rect 3375 17493 3387 17527
rect 3329 17487 3387 17493
rect 3418 17484 3424 17536
rect 3476 17524 3482 17536
rect 4157 17527 4215 17533
rect 4157 17524 4169 17527
rect 3476 17496 4169 17524
rect 3476 17484 3482 17496
rect 4157 17493 4169 17496
rect 4203 17493 4215 17527
rect 4157 17487 4215 17493
rect 4338 17484 4344 17536
rect 4396 17524 4402 17536
rect 6086 17524 6092 17536
rect 4396 17496 6092 17524
rect 4396 17484 4402 17496
rect 6086 17484 6092 17496
rect 6144 17484 6150 17536
rect 7116 17524 7144 17700
rect 9122 17688 9128 17740
rect 9180 17728 9186 17740
rect 9876 17728 9904 17756
rect 9180 17700 9904 17728
rect 10520 17728 10548 17836
rect 11882 17824 11888 17876
rect 11940 17824 11946 17876
rect 14550 17824 14556 17876
rect 14608 17864 14614 17876
rect 15105 17867 15163 17873
rect 15105 17864 15117 17867
rect 14608 17836 15117 17864
rect 14608 17824 14614 17836
rect 15105 17833 15117 17836
rect 15151 17833 15163 17867
rect 17681 17867 17739 17873
rect 15105 17827 15163 17833
rect 16776 17836 17632 17864
rect 10873 17799 10931 17805
rect 10873 17765 10885 17799
rect 10919 17796 10931 17799
rect 11900 17796 11928 17824
rect 16776 17796 16804 17836
rect 10919 17768 11468 17796
rect 11900 17768 12020 17796
rect 10919 17765 10931 17768
rect 10873 17759 10931 17765
rect 11440 17728 11468 17768
rect 11885 17731 11943 17737
rect 11885 17728 11897 17731
rect 10520 17700 11284 17728
rect 11440 17700 11897 17728
rect 9180 17688 9186 17700
rect 7190 17620 7196 17672
rect 7248 17620 7254 17672
rect 7374 17620 7380 17672
rect 7432 17660 7438 17672
rect 7467 17663 7525 17669
rect 7467 17660 7479 17663
rect 7432 17632 7479 17660
rect 7432 17620 7438 17632
rect 7467 17629 7479 17632
rect 7513 17629 7525 17663
rect 7467 17623 7525 17629
rect 7484 17592 7512 17623
rect 8018 17620 8024 17672
rect 8076 17660 8082 17672
rect 8938 17660 8944 17672
rect 8076 17632 8944 17660
rect 8076 17620 8082 17632
rect 8938 17620 8944 17632
rect 8996 17620 9002 17672
rect 9306 17620 9312 17672
rect 9364 17660 9370 17672
rect 10134 17669 10140 17672
rect 9861 17663 9919 17669
rect 9861 17660 9873 17663
rect 9364 17632 9873 17660
rect 9364 17620 9370 17632
rect 9861 17629 9873 17632
rect 9907 17660 9919 17663
rect 10103 17663 10140 17669
rect 9907 17632 9996 17660
rect 9907 17629 9919 17632
rect 9861 17623 9919 17629
rect 9968 17592 9996 17632
rect 10103 17629 10115 17663
rect 10103 17623 10140 17629
rect 10134 17620 10140 17623
rect 10192 17620 10198 17672
rect 10594 17620 10600 17672
rect 10652 17620 10658 17672
rect 11146 17620 11152 17672
rect 11204 17620 11210 17672
rect 11256 17669 11284 17700
rect 11885 17697 11897 17700
rect 11931 17697 11943 17731
rect 11992 17728 12020 17768
rect 14844 17768 16804 17796
rect 12161 17731 12219 17737
rect 12161 17728 12173 17731
rect 11992 17700 12173 17728
rect 11885 17691 11943 17697
rect 12161 17697 12173 17700
rect 12207 17697 12219 17731
rect 12161 17691 12219 17697
rect 11241 17663 11299 17669
rect 11241 17629 11253 17663
rect 11287 17629 11299 17663
rect 11241 17623 11299 17629
rect 11425 17663 11483 17669
rect 11425 17629 11437 17663
rect 11471 17629 11483 17663
rect 11425 17623 11483 17629
rect 10612 17592 10640 17620
rect 7484 17564 9812 17592
rect 9968 17564 10640 17592
rect 11164 17592 11192 17620
rect 11440 17592 11468 17623
rect 12250 17620 12256 17672
rect 12308 17669 12314 17672
rect 12308 17663 12336 17669
rect 12324 17629 12336 17663
rect 12308 17623 12336 17629
rect 12308 17620 12314 17623
rect 12434 17620 12440 17672
rect 12492 17620 12498 17672
rect 13814 17620 13820 17672
rect 13872 17660 13878 17672
rect 14093 17663 14151 17669
rect 14093 17660 14105 17663
rect 13872 17632 14105 17660
rect 13872 17620 13878 17632
rect 14093 17629 14105 17632
rect 14139 17629 14151 17663
rect 14093 17623 14151 17629
rect 14367 17663 14425 17669
rect 14367 17629 14379 17663
rect 14413 17660 14425 17663
rect 14734 17660 14740 17672
rect 14413 17632 14740 17660
rect 14413 17629 14425 17632
rect 14367 17623 14425 17629
rect 14734 17620 14740 17632
rect 14792 17620 14798 17672
rect 11164 17564 11468 17592
rect 13081 17595 13139 17601
rect 7650 17524 7656 17536
rect 7116 17496 7656 17524
rect 7650 17484 7656 17496
rect 7708 17484 7714 17536
rect 8110 17484 8116 17536
rect 8168 17524 8174 17536
rect 8205 17527 8263 17533
rect 8205 17524 8217 17527
rect 8168 17496 8217 17524
rect 8168 17484 8174 17496
rect 8205 17493 8217 17496
rect 8251 17493 8263 17527
rect 9784 17524 9812 17564
rect 13081 17561 13093 17595
rect 13127 17592 13139 17595
rect 14844 17592 14872 17768
rect 16482 17688 16488 17740
rect 16540 17728 16546 17740
rect 16669 17731 16727 17737
rect 16669 17728 16681 17731
rect 16540 17700 16681 17728
rect 16540 17688 16546 17700
rect 16669 17697 16681 17700
rect 16715 17697 16727 17731
rect 16669 17691 16727 17697
rect 15562 17620 15568 17672
rect 15620 17660 15626 17672
rect 15749 17663 15807 17669
rect 15749 17660 15761 17663
rect 15620 17632 15761 17660
rect 15620 17620 15626 17632
rect 15749 17629 15761 17632
rect 15795 17629 15807 17663
rect 16942 17660 16948 17672
rect 15749 17623 15807 17629
rect 15856 17632 16948 17660
rect 13127 17564 14872 17592
rect 13127 17561 13139 17564
rect 13081 17555 13139 17561
rect 11146 17524 11152 17536
rect 9784 17496 11152 17524
rect 8205 17487 8263 17493
rect 11146 17484 11152 17496
rect 11204 17484 11210 17536
rect 11882 17484 11888 17536
rect 11940 17524 11946 17536
rect 15856 17524 15884 17632
rect 16942 17620 16948 17632
rect 17000 17620 17006 17672
rect 17604 17592 17632 17836
rect 17681 17833 17693 17867
rect 17727 17864 17739 17867
rect 17862 17864 17868 17876
rect 17727 17836 17868 17864
rect 17727 17833 17739 17836
rect 17681 17827 17739 17833
rect 17862 17824 17868 17836
rect 17920 17824 17926 17876
rect 22370 17864 22376 17876
rect 22020 17836 22376 17864
rect 22020 17796 22048 17836
rect 22370 17824 22376 17836
rect 22428 17824 22434 17876
rect 24121 17867 24179 17873
rect 24121 17833 24133 17867
rect 24167 17864 24179 17867
rect 24872 17864 24900 18028
rect 24167 17836 24900 17864
rect 24167 17833 24179 17836
rect 24121 17827 24179 17833
rect 21468 17768 22048 17796
rect 23753 17799 23811 17805
rect 21468 17740 21496 17768
rect 23753 17765 23765 17799
rect 23799 17796 23811 17799
rect 24854 17796 24860 17808
rect 23799 17768 24860 17796
rect 23799 17765 23811 17768
rect 23753 17759 23811 17765
rect 24854 17756 24860 17768
rect 24912 17756 24918 17808
rect 21450 17688 21456 17740
rect 21508 17688 21514 17740
rect 17954 17620 17960 17672
rect 18012 17660 18018 17672
rect 19150 17660 19156 17672
rect 18012 17632 19156 17660
rect 18012 17620 18018 17632
rect 19150 17620 19156 17632
rect 19208 17660 19214 17672
rect 19521 17663 19579 17669
rect 19521 17660 19533 17663
rect 19208 17632 19533 17660
rect 19208 17620 19214 17632
rect 19521 17629 19533 17632
rect 19567 17629 19579 17663
rect 19521 17623 19579 17629
rect 20441 17663 20499 17669
rect 20441 17629 20453 17663
rect 20487 17660 20499 17663
rect 22002 17660 22008 17672
rect 20487 17632 22008 17660
rect 20487 17629 20499 17632
rect 20441 17623 20499 17629
rect 22002 17620 22008 17632
rect 22060 17620 22066 17672
rect 23569 17663 23627 17669
rect 23569 17629 23581 17663
rect 23615 17660 23627 17663
rect 23842 17660 23848 17672
rect 23615 17632 23848 17660
rect 23615 17629 23627 17632
rect 23569 17623 23627 17629
rect 23842 17620 23848 17632
rect 23900 17620 23906 17672
rect 23937 17663 23995 17669
rect 23937 17629 23949 17663
rect 23983 17660 23995 17663
rect 24210 17660 24216 17672
rect 23983 17632 24216 17660
rect 23983 17629 23995 17632
rect 23937 17623 23995 17629
rect 24210 17620 24216 17632
rect 24268 17620 24274 17672
rect 20714 17601 20720 17604
rect 20686 17595 20720 17601
rect 20686 17592 20698 17595
rect 17604 17564 20698 17592
rect 20686 17561 20698 17564
rect 20686 17555 20720 17561
rect 20714 17552 20720 17555
rect 20772 17552 20778 17604
rect 20806 17552 20812 17604
rect 20864 17592 20870 17604
rect 22272 17595 22330 17601
rect 22272 17592 22284 17595
rect 20864 17564 22284 17592
rect 20864 17552 20870 17564
rect 22272 17561 22284 17564
rect 22318 17592 22330 17595
rect 22318 17564 22784 17592
rect 22318 17561 22330 17564
rect 22272 17555 22330 17561
rect 22756 17536 22784 17564
rect 11940 17496 15884 17524
rect 11940 17484 11946 17496
rect 19334 17484 19340 17536
rect 19392 17484 19398 17536
rect 20070 17484 20076 17536
rect 20128 17524 20134 17536
rect 21450 17524 21456 17536
rect 20128 17496 21456 17524
rect 20128 17484 20134 17496
rect 21450 17484 21456 17496
rect 21508 17484 21514 17536
rect 21818 17484 21824 17536
rect 21876 17484 21882 17536
rect 22738 17484 22744 17536
rect 22796 17484 22802 17536
rect 23382 17484 23388 17536
rect 23440 17484 23446 17536
rect 1104 17434 24723 17456
rect 1104 17382 6814 17434
rect 6866 17382 6878 17434
rect 6930 17382 6942 17434
rect 6994 17382 7006 17434
rect 7058 17382 7070 17434
rect 7122 17382 12679 17434
rect 12731 17382 12743 17434
rect 12795 17382 12807 17434
rect 12859 17382 12871 17434
rect 12923 17382 12935 17434
rect 12987 17382 18544 17434
rect 18596 17382 18608 17434
rect 18660 17382 18672 17434
rect 18724 17382 18736 17434
rect 18788 17382 18800 17434
rect 18852 17382 24409 17434
rect 24461 17382 24473 17434
rect 24525 17382 24537 17434
rect 24589 17382 24601 17434
rect 24653 17382 24665 17434
rect 24717 17382 24723 17434
rect 1104 17360 24723 17382
rect 2590 17280 2596 17332
rect 2648 17320 2654 17332
rect 4338 17320 4344 17332
rect 2648 17292 4344 17320
rect 2648 17280 2654 17292
rect 4338 17280 4344 17292
rect 4396 17280 4402 17332
rect 4614 17280 4620 17332
rect 4672 17320 4678 17332
rect 4672 17292 5120 17320
rect 4672 17280 4678 17292
rect 3050 17252 3056 17264
rect 1964 17224 3056 17252
rect 1486 17144 1492 17196
rect 1544 17144 1550 17196
rect 1964 17193 1992 17224
rect 3050 17212 3056 17224
rect 3108 17252 3114 17264
rect 5092 17252 5120 17292
rect 5166 17280 5172 17332
rect 5224 17320 5230 17332
rect 7282 17320 7288 17332
rect 5224 17292 7288 17320
rect 5224 17280 5230 17292
rect 7282 17280 7288 17292
rect 7340 17320 7346 17332
rect 7929 17323 7987 17329
rect 7929 17320 7941 17323
rect 7340 17292 7941 17320
rect 7340 17280 7346 17292
rect 7929 17289 7941 17292
rect 7975 17289 7987 17323
rect 8294 17320 8300 17332
rect 7929 17283 7987 17289
rect 8018 17292 8300 17320
rect 3108 17224 4752 17252
rect 5092 17224 5178 17252
rect 3108 17212 3114 17224
rect 1949 17187 2007 17193
rect 1949 17153 1961 17187
rect 1995 17153 2007 17187
rect 2222 17184 2228 17196
rect 2183 17156 2228 17184
rect 1949 17147 2007 17153
rect 2222 17144 2228 17156
rect 2280 17144 2286 17196
rect 3160 17116 3188 17224
rect 3234 17144 3240 17196
rect 3292 17184 3298 17196
rect 3603 17187 3661 17193
rect 3603 17184 3615 17187
rect 3292 17156 3615 17184
rect 3292 17144 3298 17156
rect 3603 17153 3615 17156
rect 3649 17184 3661 17187
rect 4062 17184 4068 17196
rect 3649 17156 4068 17184
rect 3649 17153 3661 17156
rect 3603 17147 3661 17153
rect 4062 17144 4068 17156
rect 4120 17144 4126 17196
rect 4724 17128 4752 17224
rect 5150 17223 5178 17224
rect 6638 17223 6644 17264
rect 5150 17217 5209 17223
rect 5150 17186 5163 17217
rect 5151 17183 5163 17186
rect 5197 17183 5209 17217
rect 6623 17217 6644 17223
rect 5151 17177 5209 17183
rect 5902 17144 5908 17196
rect 5960 17184 5966 17196
rect 6362 17184 6368 17196
rect 5960 17156 6368 17184
rect 5960 17144 5966 17156
rect 6362 17144 6368 17156
rect 6420 17144 6426 17196
rect 6623 17183 6635 17217
rect 6696 17212 6702 17264
rect 7098 17212 7104 17264
rect 7156 17252 7162 17264
rect 8018 17252 8046 17292
rect 8294 17280 8300 17292
rect 8352 17280 8358 17332
rect 8846 17280 8852 17332
rect 8904 17320 8910 17332
rect 10410 17320 10416 17332
rect 8904 17292 10416 17320
rect 8904 17280 8910 17292
rect 10410 17280 10416 17292
rect 10468 17280 10474 17332
rect 12250 17320 12256 17332
rect 11072 17292 12256 17320
rect 9033 17255 9091 17261
rect 7156 17224 8046 17252
rect 8312 17224 8892 17252
rect 7156 17212 7162 17224
rect 6669 17186 6684 17212
rect 6669 17183 6681 17186
rect 6623 17177 6681 17183
rect 8018 17144 8024 17196
rect 8076 17184 8082 17196
rect 8312 17193 8340 17224
rect 8864 17196 8892 17224
rect 9033 17221 9045 17255
rect 9079 17221 9091 17255
rect 9033 17215 9091 17221
rect 8205 17187 8263 17193
rect 8205 17184 8217 17187
rect 8076 17156 8217 17184
rect 8076 17144 8082 17156
rect 8205 17153 8217 17156
rect 8251 17153 8263 17187
rect 8205 17147 8263 17153
rect 8297 17187 8355 17193
rect 8297 17153 8309 17187
rect 8343 17153 8355 17187
rect 8297 17147 8355 17153
rect 8570 17144 8576 17196
rect 8628 17184 8634 17196
rect 8665 17187 8723 17193
rect 8665 17184 8677 17187
rect 8628 17156 8677 17184
rect 8628 17144 8634 17156
rect 8665 17153 8677 17156
rect 8711 17153 8723 17187
rect 8665 17147 8723 17153
rect 8846 17144 8852 17196
rect 8904 17144 8910 17196
rect 3329 17119 3387 17125
rect 3329 17116 3341 17119
rect 3160 17088 3341 17116
rect 3329 17085 3341 17088
rect 3375 17085 3387 17119
rect 3329 17079 3387 17085
rect 4706 17076 4712 17128
rect 4764 17116 4770 17128
rect 4893 17119 4951 17125
rect 4893 17116 4905 17119
rect 4764 17088 4905 17116
rect 4764 17076 4770 17088
rect 4893 17085 4905 17088
rect 4939 17085 4951 17119
rect 4893 17079 4951 17085
rect 8110 17076 8116 17128
rect 8168 17076 8174 17128
rect 6178 17048 6184 17060
rect 5828 17020 6184 17048
rect 842 16940 848 16992
rect 900 16980 906 16992
rect 1581 16983 1639 16989
rect 1581 16980 1593 16983
rect 900 16952 1593 16980
rect 900 16940 906 16952
rect 1581 16949 1593 16952
rect 1627 16949 1639 16983
rect 1581 16943 1639 16949
rect 2961 16983 3019 16989
rect 2961 16949 2973 16983
rect 3007 16980 3019 16983
rect 3602 16980 3608 16992
rect 3007 16952 3608 16980
rect 3007 16949 3019 16952
rect 2961 16943 3019 16949
rect 3602 16940 3608 16952
rect 3660 16940 3666 16992
rect 4341 16983 4399 16989
rect 4341 16949 4353 16983
rect 4387 16980 4399 16983
rect 4430 16980 4436 16992
rect 4387 16952 4436 16980
rect 4387 16949 4399 16952
rect 4341 16943 4399 16949
rect 4430 16940 4436 16952
rect 4488 16940 4494 16992
rect 5350 16940 5356 16992
rect 5408 16980 5414 16992
rect 5828 16980 5856 17020
rect 6178 17008 6184 17020
rect 6236 17008 6242 17060
rect 7190 17008 7196 17060
rect 7248 17048 7254 17060
rect 9048 17048 9076 17215
rect 9122 17212 9128 17264
rect 9180 17252 9186 17264
rect 11072 17252 11100 17292
rect 12250 17280 12256 17292
rect 12308 17280 12314 17332
rect 12434 17280 12440 17332
rect 12492 17320 12498 17332
rect 12529 17323 12587 17329
rect 12529 17320 12541 17323
rect 12492 17292 12541 17320
rect 12492 17280 12498 17292
rect 12529 17289 12541 17292
rect 12575 17289 12587 17323
rect 15286 17320 15292 17332
rect 12529 17283 12587 17289
rect 14844 17292 15292 17320
rect 9180 17224 11100 17252
rect 9180 17212 9186 17224
rect 11146 17212 11152 17264
rect 11204 17252 11210 17264
rect 14844 17252 14872 17292
rect 15286 17280 15292 17292
rect 15344 17280 15350 17332
rect 16298 17280 16304 17332
rect 16356 17320 16362 17332
rect 16574 17320 16580 17332
rect 16356 17292 16580 17320
rect 16356 17280 16362 17292
rect 16574 17280 16580 17292
rect 16632 17280 16638 17332
rect 17310 17280 17316 17332
rect 17368 17320 17374 17332
rect 17681 17323 17739 17329
rect 17681 17320 17693 17323
rect 17368 17292 17693 17320
rect 17368 17280 17374 17292
rect 17681 17289 17693 17292
rect 17727 17289 17739 17323
rect 17681 17283 17739 17289
rect 21818 17280 21824 17332
rect 21876 17280 21882 17332
rect 22557 17323 22615 17329
rect 22557 17289 22569 17323
rect 22603 17289 22615 17323
rect 22557 17283 22615 17289
rect 19150 17261 19156 17264
rect 19144 17252 19156 17261
rect 11204 17224 14872 17252
rect 19111 17224 19156 17252
rect 11204 17212 11210 17224
rect 19144 17215 19156 17224
rect 19150 17212 19156 17215
rect 19208 17212 19214 17264
rect 9306 17144 9312 17196
rect 9364 17184 9370 17196
rect 9735 17187 9793 17193
rect 9735 17184 9747 17187
rect 9364 17156 9747 17184
rect 9364 17144 9370 17156
rect 9735 17153 9747 17156
rect 9781 17153 9793 17187
rect 9735 17147 9793 17153
rect 9858 17144 9864 17196
rect 9916 17184 9922 17196
rect 11759 17187 11817 17193
rect 11759 17184 11771 17187
rect 9916 17156 11771 17184
rect 9916 17144 9922 17156
rect 11759 17153 11771 17156
rect 11805 17153 11817 17187
rect 11759 17147 11817 17153
rect 13446 17144 13452 17196
rect 13504 17184 13510 17196
rect 14829 17187 14887 17193
rect 14829 17184 14841 17187
rect 13504 17156 14841 17184
rect 13504 17144 13510 17156
rect 14829 17153 14841 17156
rect 14875 17153 14887 17187
rect 14829 17147 14887 17153
rect 15010 17144 15016 17196
rect 15068 17144 15074 17196
rect 15562 17144 15568 17196
rect 15620 17144 15626 17196
rect 16482 17144 16488 17196
rect 16540 17144 16546 17196
rect 16574 17144 16580 17196
rect 16632 17184 16638 17196
rect 16911 17187 16969 17193
rect 16911 17184 16923 17187
rect 16632 17156 16923 17184
rect 16632 17144 16638 17156
rect 16911 17153 16923 17156
rect 16957 17153 16969 17187
rect 16911 17147 16969 17153
rect 19610 17144 19616 17196
rect 19668 17184 19674 17196
rect 20591 17187 20649 17193
rect 20591 17184 20603 17187
rect 19668 17156 20603 17184
rect 19668 17144 19674 17156
rect 20591 17153 20603 17156
rect 20637 17153 20649 17187
rect 20591 17147 20649 17153
rect 20714 17144 20720 17196
rect 20772 17184 20778 17196
rect 21836 17184 21864 17280
rect 22005 17187 22063 17193
rect 22005 17184 22017 17187
rect 20772 17156 21036 17184
rect 21836 17156 22017 17184
rect 20772 17144 20778 17156
rect 9493 17119 9551 17125
rect 9493 17085 9505 17119
rect 9539 17085 9551 17119
rect 9493 17079 9551 17085
rect 9508 17048 9536 17079
rect 10594 17076 10600 17128
rect 10652 17116 10658 17128
rect 11517 17119 11575 17125
rect 11517 17116 11529 17119
rect 10652 17088 11529 17116
rect 10652 17076 10658 17088
rect 11517 17085 11529 17088
rect 11563 17085 11575 17119
rect 11517 17079 11575 17085
rect 7248 17020 7972 17048
rect 9048 17020 9444 17048
rect 9508 17020 9628 17048
rect 7248 17008 7254 17020
rect 7944 16992 7972 17020
rect 5408 16952 5856 16980
rect 5408 16940 5414 16952
rect 5902 16940 5908 16992
rect 5960 16940 5966 16992
rect 6086 16940 6092 16992
rect 6144 16980 6150 16992
rect 7098 16980 7104 16992
rect 6144 16952 7104 16980
rect 6144 16940 6150 16952
rect 7098 16940 7104 16952
rect 7156 16940 7162 16992
rect 7374 16940 7380 16992
rect 7432 16940 7438 16992
rect 7926 16940 7932 16992
rect 7984 16940 7990 16992
rect 9214 16940 9220 16992
rect 9272 16940 9278 16992
rect 9416 16980 9444 17020
rect 9600 16992 9628 17020
rect 9490 16980 9496 16992
rect 9416 16952 9496 16980
rect 9490 16940 9496 16952
rect 9548 16940 9554 16992
rect 9582 16940 9588 16992
rect 9640 16940 9646 16992
rect 10226 16940 10232 16992
rect 10284 16980 10290 16992
rect 10505 16983 10563 16989
rect 10505 16980 10517 16983
rect 10284 16952 10517 16980
rect 10284 16940 10290 16952
rect 10505 16949 10517 16952
rect 10551 16949 10563 16983
rect 11520 16980 11548 17079
rect 14366 17076 14372 17128
rect 14424 17116 14430 17128
rect 14645 17119 14703 17125
rect 14645 17116 14657 17119
rect 14424 17088 14657 17116
rect 14424 17076 14430 17088
rect 14645 17085 14657 17088
rect 14691 17085 14703 17119
rect 14645 17079 14703 17085
rect 14734 17076 14740 17128
rect 14792 17116 14798 17128
rect 15028 17116 15056 17144
rect 15682 17119 15740 17125
rect 15682 17116 15694 17119
rect 14792 17088 15694 17116
rect 14792 17076 14798 17088
rect 15682 17085 15694 17088
rect 15728 17085 15740 17119
rect 15682 17079 15740 17085
rect 15841 17119 15899 17125
rect 15841 17085 15853 17119
rect 15887 17116 15899 17119
rect 16022 17116 16028 17128
rect 15887 17088 16028 17116
rect 15887 17085 15899 17088
rect 15841 17079 15899 17085
rect 16022 17076 16028 17088
rect 16080 17076 16086 17128
rect 16500 17116 16528 17144
rect 16669 17119 16727 17125
rect 16669 17116 16681 17119
rect 16500 17088 16681 17116
rect 16669 17085 16681 17088
rect 16715 17085 16727 17119
rect 16669 17079 16727 17085
rect 17954 17076 17960 17128
rect 18012 17116 18018 17128
rect 18874 17116 18880 17128
rect 18012 17088 18880 17116
rect 18012 17076 18018 17088
rect 18874 17076 18880 17088
rect 18932 17076 18938 17128
rect 20346 17076 20352 17128
rect 20404 17076 20410 17128
rect 21008 17116 21036 17156
rect 22005 17153 22017 17156
rect 22051 17153 22063 17187
rect 22005 17147 22063 17153
rect 22281 17187 22339 17193
rect 22281 17153 22293 17187
rect 22327 17184 22339 17187
rect 22572 17184 22600 17283
rect 23382 17280 23388 17332
rect 23440 17280 23446 17332
rect 23400 17252 23428 17280
rect 24029 17255 24087 17261
rect 24029 17252 24041 17255
rect 23032 17224 23428 17252
rect 23584 17224 24041 17252
rect 22327 17156 22600 17184
rect 22327 17153 22339 17156
rect 22281 17147 22339 17153
rect 22738 17144 22744 17196
rect 22796 17144 22802 17196
rect 23032 17193 23060 17224
rect 23017 17187 23075 17193
rect 23017 17153 23029 17187
rect 23063 17153 23075 17187
rect 23017 17147 23075 17153
rect 23293 17187 23351 17193
rect 23293 17153 23305 17187
rect 23339 17184 23351 17187
rect 23584 17184 23612 17224
rect 24029 17221 24041 17224
rect 24075 17221 24087 17255
rect 24029 17215 24087 17221
rect 23339 17156 23612 17184
rect 23339 17153 23351 17156
rect 23293 17147 23351 17153
rect 23750 17144 23756 17196
rect 23808 17144 23814 17196
rect 23842 17144 23848 17196
rect 23900 17144 23906 17196
rect 23860 17116 23888 17144
rect 21008 17088 23888 17116
rect 24029 17119 24087 17125
rect 24029 17085 24041 17119
rect 24075 17116 24087 17119
rect 24075 17088 24164 17116
rect 24075 17085 24087 17088
rect 24029 17079 24087 17085
rect 15286 17008 15292 17060
rect 15344 17008 15350 17060
rect 23845 17051 23903 17057
rect 23845 17048 23857 17051
rect 22756 17020 23857 17048
rect 12250 16980 12256 16992
rect 11520 16952 12256 16980
rect 10505 16943 10563 16949
rect 12250 16940 12256 16952
rect 12308 16940 12314 16992
rect 16482 16940 16488 16992
rect 16540 16940 16546 16992
rect 20257 16983 20315 16989
rect 20257 16949 20269 16983
rect 20303 16980 20315 16983
rect 20714 16980 20720 16992
rect 20303 16952 20720 16980
rect 20303 16949 20315 16952
rect 20257 16943 20315 16949
rect 20714 16940 20720 16952
rect 20772 16940 20778 16992
rect 21082 16940 21088 16992
rect 21140 16980 21146 16992
rect 21361 16983 21419 16989
rect 21361 16980 21373 16983
rect 21140 16952 21373 16980
rect 21140 16940 21146 16952
rect 21361 16949 21373 16952
rect 21407 16949 21419 16983
rect 21361 16943 21419 16949
rect 21821 16983 21879 16989
rect 21821 16949 21833 16983
rect 21867 16980 21879 16983
rect 22278 16980 22284 16992
rect 21867 16952 22284 16980
rect 21867 16949 21879 16952
rect 21821 16943 21879 16949
rect 22278 16940 22284 16952
rect 22336 16940 22342 16992
rect 22373 16983 22431 16989
rect 22373 16949 22385 16983
rect 22419 16980 22431 16983
rect 22756 16980 22784 17020
rect 23845 17017 23857 17020
rect 23891 17017 23903 17051
rect 23845 17011 23903 17017
rect 24136 16992 24164 17088
rect 22419 16952 22784 16980
rect 22833 16983 22891 16989
rect 22419 16949 22431 16952
rect 22373 16943 22431 16949
rect 22833 16949 22845 16983
rect 22879 16980 22891 16983
rect 23474 16980 23480 16992
rect 22879 16952 23480 16980
rect 22879 16949 22891 16952
rect 22833 16943 22891 16949
rect 23474 16940 23480 16952
rect 23532 16940 23538 16992
rect 23566 16940 23572 16992
rect 23624 16940 23630 16992
rect 24118 16940 24124 16992
rect 24176 16940 24182 16992
rect 1104 16890 24564 16912
rect 1104 16838 3882 16890
rect 3934 16838 3946 16890
rect 3998 16838 4010 16890
rect 4062 16838 4074 16890
rect 4126 16838 4138 16890
rect 4190 16838 9747 16890
rect 9799 16838 9811 16890
rect 9863 16838 9875 16890
rect 9927 16838 9939 16890
rect 9991 16838 10003 16890
rect 10055 16838 15612 16890
rect 15664 16838 15676 16890
rect 15728 16838 15740 16890
rect 15792 16838 15804 16890
rect 15856 16838 15868 16890
rect 15920 16838 21477 16890
rect 21529 16838 21541 16890
rect 21593 16838 21605 16890
rect 21657 16838 21669 16890
rect 21721 16838 21733 16890
rect 21785 16838 24564 16890
rect 1104 16816 24564 16838
rect 5534 16776 5540 16788
rect 2332 16748 4752 16776
rect 1762 16708 1768 16720
rect 1596 16680 1768 16708
rect 1596 16649 1624 16680
rect 1762 16668 1768 16680
rect 1820 16668 1826 16720
rect 1854 16668 1860 16720
rect 1912 16708 1918 16720
rect 2225 16711 2283 16717
rect 2225 16708 2237 16711
rect 1912 16680 2237 16708
rect 1912 16668 1918 16680
rect 2225 16677 2237 16680
rect 2271 16677 2283 16711
rect 2225 16671 2283 16677
rect 2332 16652 2360 16748
rect 4614 16708 4620 16720
rect 3344 16680 4620 16708
rect 1581 16643 1639 16649
rect 1581 16609 1593 16643
rect 1627 16609 1639 16643
rect 1581 16603 1639 16609
rect 2314 16600 2320 16652
rect 2372 16640 2378 16652
rect 2501 16643 2559 16649
rect 2501 16640 2513 16643
rect 2372 16612 2513 16640
rect 2372 16600 2378 16612
rect 2501 16609 2513 16612
rect 2547 16609 2559 16643
rect 2501 16603 2559 16609
rect 2590 16600 2596 16652
rect 2648 16649 2654 16652
rect 2648 16643 2676 16649
rect 2664 16609 2676 16643
rect 2648 16603 2676 16609
rect 2648 16600 2654 16603
rect 2958 16600 2964 16652
rect 3016 16640 3022 16652
rect 3344 16640 3372 16680
rect 4614 16668 4620 16680
rect 4672 16668 4678 16720
rect 3016 16612 3372 16640
rect 3016 16600 3022 16612
rect 3418 16600 3424 16652
rect 3476 16600 3482 16652
rect 4724 16640 4752 16748
rect 4908 16748 5540 16776
rect 4908 16717 4936 16748
rect 5534 16736 5540 16748
rect 5592 16736 5598 16788
rect 5902 16736 5908 16788
rect 5960 16736 5966 16788
rect 7374 16776 7380 16788
rect 6840 16748 7380 16776
rect 4893 16711 4951 16717
rect 4893 16677 4905 16711
rect 4939 16677 4951 16711
rect 4893 16671 4951 16677
rect 5166 16640 5172 16652
rect 4724 16612 5172 16640
rect 5166 16600 5172 16612
rect 5224 16600 5230 16652
rect 5350 16649 5356 16652
rect 5307 16643 5356 16649
rect 5307 16609 5319 16643
rect 5353 16609 5356 16643
rect 5307 16603 5356 16609
rect 5350 16600 5356 16603
rect 5408 16600 5414 16652
rect 5445 16643 5503 16649
rect 5445 16609 5457 16643
rect 5491 16640 5503 16643
rect 5920 16640 5948 16736
rect 6840 16717 6868 16748
rect 7374 16736 7380 16748
rect 7432 16736 7438 16788
rect 7926 16736 7932 16788
rect 7984 16776 7990 16788
rect 9582 16776 9588 16788
rect 7984 16748 9588 16776
rect 7984 16736 7990 16748
rect 9582 16736 9588 16748
rect 9640 16776 9646 16788
rect 12250 16776 12256 16788
rect 9640 16748 11652 16776
rect 9640 16736 9646 16748
rect 6825 16711 6883 16717
rect 6104 16680 6408 16708
rect 6104 16652 6132 16680
rect 5491 16612 5948 16640
rect 5491 16609 5503 16612
rect 5445 16603 5503 16609
rect 6086 16600 6092 16652
rect 6144 16600 6150 16652
rect 6178 16600 6184 16652
rect 6236 16600 6242 16652
rect 6380 16649 6408 16680
rect 6825 16677 6837 16711
rect 6871 16677 6883 16711
rect 6825 16671 6883 16677
rect 6365 16643 6423 16649
rect 6365 16609 6377 16643
rect 6411 16609 6423 16643
rect 6730 16640 6736 16652
rect 6365 16603 6423 16609
rect 6472 16612 6736 16640
rect 1765 16575 1823 16581
rect 1765 16541 1777 16575
rect 1811 16572 1823 16575
rect 1946 16572 1952 16584
rect 1811 16544 1952 16572
rect 1811 16541 1823 16544
rect 1765 16535 1823 16541
rect 1946 16532 1952 16544
rect 2004 16532 2010 16584
rect 2774 16532 2780 16584
rect 2832 16532 2838 16584
rect 3786 16532 3792 16584
rect 3844 16532 3850 16584
rect 3878 16532 3884 16584
rect 3936 16572 3942 16584
rect 4249 16575 4307 16581
rect 4249 16572 4261 16575
rect 3936 16544 4261 16572
rect 3936 16532 3942 16544
rect 4249 16541 4261 16544
rect 4295 16541 4307 16575
rect 4249 16535 4307 16541
rect 4338 16532 4344 16584
rect 4396 16572 4402 16584
rect 4433 16575 4491 16581
rect 4433 16572 4445 16575
rect 4396 16544 4445 16572
rect 4396 16532 4402 16544
rect 4433 16541 4445 16544
rect 4479 16541 4491 16575
rect 4433 16535 4491 16541
rect 6270 16532 6276 16584
rect 6328 16572 6334 16584
rect 6472 16572 6500 16612
rect 6730 16600 6736 16612
rect 6788 16640 6794 16652
rect 7218 16643 7276 16649
rect 7218 16640 7230 16643
rect 6788 16612 7230 16640
rect 6788 16600 6794 16612
rect 7218 16609 7230 16612
rect 7264 16609 7276 16643
rect 7218 16603 7276 16609
rect 8018 16600 8024 16652
rect 8076 16640 8082 16652
rect 9674 16640 9680 16652
rect 8076 16612 9680 16640
rect 8076 16600 8082 16612
rect 9646 16600 9680 16612
rect 9732 16600 9738 16652
rect 10152 16649 10180 16748
rect 10870 16668 10876 16720
rect 10928 16708 10934 16720
rect 11149 16711 11207 16717
rect 11149 16708 11161 16711
rect 10928 16680 11161 16708
rect 10928 16668 10934 16680
rect 11149 16677 11161 16680
rect 11195 16677 11207 16711
rect 11149 16671 11207 16677
rect 11624 16652 11652 16748
rect 11900 16748 12256 16776
rect 10137 16643 10195 16649
rect 10137 16609 10149 16643
rect 10183 16609 10195 16643
rect 10137 16603 10195 16609
rect 11606 16600 11612 16652
rect 11664 16600 11670 16652
rect 11900 16649 11928 16748
rect 12250 16736 12256 16748
rect 12308 16736 12314 16788
rect 15286 16736 15292 16788
rect 15344 16776 15350 16788
rect 15381 16779 15439 16785
rect 15381 16776 15393 16779
rect 15344 16748 15393 16776
rect 15344 16736 15350 16748
rect 15381 16745 15393 16748
rect 15427 16745 15439 16779
rect 18693 16779 18751 16785
rect 15381 16739 15439 16745
rect 16960 16748 18000 16776
rect 16960 16649 16988 16748
rect 17972 16652 18000 16748
rect 18693 16745 18705 16779
rect 18739 16776 18751 16779
rect 21450 16776 21456 16788
rect 18739 16748 21456 16776
rect 18739 16745 18751 16748
rect 18693 16739 18751 16745
rect 21450 16736 21456 16748
rect 21508 16736 21514 16788
rect 21821 16779 21879 16785
rect 21821 16745 21833 16779
rect 21867 16776 21879 16779
rect 22189 16779 22247 16785
rect 22189 16776 22201 16779
rect 21867 16748 22201 16776
rect 21867 16745 21879 16748
rect 21821 16739 21879 16745
rect 22189 16745 22201 16748
rect 22235 16745 22247 16779
rect 22189 16739 22247 16745
rect 22278 16736 22284 16788
rect 22336 16776 22342 16788
rect 22336 16748 22582 16776
rect 22336 16736 22342 16748
rect 18601 16711 18659 16717
rect 18601 16677 18613 16711
rect 18647 16708 18659 16711
rect 18969 16711 19027 16717
rect 18969 16708 18981 16711
rect 18647 16680 18981 16708
rect 18647 16677 18659 16680
rect 18601 16671 18659 16677
rect 18969 16677 18981 16680
rect 19015 16677 19027 16711
rect 19613 16711 19671 16717
rect 19613 16708 19625 16711
rect 18969 16671 19027 16677
rect 19168 16680 19625 16708
rect 11885 16643 11943 16649
rect 11885 16609 11897 16643
rect 11931 16609 11943 16643
rect 16945 16643 17003 16649
rect 11885 16603 11943 16609
rect 12544 16612 14136 16640
rect 6328 16544 6500 16572
rect 6328 16532 6334 16544
rect 7098 16532 7104 16584
rect 7156 16532 7162 16584
rect 7372 16532 7378 16584
rect 7430 16532 7436 16584
rect 9646 16572 9674 16600
rect 10042 16572 10048 16584
rect 9646 16544 10048 16572
rect 10042 16532 10048 16544
rect 10100 16572 10106 16584
rect 10379 16575 10437 16581
rect 10379 16572 10391 16575
rect 10100 16544 10391 16572
rect 10100 16532 10106 16544
rect 10379 16541 10391 16544
rect 10425 16541 10437 16575
rect 10379 16535 10437 16541
rect 12159 16575 12217 16581
rect 12159 16541 12171 16575
rect 12205 16572 12217 16575
rect 12544 16572 12572 16612
rect 14108 16584 14136 16612
rect 16945 16609 16957 16643
rect 16991 16609 17003 16643
rect 16945 16603 17003 16609
rect 17954 16600 17960 16652
rect 18012 16600 18018 16652
rect 18785 16643 18843 16649
rect 18785 16609 18797 16643
rect 18831 16640 18843 16643
rect 19168 16640 19196 16680
rect 19613 16677 19625 16680
rect 19659 16677 19671 16711
rect 20990 16708 20996 16720
rect 19613 16671 19671 16677
rect 20548 16680 20996 16708
rect 18831 16612 19196 16640
rect 18831 16609 18843 16612
rect 18785 16603 18843 16609
rect 19334 16600 19340 16652
rect 19392 16640 19398 16652
rect 20073 16643 20131 16649
rect 19392 16612 20024 16640
rect 19392 16600 19398 16612
rect 12205 16544 12572 16572
rect 12205 16541 12217 16544
rect 12159 16535 12217 16541
rect 9122 16504 9128 16516
rect 3896 16476 4476 16504
rect 842 16396 848 16448
rect 900 16436 906 16448
rect 1210 16436 1216 16448
rect 900 16408 1216 16436
rect 900 16396 906 16408
rect 1210 16396 1216 16408
rect 1268 16396 1274 16448
rect 1670 16396 1676 16448
rect 1728 16436 1734 16448
rect 3896 16436 3924 16476
rect 1728 16408 3924 16436
rect 3973 16439 4031 16445
rect 1728 16396 1734 16408
rect 3973 16405 3985 16439
rect 4019 16436 4031 16439
rect 4246 16436 4252 16448
rect 4019 16408 4252 16436
rect 4019 16405 4031 16408
rect 3973 16399 4031 16405
rect 4246 16396 4252 16408
rect 4304 16396 4310 16448
rect 4448 16436 4476 16476
rect 7944 16476 9128 16504
rect 5902 16436 5908 16448
rect 4448 16408 5908 16436
rect 5902 16396 5908 16408
rect 5960 16396 5966 16448
rect 6089 16439 6147 16445
rect 6089 16405 6101 16439
rect 6135 16436 6147 16439
rect 6178 16436 6184 16448
rect 6135 16408 6184 16436
rect 6135 16405 6147 16408
rect 6089 16399 6147 16405
rect 6178 16396 6184 16408
rect 6236 16396 6242 16448
rect 6546 16396 6552 16448
rect 6604 16436 6610 16448
rect 7944 16436 7972 16476
rect 9122 16464 9128 16476
rect 9180 16464 9186 16516
rect 9398 16464 9404 16516
rect 9456 16504 9462 16516
rect 9456 16476 11560 16504
rect 9456 16464 9462 16476
rect 6604 16408 7972 16436
rect 6604 16396 6610 16408
rect 8018 16396 8024 16448
rect 8076 16396 8082 16448
rect 9490 16396 9496 16448
rect 9548 16436 9554 16448
rect 11422 16436 11428 16448
rect 9548 16408 11428 16436
rect 9548 16396 9554 16408
rect 11422 16396 11428 16408
rect 11480 16396 11486 16448
rect 11532 16436 11560 16476
rect 11974 16464 11980 16516
rect 12032 16504 12038 16516
rect 12174 16504 12202 16535
rect 13354 16532 13360 16584
rect 13412 16572 13418 16584
rect 13633 16575 13691 16581
rect 13633 16572 13645 16575
rect 13412 16544 13645 16572
rect 13412 16532 13418 16544
rect 13633 16541 13645 16544
rect 13679 16541 13691 16575
rect 13633 16535 13691 16541
rect 14090 16532 14096 16584
rect 14148 16532 14154 16584
rect 14369 16575 14427 16581
rect 14369 16541 14381 16575
rect 14415 16541 14427 16575
rect 14643 16575 14701 16581
rect 14643 16572 14655 16575
rect 14369 16535 14427 16541
rect 14642 16541 14655 16572
rect 14689 16541 14701 16575
rect 14642 16535 14701 16541
rect 12032 16476 12202 16504
rect 12032 16464 12038 16476
rect 14384 16448 14412 16535
rect 14550 16464 14556 16516
rect 14608 16504 14614 16516
rect 14642 16504 14670 16535
rect 16482 16532 16488 16584
rect 16540 16572 16546 16584
rect 17201 16575 17259 16581
rect 17201 16572 17213 16575
rect 16540 16544 17213 16572
rect 16540 16532 16546 16544
rect 17201 16541 17213 16544
rect 17247 16541 17259 16575
rect 17201 16535 17259 16541
rect 18414 16532 18420 16584
rect 18472 16572 18478 16584
rect 18509 16575 18567 16581
rect 18509 16572 18521 16575
rect 18472 16544 18521 16572
rect 18472 16532 18478 16544
rect 18509 16541 18521 16544
rect 18555 16541 18567 16575
rect 18509 16535 18567 16541
rect 18874 16532 18880 16584
rect 18932 16532 18938 16584
rect 19429 16575 19487 16581
rect 19429 16572 19441 16575
rect 18984 16544 19441 16572
rect 18984 16504 19012 16544
rect 19429 16541 19441 16544
rect 19475 16541 19487 16575
rect 19429 16535 19487 16541
rect 19518 16532 19524 16584
rect 19576 16532 19582 16584
rect 19996 16581 20024 16612
rect 20073 16609 20085 16643
rect 20119 16640 20131 16643
rect 20441 16643 20499 16649
rect 20441 16640 20453 16643
rect 20119 16612 20453 16640
rect 20119 16609 20131 16612
rect 20073 16603 20131 16609
rect 20441 16609 20453 16612
rect 20487 16609 20499 16643
rect 20441 16603 20499 16609
rect 19705 16575 19763 16581
rect 19705 16541 19717 16575
rect 19751 16541 19763 16575
rect 19705 16535 19763 16541
rect 19981 16575 20039 16581
rect 19981 16541 19993 16575
rect 20027 16541 20039 16575
rect 19981 16535 20039 16541
rect 20349 16575 20407 16581
rect 20349 16541 20361 16575
rect 20395 16572 20407 16575
rect 20548 16572 20576 16680
rect 20990 16668 20996 16680
rect 21048 16668 21054 16720
rect 20625 16643 20683 16649
rect 20625 16609 20637 16643
rect 20671 16640 20683 16643
rect 21085 16643 21143 16649
rect 21085 16640 21097 16643
rect 20671 16612 21097 16640
rect 20671 16609 20683 16612
rect 20625 16603 20683 16609
rect 21085 16609 21097 16612
rect 21131 16609 21143 16643
rect 21085 16603 21143 16609
rect 22005 16643 22063 16649
rect 22005 16609 22017 16643
rect 22051 16640 22063 16643
rect 22465 16643 22523 16649
rect 22465 16640 22477 16643
rect 22051 16612 22477 16640
rect 22051 16609 22063 16612
rect 22005 16603 22063 16609
rect 22465 16609 22477 16612
rect 22511 16609 22523 16643
rect 22465 16603 22523 16609
rect 20395 16544 20576 16572
rect 20395 16541 20407 16544
rect 20349 16535 20407 16541
rect 19720 16504 19748 16535
rect 20714 16532 20720 16584
rect 20772 16572 20778 16584
rect 20901 16575 20959 16581
rect 20901 16572 20913 16575
rect 20772 16544 20913 16572
rect 20772 16532 20778 16544
rect 20901 16541 20913 16544
rect 20947 16541 20959 16575
rect 20901 16535 20959 16541
rect 20990 16532 20996 16584
rect 21048 16532 21054 16584
rect 21177 16575 21235 16581
rect 21177 16541 21189 16575
rect 21223 16541 21235 16575
rect 21177 16535 21235 16541
rect 21729 16575 21787 16581
rect 21729 16541 21741 16575
rect 21775 16541 21787 16575
rect 21729 16535 21787 16541
rect 14608 16476 14670 16504
rect 18340 16476 19012 16504
rect 19260 16476 19748 16504
rect 14608 16464 14614 16476
rect 12434 16436 12440 16448
rect 11532 16408 12440 16436
rect 12434 16396 12440 16408
rect 12492 16396 12498 16448
rect 12897 16439 12955 16445
rect 12897 16405 12909 16439
rect 12943 16436 12955 16439
rect 13078 16436 13084 16448
rect 12943 16408 13084 16436
rect 12943 16405 12955 16408
rect 12897 16399 12955 16405
rect 13078 16396 13084 16408
rect 13136 16396 13142 16448
rect 14366 16396 14372 16448
rect 14424 16436 14430 16448
rect 15102 16436 15108 16448
rect 14424 16408 15108 16436
rect 14424 16396 14430 16408
rect 15102 16396 15108 16408
rect 15160 16396 15166 16448
rect 18340 16445 18368 16476
rect 19260 16445 19288 16476
rect 20622 16464 20628 16516
rect 20680 16464 20686 16516
rect 21192 16504 21220 16535
rect 20732 16476 21220 16504
rect 21744 16504 21772 16535
rect 22094 16532 22100 16584
rect 22152 16532 22158 16584
rect 22554 16581 22582 16748
rect 23474 16736 23480 16788
rect 23532 16736 23538 16788
rect 23661 16779 23719 16785
rect 23661 16745 23673 16779
rect 23707 16776 23719 16779
rect 23750 16776 23756 16788
rect 23707 16748 23756 16776
rect 23707 16745 23719 16748
rect 23661 16739 23719 16745
rect 23750 16736 23756 16748
rect 23808 16736 23814 16788
rect 24118 16736 24124 16788
rect 24176 16736 24182 16788
rect 23492 16640 23520 16736
rect 23492 16612 23704 16640
rect 22373 16575 22431 16581
rect 22373 16541 22385 16575
rect 22419 16541 22431 16575
rect 22554 16575 22615 16581
rect 22554 16544 22569 16575
rect 22373 16535 22431 16541
rect 22557 16541 22569 16544
rect 22603 16541 22615 16575
rect 22557 16535 22615 16541
rect 22649 16575 22707 16581
rect 22649 16541 22661 16575
rect 22695 16541 22707 16575
rect 22649 16535 22707 16541
rect 22907 16545 22965 16551
rect 22394 16504 22422 16535
rect 22462 16504 22468 16516
rect 21744 16476 22468 16504
rect 20732 16445 20760 16476
rect 22462 16464 22468 16476
rect 22520 16464 22526 16516
rect 18325 16439 18383 16445
rect 18325 16405 18337 16439
rect 18371 16405 18383 16439
rect 18325 16399 18383 16405
rect 19245 16439 19303 16445
rect 19245 16405 19257 16439
rect 19291 16405 19303 16439
rect 19245 16399 19303 16405
rect 20717 16439 20775 16445
rect 20717 16405 20729 16439
rect 20763 16405 20775 16439
rect 20717 16399 20775 16405
rect 22005 16439 22063 16445
rect 22005 16405 22017 16439
rect 22051 16436 22063 16439
rect 22094 16436 22100 16448
rect 22051 16408 22100 16436
rect 22051 16405 22063 16408
rect 22005 16399 22063 16405
rect 22094 16396 22100 16408
rect 22152 16396 22158 16448
rect 22186 16396 22192 16448
rect 22244 16436 22250 16448
rect 22664 16436 22692 16535
rect 22907 16511 22919 16545
rect 22953 16511 22965 16545
rect 22907 16505 22965 16511
rect 22244 16408 22692 16436
rect 22244 16396 22250 16408
rect 22830 16396 22836 16448
rect 22888 16436 22894 16448
rect 22922 16436 22950 16505
rect 23676 16504 23704 16612
rect 23768 16572 23796 16736
rect 24029 16575 24087 16581
rect 24029 16572 24041 16575
rect 23768 16544 24041 16572
rect 24029 16541 24041 16544
rect 24075 16541 24087 16575
rect 24029 16535 24087 16541
rect 24213 16575 24271 16581
rect 24213 16541 24225 16575
rect 24259 16541 24271 16575
rect 24213 16535 24271 16541
rect 24228 16504 24256 16535
rect 23676 16476 24256 16504
rect 22888 16408 22950 16436
rect 22888 16396 22894 16408
rect 1104 16346 24723 16368
rect 1104 16294 6814 16346
rect 6866 16294 6878 16346
rect 6930 16294 6942 16346
rect 6994 16294 7006 16346
rect 7058 16294 7070 16346
rect 7122 16294 12679 16346
rect 12731 16294 12743 16346
rect 12795 16294 12807 16346
rect 12859 16294 12871 16346
rect 12923 16294 12935 16346
rect 12987 16294 18544 16346
rect 18596 16294 18608 16346
rect 18660 16294 18672 16346
rect 18724 16294 18736 16346
rect 18788 16294 18800 16346
rect 18852 16294 24409 16346
rect 24461 16294 24473 16346
rect 24525 16294 24537 16346
rect 24589 16294 24601 16346
rect 24653 16294 24665 16346
rect 24717 16294 24723 16346
rect 1104 16272 24723 16294
rect 2038 16192 2044 16244
rect 2096 16232 2102 16244
rect 2222 16232 2228 16244
rect 2096 16204 2228 16232
rect 2096 16192 2102 16204
rect 2222 16192 2228 16204
rect 2280 16192 2286 16244
rect 2685 16235 2743 16241
rect 2685 16201 2697 16235
rect 2731 16232 2743 16235
rect 2774 16232 2780 16244
rect 2731 16204 2780 16232
rect 2731 16201 2743 16204
rect 2685 16195 2743 16201
rect 2774 16192 2780 16204
rect 2832 16192 2838 16244
rect 4338 16232 4344 16244
rect 3436 16204 4344 16232
rect 2958 16164 2964 16176
rect 1962 16136 2964 16164
rect 1962 16135 1990 16136
rect 1931 16129 1990 16135
rect 1931 16095 1943 16129
rect 1977 16098 1990 16129
rect 2958 16124 2964 16136
rect 3016 16124 3022 16176
rect 1977 16095 1989 16098
rect 1931 16089 1989 16095
rect 2314 16056 2320 16108
rect 2372 16096 2378 16108
rect 3436 16105 3464 16204
rect 4338 16192 4344 16204
rect 4396 16192 4402 16244
rect 5902 16192 5908 16244
rect 5960 16192 5966 16244
rect 7374 16192 7380 16244
rect 7432 16232 7438 16244
rect 7653 16235 7711 16241
rect 7653 16232 7665 16235
rect 7432 16204 7665 16232
rect 7432 16192 7438 16204
rect 7653 16201 7665 16204
rect 7699 16201 7711 16235
rect 7653 16195 7711 16201
rect 8846 16192 8852 16244
rect 8904 16232 8910 16244
rect 9033 16235 9091 16241
rect 9033 16232 9045 16235
rect 8904 16204 9045 16232
rect 8904 16192 8910 16204
rect 9033 16201 9045 16204
rect 9079 16201 9091 16235
rect 12069 16235 12127 16241
rect 12069 16232 12081 16235
rect 9033 16195 9091 16201
rect 9140 16204 12081 16232
rect 5920 16164 5948 16192
rect 9140 16164 9168 16204
rect 12069 16201 12081 16204
rect 12115 16232 12127 16235
rect 12115 16204 12434 16232
rect 12115 16201 12127 16204
rect 12069 16195 12127 16201
rect 5920 16136 9168 16164
rect 3421 16099 3479 16105
rect 3421 16096 3433 16099
rect 2372 16068 3433 16096
rect 2372 16056 2378 16068
rect 3421 16065 3433 16068
rect 3467 16065 3479 16099
rect 3421 16059 3479 16065
rect 4154 16056 4160 16108
rect 4212 16056 4218 16108
rect 4430 16056 4436 16108
rect 4488 16056 4494 16108
rect 5258 16056 5264 16108
rect 5316 16096 5322 16108
rect 6086 16096 6092 16108
rect 5316 16068 6092 16096
rect 5316 16056 5322 16068
rect 6086 16056 6092 16068
rect 6144 16056 6150 16108
rect 6362 16056 6368 16108
rect 6420 16096 6426 16108
rect 6641 16099 6699 16105
rect 6641 16096 6653 16099
rect 6420 16068 6653 16096
rect 6420 16056 6426 16068
rect 6641 16065 6653 16068
rect 6687 16065 6699 16099
rect 6641 16059 6699 16065
rect 6822 16056 6828 16108
rect 6880 16096 6886 16108
rect 6915 16099 6973 16105
rect 6915 16096 6927 16099
rect 6880 16068 6927 16096
rect 6880 16056 6886 16068
rect 6915 16065 6927 16068
rect 6961 16065 6973 16099
rect 6915 16059 6973 16065
rect 7926 16056 7932 16108
rect 7984 16096 7990 16108
rect 8021 16099 8079 16105
rect 8021 16096 8033 16099
rect 7984 16068 8033 16096
rect 7984 16056 7990 16068
rect 8021 16065 8033 16068
rect 8067 16065 8079 16099
rect 8294 16096 8300 16108
rect 8255 16068 8300 16096
rect 8021 16059 8079 16065
rect 8294 16056 8300 16068
rect 8352 16056 8358 16108
rect 9490 16056 9496 16108
rect 9548 16056 9554 16108
rect 12406 16096 12434 16204
rect 12986 16192 12992 16244
rect 13044 16232 13050 16244
rect 13170 16232 13176 16244
rect 13044 16204 13176 16232
rect 13044 16192 13050 16204
rect 13170 16192 13176 16204
rect 13228 16192 13234 16244
rect 13446 16192 13452 16244
rect 13504 16232 13510 16244
rect 13630 16232 13636 16244
rect 13504 16204 13636 16232
rect 13504 16192 13510 16204
rect 13630 16192 13636 16204
rect 13688 16192 13694 16244
rect 14090 16192 14096 16244
rect 14148 16232 14154 16244
rect 14148 16204 15725 16232
rect 14148 16192 14154 16204
rect 15194 16164 15200 16176
rect 14198 16136 15200 16164
rect 12621 16099 12679 16105
rect 12621 16096 12633 16099
rect 12406 16068 12633 16096
rect 12621 16065 12633 16068
rect 12667 16065 12679 16099
rect 12621 16059 12679 16065
rect 13354 16056 13360 16108
rect 13412 16056 13418 16108
rect 13630 16056 13636 16108
rect 13688 16056 13694 16108
rect 1394 15988 1400 16040
rect 1452 16028 1458 16040
rect 1673 16031 1731 16037
rect 1673 16028 1685 16031
rect 1452 16000 1685 16028
rect 1452 15988 1458 16000
rect 1673 15997 1685 16000
rect 1719 15997 1731 16031
rect 1673 15991 1731 15997
rect 3237 16031 3295 16037
rect 3237 15997 3249 16031
rect 3283 15997 3295 16031
rect 3237 15991 3295 15997
rect 3252 15960 3280 15991
rect 3602 15988 3608 16040
rect 3660 16028 3666 16040
rect 3881 16031 3939 16037
rect 3881 16028 3893 16031
rect 3660 16000 3893 16028
rect 3660 15988 3666 16000
rect 3881 15997 3893 16000
rect 3927 15997 3939 16031
rect 3881 15991 3939 15997
rect 4295 16031 4353 16037
rect 4295 15997 4307 16031
rect 4341 16028 4353 16031
rect 6270 16028 6276 16040
rect 4341 16000 6276 16028
rect 4341 15997 4353 16000
rect 4295 15991 4353 15997
rect 6270 15988 6276 16000
rect 6328 15988 6334 16040
rect 7650 15988 7656 16040
rect 7708 15988 7714 16040
rect 9582 16028 9588 16040
rect 8680 16000 9588 16028
rect 3252 15932 3832 15960
rect 1762 15852 1768 15904
rect 1820 15892 1826 15904
rect 2774 15892 2780 15904
rect 1820 15864 2780 15892
rect 1820 15852 1826 15864
rect 2774 15852 2780 15864
rect 2832 15892 2838 15904
rect 3252 15892 3280 15932
rect 3804 15904 3832 15932
rect 2832 15864 3280 15892
rect 2832 15852 2838 15864
rect 3786 15852 3792 15904
rect 3844 15852 3850 15904
rect 4246 15852 4252 15904
rect 4304 15892 4310 15904
rect 5077 15895 5135 15901
rect 5077 15892 5089 15895
rect 4304 15864 5089 15892
rect 4304 15852 4310 15864
rect 5077 15861 5089 15864
rect 5123 15861 5135 15895
rect 7668 15892 7696 15988
rect 8680 15892 8708 16000
rect 9582 15988 9588 16000
rect 9640 16028 9646 16040
rect 9677 16031 9735 16037
rect 9677 16028 9689 16031
rect 9640 16000 9689 16028
rect 9640 15988 9646 16000
rect 9677 15997 9689 16000
rect 9723 15997 9735 16031
rect 9677 15991 9735 15997
rect 10042 15988 10048 16040
rect 10100 15988 10106 16040
rect 10134 15988 10140 16040
rect 10192 15988 10198 16040
rect 10413 16031 10471 16037
rect 10413 16028 10425 16031
rect 10244 16000 10425 16028
rect 10060 15960 10088 15988
rect 10244 15960 10272 16000
rect 10413 15997 10425 16000
rect 10459 15997 10471 16031
rect 10413 15991 10471 15997
rect 10548 15988 10554 16040
rect 10606 15988 10612 16040
rect 10689 16031 10747 16037
rect 10689 15997 10701 16031
rect 10735 16028 10747 16031
rect 10870 16028 10876 16040
rect 10735 16000 10876 16028
rect 10735 15997 10747 16000
rect 10689 15991 10747 15997
rect 10870 15988 10876 16000
rect 10928 15988 10934 16040
rect 12434 15988 12440 16040
rect 12492 15988 12498 16040
rect 13078 15988 13084 16040
rect 13136 15988 13142 16040
rect 13495 16031 13553 16037
rect 13495 16028 13507 16031
rect 13188 16000 13507 16028
rect 10060 15932 10272 15960
rect 12342 15920 12348 15972
rect 12400 15960 12406 15972
rect 13188 15960 13216 16000
rect 13495 15997 13507 16000
rect 13541 16028 13553 16031
rect 14198 16028 14226 16136
rect 15194 16124 15200 16136
rect 15252 16124 15258 16176
rect 15286 16056 15292 16108
rect 15344 16096 15350 16108
rect 15379 16099 15437 16105
rect 15379 16096 15391 16099
rect 15344 16068 15391 16096
rect 15344 16056 15350 16068
rect 15379 16065 15391 16068
rect 15425 16065 15437 16099
rect 15379 16059 15437 16065
rect 13541 16000 14226 16028
rect 13541 15997 13553 16000
rect 13495 15991 13553 15997
rect 15102 15988 15108 16040
rect 15160 15988 15166 16040
rect 15697 16028 15725 16204
rect 16022 16192 16028 16244
rect 16080 16232 16086 16244
rect 16117 16235 16175 16241
rect 16117 16232 16129 16235
rect 16080 16204 16129 16232
rect 16080 16192 16086 16204
rect 16117 16201 16129 16204
rect 16163 16201 16175 16235
rect 16117 16195 16175 16201
rect 16482 16192 16488 16244
rect 16540 16192 16546 16244
rect 17405 16235 17463 16241
rect 17405 16201 17417 16235
rect 17451 16201 17463 16235
rect 17405 16195 17463 16201
rect 16500 16096 16528 16192
rect 17420 16164 17448 16195
rect 18414 16192 18420 16244
rect 18472 16232 18478 16244
rect 18785 16235 18843 16241
rect 18785 16232 18797 16235
rect 18472 16204 18797 16232
rect 18472 16192 18478 16204
rect 18785 16201 18797 16204
rect 18831 16232 18843 16235
rect 19518 16232 19524 16244
rect 18831 16204 19524 16232
rect 18831 16201 18843 16204
rect 18785 16195 18843 16201
rect 19518 16192 19524 16204
rect 19576 16192 19582 16244
rect 22094 16192 22100 16244
rect 22152 16232 22158 16244
rect 22152 16204 22416 16232
rect 22152 16192 22158 16204
rect 18874 16164 18880 16176
rect 17420 16136 18880 16164
rect 18874 16124 18880 16136
rect 18932 16124 18938 16176
rect 21450 16124 21456 16176
rect 21508 16164 21514 16176
rect 22388 16164 22416 16204
rect 22462 16192 22468 16244
rect 22520 16232 22526 16244
rect 22833 16235 22891 16241
rect 22833 16232 22845 16235
rect 22520 16204 22845 16232
rect 22520 16192 22526 16204
rect 22833 16201 22845 16204
rect 22879 16201 22891 16235
rect 22833 16195 22891 16201
rect 24121 16235 24179 16241
rect 24121 16201 24133 16235
rect 24167 16232 24179 16235
rect 24854 16232 24860 16244
rect 24167 16204 24860 16232
rect 24167 16201 24179 16204
rect 24121 16195 24179 16201
rect 24854 16192 24860 16204
rect 24912 16192 24918 16244
rect 21508 16136 22324 16164
rect 22388 16136 23980 16164
rect 21508 16124 21514 16136
rect 17589 16099 17647 16105
rect 17589 16096 17601 16099
rect 16500 16068 17601 16096
rect 17589 16065 17601 16068
rect 17635 16065 17647 16099
rect 18015 16099 18073 16105
rect 18015 16096 18027 16099
rect 17589 16059 17647 16065
rect 17676 16068 18027 16096
rect 17676 16028 17704 16068
rect 18015 16065 18027 16068
rect 18061 16065 18073 16099
rect 18015 16059 18073 16065
rect 18506 16056 18512 16108
rect 18564 16096 18570 16108
rect 22296 16106 22324 16136
rect 22063 16099 22121 16105
rect 22063 16096 22075 16099
rect 18564 16068 22075 16096
rect 18564 16056 18570 16068
rect 22063 16065 22075 16068
rect 22109 16065 22121 16099
rect 22296 16096 22508 16106
rect 23952 16105 23980 16136
rect 23569 16099 23627 16105
rect 23569 16096 23581 16099
rect 22296 16078 23581 16096
rect 22480 16068 23581 16078
rect 22063 16059 22121 16065
rect 23569 16065 23581 16068
rect 23615 16065 23627 16099
rect 23569 16059 23627 16065
rect 23937 16099 23995 16105
rect 23937 16065 23949 16099
rect 23983 16065 23995 16099
rect 23937 16059 23995 16065
rect 15697 16000 17704 16028
rect 17773 16031 17831 16037
rect 17773 15997 17785 16031
rect 17819 15997 17831 16031
rect 17773 15991 17831 15997
rect 17788 15960 17816 15991
rect 20346 15988 20352 16040
rect 20404 16028 20410 16040
rect 21821 16031 21879 16037
rect 21821 16028 21833 16031
rect 20404 16000 21833 16028
rect 20404 15988 20410 16000
rect 21821 15997 21833 16000
rect 21867 15997 21879 16031
rect 21821 15991 21879 15997
rect 12400 15932 13216 15960
rect 17696 15932 17816 15960
rect 12400 15920 12406 15932
rect 17696 15904 17724 15932
rect 7668 15864 8708 15892
rect 5077 15855 5135 15861
rect 9122 15852 9128 15904
rect 9180 15892 9186 15904
rect 11333 15895 11391 15901
rect 11333 15892 11345 15895
rect 9180 15864 11345 15892
rect 9180 15852 9186 15864
rect 11333 15861 11345 15864
rect 11379 15861 11391 15895
rect 11333 15855 11391 15861
rect 14277 15895 14335 15901
rect 14277 15861 14289 15895
rect 14323 15892 14335 15895
rect 16574 15892 16580 15904
rect 14323 15864 16580 15892
rect 14323 15861 14335 15864
rect 14277 15855 14335 15861
rect 16574 15852 16580 15864
rect 16632 15852 16638 15904
rect 17678 15852 17684 15904
rect 17736 15852 17742 15904
rect 21836 15892 21864 15991
rect 22186 15892 22192 15904
rect 21836 15864 22192 15892
rect 22186 15852 22192 15864
rect 22244 15852 22250 15904
rect 23750 15852 23756 15904
rect 23808 15852 23814 15904
rect 1104 15802 24564 15824
rect 1104 15750 3882 15802
rect 3934 15750 3946 15802
rect 3998 15750 4010 15802
rect 4062 15750 4074 15802
rect 4126 15750 4138 15802
rect 4190 15750 9747 15802
rect 9799 15750 9811 15802
rect 9863 15750 9875 15802
rect 9927 15750 9939 15802
rect 9991 15750 10003 15802
rect 10055 15750 15612 15802
rect 15664 15750 15676 15802
rect 15728 15750 15740 15802
rect 15792 15750 15804 15802
rect 15856 15750 15868 15802
rect 15920 15750 21477 15802
rect 21529 15750 21541 15802
rect 21593 15750 21605 15802
rect 21657 15750 21669 15802
rect 21721 15750 21733 15802
rect 21785 15750 24564 15802
rect 1104 15728 24564 15750
rect 1118 15648 1124 15700
rect 1176 15688 1182 15700
rect 2133 15691 2191 15697
rect 2133 15688 2145 15691
rect 1176 15660 2145 15688
rect 1176 15648 1182 15660
rect 2133 15657 2145 15660
rect 2179 15657 2191 15691
rect 3237 15691 3295 15697
rect 3237 15688 3249 15691
rect 2133 15651 2191 15657
rect 2746 15660 3249 15688
rect 1210 15580 1216 15632
rect 1268 15620 1274 15632
rect 2746 15620 2774 15660
rect 3237 15657 3249 15660
rect 3283 15657 3295 15691
rect 3237 15651 3295 15657
rect 3326 15648 3332 15700
rect 3384 15688 3390 15700
rect 3973 15691 4031 15697
rect 3973 15688 3985 15691
rect 3384 15660 3985 15688
rect 3384 15648 3390 15660
rect 3973 15657 3985 15660
rect 4019 15657 4031 15691
rect 3973 15651 4031 15657
rect 4080 15660 5212 15688
rect 1268 15592 2774 15620
rect 1268 15580 1274 15592
rect 4080 15552 4108 15660
rect 5184 15620 5212 15660
rect 5534 15648 5540 15700
rect 5592 15648 5598 15700
rect 11330 15648 11336 15700
rect 11388 15688 11394 15700
rect 12250 15688 12256 15700
rect 11388 15660 12256 15688
rect 11388 15648 11394 15660
rect 12250 15648 12256 15660
rect 12308 15688 12314 15700
rect 12308 15660 13308 15688
rect 12308 15648 12314 15660
rect 5184 15592 7328 15620
rect 2746 15524 4108 15552
rect 1673 15487 1731 15493
rect 1673 15453 1685 15487
rect 1719 15484 1731 15487
rect 2041 15487 2099 15493
rect 2041 15484 2053 15487
rect 1719 15456 2053 15484
rect 1719 15453 1731 15456
rect 1673 15447 1731 15453
rect 2041 15453 2053 15456
rect 2087 15484 2099 15487
rect 2746 15484 2774 15524
rect 7300 15496 7328 15592
rect 9582 15580 9588 15632
rect 9640 15620 9646 15632
rect 11606 15620 11612 15632
rect 9640 15592 11612 15620
rect 9640 15580 9646 15592
rect 11606 15580 11612 15592
rect 11664 15620 11670 15632
rect 12158 15620 12164 15632
rect 11664 15592 12164 15620
rect 11664 15580 11670 15592
rect 12158 15580 12164 15592
rect 12216 15580 12222 15632
rect 12710 15620 12738 15660
rect 12636 15592 12738 15620
rect 13280 15620 13308 15660
rect 13630 15648 13636 15700
rect 13688 15648 13694 15700
rect 15930 15688 15936 15700
rect 14568 15660 15936 15688
rect 13280 15592 14412 15620
rect 12636 15561 12664 15592
rect 14384 15564 14412 15592
rect 12621 15555 12679 15561
rect 12621 15521 12633 15555
rect 12667 15521 12679 15555
rect 12621 15515 12679 15521
rect 14366 15512 14372 15564
rect 14424 15512 14430 15564
rect 2087 15456 2774 15484
rect 3145 15487 3203 15493
rect 2087 15453 2099 15456
rect 2041 15447 2099 15453
rect 3145 15453 3157 15487
rect 3191 15453 3203 15487
rect 3145 15447 3203 15453
rect 4525 15487 4583 15493
rect 4525 15453 4537 15487
rect 4571 15484 4583 15487
rect 4706 15484 4712 15496
rect 4571 15456 4712 15484
rect 4571 15453 4583 15456
rect 4525 15447 4583 15453
rect 1302 15376 1308 15428
rect 1360 15416 1366 15428
rect 2593 15419 2651 15425
rect 1360 15388 1716 15416
rect 1360 15376 1366 15388
rect 1688 15348 1716 15388
rect 2593 15385 2605 15419
rect 2639 15416 2651 15419
rect 2958 15416 2964 15428
rect 2639 15388 2964 15416
rect 2639 15385 2651 15388
rect 2593 15379 2651 15385
rect 2958 15376 2964 15388
rect 3016 15376 3022 15428
rect 2685 15351 2743 15357
rect 2685 15348 2697 15351
rect 1688 15320 2697 15348
rect 2685 15317 2697 15320
rect 2731 15317 2743 15351
rect 3160 15348 3188 15447
rect 4706 15444 4712 15456
rect 4764 15444 4770 15496
rect 4798 15444 4804 15496
rect 4856 15484 4862 15496
rect 7190 15484 7196 15496
rect 4856 15456 7196 15484
rect 4856 15444 4862 15456
rect 7190 15444 7196 15456
rect 7248 15444 7254 15496
rect 7282 15444 7288 15496
rect 7340 15444 7346 15496
rect 8018 15444 8024 15496
rect 8076 15444 8082 15496
rect 9398 15444 9404 15496
rect 9456 15484 9462 15496
rect 9677 15487 9735 15493
rect 9677 15484 9689 15487
rect 9456 15456 9689 15484
rect 9456 15444 9462 15456
rect 9677 15453 9689 15456
rect 9723 15453 9735 15487
rect 9677 15447 9735 15453
rect 10134 15444 10140 15496
rect 10192 15484 10198 15496
rect 10502 15484 10508 15496
rect 10192 15456 10508 15484
rect 10192 15444 10198 15456
rect 10502 15444 10508 15456
rect 10560 15444 10566 15496
rect 12895 15487 12953 15493
rect 12895 15453 12907 15487
rect 12941 15484 12953 15487
rect 12941 15456 13492 15484
rect 12941 15453 12953 15456
rect 12895 15447 12953 15453
rect 3881 15419 3939 15425
rect 3881 15385 3893 15419
rect 3927 15416 3939 15419
rect 8036 15416 8064 15444
rect 3927 15388 8064 15416
rect 3927 15385 3939 15388
rect 3881 15379 3939 15385
rect 11238 15376 11244 15428
rect 11296 15416 11302 15428
rect 12910 15416 12938 15447
rect 11296 15388 12938 15416
rect 13464 15416 13492 15456
rect 14090 15444 14096 15496
rect 14148 15484 14154 15496
rect 14568 15493 14596 15660
rect 15930 15648 15936 15660
rect 15988 15648 15994 15700
rect 16206 15580 16212 15632
rect 16264 15620 16270 15632
rect 16264 15592 19334 15620
rect 16264 15580 16270 15592
rect 15145 15524 18552 15552
rect 14553 15487 14611 15493
rect 14553 15484 14565 15487
rect 14148 15456 14565 15484
rect 14148 15444 14154 15456
rect 14553 15453 14565 15456
rect 14599 15453 14611 15487
rect 14826 15484 14832 15496
rect 14787 15456 14832 15484
rect 14553 15447 14611 15453
rect 14826 15444 14832 15456
rect 14884 15444 14890 15496
rect 15145 15484 15173 15524
rect 18524 15496 18552 15524
rect 14936 15456 15173 15484
rect 14734 15416 14740 15428
rect 13464 15388 14740 15416
rect 11296 15376 11302 15388
rect 14734 15376 14740 15388
rect 14792 15416 14798 15428
rect 14936 15416 14964 15456
rect 16574 15444 16580 15496
rect 16632 15484 16638 15496
rect 17681 15487 17739 15493
rect 17681 15484 17693 15487
rect 16632 15456 17693 15484
rect 16632 15444 16638 15456
rect 17681 15453 17693 15456
rect 17727 15453 17739 15487
rect 17681 15447 17739 15453
rect 18506 15444 18512 15496
rect 18564 15444 18570 15496
rect 14792 15388 14964 15416
rect 14792 15376 14798 15388
rect 15102 15376 15108 15428
rect 15160 15416 15166 15428
rect 17218 15416 17224 15428
rect 15160 15388 17224 15416
rect 15160 15376 15166 15388
rect 17218 15376 17224 15388
rect 17276 15376 17282 15428
rect 19306 15416 19334 15592
rect 19797 15487 19855 15493
rect 19797 15453 19809 15487
rect 19843 15484 19855 15487
rect 19978 15484 19984 15496
rect 19843 15456 19984 15484
rect 19843 15453 19855 15456
rect 19797 15447 19855 15453
rect 19978 15444 19984 15456
rect 20036 15444 20042 15496
rect 23842 15444 23848 15496
rect 23900 15444 23906 15496
rect 22646 15416 22652 15428
rect 19306 15388 22652 15416
rect 22646 15376 22652 15388
rect 22704 15376 22710 15428
rect 24213 15419 24271 15425
rect 24213 15385 24225 15419
rect 24259 15416 24271 15419
rect 24854 15416 24860 15428
rect 24259 15388 24860 15416
rect 24259 15385 24271 15388
rect 24213 15379 24271 15385
rect 24854 15376 24860 15388
rect 24912 15376 24918 15428
rect 5534 15348 5540 15360
rect 3160 15320 5540 15348
rect 2685 15311 2743 15317
rect 5534 15308 5540 15320
rect 5592 15308 5598 15360
rect 11422 15308 11428 15360
rect 11480 15348 11486 15360
rect 13446 15348 13452 15360
rect 11480 15320 13452 15348
rect 11480 15308 11486 15320
rect 13446 15308 13452 15320
rect 13504 15308 13510 15360
rect 13906 15308 13912 15360
rect 13964 15348 13970 15360
rect 14274 15348 14280 15360
rect 13964 15320 14280 15348
rect 13964 15308 13970 15320
rect 14274 15308 14280 15320
rect 14332 15308 14338 15360
rect 14826 15308 14832 15360
rect 14884 15348 14890 15360
rect 15010 15348 15016 15360
rect 14884 15320 15016 15348
rect 14884 15308 14890 15320
rect 15010 15308 15016 15320
rect 15068 15308 15074 15360
rect 15470 15308 15476 15360
rect 15528 15348 15534 15360
rect 15565 15351 15623 15357
rect 15565 15348 15577 15351
rect 15528 15320 15577 15348
rect 15528 15308 15534 15320
rect 15565 15317 15577 15320
rect 15611 15317 15623 15351
rect 15565 15311 15623 15317
rect 17497 15351 17555 15357
rect 17497 15317 17509 15351
rect 17543 15348 17555 15351
rect 18046 15348 18052 15360
rect 17543 15320 18052 15348
rect 17543 15317 17555 15320
rect 17497 15311 17555 15317
rect 18046 15308 18052 15320
rect 18104 15308 18110 15360
rect 19613 15351 19671 15357
rect 19613 15317 19625 15351
rect 19659 15348 19671 15351
rect 20346 15348 20352 15360
rect 19659 15320 20352 15348
rect 19659 15317 19671 15320
rect 19613 15311 19671 15317
rect 20346 15308 20352 15320
rect 20404 15308 20410 15360
rect 20806 15308 20812 15360
rect 20864 15348 20870 15360
rect 21358 15348 21364 15360
rect 20864 15320 21364 15348
rect 20864 15308 20870 15320
rect 21358 15308 21364 15320
rect 21416 15308 21422 15360
rect 1104 15258 24723 15280
rect 1104 15206 6814 15258
rect 6866 15206 6878 15258
rect 6930 15206 6942 15258
rect 6994 15206 7006 15258
rect 7058 15206 7070 15258
rect 7122 15206 12679 15258
rect 12731 15206 12743 15258
rect 12795 15206 12807 15258
rect 12859 15206 12871 15258
rect 12923 15206 12935 15258
rect 12987 15206 18544 15258
rect 18596 15206 18608 15258
rect 18660 15206 18672 15258
rect 18724 15206 18736 15258
rect 18788 15206 18800 15258
rect 18852 15206 24409 15258
rect 24461 15206 24473 15258
rect 24525 15206 24537 15258
rect 24589 15206 24601 15258
rect 24653 15206 24665 15258
rect 24717 15206 24723 15258
rect 1104 15184 24723 15206
rect 1302 15104 1308 15156
rect 1360 15144 1366 15156
rect 3145 15147 3203 15153
rect 3145 15144 3157 15147
rect 1360 15116 3157 15144
rect 1360 15104 1366 15116
rect 3145 15113 3157 15116
rect 3191 15113 3203 15147
rect 3145 15107 3203 15113
rect 3694 15104 3700 15156
rect 3752 15104 3758 15156
rect 4430 15104 4436 15156
rect 4488 15144 4494 15156
rect 7190 15144 7196 15156
rect 4488 15116 7196 15144
rect 4488 15104 4494 15116
rect 7190 15104 7196 15116
rect 7248 15104 7254 15156
rect 8018 15104 8024 15156
rect 8076 15144 8082 15156
rect 10321 15147 10379 15153
rect 8076 15116 10272 15144
rect 8076 15104 8082 15116
rect 658 15036 664 15088
rect 716 15036 722 15088
rect 4338 15076 4344 15088
rect 2976 15048 4344 15076
rect 676 15008 704 15036
rect 1639 15011 1697 15017
rect 1639 15008 1651 15011
rect 676 14980 1651 15008
rect 1639 14977 1651 14980
rect 1685 15008 1697 15011
rect 2976 15008 3004 15048
rect 4338 15036 4344 15048
rect 4396 15036 4402 15088
rect 4522 15076 4528 15088
rect 4448 15048 4528 15076
rect 1685 14980 3004 15008
rect 3053 15011 3111 15017
rect 1685 14977 1697 14980
rect 1639 14971 1697 14977
rect 3053 14977 3065 15011
rect 3099 14977 3111 15011
rect 3053 14971 3111 14977
rect 3605 15011 3663 15017
rect 3605 14977 3617 15011
rect 3651 14977 3663 15011
rect 3605 14971 3663 14977
rect 1394 14900 1400 14952
rect 1452 14900 1458 14952
rect 2222 14764 2228 14816
rect 2280 14804 2286 14816
rect 2409 14807 2467 14813
rect 2409 14804 2421 14807
rect 2280 14776 2421 14804
rect 2280 14764 2286 14776
rect 2409 14773 2421 14776
rect 2455 14773 2467 14807
rect 3068 14804 3096 14971
rect 3620 14940 3648 14971
rect 3694 14968 3700 15020
rect 3752 15008 3758 15020
rect 4448 15008 4476 15048
rect 4522 15036 4528 15048
rect 4580 15076 4586 15088
rect 10244 15076 10272 15116
rect 10321 15113 10333 15147
rect 10367 15144 10379 15147
rect 10367 15116 17264 15144
rect 10367 15113 10379 15116
rect 10321 15107 10379 15113
rect 4580 15048 4844 15076
rect 10244 15048 13308 15076
rect 4580 15036 4586 15048
rect 4816 15038 4844 15048
rect 4875 15041 4933 15047
rect 4875 15038 4887 15041
rect 4816 15010 4887 15038
rect 3752 14980 4476 15008
rect 4875 15007 4887 15010
rect 4921 15007 4933 15041
rect 4875 15001 4933 15007
rect 7375 15011 7433 15017
rect 3752 14968 3758 14980
rect 7375 14977 7387 15011
rect 7421 15008 7433 15011
rect 7466 15008 7472 15020
rect 7421 14980 7472 15008
rect 7421 14977 7433 14980
rect 7375 14971 7433 14977
rect 7466 14968 7472 14980
rect 7524 14968 7530 15020
rect 8478 14968 8484 15020
rect 8536 14968 8542 15020
rect 9398 14968 9404 15020
rect 9456 14968 9462 15020
rect 4522 14940 4528 14952
rect 3620 14912 4528 14940
rect 4522 14900 4528 14912
rect 4580 14900 4586 14952
rect 4617 14943 4675 14949
rect 4617 14909 4629 14943
rect 4663 14909 4675 14943
rect 4617 14903 4675 14909
rect 3786 14832 3792 14884
rect 3844 14872 3850 14884
rect 4154 14872 4160 14884
rect 3844 14844 4160 14872
rect 3844 14832 3850 14844
rect 4154 14832 4160 14844
rect 4212 14872 4218 14884
rect 4632 14872 4660 14903
rect 7098 14900 7104 14952
rect 7156 14900 7162 14952
rect 8294 14900 8300 14952
rect 8352 14940 8358 14952
rect 8665 14943 8723 14949
rect 8665 14940 8677 14943
rect 8352 14912 8677 14940
rect 8352 14900 8358 14912
rect 8665 14909 8677 14912
rect 8711 14909 8723 14943
rect 8665 14903 8723 14909
rect 9030 14900 9036 14952
rect 9088 14940 9094 14952
rect 9518 14943 9576 14949
rect 9518 14940 9530 14943
rect 9088 14912 9530 14940
rect 9088 14900 9094 14912
rect 9518 14909 9530 14912
rect 9564 14909 9576 14943
rect 9518 14903 9576 14909
rect 9677 14943 9735 14949
rect 9677 14909 9689 14943
rect 9723 14940 9735 14943
rect 9723 14912 10180 14940
rect 9723 14909 9735 14912
rect 9677 14903 9735 14909
rect 10152 14884 10180 14912
rect 10226 14900 10232 14952
rect 10284 14940 10290 14952
rect 11974 14940 11980 14952
rect 10284 14912 11980 14940
rect 10284 14900 10290 14912
rect 11974 14900 11980 14912
rect 12032 14900 12038 14952
rect 13170 14900 13176 14952
rect 13228 14900 13234 14952
rect 13280 14940 13308 15048
rect 16574 15036 16580 15088
rect 16632 15036 16638 15088
rect 17236 15076 17264 15116
rect 18138 15104 18144 15156
rect 18196 15144 18202 15156
rect 18966 15144 18972 15156
rect 18196 15116 18972 15144
rect 18196 15104 18202 15116
rect 18966 15104 18972 15116
rect 19024 15104 19030 15156
rect 20901 15147 20959 15153
rect 20901 15113 20913 15147
rect 20947 15144 20959 15147
rect 20947 15116 23980 15144
rect 20947 15113 20959 15116
rect 20901 15107 20959 15113
rect 17236 15048 22508 15076
rect 14277 15011 14335 15017
rect 14277 14977 14289 15011
rect 14323 15008 14335 15011
rect 14323 14980 14688 15008
rect 14323 14977 14335 14980
rect 14277 14971 14335 14977
rect 13280 14912 14320 14940
rect 8113 14875 8171 14881
rect 4212 14844 4660 14872
rect 5460 14844 7236 14872
rect 4212 14832 4218 14844
rect 5460 14804 5488 14844
rect 3068 14776 5488 14804
rect 2409 14767 2467 14773
rect 5534 14764 5540 14816
rect 5592 14804 5598 14816
rect 5629 14807 5687 14813
rect 5629 14804 5641 14807
rect 5592 14776 5641 14804
rect 5592 14764 5598 14776
rect 5629 14773 5641 14776
rect 5675 14773 5687 14807
rect 7208 14804 7236 14844
rect 8113 14841 8125 14875
rect 8159 14872 8171 14875
rect 9125 14875 9183 14881
rect 9125 14872 9137 14875
rect 8159 14844 9137 14872
rect 8159 14841 8171 14844
rect 8113 14835 8171 14841
rect 9125 14841 9137 14844
rect 9171 14841 9183 14875
rect 9125 14835 9183 14841
rect 10134 14832 10140 14884
rect 10192 14832 10198 14884
rect 10594 14804 10600 14816
rect 7208 14776 10600 14804
rect 5629 14767 5687 14773
rect 10594 14764 10600 14776
rect 10652 14764 10658 14816
rect 13188 14804 13216 14900
rect 14292 14884 14320 14912
rect 14458 14900 14464 14952
rect 14516 14900 14522 14952
rect 14660 14940 14688 14980
rect 15470 14968 15476 15020
rect 15528 14968 15534 15020
rect 16298 14968 16304 15020
rect 16356 14968 16362 15020
rect 16592 15008 16620 15036
rect 17201 15011 17259 15017
rect 17201 15008 17213 15011
rect 16592 14980 17213 15008
rect 17201 14977 17213 14980
rect 17247 14977 17259 15011
rect 17201 14971 17259 14977
rect 18690 14968 18696 15020
rect 18748 14968 18754 15020
rect 18874 14968 18880 15020
rect 18932 14968 18938 15020
rect 19420 15011 19478 15017
rect 19420 14977 19432 15011
rect 19466 15008 19478 15011
rect 19978 15008 19984 15020
rect 19466 14980 19984 15008
rect 19466 14977 19478 14980
rect 19420 14971 19478 14977
rect 19978 14968 19984 14980
rect 20036 14968 20042 15020
rect 20622 14968 20628 15020
rect 20680 14968 20686 15020
rect 21177 15011 21235 15017
rect 21177 15008 21189 15011
rect 20824 14980 21189 15008
rect 14826 14940 14832 14952
rect 14660 14912 14832 14940
rect 14826 14900 14832 14912
rect 14884 14900 14890 14952
rect 15194 14900 15200 14952
rect 15252 14900 15258 14952
rect 15335 14943 15393 14949
rect 15335 14909 15347 14943
rect 15381 14940 15393 14943
rect 16316 14940 16344 14968
rect 15381 14912 16344 14940
rect 16945 14943 17003 14949
rect 15381 14909 15393 14912
rect 15335 14903 15393 14909
rect 16945 14909 16957 14943
rect 16991 14909 17003 14943
rect 19153 14943 19211 14949
rect 19153 14940 19165 14943
rect 16945 14903 17003 14909
rect 17972 14912 19165 14940
rect 14274 14832 14280 14884
rect 14332 14832 14338 14884
rect 14918 14832 14924 14884
rect 14976 14832 14982 14884
rect 16117 14807 16175 14813
rect 16117 14804 16129 14807
rect 13188 14776 16129 14804
rect 16117 14773 16129 14776
rect 16163 14773 16175 14807
rect 16960 14804 16988 14903
rect 17972 14816 18000 14912
rect 19153 14909 19165 14912
rect 19199 14909 19211 14943
rect 20824 14940 20852 14980
rect 21177 14977 21189 14980
rect 21223 14977 21235 15011
rect 21177 14971 21235 14977
rect 22002 14968 22008 15020
rect 22060 15008 22066 15020
rect 22281 15011 22339 15017
rect 22281 15008 22293 15011
rect 22060 14980 22293 15008
rect 22060 14968 22066 14980
rect 22281 14977 22293 14980
rect 22327 14977 22339 15011
rect 22480 15008 22508 15048
rect 22548 15011 22606 15017
rect 22548 15008 22560 15011
rect 22480 14980 22560 15008
rect 22281 14971 22339 14977
rect 22548 14977 22560 14980
rect 22594 15008 22606 15011
rect 23014 15008 23020 15020
rect 22594 14980 23020 15008
rect 22594 14977 22606 14980
rect 22548 14971 22606 14977
rect 23014 14968 23020 14980
rect 23072 14968 23078 15020
rect 23952 15017 23980 15116
rect 23937 15011 23995 15017
rect 23937 14977 23949 15011
rect 23983 14977 23995 15011
rect 23937 14971 23995 14977
rect 19153 14903 19211 14909
rect 20548 14912 20852 14940
rect 20901 14943 20959 14949
rect 20548 14881 20576 14912
rect 20901 14909 20913 14943
rect 20947 14940 20959 14943
rect 20947 14912 21404 14940
rect 20947 14909 20959 14912
rect 20901 14903 20959 14909
rect 20533 14875 20591 14881
rect 20533 14841 20545 14875
rect 20579 14841 20591 14875
rect 20533 14835 20591 14841
rect 20717 14875 20775 14881
rect 20717 14841 20729 14875
rect 20763 14872 20775 14875
rect 21082 14872 21088 14884
rect 20763 14844 21088 14872
rect 20763 14841 20775 14844
rect 20717 14835 20775 14841
rect 21082 14832 21088 14844
rect 21140 14832 21146 14884
rect 21376 14816 21404 14912
rect 17954 14804 17960 14816
rect 16960 14776 17960 14804
rect 16117 14767 16175 14773
rect 17954 14764 17960 14776
rect 18012 14764 18018 14816
rect 18322 14764 18328 14816
rect 18380 14764 18386 14816
rect 18782 14764 18788 14816
rect 18840 14764 18846 14816
rect 19150 14764 19156 14816
rect 19208 14804 19214 14816
rect 20806 14804 20812 14816
rect 19208 14776 20812 14804
rect 19208 14764 19214 14776
rect 20806 14764 20812 14776
rect 20864 14764 20870 14816
rect 20990 14764 20996 14816
rect 21048 14764 21054 14816
rect 21358 14764 21364 14816
rect 21416 14764 21422 14816
rect 23290 14764 23296 14816
rect 23348 14804 23354 14816
rect 23661 14807 23719 14813
rect 23661 14804 23673 14807
rect 23348 14776 23673 14804
rect 23348 14764 23354 14776
rect 23661 14773 23673 14776
rect 23707 14773 23719 14807
rect 23661 14767 23719 14773
rect 24118 14764 24124 14816
rect 24176 14764 24182 14816
rect 1104 14714 24564 14736
rect 1104 14662 3882 14714
rect 3934 14662 3946 14714
rect 3998 14662 4010 14714
rect 4062 14662 4074 14714
rect 4126 14662 4138 14714
rect 4190 14662 9747 14714
rect 9799 14662 9811 14714
rect 9863 14662 9875 14714
rect 9927 14662 9939 14714
rect 9991 14662 10003 14714
rect 10055 14662 15612 14714
rect 15664 14662 15676 14714
rect 15728 14662 15740 14714
rect 15792 14662 15804 14714
rect 15856 14662 15868 14714
rect 15920 14662 21477 14714
rect 21529 14662 21541 14714
rect 21593 14662 21605 14714
rect 21657 14662 21669 14714
rect 21721 14662 21733 14714
rect 21785 14662 24564 14714
rect 1104 14640 24564 14662
rect 1578 14560 1584 14612
rect 1636 14560 1642 14612
rect 3053 14603 3111 14609
rect 3053 14600 3065 14603
rect 2746 14572 3065 14600
rect 1118 14492 1124 14544
rect 1176 14532 1182 14544
rect 2746 14532 2774 14572
rect 3053 14569 3065 14572
rect 3099 14569 3111 14603
rect 3053 14563 3111 14569
rect 3970 14560 3976 14612
rect 4028 14560 4034 14612
rect 7098 14560 7104 14612
rect 7156 14600 7162 14612
rect 9953 14603 10011 14609
rect 7156 14572 9674 14600
rect 7156 14560 7162 14572
rect 1176 14504 2774 14532
rect 1176 14492 1182 14504
rect 4154 14492 4160 14544
rect 4212 14532 4218 14544
rect 4212 14504 5120 14532
rect 4212 14492 4218 14504
rect 290 14424 296 14476
rect 348 14464 354 14476
rect 934 14464 940 14476
rect 348 14436 940 14464
rect 348 14424 354 14436
rect 934 14424 940 14436
rect 992 14464 998 14476
rect 4525 14467 4583 14473
rect 4525 14464 4537 14467
rect 992 14436 4537 14464
rect 992 14424 998 14436
rect 4525 14433 4537 14436
rect 4571 14433 4583 14467
rect 4525 14427 4583 14433
rect 4982 14424 4988 14476
rect 5040 14424 5046 14476
rect 5092 14464 5120 14504
rect 5258 14464 5264 14476
rect 5092 14436 5264 14464
rect 5258 14424 5264 14436
rect 5316 14424 5322 14476
rect 5534 14424 5540 14476
rect 5592 14424 5598 14476
rect 6362 14424 6368 14476
rect 6420 14464 6426 14476
rect 8956 14473 8984 14572
rect 9646 14532 9674 14572
rect 9953 14569 9965 14603
rect 9999 14600 10011 14603
rect 10134 14600 10140 14612
rect 9999 14572 10140 14600
rect 9999 14569 10011 14572
rect 9953 14563 10011 14569
rect 10134 14560 10140 14572
rect 10192 14560 10198 14612
rect 11330 14560 11336 14612
rect 11388 14560 11394 14612
rect 13078 14600 13084 14612
rect 12084 14572 13084 14600
rect 11348 14532 11376 14560
rect 9646 14504 11376 14532
rect 11882 14492 11888 14544
rect 11940 14492 11946 14544
rect 11974 14492 11980 14544
rect 12032 14532 12038 14544
rect 12084 14532 12112 14572
rect 13078 14560 13084 14572
rect 13136 14560 13142 14612
rect 14918 14560 14924 14612
rect 14976 14600 14982 14612
rect 15105 14603 15163 14609
rect 15105 14600 15117 14603
rect 14976 14572 15117 14600
rect 14976 14560 14982 14572
rect 15105 14569 15117 14572
rect 15151 14569 15163 14603
rect 15105 14563 15163 14569
rect 15194 14560 15200 14612
rect 15252 14600 15258 14612
rect 15930 14600 15936 14612
rect 15252 14572 15936 14600
rect 15252 14560 15258 14572
rect 15930 14560 15936 14572
rect 15988 14560 15994 14612
rect 16574 14560 16580 14612
rect 16632 14600 16638 14612
rect 17402 14600 17408 14612
rect 16632 14572 17408 14600
rect 16632 14560 16638 14572
rect 17402 14560 17408 14572
rect 17460 14560 17466 14612
rect 18690 14560 18696 14612
rect 18748 14560 18754 14612
rect 18782 14560 18788 14612
rect 18840 14560 18846 14612
rect 20622 14560 20628 14612
rect 20680 14560 20686 14612
rect 20990 14560 20996 14612
rect 21048 14560 21054 14612
rect 21082 14560 21088 14612
rect 21140 14560 21146 14612
rect 21358 14560 21364 14612
rect 21416 14560 21422 14612
rect 23750 14600 23756 14612
rect 22296 14572 23756 14600
rect 12032 14504 12112 14532
rect 12032 14492 12038 14504
rect 7377 14467 7435 14473
rect 7377 14464 7389 14467
rect 6420 14436 7389 14464
rect 6420 14424 6426 14436
rect 7377 14433 7389 14436
rect 7423 14433 7435 14467
rect 7377 14427 7435 14433
rect 8941 14467 8999 14473
rect 8941 14433 8953 14467
rect 8987 14433 8999 14467
rect 8941 14427 8999 14433
rect 10870 14424 10876 14476
rect 10928 14424 10934 14476
rect 11900 14464 11928 14492
rect 12084 14473 12112 14504
rect 12069 14467 12127 14473
rect 11900 14436 12020 14464
rect 2593 14399 2651 14405
rect 2593 14365 2605 14399
rect 2639 14396 2651 14399
rect 2682 14396 2688 14408
rect 2639 14368 2688 14396
rect 2639 14365 2651 14368
rect 2593 14359 2651 14365
rect 2682 14356 2688 14368
rect 2740 14396 2746 14408
rect 2961 14399 3019 14405
rect 2961 14396 2973 14399
rect 2740 14368 2973 14396
rect 2740 14356 2746 14368
rect 2961 14365 2973 14368
rect 3007 14365 3019 14399
rect 2961 14359 3019 14365
rect 4341 14399 4399 14405
rect 4341 14365 4353 14399
rect 4387 14396 4399 14399
rect 4430 14396 4436 14408
rect 4387 14368 4436 14396
rect 4387 14365 4399 14368
rect 4341 14359 4399 14365
rect 4430 14356 4436 14368
rect 4488 14356 4494 14408
rect 5442 14405 5448 14408
rect 5399 14399 5448 14405
rect 5399 14365 5411 14399
rect 5445 14365 5448 14399
rect 5399 14359 5448 14365
rect 5442 14356 5448 14359
rect 5500 14356 5506 14408
rect 7558 14356 7564 14408
rect 7616 14396 7622 14408
rect 7651 14399 7709 14405
rect 7651 14396 7663 14399
rect 7616 14368 7663 14396
rect 7616 14356 7622 14368
rect 7651 14365 7663 14368
rect 7697 14396 7709 14399
rect 8018 14396 8024 14408
rect 7697 14368 8024 14396
rect 7697 14365 7709 14368
rect 7651 14359 7709 14365
rect 8018 14356 8024 14368
rect 8076 14356 8082 14408
rect 8754 14356 8760 14408
rect 8812 14396 8818 14408
rect 9183 14399 9241 14405
rect 9183 14396 9195 14399
rect 8812 14368 9195 14396
rect 8812 14356 8818 14368
rect 9183 14365 9195 14368
rect 9229 14365 9241 14399
rect 9183 14359 9241 14365
rect 1486 14288 1492 14340
rect 1544 14288 1550 14340
rect 3881 14331 3939 14337
rect 3881 14297 3893 14331
rect 3927 14328 3939 14331
rect 4522 14328 4528 14340
rect 3927 14300 4528 14328
rect 3927 14297 3939 14300
rect 3881 14291 3939 14297
rect 4522 14288 4528 14300
rect 4580 14288 4586 14340
rect 7190 14288 7196 14340
rect 7248 14328 7254 14340
rect 10888 14328 10916 14424
rect 11885 14399 11943 14405
rect 11885 14365 11897 14399
rect 11931 14365 11943 14399
rect 11992 14396 12020 14436
rect 12069 14433 12081 14467
rect 12115 14433 12127 14467
rect 12069 14427 12127 14433
rect 12311 14399 12369 14405
rect 12311 14396 12323 14399
rect 11992 14368 12323 14396
rect 11885 14359 11943 14365
rect 12311 14365 12323 14368
rect 12357 14365 12369 14399
rect 12311 14359 12369 14365
rect 7248 14300 10916 14328
rect 7248 14288 7254 14300
rect 2314 14220 2320 14272
rect 2372 14260 2378 14272
rect 4890 14260 4896 14272
rect 2372 14232 4896 14260
rect 2372 14220 2378 14232
rect 4890 14220 4896 14232
rect 4948 14220 4954 14272
rect 5074 14220 5080 14272
rect 5132 14260 5138 14272
rect 6181 14263 6239 14269
rect 6181 14260 6193 14263
rect 5132 14232 6193 14260
rect 5132 14220 5138 14232
rect 6181 14229 6193 14232
rect 6227 14229 6239 14263
rect 6181 14223 6239 14229
rect 8294 14220 8300 14272
rect 8352 14260 8358 14272
rect 8389 14263 8447 14269
rect 8389 14260 8401 14263
rect 8352 14232 8401 14260
rect 8352 14220 8358 14232
rect 8389 14229 8401 14232
rect 8435 14229 8447 14263
rect 11900 14260 11928 14359
rect 14090 14356 14096 14408
rect 14148 14356 14154 14408
rect 14335 14399 14393 14405
rect 14335 14396 14347 14399
rect 14200 14368 14347 14396
rect 14200 14340 14228 14368
rect 14335 14365 14347 14368
rect 14381 14396 14393 14399
rect 15194 14396 15200 14408
rect 14381 14368 15200 14396
rect 14381 14365 14393 14368
rect 14335 14359 14393 14365
rect 15194 14356 15200 14368
rect 15252 14356 15258 14408
rect 17494 14356 17500 14408
rect 17552 14356 17558 14408
rect 17678 14356 17684 14408
rect 17736 14356 17742 14408
rect 18708 14396 18736 14560
rect 18800 14464 18828 14560
rect 19521 14467 19579 14473
rect 19521 14464 19533 14467
rect 18800 14436 19533 14464
rect 19521 14433 19533 14436
rect 19567 14433 19579 14467
rect 20640 14464 20668 14560
rect 21008 14532 21036 14560
rect 21008 14504 21496 14532
rect 21000 14464 21119 14472
rect 20640 14444 21119 14464
rect 20640 14436 21028 14444
rect 19521 14427 19579 14433
rect 19245 14399 19303 14405
rect 19245 14396 19257 14399
rect 17788 14395 17982 14396
rect 17788 14389 18013 14395
rect 17788 14368 17967 14389
rect 14182 14288 14188 14340
rect 14240 14288 14246 14340
rect 17512 14328 17540 14356
rect 17788 14328 17816 14368
rect 17954 14358 17967 14368
rect 17955 14355 17967 14358
rect 18001 14355 18013 14389
rect 18708 14368 19257 14396
rect 19245 14365 19257 14368
rect 19291 14365 19303 14399
rect 19245 14359 19303 14365
rect 19337 14399 19395 14405
rect 19337 14365 19349 14399
rect 19383 14365 19395 14399
rect 19613 14399 19671 14405
rect 19613 14396 19625 14399
rect 19337 14359 19395 14365
rect 19444 14368 19625 14396
rect 17955 14349 18013 14355
rect 17512 14300 17816 14328
rect 18138 14288 18144 14340
rect 18196 14328 18202 14340
rect 19352 14328 19380 14359
rect 18196 14300 19380 14328
rect 18196 14288 18202 14300
rect 12434 14260 12440 14272
rect 11900 14232 12440 14260
rect 8389 14223 8447 14229
rect 12434 14220 12440 14232
rect 12492 14220 12498 14272
rect 13078 14220 13084 14272
rect 13136 14220 13142 14272
rect 13446 14220 13452 14272
rect 13504 14260 13510 14272
rect 14734 14260 14740 14272
rect 13504 14232 14740 14260
rect 13504 14220 13510 14232
rect 14734 14220 14740 14232
rect 14792 14220 14798 14272
rect 15010 14220 15016 14272
rect 15068 14260 15074 14272
rect 16206 14260 16212 14272
rect 15068 14232 16212 14260
rect 15068 14220 15074 14232
rect 16206 14220 16212 14232
rect 16264 14220 16270 14272
rect 17678 14220 17684 14272
rect 17736 14260 17742 14272
rect 19444 14260 19472 14368
rect 19613 14365 19625 14368
rect 19659 14365 19671 14399
rect 19613 14359 19671 14365
rect 19887 14399 19945 14405
rect 19887 14365 19899 14399
rect 19933 14396 19945 14399
rect 19978 14396 19984 14408
rect 19933 14368 19984 14396
rect 19933 14365 19945 14368
rect 19887 14359 19945 14365
rect 19978 14356 19984 14368
rect 20036 14356 20042 14408
rect 20346 14356 20352 14408
rect 20404 14396 20410 14408
rect 20993 14399 21051 14405
rect 20404 14392 20944 14396
rect 20993 14392 21005 14399
rect 20404 14368 21005 14392
rect 20404 14356 20410 14368
rect 20916 14365 21005 14368
rect 21039 14365 21051 14399
rect 21091 14396 21119 14444
rect 21468 14405 21496 14504
rect 22296 14405 22324 14572
rect 23750 14560 23756 14572
rect 23808 14560 23814 14612
rect 22557 14535 22615 14541
rect 22557 14501 22569 14535
rect 22603 14501 22615 14535
rect 22557 14495 22615 14501
rect 21269 14399 21327 14405
rect 21269 14396 21281 14399
rect 21091 14368 21281 14396
rect 20916 14364 21051 14365
rect 20993 14359 21051 14364
rect 21269 14365 21281 14368
rect 21315 14365 21327 14399
rect 21269 14359 21327 14365
rect 21453 14399 21511 14405
rect 21453 14365 21465 14399
rect 21499 14365 21511 14399
rect 21453 14359 21511 14365
rect 22281 14399 22339 14405
rect 22281 14365 22293 14399
rect 22327 14365 22339 14399
rect 22281 14359 22339 14365
rect 22465 14399 22523 14405
rect 22465 14365 22477 14399
rect 22511 14396 22523 14399
rect 22572 14396 22600 14495
rect 22830 14492 22836 14544
rect 22888 14492 22894 14544
rect 23290 14492 23296 14544
rect 23348 14492 23354 14544
rect 23584 14504 24072 14532
rect 23308 14464 23336 14492
rect 22756 14436 23336 14464
rect 22756 14405 22784 14436
rect 22511 14368 22600 14396
rect 22741 14399 22799 14405
rect 22511 14365 22523 14368
rect 22465 14359 22523 14365
rect 22741 14365 22753 14399
rect 22787 14365 22799 14399
rect 22741 14359 22799 14365
rect 23014 14356 23020 14408
rect 23072 14356 23078 14408
rect 23584 14396 23612 14504
rect 24044 14473 24072 14504
rect 24029 14467 24087 14473
rect 24029 14433 24041 14467
rect 24075 14433 24087 14467
rect 24029 14427 24087 14433
rect 23216 14368 23612 14396
rect 19521 14331 19579 14337
rect 19521 14297 19533 14331
rect 19567 14328 19579 14331
rect 20806 14328 20812 14340
rect 19567 14300 20812 14328
rect 19567 14297 19579 14300
rect 19521 14291 19579 14297
rect 20806 14288 20812 14300
rect 20864 14288 20870 14340
rect 22373 14331 22431 14337
rect 22373 14297 22385 14331
rect 22419 14328 22431 14331
rect 23216 14328 23244 14368
rect 23750 14356 23756 14408
rect 23808 14356 23814 14408
rect 23842 14356 23848 14408
rect 23900 14356 23906 14408
rect 22419 14300 23244 14328
rect 23293 14331 23351 14337
rect 22419 14297 22431 14300
rect 22373 14291 22431 14297
rect 23293 14297 23305 14331
rect 23339 14328 23351 14331
rect 24029 14331 24087 14337
rect 24029 14328 24041 14331
rect 23339 14300 24041 14328
rect 23339 14297 23351 14300
rect 23293 14291 23351 14297
rect 24029 14297 24041 14300
rect 24075 14297 24087 14331
rect 24029 14291 24087 14297
rect 19794 14260 19800 14272
rect 17736 14232 19800 14260
rect 17736 14220 17742 14232
rect 19794 14220 19800 14232
rect 19852 14220 19858 14272
rect 21174 14220 21180 14272
rect 21232 14260 21238 14272
rect 23014 14260 23020 14272
rect 21232 14232 23020 14260
rect 21232 14220 21238 14232
rect 23014 14220 23020 14232
rect 23072 14220 23078 14272
rect 23569 14263 23627 14269
rect 23569 14229 23581 14263
rect 23615 14260 23627 14263
rect 24854 14260 24860 14272
rect 23615 14232 24860 14260
rect 23615 14229 23627 14232
rect 23569 14223 23627 14229
rect 24854 14220 24860 14232
rect 24912 14220 24918 14272
rect 1104 14170 24723 14192
rect 1104 14118 6814 14170
rect 6866 14118 6878 14170
rect 6930 14118 6942 14170
rect 6994 14118 7006 14170
rect 7058 14118 7070 14170
rect 7122 14118 12679 14170
rect 12731 14118 12743 14170
rect 12795 14118 12807 14170
rect 12859 14118 12871 14170
rect 12923 14118 12935 14170
rect 12987 14118 18544 14170
rect 18596 14118 18608 14170
rect 18660 14118 18672 14170
rect 18724 14118 18736 14170
rect 18788 14118 18800 14170
rect 18852 14118 24409 14170
rect 24461 14118 24473 14170
rect 24525 14118 24537 14170
rect 24589 14118 24601 14170
rect 24653 14118 24665 14170
rect 24717 14118 24723 14170
rect 1104 14096 24723 14118
rect 1486 14016 1492 14068
rect 1544 14056 1550 14068
rect 7650 14056 7656 14068
rect 1544 14028 7656 14056
rect 1544 14016 1550 14028
rect 7650 14016 7656 14028
rect 7708 14016 7714 14068
rect 7742 14016 7748 14068
rect 7800 14056 7806 14068
rect 8941 14059 8999 14065
rect 8941 14056 8953 14059
rect 7800 14028 8953 14056
rect 7800 14016 7806 14028
rect 8941 14025 8953 14028
rect 8987 14025 8999 14059
rect 12066 14056 12072 14068
rect 8941 14019 8999 14025
rect 10318 14028 12072 14056
rect 1670 13988 1676 14000
rect 1504 13960 1676 13988
rect 1504 13864 1532 13960
rect 1670 13948 1676 13960
rect 1728 13948 1734 14000
rect 6362 13988 6368 14000
rect 4908 13960 6368 13988
rect 3679 13953 3737 13959
rect 2406 13880 2412 13932
rect 2464 13880 2470 13932
rect 2590 13929 2596 13932
rect 2547 13923 2596 13929
rect 2547 13889 2559 13923
rect 2593 13889 2596 13923
rect 2547 13883 2596 13889
rect 2590 13880 2596 13883
rect 2648 13880 2654 13932
rect 3679 13920 3691 13953
rect 3252 13919 3691 13920
rect 3725 13950 3737 13953
rect 3725 13919 3740 13950
rect 4908 13929 4936 13960
rect 6362 13948 6368 13960
rect 6420 13948 6426 14000
rect 10318 13959 10346 14028
rect 12066 14016 12072 14028
rect 12124 14016 12130 14068
rect 12158 14016 12164 14068
rect 12216 14056 12222 14068
rect 13354 14056 13360 14068
rect 12216 14028 13360 14056
rect 12216 14016 12222 14028
rect 13354 14016 13360 14028
rect 13412 14056 13418 14068
rect 13633 14059 13691 14065
rect 13633 14056 13645 14059
rect 13412 14028 13645 14056
rect 13412 14016 13418 14028
rect 13633 14025 13645 14028
rect 13679 14025 13691 14059
rect 13633 14019 13691 14025
rect 14016 14028 17354 14056
rect 14016 13988 14044 14028
rect 11072 13960 11744 13988
rect 10303 13953 10361 13959
rect 3252 13892 3740 13919
rect 4893 13923 4951 13929
rect 1486 13812 1492 13864
rect 1544 13812 1550 13864
rect 1673 13855 1731 13861
rect 1673 13821 1685 13855
rect 1719 13852 1731 13855
rect 2133 13855 2191 13861
rect 1719 13824 1900 13852
rect 1719 13821 1731 13824
rect 1673 13815 1731 13821
rect 1872 13796 1900 13824
rect 2133 13821 2145 13855
rect 2179 13852 2191 13855
rect 2222 13852 2228 13864
rect 2179 13824 2228 13852
rect 2179 13821 2191 13824
rect 2133 13815 2191 13821
rect 2222 13812 2228 13824
rect 2280 13812 2286 13864
rect 2682 13812 2688 13864
rect 2740 13812 2746 13864
rect 2866 13812 2872 13864
rect 2924 13852 2930 13864
rect 3252 13852 3280 13892
rect 4893 13889 4905 13923
rect 4939 13889 4951 13923
rect 5166 13920 5172 13932
rect 5127 13892 5172 13920
rect 4893 13883 4951 13889
rect 5166 13880 5172 13892
rect 5224 13880 5230 13932
rect 5534 13880 5540 13932
rect 5592 13920 5598 13932
rect 6546 13920 6552 13932
rect 5592 13892 6552 13920
rect 5592 13880 5598 13892
rect 6546 13880 6552 13892
rect 6604 13920 6610 13932
rect 7285 13923 7343 13929
rect 7285 13920 7297 13923
rect 6604 13892 7297 13920
rect 6604 13880 6610 13892
rect 7285 13889 7297 13892
rect 7331 13889 7343 13923
rect 7285 13883 7343 13889
rect 7466 13880 7472 13932
rect 7524 13880 7530 13932
rect 8294 13880 8300 13932
rect 8352 13880 8358 13932
rect 9306 13880 9312 13932
rect 9364 13880 9370 13932
rect 10303 13919 10315 13953
rect 10349 13919 10361 13953
rect 10303 13913 10361 13919
rect 2924 13824 3280 13852
rect 3421 13855 3479 13861
rect 2924 13812 2930 13824
rect 3421 13821 3433 13855
rect 3467 13821 3479 13855
rect 3421 13815 3479 13821
rect 1854 13744 1860 13796
rect 1912 13744 1918 13796
rect 1946 13676 1952 13728
rect 2004 13716 2010 13728
rect 2866 13716 2872 13728
rect 2004 13688 2872 13716
rect 2004 13676 2010 13688
rect 2866 13676 2872 13688
rect 2924 13676 2930 13728
rect 3234 13676 3240 13728
rect 3292 13716 3298 13728
rect 3329 13719 3387 13725
rect 3329 13716 3341 13719
rect 3292 13688 3341 13716
rect 3292 13676 3298 13688
rect 3329 13685 3341 13688
rect 3375 13685 3387 13719
rect 3436 13716 3464 13815
rect 6454 13812 6460 13864
rect 6512 13852 6518 13864
rect 6730 13852 6736 13864
rect 6512 13824 6736 13852
rect 6512 13812 6518 13824
rect 6730 13812 6736 13824
rect 6788 13812 6794 13864
rect 7101 13855 7159 13861
rect 7101 13821 7113 13855
rect 7147 13852 7159 13855
rect 7190 13852 7196 13864
rect 7147 13824 7196 13852
rect 7147 13821 7159 13824
rect 7101 13815 7159 13821
rect 7190 13812 7196 13824
rect 7248 13852 7254 13864
rect 7484 13852 7512 13880
rect 7248 13824 7512 13852
rect 7248 13812 7254 13824
rect 8018 13812 8024 13864
rect 8076 13812 8082 13864
rect 8202 13861 8208 13864
rect 8159 13855 8208 13861
rect 8159 13821 8171 13855
rect 8205 13821 8208 13855
rect 8159 13815 8208 13821
rect 8202 13812 8208 13815
rect 8260 13852 8266 13864
rect 9324 13852 9352 13880
rect 8260 13824 9352 13852
rect 10045 13855 10103 13861
rect 8260 13812 8266 13824
rect 10045 13821 10057 13855
rect 10091 13821 10103 13855
rect 10045 13815 10103 13821
rect 7466 13784 7472 13796
rect 5828 13756 7472 13784
rect 3786 13716 3792 13728
rect 3436 13688 3792 13716
rect 3329 13679 3387 13685
rect 3786 13676 3792 13688
rect 3844 13676 3850 13728
rect 4430 13676 4436 13728
rect 4488 13676 4494 13728
rect 4614 13676 4620 13728
rect 4672 13716 4678 13728
rect 5828 13716 5856 13756
rect 7466 13744 7472 13756
rect 7524 13744 7530 13796
rect 7742 13744 7748 13796
rect 7800 13744 7806 13796
rect 10060 13784 10088 13815
rect 11072 13793 11100 13960
rect 11517 13923 11575 13929
rect 11517 13889 11529 13923
rect 11563 13889 11575 13923
rect 11716 13920 11744 13960
rect 13832 13960 14044 13988
rect 11716 13892 11834 13920
rect 11517 13883 11575 13889
rect 9048 13756 10088 13784
rect 9048 13728 9076 13756
rect 4672 13688 5856 13716
rect 4672 13676 4678 13688
rect 5902 13676 5908 13728
rect 5960 13676 5966 13728
rect 9030 13676 9036 13728
rect 9088 13676 9094 13728
rect 10060 13716 10088 13756
rect 11057 13787 11115 13793
rect 11057 13753 11069 13787
rect 11103 13753 11115 13787
rect 11057 13747 11115 13753
rect 11330 13744 11336 13796
rect 11388 13784 11394 13796
rect 11520 13784 11548 13883
rect 11606 13812 11612 13864
rect 11664 13852 11670 13864
rect 11701 13855 11759 13861
rect 11701 13852 11713 13855
rect 11664 13824 11713 13852
rect 11664 13812 11670 13824
rect 11701 13821 11713 13824
rect 11747 13821 11759 13855
rect 11806 13852 11834 13892
rect 12434 13880 12440 13932
rect 12492 13880 12498 13932
rect 12710 13880 12716 13932
rect 12768 13880 12774 13932
rect 13357 13923 13415 13929
rect 13357 13889 13369 13923
rect 13403 13920 13415 13923
rect 13832 13920 13860 13960
rect 14734 13948 14740 14000
rect 14792 13948 14798 14000
rect 15286 13948 15292 14000
rect 15344 13988 15350 14000
rect 15562 13988 15568 14000
rect 15344 13960 15568 13988
rect 15344 13948 15350 13960
rect 15562 13948 15568 13960
rect 15620 13988 15626 14000
rect 15620 13960 16954 13988
rect 15620 13948 15626 13960
rect 13403 13892 13860 13920
rect 13403 13889 13415 13892
rect 13357 13883 13415 13889
rect 13906 13880 13912 13932
rect 13964 13880 13970 13932
rect 13998 13880 14004 13932
rect 14056 13880 14062 13932
rect 14182 13880 14188 13932
rect 14240 13920 14246 13932
rect 14369 13923 14427 13929
rect 14369 13920 14381 13923
rect 14240 13892 14381 13920
rect 14240 13880 14246 13892
rect 14369 13889 14381 13892
rect 14415 13889 14427 13923
rect 14369 13883 14427 13889
rect 14550 13880 14556 13932
rect 14608 13920 14614 13932
rect 16926 13929 16954 13960
rect 15439 13923 15497 13929
rect 15439 13920 15451 13923
rect 14608 13892 15451 13920
rect 14608 13880 14614 13892
rect 15439 13889 15451 13892
rect 15485 13889 15497 13923
rect 15439 13883 15497 13889
rect 16911 13923 16969 13929
rect 16911 13889 16923 13923
rect 16957 13889 16969 13923
rect 16911 13883 16969 13889
rect 12161 13855 12219 13861
rect 12161 13852 12173 13855
rect 11806 13824 12173 13852
rect 11701 13815 11759 13821
rect 12161 13821 12173 13824
rect 12207 13821 12219 13855
rect 12575 13855 12633 13861
rect 12575 13852 12587 13855
rect 12161 13815 12219 13821
rect 12250 13824 12587 13852
rect 11790 13784 11796 13796
rect 11388 13756 11796 13784
rect 11388 13744 11394 13756
rect 11790 13744 11796 13756
rect 11848 13744 11854 13796
rect 10870 13716 10876 13728
rect 10060 13688 10876 13716
rect 10870 13676 10876 13688
rect 10928 13676 10934 13728
rect 11606 13676 11612 13728
rect 11664 13716 11670 13728
rect 12250 13716 12278 13824
rect 12575 13821 12587 13824
rect 12621 13821 12633 13855
rect 12575 13815 12633 13821
rect 13078 13812 13084 13864
rect 13136 13852 13142 13864
rect 13136 13824 13478 13852
rect 13136 13812 13142 13824
rect 15010 13812 15016 13864
rect 15068 13852 15074 13864
rect 15197 13855 15255 13861
rect 15197 13852 15209 13855
rect 15068 13824 15209 13852
rect 15068 13812 15074 13824
rect 15197 13821 15209 13824
rect 15243 13821 15255 13855
rect 15197 13815 15255 13821
rect 16206 13812 16212 13864
rect 16264 13852 16270 13864
rect 16669 13855 16727 13861
rect 16669 13852 16681 13855
rect 16264 13824 16681 13852
rect 16264 13812 16270 13824
rect 16669 13821 16681 13824
rect 16715 13821 16727 13855
rect 17326 13852 17354 14028
rect 18046 14016 18052 14068
rect 18104 14016 18110 14068
rect 18138 14016 18144 14068
rect 18196 14016 18202 14068
rect 18322 14016 18328 14068
rect 18380 14016 18386 14068
rect 18601 14059 18659 14065
rect 18601 14025 18613 14059
rect 18647 14056 18659 14059
rect 18874 14056 18880 14068
rect 18647 14028 18880 14056
rect 18647 14025 18659 14028
rect 18601 14019 18659 14025
rect 18874 14016 18880 14028
rect 18932 14016 18938 14068
rect 19886 14016 19892 14068
rect 19944 14056 19950 14068
rect 20162 14056 20168 14068
rect 19944 14028 20168 14056
rect 19944 14016 19950 14028
rect 20162 14016 20168 14028
rect 20220 14016 20226 14068
rect 22278 14016 22284 14068
rect 22336 14056 22342 14068
rect 22373 14059 22431 14065
rect 22373 14056 22385 14059
rect 22336 14028 22385 14056
rect 22336 14016 22342 14028
rect 22373 14025 22385 14028
rect 22419 14025 22431 14059
rect 22373 14019 22431 14025
rect 22741 14059 22799 14065
rect 22741 14025 22753 14059
rect 22787 14056 22799 14059
rect 23842 14056 23848 14068
rect 22787 14028 23848 14056
rect 22787 14025 22799 14028
rect 22741 14019 22799 14025
rect 23842 14016 23848 14028
rect 23900 14016 23906 14068
rect 23937 14059 23995 14065
rect 23937 14025 23949 14059
rect 23983 14025 23995 14059
rect 23937 14019 23995 14025
rect 18064 13929 18092 14016
rect 18049 13923 18107 13929
rect 18049 13889 18061 13923
rect 18095 13889 18107 13923
rect 18340 13920 18368 14016
rect 18966 13948 18972 14000
rect 19024 13988 19030 14000
rect 21174 13988 21180 14000
rect 19024 13960 21180 13988
rect 19024 13948 19030 13960
rect 21174 13948 21180 13960
rect 21232 13948 21238 14000
rect 22186 13988 22192 14000
rect 21468 13960 22192 13988
rect 18785 13923 18843 13929
rect 18785 13920 18797 13923
rect 18340 13892 18797 13920
rect 18049 13883 18107 13889
rect 18785 13889 18797 13892
rect 18831 13889 18843 13923
rect 18785 13883 18843 13889
rect 19794 13880 19800 13932
rect 19852 13920 19858 13932
rect 21468 13920 21496 13960
rect 22186 13948 22192 13960
rect 22244 13988 22250 14000
rect 22244 13960 22968 13988
rect 22244 13948 22250 13960
rect 19852 13892 21496 13920
rect 21545 13923 21603 13929
rect 19852 13880 19858 13892
rect 21545 13889 21557 13923
rect 21591 13889 21603 13923
rect 21545 13883 21603 13889
rect 21082 13852 21088 13864
rect 17326 13824 21088 13852
rect 16669 13815 16727 13821
rect 15948 13756 16528 13784
rect 11664 13688 12278 13716
rect 11664 13676 11670 13688
rect 13078 13676 13084 13728
rect 13136 13716 13142 13728
rect 13538 13716 13544 13728
rect 13136 13688 13544 13716
rect 13136 13676 13142 13688
rect 13538 13676 13544 13688
rect 13596 13676 13602 13728
rect 14826 13676 14832 13728
rect 14884 13716 14890 13728
rect 14921 13719 14979 13725
rect 14921 13716 14933 13719
rect 14884 13688 14933 13716
rect 14884 13676 14890 13688
rect 14921 13685 14933 13688
rect 14967 13716 14979 13719
rect 15948 13716 15976 13756
rect 16500 13728 16528 13756
rect 14967 13688 15976 13716
rect 14967 13685 14979 13688
rect 14921 13679 14979 13685
rect 16206 13676 16212 13728
rect 16264 13676 16270 13728
rect 16482 13676 16488 13728
rect 16540 13676 16546 13728
rect 16684 13716 16712 13815
rect 21082 13812 21088 13824
rect 21140 13852 21146 13864
rect 21560 13852 21588 13883
rect 22094 13880 22100 13932
rect 22152 13880 22158 13932
rect 22278 13880 22284 13932
rect 22336 13880 22342 13932
rect 22554 13880 22560 13932
rect 22612 13880 22618 13932
rect 22940 13929 22968 13960
rect 23014 13948 23020 14000
rect 23072 13988 23078 14000
rect 23072 13960 23152 13988
rect 23072 13948 23078 13960
rect 23124 13950 23152 13960
rect 23183 13953 23241 13959
rect 23183 13950 23195 13953
rect 22925 13923 22983 13929
rect 22673 13913 22731 13919
rect 22673 13879 22685 13913
rect 22719 13910 22731 13913
rect 22719 13879 22750 13910
rect 22925 13889 22937 13923
rect 22971 13889 22983 13923
rect 23124 13922 23195 13950
rect 23183 13919 23195 13922
rect 23229 13919 23241 13953
rect 23750 13948 23756 14000
rect 23808 13988 23814 14000
rect 23952 13988 23980 14019
rect 23808 13960 23980 13988
rect 23808 13948 23814 13960
rect 23183 13913 23241 13919
rect 22925 13883 22983 13889
rect 22673 13873 22750 13879
rect 21140 13824 21588 13852
rect 22722 13852 22750 13873
rect 22830 13852 22836 13864
rect 22722 13824 22836 13852
rect 21140 13812 21146 13824
rect 22830 13812 22836 13824
rect 22888 13812 22894 13864
rect 18322 13784 18328 13796
rect 17326 13756 18328 13784
rect 17326 13716 17354 13756
rect 18322 13744 18328 13756
rect 18380 13784 18386 13796
rect 19150 13784 19156 13796
rect 18380 13756 19156 13784
rect 18380 13744 18386 13756
rect 19150 13744 19156 13756
rect 19208 13744 19214 13796
rect 20346 13744 20352 13796
rect 20404 13784 20410 13796
rect 20404 13756 22692 13784
rect 20404 13744 20410 13756
rect 22664 13728 22692 13756
rect 16684 13688 17354 13716
rect 17678 13676 17684 13728
rect 17736 13676 17742 13728
rect 21358 13676 21364 13728
rect 21416 13676 21422 13728
rect 22186 13676 22192 13728
rect 22244 13676 22250 13728
rect 22646 13676 22652 13728
rect 22704 13676 22710 13728
rect 1104 13626 24564 13648
rect 1104 13574 3882 13626
rect 3934 13574 3946 13626
rect 3998 13574 4010 13626
rect 4062 13574 4074 13626
rect 4126 13574 4138 13626
rect 4190 13574 9747 13626
rect 9799 13574 9811 13626
rect 9863 13574 9875 13626
rect 9927 13574 9939 13626
rect 9991 13574 10003 13626
rect 10055 13574 15612 13626
rect 15664 13574 15676 13626
rect 15728 13574 15740 13626
rect 15792 13574 15804 13626
rect 15856 13574 15868 13626
rect 15920 13574 21477 13626
rect 21529 13574 21541 13626
rect 21593 13574 21605 13626
rect 21657 13574 21669 13626
rect 21721 13574 21733 13626
rect 21785 13574 24564 13626
rect 1104 13552 24564 13574
rect 2501 13515 2559 13521
rect 2501 13481 2513 13515
rect 2547 13512 2559 13515
rect 2682 13512 2688 13524
rect 2547 13484 2688 13512
rect 2547 13481 2559 13484
rect 2501 13475 2559 13481
rect 2682 13472 2688 13484
rect 2740 13472 2746 13524
rect 4982 13472 4988 13524
rect 5040 13512 5046 13524
rect 5077 13515 5135 13521
rect 5077 13512 5089 13515
rect 5040 13484 5089 13512
rect 5040 13472 5046 13484
rect 5077 13481 5089 13484
rect 5123 13481 5135 13515
rect 5077 13475 5135 13481
rect 7650 13472 7656 13524
rect 7708 13472 7714 13524
rect 11882 13512 11888 13524
rect 7760 13484 11888 13512
rect 5902 13404 5908 13456
rect 5960 13444 5966 13456
rect 6457 13447 6515 13453
rect 6457 13444 6469 13447
rect 5960 13416 6469 13444
rect 5960 13404 5966 13416
rect 6457 13413 6469 13416
rect 6503 13413 6515 13447
rect 6457 13407 6515 13413
rect 3694 13336 3700 13388
rect 3752 13336 3758 13388
rect 3786 13336 3792 13388
rect 3844 13376 3850 13388
rect 4065 13379 4123 13385
rect 4065 13376 4077 13379
rect 3844 13348 4077 13376
rect 3844 13336 3850 13348
rect 4065 13345 4077 13348
rect 4111 13345 4123 13379
rect 4065 13339 4123 13345
rect 4890 13336 4896 13388
rect 4948 13376 4954 13388
rect 5166 13376 5172 13388
rect 4948 13348 5172 13376
rect 4948 13336 4954 13348
rect 5166 13336 5172 13348
rect 5224 13336 5230 13388
rect 6086 13336 6092 13388
rect 6144 13376 6150 13388
rect 6850 13379 6908 13385
rect 6850 13376 6862 13379
rect 6144 13348 6862 13376
rect 6144 13336 6150 13348
rect 6850 13345 6862 13348
rect 6896 13345 6908 13379
rect 7374 13376 7380 13388
rect 6850 13339 6908 13345
rect 7024 13348 7380 13376
rect 1394 13268 1400 13320
rect 1452 13308 1458 13320
rect 1489 13311 1547 13317
rect 1489 13308 1501 13311
rect 1452 13280 1501 13308
rect 1452 13268 1458 13280
rect 1489 13277 1501 13280
rect 1535 13277 1547 13311
rect 1489 13271 1547 13277
rect 1763 13311 1821 13317
rect 1763 13277 1775 13311
rect 1809 13308 1821 13311
rect 3712 13308 3740 13336
rect 1809 13280 3740 13308
rect 4338 13287 4344 13320
rect 4323 13281 4344 13287
rect 1809 13277 1821 13280
rect 1763 13271 1821 13277
rect 1504 13240 1532 13271
rect 1946 13240 1952 13252
rect 1504 13212 1952 13240
rect 1946 13200 1952 13212
rect 2004 13200 2010 13252
rect 2038 13200 2044 13252
rect 2096 13240 2102 13252
rect 2590 13240 2596 13252
rect 2096 13212 2596 13240
rect 2096 13200 2102 13212
rect 2590 13200 2596 13212
rect 2648 13200 2654 13252
rect 2682 13200 2688 13252
rect 2740 13240 2746 13252
rect 3694 13240 3700 13252
rect 2740 13212 3700 13240
rect 2740 13200 2746 13212
rect 3694 13200 3700 13212
rect 3752 13200 3758 13252
rect 4323 13247 4335 13281
rect 4396 13268 4402 13320
rect 5718 13268 5724 13320
rect 5776 13308 5782 13320
rect 5813 13311 5871 13317
rect 5813 13308 5825 13311
rect 5776 13280 5825 13308
rect 5776 13268 5782 13280
rect 5813 13277 5825 13280
rect 5859 13277 5871 13311
rect 5813 13271 5871 13277
rect 5997 13311 6055 13317
rect 5997 13277 6009 13311
rect 6043 13277 6055 13311
rect 5997 13271 6055 13277
rect 4369 13250 4382 13268
rect 4369 13247 4381 13250
rect 4323 13241 4381 13247
rect 5166 13200 5172 13252
rect 5224 13240 5230 13252
rect 6012 13240 6040 13271
rect 6730 13268 6736 13320
rect 6788 13268 6794 13320
rect 7024 13317 7052 13348
rect 7374 13336 7380 13348
rect 7432 13336 7438 13388
rect 7650 13336 7656 13388
rect 7708 13376 7714 13388
rect 7760 13376 7788 13484
rect 11882 13472 11888 13484
rect 11940 13472 11946 13524
rect 11977 13515 12035 13521
rect 11977 13481 11989 13515
rect 12023 13512 12035 13515
rect 12710 13512 12716 13524
rect 12023 13484 12716 13512
rect 12023 13481 12035 13484
rect 11977 13475 12035 13481
rect 12710 13472 12716 13484
rect 12768 13472 12774 13524
rect 13633 13515 13691 13521
rect 13633 13481 13645 13515
rect 13679 13512 13691 13515
rect 13998 13512 14004 13524
rect 13679 13484 14004 13512
rect 13679 13481 13691 13484
rect 13633 13475 13691 13481
rect 13998 13472 14004 13484
rect 14056 13472 14062 13524
rect 14366 13472 14372 13524
rect 14424 13512 14430 13524
rect 16022 13512 16028 13524
rect 14424 13484 16028 13512
rect 14424 13472 14430 13484
rect 16022 13472 16028 13484
rect 16080 13472 16086 13524
rect 16482 13472 16488 13524
rect 16540 13512 16546 13524
rect 17034 13512 17040 13524
rect 16540 13484 17040 13512
rect 16540 13472 16546 13484
rect 17034 13472 17040 13484
rect 17092 13472 17098 13524
rect 22189 13515 22247 13521
rect 22189 13481 22201 13515
rect 22235 13512 22247 13515
rect 22554 13512 22560 13524
rect 22235 13484 22560 13512
rect 22235 13481 22247 13484
rect 22189 13475 22247 13481
rect 22554 13472 22560 13484
rect 22612 13472 22618 13524
rect 24118 13472 24124 13524
rect 24176 13472 24182 13524
rect 16117 13447 16175 13453
rect 16117 13413 16129 13447
rect 16163 13444 16175 13447
rect 16206 13444 16212 13456
rect 16163 13416 16212 13444
rect 16163 13413 16175 13416
rect 16117 13407 16175 13413
rect 16206 13404 16212 13416
rect 16264 13404 16270 13456
rect 7708 13348 7788 13376
rect 7708 13336 7714 13348
rect 8662 13336 8668 13388
rect 8720 13376 8726 13388
rect 8941 13379 8999 13385
rect 8941 13376 8953 13379
rect 8720 13348 8953 13376
rect 8720 13336 8726 13348
rect 8941 13345 8953 13348
rect 8987 13345 8999 13379
rect 8941 13339 8999 13345
rect 10870 13336 10876 13388
rect 10928 13376 10934 13388
rect 10928 13348 11008 13376
rect 10928 13336 10934 13348
rect 7009 13311 7067 13317
rect 7009 13277 7021 13311
rect 7055 13277 7067 13311
rect 7009 13271 7067 13277
rect 9215 13311 9273 13317
rect 9215 13277 9227 13311
rect 9261 13308 9273 13311
rect 10226 13308 10232 13320
rect 9261 13280 10232 13308
rect 9261 13277 9273 13280
rect 9215 13271 9273 13277
rect 10226 13268 10232 13280
rect 10284 13268 10290 13320
rect 10502 13268 10508 13320
rect 10560 13268 10566 13320
rect 10980 13317 11008 13348
rect 11974 13336 11980 13388
rect 12032 13376 12038 13388
rect 12621 13379 12679 13385
rect 12621 13376 12633 13379
rect 12032 13348 12633 13376
rect 12032 13336 12038 13348
rect 12621 13345 12633 13348
rect 12667 13345 12679 13379
rect 12621 13339 12679 13345
rect 14458 13336 14464 13388
rect 14516 13376 14522 13388
rect 15657 13379 15715 13385
rect 15657 13376 15669 13379
rect 14516 13348 15669 13376
rect 14516 13336 14522 13348
rect 15657 13345 15669 13348
rect 15703 13345 15715 13379
rect 15657 13339 15715 13345
rect 10965 13311 11023 13317
rect 10965 13277 10977 13311
rect 11011 13277 11023 13311
rect 10965 13271 11023 13277
rect 11239 13311 11297 13317
rect 11239 13277 11251 13311
rect 11285 13308 11297 13311
rect 11698 13308 11704 13320
rect 11285 13280 11704 13308
rect 11285 13277 11297 13280
rect 11239 13271 11297 13277
rect 5224 13212 6040 13240
rect 5224 13200 5230 13212
rect 8570 13200 8576 13252
rect 8628 13240 8634 13252
rect 10980 13240 11008 13271
rect 11698 13268 11704 13280
rect 11756 13268 11762 13320
rect 11992 13240 12020 13336
rect 12895 13311 12953 13317
rect 12895 13277 12907 13311
rect 12941 13308 12953 13311
rect 14274 13308 14280 13320
rect 12941 13280 14280 13308
rect 12941 13277 12953 13280
rect 12895 13271 12953 13277
rect 14274 13268 14280 13280
rect 14332 13268 14338 13320
rect 15286 13268 15292 13320
rect 15344 13308 15350 13320
rect 15473 13311 15531 13317
rect 15473 13308 15485 13311
rect 15344 13280 15485 13308
rect 15344 13268 15350 13280
rect 15473 13277 15485 13280
rect 15519 13277 15531 13311
rect 15473 13271 15531 13277
rect 8628 13212 10088 13240
rect 10980 13212 12020 13240
rect 8628 13200 8634 13212
rect 2222 13132 2228 13184
rect 2280 13172 2286 13184
rect 6178 13172 6184 13184
rect 2280 13144 6184 13172
rect 2280 13132 2286 13144
rect 6178 13132 6184 13144
rect 6236 13132 6242 13184
rect 9950 13132 9956 13184
rect 10008 13132 10014 13184
rect 10060 13172 10088 13212
rect 12066 13200 12072 13252
rect 12124 13240 12130 13252
rect 13998 13240 14004 13252
rect 12124 13212 14004 13240
rect 12124 13200 12130 13212
rect 13998 13200 14004 13212
rect 14056 13200 14062 13252
rect 11606 13172 11612 13184
rect 10060 13144 11612 13172
rect 11606 13132 11612 13144
rect 11664 13132 11670 13184
rect 11974 13132 11980 13184
rect 12032 13172 12038 13184
rect 13354 13172 13360 13184
rect 12032 13144 13360 13172
rect 12032 13132 12038 13144
rect 13354 13132 13360 13144
rect 13412 13172 13418 13184
rect 14182 13172 14188 13184
rect 13412 13144 14188 13172
rect 13412 13132 13418 13144
rect 14182 13132 14188 13144
rect 14240 13132 14246 13184
rect 15672 13172 15700 13339
rect 16390 13336 16396 13388
rect 16448 13336 16454 13388
rect 16482 13336 16488 13388
rect 16540 13385 16546 13388
rect 16540 13379 16568 13385
rect 16556 13345 16568 13379
rect 16540 13339 16568 13345
rect 16669 13379 16727 13385
rect 16669 13345 16681 13379
rect 16715 13376 16727 13379
rect 17678 13376 17684 13388
rect 16715 13348 17684 13376
rect 16715 13345 16727 13348
rect 16669 13339 16727 13345
rect 16540 13336 16546 13339
rect 17678 13336 17684 13348
rect 17736 13336 17742 13388
rect 22002 13336 22008 13388
rect 22060 13336 22066 13388
rect 20809 13311 20867 13317
rect 20809 13277 20821 13311
rect 20855 13308 20867 13311
rect 22020 13308 22048 13336
rect 20855 13280 22048 13308
rect 22281 13311 22339 13317
rect 20855 13277 20867 13280
rect 20809 13271 20867 13277
rect 21192 13252 21220 13280
rect 22281 13277 22293 13311
rect 22327 13308 22339 13311
rect 22327 13280 22416 13308
rect 22554 13307 22560 13320
rect 22327 13277 22339 13280
rect 22281 13271 22339 13277
rect 22388 13252 22416 13280
rect 22523 13301 22560 13307
rect 22523 13267 22535 13301
rect 22612 13268 22618 13320
rect 23937 13311 23995 13317
rect 23937 13277 23949 13311
rect 23983 13277 23995 13311
rect 23937 13271 23995 13277
rect 22569 13267 22581 13268
rect 22523 13261 22581 13267
rect 21082 13249 21088 13252
rect 21076 13240 21088 13249
rect 21043 13212 21088 13240
rect 21076 13203 21088 13212
rect 21082 13200 21088 13203
rect 21140 13200 21146 13252
rect 21174 13200 21180 13252
rect 21232 13200 21238 13252
rect 22370 13200 22376 13252
rect 22428 13200 22434 13252
rect 22830 13200 22836 13252
rect 22888 13240 22894 13252
rect 23952 13240 23980 13271
rect 22888 13212 23980 13240
rect 22888 13200 22894 13212
rect 16390 13172 16396 13184
rect 15672 13144 16396 13172
rect 16390 13132 16396 13144
rect 16448 13132 16454 13184
rect 17310 13132 17316 13184
rect 17368 13132 17374 13184
rect 22278 13132 22284 13184
rect 22336 13172 22342 13184
rect 23293 13175 23351 13181
rect 23293 13172 23305 13175
rect 22336 13144 23305 13172
rect 22336 13132 22342 13144
rect 23293 13141 23305 13144
rect 23339 13141 23351 13175
rect 23293 13135 23351 13141
rect 1104 13082 24723 13104
rect 1104 13030 6814 13082
rect 6866 13030 6878 13082
rect 6930 13030 6942 13082
rect 6994 13030 7006 13082
rect 7058 13030 7070 13082
rect 7122 13030 12679 13082
rect 12731 13030 12743 13082
rect 12795 13030 12807 13082
rect 12859 13030 12871 13082
rect 12923 13030 12935 13082
rect 12987 13030 18544 13082
rect 18596 13030 18608 13082
rect 18660 13030 18672 13082
rect 18724 13030 18736 13082
rect 18788 13030 18800 13082
rect 18852 13030 24409 13082
rect 24461 13030 24473 13082
rect 24525 13030 24537 13082
rect 24589 13030 24601 13082
rect 24653 13030 24665 13082
rect 24717 13030 24723 13082
rect 1104 13008 24723 13030
rect 1210 12928 1216 12980
rect 1268 12968 1274 12980
rect 2317 12971 2375 12977
rect 2317 12968 2329 12971
rect 1268 12940 2329 12968
rect 1268 12928 1274 12940
rect 2317 12937 2329 12940
rect 2363 12937 2375 12971
rect 2317 12931 2375 12937
rect 3602 12928 3608 12980
rect 3660 12968 3666 12980
rect 4801 12971 4859 12977
rect 4801 12968 4813 12971
rect 3660 12940 4813 12968
rect 3660 12928 3666 12940
rect 4801 12937 4813 12940
rect 4847 12937 4859 12971
rect 4801 12931 4859 12937
rect 6178 12928 6184 12980
rect 6236 12968 6242 12980
rect 6730 12968 6736 12980
rect 6236 12940 6736 12968
rect 6236 12928 6242 12940
rect 6730 12928 6736 12940
rect 6788 12928 6794 12980
rect 7742 12928 7748 12980
rect 7800 12968 7806 12980
rect 7837 12971 7895 12977
rect 7837 12968 7849 12971
rect 7800 12940 7849 12968
rect 7800 12928 7806 12940
rect 7837 12937 7849 12940
rect 7883 12937 7895 12971
rect 17310 12968 17316 12980
rect 7837 12931 7895 12937
rect 8588 12940 17316 12968
rect 1673 12903 1731 12909
rect 1673 12869 1685 12903
rect 1719 12900 1731 12903
rect 2130 12900 2136 12912
rect 1719 12872 2136 12900
rect 1719 12869 1731 12872
rect 1673 12863 1731 12869
rect 2130 12860 2136 12872
rect 2188 12860 2194 12912
rect 2222 12860 2228 12912
rect 2280 12860 2286 12912
rect 4709 12903 4767 12909
rect 4709 12869 4721 12903
rect 4755 12900 4767 12903
rect 8588 12900 8616 12940
rect 17310 12928 17316 12940
rect 17368 12928 17374 12980
rect 18966 12928 18972 12980
rect 19024 12968 19030 12980
rect 19024 12940 20852 12968
rect 19024 12928 19030 12940
rect 4755 12872 8616 12900
rect 4755 12869 4767 12872
rect 4709 12863 4767 12869
rect 9490 12860 9496 12912
rect 9548 12860 9554 12912
rect 9769 12903 9827 12909
rect 9769 12869 9781 12903
rect 9815 12900 9827 12903
rect 10502 12900 10508 12912
rect 9815 12872 10508 12900
rect 9815 12869 9827 12872
rect 9769 12863 9827 12869
rect 10502 12860 10508 12872
rect 10560 12860 10566 12912
rect 10594 12860 10600 12912
rect 10652 12860 10658 12912
rect 11330 12860 11336 12912
rect 11388 12860 11394 12912
rect 11606 12860 11612 12912
rect 11664 12900 11670 12912
rect 19889 12903 19947 12909
rect 19889 12900 19901 12903
rect 11664 12872 19901 12900
rect 11664 12860 11670 12872
rect 19889 12869 19901 12872
rect 19935 12869 19947 12903
rect 20714 12900 20720 12912
rect 19889 12863 19947 12869
rect 19996 12872 20720 12900
rect 2406 12792 2412 12844
rect 2464 12792 2470 12844
rect 2682 12792 2688 12844
rect 2740 12792 2746 12844
rect 2866 12792 2872 12844
rect 2924 12792 2930 12844
rect 3694 12792 3700 12844
rect 3752 12841 3758 12844
rect 3752 12835 3780 12841
rect 3768 12801 3780 12835
rect 3752 12795 3780 12801
rect 3752 12792 3758 12795
rect 6362 12792 6368 12844
rect 6420 12832 6426 12844
rect 6730 12832 6736 12844
rect 6420 12804 6736 12832
rect 6420 12792 6426 12804
rect 6730 12792 6736 12804
rect 6788 12832 6794 12844
rect 6825 12835 6883 12841
rect 6825 12832 6837 12835
rect 6788 12804 6837 12832
rect 6788 12792 6794 12804
rect 6825 12801 6837 12804
rect 6871 12801 6883 12835
rect 6825 12795 6883 12801
rect 7099 12835 7157 12841
rect 7099 12801 7111 12835
rect 7145 12832 7157 12835
rect 7650 12832 7656 12844
rect 7145 12804 7656 12832
rect 7145 12801 7157 12804
rect 7099 12795 7157 12801
rect 7650 12792 7656 12804
rect 7708 12792 7714 12844
rect 9861 12835 9919 12841
rect 9861 12801 9873 12835
rect 9907 12832 9919 12835
rect 10134 12832 10140 12844
rect 9907 12804 10140 12832
rect 9907 12801 9919 12804
rect 9861 12795 9919 12801
rect 10134 12792 10140 12804
rect 10192 12792 10198 12844
rect 10229 12835 10287 12841
rect 10229 12801 10241 12835
rect 10275 12832 10287 12835
rect 11348 12832 11376 12860
rect 11759 12835 11817 12841
rect 11759 12832 11771 12835
rect 10275 12804 11376 12832
rect 11440 12804 11771 12832
rect 10275 12801 10287 12804
rect 10229 12795 10287 12801
rect 2424 12764 2452 12792
rect 3605 12767 3663 12773
rect 3605 12764 3617 12767
rect 2424 12736 3617 12764
rect 3605 12733 3617 12736
rect 3651 12733 3663 12767
rect 3605 12727 3663 12733
rect 3881 12767 3939 12773
rect 3881 12733 3893 12767
rect 3927 12764 3939 12767
rect 4430 12764 4436 12776
rect 3927 12736 4436 12764
rect 3927 12733 3939 12736
rect 3881 12727 3939 12733
rect 4430 12724 4436 12736
rect 4488 12724 4494 12776
rect 4522 12724 4528 12776
rect 4580 12764 4586 12776
rect 6270 12764 6276 12776
rect 4580 12736 6276 12764
rect 4580 12724 4586 12736
rect 6270 12724 6276 12736
rect 6328 12724 6334 12776
rect 9950 12724 9956 12776
rect 10008 12724 10014 12776
rect 10778 12724 10784 12776
rect 10836 12724 10842 12776
rect 11146 12724 11152 12776
rect 11204 12764 11210 12776
rect 11440 12764 11468 12804
rect 11759 12801 11771 12804
rect 11805 12801 11817 12835
rect 11759 12795 11817 12801
rect 11882 12792 11888 12844
rect 11940 12832 11946 12844
rect 14795 12835 14853 12841
rect 14795 12832 14807 12835
rect 11940 12804 14807 12832
rect 11940 12792 11946 12804
rect 14795 12801 14807 12804
rect 14841 12801 14853 12835
rect 14795 12795 14853 12801
rect 15930 12792 15936 12844
rect 15988 12832 15994 12844
rect 16114 12832 16120 12844
rect 15988 12804 16120 12832
rect 15988 12792 15994 12804
rect 16114 12792 16120 12804
rect 16172 12792 16178 12844
rect 17311 12835 17369 12841
rect 17311 12801 17323 12835
rect 17357 12832 17369 12835
rect 17402 12832 17408 12844
rect 17357 12804 17408 12832
rect 17357 12801 17369 12804
rect 17311 12795 17369 12801
rect 17402 12792 17408 12804
rect 17460 12792 17466 12844
rect 19610 12792 19616 12844
rect 19668 12792 19674 12844
rect 19996 12841 20024 12872
rect 20714 12860 20720 12872
rect 20772 12860 20778 12912
rect 19981 12835 20039 12841
rect 19981 12801 19993 12835
rect 20027 12801 20039 12835
rect 19981 12795 20039 12801
rect 20346 12792 20352 12844
rect 20404 12792 20410 12844
rect 20591 12835 20649 12841
rect 20591 12801 20603 12835
rect 20637 12832 20649 12835
rect 20824 12832 20852 12940
rect 21358 12928 21364 12980
rect 21416 12928 21422 12980
rect 22741 12971 22799 12977
rect 22741 12937 22753 12971
rect 22787 12968 22799 12971
rect 23290 12968 23296 12980
rect 22787 12940 23296 12968
rect 22787 12937 22799 12940
rect 22741 12931 22799 12937
rect 23290 12928 23296 12940
rect 23348 12928 23354 12980
rect 23385 12971 23443 12977
rect 23385 12937 23397 12971
rect 23431 12968 23443 12971
rect 24854 12968 24860 12980
rect 23431 12940 24860 12968
rect 23431 12937 23443 12940
rect 23385 12931 23443 12937
rect 24854 12928 24860 12940
rect 24912 12928 24918 12980
rect 20637 12804 20852 12832
rect 21376 12832 21404 12928
rect 21450 12860 21456 12912
rect 21508 12900 21514 12912
rect 23661 12903 23719 12909
rect 23661 12900 23673 12903
rect 21508 12872 23673 12900
rect 21508 12860 21514 12872
rect 23661 12869 23673 12872
rect 23707 12869 23719 12903
rect 23661 12863 23719 12869
rect 22005 12835 22063 12841
rect 22005 12832 22017 12835
rect 21376 12804 22017 12832
rect 20637 12801 20649 12804
rect 20591 12795 20649 12801
rect 22005 12801 22017 12804
rect 22051 12801 22063 12835
rect 22005 12795 22063 12801
rect 22186 12792 22192 12844
rect 22244 12792 22250 12844
rect 22278 12792 22284 12844
rect 22336 12832 22342 12844
rect 22465 12835 22523 12841
rect 22465 12832 22477 12835
rect 22336 12804 22477 12832
rect 22336 12792 22342 12804
rect 22465 12801 22477 12804
rect 22511 12801 22523 12835
rect 22465 12795 22523 12801
rect 22646 12792 22652 12844
rect 22704 12832 22710 12844
rect 22925 12835 22983 12841
rect 22925 12832 22937 12835
rect 22704 12804 22937 12832
rect 22704 12792 22710 12804
rect 22925 12801 22937 12804
rect 22971 12801 22983 12835
rect 22925 12795 22983 12801
rect 23201 12835 23259 12841
rect 23201 12801 23213 12835
rect 23247 12801 23259 12835
rect 23201 12795 23259 12801
rect 11204 12736 11468 12764
rect 11204 12724 11210 12736
rect 3326 12656 3332 12708
rect 3384 12656 3390 12708
rect 4338 12656 4344 12708
rect 4396 12656 4402 12708
rect 1394 12588 1400 12640
rect 1452 12628 1458 12640
rect 1765 12631 1823 12637
rect 1765 12628 1777 12631
rect 1452 12600 1777 12628
rect 1452 12588 1458 12600
rect 1765 12597 1777 12600
rect 1811 12597 1823 12631
rect 1765 12591 1823 12597
rect 2866 12588 2872 12640
rect 2924 12628 2930 12640
rect 4356 12628 4384 12656
rect 2924 12600 4384 12628
rect 2924 12588 2930 12600
rect 4522 12588 4528 12640
rect 4580 12588 4586 12640
rect 10796 12637 10824 12724
rect 10781 12631 10839 12637
rect 10781 12597 10793 12631
rect 10827 12597 10839 12631
rect 11440 12628 11468 12736
rect 11514 12724 11520 12776
rect 11572 12724 11578 12776
rect 12434 12724 12440 12776
rect 12492 12764 12498 12776
rect 12986 12764 12992 12776
rect 12492 12736 12992 12764
rect 12492 12724 12498 12736
rect 12986 12724 12992 12736
rect 13044 12724 13050 12776
rect 14274 12724 14280 12776
rect 14332 12764 14338 12776
rect 14553 12767 14611 12773
rect 14553 12764 14565 12767
rect 14332 12736 14565 12764
rect 14332 12724 14338 12736
rect 14553 12733 14565 12736
rect 14599 12733 14611 12767
rect 14553 12727 14611 12733
rect 17037 12767 17095 12773
rect 17037 12733 17049 12767
rect 17083 12733 17095 12767
rect 17037 12727 17095 12733
rect 19797 12767 19855 12773
rect 19797 12733 19809 12767
rect 19843 12764 19855 12767
rect 20254 12764 20260 12776
rect 19843 12736 20260 12764
rect 19843 12733 19855 12736
rect 19797 12727 19855 12733
rect 12406 12668 13584 12696
rect 12406 12628 12434 12668
rect 13556 12640 13584 12668
rect 17052 12640 17080 12727
rect 20254 12724 20260 12736
rect 20312 12724 20318 12776
rect 20364 12696 20392 12792
rect 22204 12764 22232 12792
rect 22741 12767 22799 12773
rect 22741 12764 22753 12767
rect 22204 12736 22753 12764
rect 22741 12733 22753 12736
rect 22787 12733 22799 12767
rect 22741 12727 22799 12733
rect 23216 12696 23244 12795
rect 17696 12668 20392 12696
rect 21284 12668 23244 12696
rect 11440 12600 12434 12628
rect 10781 12591 10839 12597
rect 12526 12588 12532 12640
rect 12584 12588 12590 12640
rect 13538 12588 13544 12640
rect 13596 12588 13602 12640
rect 13814 12588 13820 12640
rect 13872 12628 13878 12640
rect 14090 12628 14096 12640
rect 13872 12600 14096 12628
rect 13872 12588 13878 12600
rect 14090 12588 14096 12600
rect 14148 12588 14154 12640
rect 14826 12588 14832 12640
rect 14884 12628 14890 12640
rect 15565 12631 15623 12637
rect 15565 12628 15577 12631
rect 14884 12600 15577 12628
rect 14884 12588 14890 12600
rect 15565 12597 15577 12600
rect 15611 12597 15623 12631
rect 15565 12591 15623 12597
rect 17034 12588 17040 12640
rect 17092 12628 17098 12640
rect 17696 12628 17724 12668
rect 17092 12600 17724 12628
rect 17092 12588 17098 12600
rect 18046 12588 18052 12640
rect 18104 12588 18110 12640
rect 19150 12588 19156 12640
rect 19208 12628 19214 12640
rect 19794 12628 19800 12640
rect 19208 12600 19800 12628
rect 19208 12588 19214 12600
rect 19794 12588 19800 12600
rect 19852 12588 19858 12640
rect 20438 12588 20444 12640
rect 20496 12628 20502 12640
rect 21284 12628 21312 12668
rect 20496 12600 21312 12628
rect 20496 12588 20502 12600
rect 21358 12588 21364 12640
rect 21416 12588 21422 12640
rect 22097 12631 22155 12637
rect 22097 12597 22109 12631
rect 22143 12628 22155 12631
rect 22557 12631 22615 12637
rect 22557 12628 22569 12631
rect 22143 12600 22569 12628
rect 22143 12597 22155 12600
rect 22097 12591 22155 12597
rect 22557 12597 22569 12600
rect 22603 12597 22615 12631
rect 22557 12591 22615 12597
rect 22738 12588 22744 12640
rect 22796 12628 22802 12640
rect 23017 12631 23075 12637
rect 23017 12628 23029 12631
rect 22796 12600 23029 12628
rect 22796 12588 22802 12600
rect 23017 12597 23029 12600
rect 23063 12597 23075 12631
rect 23017 12591 23075 12597
rect 23934 12588 23940 12640
rect 23992 12588 23998 12640
rect 1104 12538 24564 12560
rect 1104 12486 3882 12538
rect 3934 12486 3946 12538
rect 3998 12486 4010 12538
rect 4062 12486 4074 12538
rect 4126 12486 4138 12538
rect 4190 12486 9747 12538
rect 9799 12486 9811 12538
rect 9863 12486 9875 12538
rect 9927 12486 9939 12538
rect 9991 12486 10003 12538
rect 10055 12486 15612 12538
rect 15664 12486 15676 12538
rect 15728 12486 15740 12538
rect 15792 12486 15804 12538
rect 15856 12486 15868 12538
rect 15920 12486 21477 12538
rect 21529 12486 21541 12538
rect 21593 12486 21605 12538
rect 21657 12486 21669 12538
rect 21721 12486 21733 12538
rect 21785 12486 24564 12538
rect 1104 12464 24564 12486
rect 1578 12384 1584 12436
rect 1636 12384 1642 12436
rect 3326 12384 3332 12436
rect 3384 12384 3390 12436
rect 3694 12384 3700 12436
rect 3752 12424 3758 12436
rect 4709 12427 4767 12433
rect 4709 12424 4721 12427
rect 3752 12396 4721 12424
rect 3752 12384 3758 12396
rect 4709 12393 4721 12396
rect 4755 12393 4767 12427
rect 4709 12387 4767 12393
rect 5166 12384 5172 12436
rect 5224 12424 5230 12436
rect 5224 12396 6776 12424
rect 5224 12384 5230 12396
rect 3786 12248 3792 12300
rect 3844 12248 3850 12300
rect 1486 12180 1492 12232
rect 1544 12180 1550 12232
rect 2317 12223 2375 12229
rect 2317 12189 2329 12223
rect 2363 12189 2375 12223
rect 2317 12183 2375 12189
rect 2332 12152 2360 12183
rect 2590 12180 2596 12232
rect 2648 12180 2654 12232
rect 3804 12152 3832 12248
rect 4706 12180 4712 12232
rect 4764 12220 4770 12232
rect 5258 12220 5264 12232
rect 4764 12192 5264 12220
rect 4764 12180 4770 12192
rect 5258 12180 5264 12192
rect 5316 12220 5322 12232
rect 5445 12223 5503 12229
rect 5445 12220 5457 12223
rect 5316 12192 5457 12220
rect 5316 12180 5322 12192
rect 5445 12189 5457 12192
rect 5491 12189 5503 12223
rect 5445 12183 5503 12189
rect 5703 12193 5761 12199
rect 2332 12124 3832 12152
rect 4065 12155 4123 12161
rect 4065 12121 4077 12155
rect 4111 12152 4123 12155
rect 4617 12155 4675 12161
rect 4111 12124 4568 12152
rect 4111 12121 4123 12124
rect 4065 12115 4123 12121
rect 3418 12044 3424 12096
rect 3476 12084 3482 12096
rect 4157 12087 4215 12093
rect 4157 12084 4169 12087
rect 3476 12056 4169 12084
rect 3476 12044 3482 12056
rect 4157 12053 4169 12056
rect 4203 12053 4215 12087
rect 4540 12084 4568 12124
rect 4617 12121 4629 12155
rect 4663 12152 4675 12155
rect 5703 12159 5715 12193
rect 5749 12190 5761 12193
rect 5749 12159 5764 12190
rect 5703 12153 5764 12159
rect 5736 12152 5764 12153
rect 4663 12124 5672 12152
rect 5736 12124 6684 12152
rect 4663 12121 4675 12124
rect 4617 12115 4675 12121
rect 5534 12084 5540 12096
rect 4540 12056 5540 12084
rect 4157 12047 4215 12053
rect 5534 12044 5540 12056
rect 5592 12044 5598 12096
rect 5644 12084 5672 12124
rect 6656 12096 6684 12124
rect 6362 12084 6368 12096
rect 5644 12056 6368 12084
rect 6362 12044 6368 12056
rect 6420 12044 6426 12096
rect 6454 12044 6460 12096
rect 6512 12044 6518 12096
rect 6638 12044 6644 12096
rect 6696 12044 6702 12096
rect 6748 12084 6776 12396
rect 10042 12384 10048 12436
rect 10100 12424 10106 12436
rect 10597 12427 10655 12433
rect 10597 12424 10609 12427
rect 10100 12396 10609 12424
rect 10100 12384 10106 12396
rect 10597 12393 10609 12396
rect 10643 12393 10655 12427
rect 10597 12387 10655 12393
rect 11882 12384 11888 12436
rect 11940 12424 11946 12436
rect 12158 12424 12164 12436
rect 11940 12396 12164 12424
rect 11940 12384 11946 12396
rect 12158 12384 12164 12396
rect 12216 12384 12222 12436
rect 12434 12384 12440 12436
rect 12492 12424 12498 12436
rect 13909 12427 13967 12433
rect 13909 12424 13921 12427
rect 12492 12396 13921 12424
rect 12492 12384 12498 12396
rect 13909 12393 13921 12396
rect 13955 12393 13967 12427
rect 13909 12387 13967 12393
rect 13998 12384 14004 12436
rect 14056 12424 14062 12436
rect 14182 12424 14188 12436
rect 14056 12396 14188 12424
rect 14056 12384 14062 12396
rect 14182 12384 14188 12396
rect 14240 12384 14246 12436
rect 18969 12427 19027 12433
rect 18969 12393 18981 12427
rect 19015 12424 19027 12427
rect 19610 12424 19616 12436
rect 19015 12396 19616 12424
rect 19015 12393 19027 12396
rect 18969 12387 19027 12393
rect 19610 12384 19616 12396
rect 19668 12384 19674 12436
rect 19702 12384 19708 12436
rect 19760 12424 19766 12436
rect 19760 12396 19930 12424
rect 19760 12384 19766 12396
rect 12342 12356 12348 12368
rect 12084 12328 12348 12356
rect 8662 12248 8668 12300
rect 8720 12288 8726 12300
rect 12084 12297 12112 12328
rect 12342 12316 12348 12328
rect 12400 12316 12406 12368
rect 12526 12316 12532 12368
rect 12584 12356 12590 12368
rect 12584 12316 12597 12356
rect 15562 12316 15568 12368
rect 15620 12356 15626 12368
rect 15930 12356 15936 12368
rect 15620 12328 15936 12356
rect 15620 12316 15626 12328
rect 15930 12316 15936 12328
rect 15988 12356 15994 12368
rect 17957 12359 18015 12365
rect 17957 12356 17969 12359
rect 15988 12328 17969 12356
rect 15988 12316 15994 12328
rect 17957 12325 17969 12328
rect 18003 12325 18015 12359
rect 17957 12319 18015 12325
rect 9585 12291 9643 12297
rect 9585 12288 9597 12291
rect 8720 12260 9597 12288
rect 8720 12248 8726 12260
rect 9585 12257 9597 12260
rect 9631 12257 9643 12291
rect 9585 12251 9643 12257
rect 12069 12291 12127 12297
rect 12069 12257 12081 12291
rect 12115 12257 12127 12291
rect 12069 12251 12127 12257
rect 12158 12248 12164 12300
rect 12216 12288 12222 12300
rect 12253 12291 12311 12297
rect 12253 12288 12265 12291
rect 12216 12260 12265 12288
rect 12216 12248 12222 12260
rect 12253 12257 12265 12260
rect 12299 12257 12311 12291
rect 12569 12288 12597 12316
rect 12713 12291 12771 12297
rect 12713 12288 12725 12291
rect 12569 12260 12725 12288
rect 12253 12251 12311 12257
rect 12713 12257 12725 12260
rect 12759 12257 12771 12291
rect 12713 12251 12771 12257
rect 12986 12248 12992 12300
rect 13044 12248 13050 12300
rect 14918 12248 14924 12300
rect 14976 12248 14982 12300
rect 15746 12248 15752 12300
rect 15804 12288 15810 12300
rect 15804 12260 18736 12288
rect 15804 12248 15810 12260
rect 9859 12223 9917 12229
rect 9859 12189 9871 12223
rect 9905 12220 9917 12223
rect 11238 12220 11244 12232
rect 9905 12192 11244 12220
rect 9905 12189 9917 12192
rect 9859 12183 9917 12189
rect 11238 12180 11244 12192
rect 11296 12180 11302 12232
rect 13078 12180 13084 12232
rect 13136 12229 13142 12232
rect 13136 12223 13164 12229
rect 13152 12189 13164 12223
rect 13136 12183 13164 12189
rect 13136 12180 13142 12183
rect 13262 12180 13268 12232
rect 13320 12180 13326 12232
rect 14734 12180 14740 12232
rect 14792 12180 14798 12232
rect 16298 12220 16304 12232
rect 15488 12214 16304 12220
rect 15470 12210 16304 12214
rect 15454 12192 16304 12210
rect 15454 12186 15516 12192
rect 15454 12182 15498 12186
rect 8754 12112 8760 12164
rect 8812 12152 8818 12164
rect 11974 12152 11980 12164
rect 8812 12124 11980 12152
rect 8812 12112 8818 12124
rect 11974 12112 11980 12124
rect 12032 12112 12038 12164
rect 13924 12124 14504 12152
rect 13924 12084 13952 12124
rect 6748 12056 13952 12084
rect 13998 12044 14004 12096
rect 14056 12084 14062 12096
rect 14366 12084 14372 12096
rect 14056 12056 14372 12084
rect 14056 12044 14062 12056
rect 14366 12044 14372 12056
rect 14424 12044 14430 12096
rect 14476 12084 14504 12124
rect 14550 12112 14556 12164
rect 14608 12152 14614 12164
rect 14645 12155 14703 12161
rect 14645 12152 14657 12155
rect 14608 12124 14657 12152
rect 14608 12112 14614 12124
rect 14645 12121 14657 12124
rect 14691 12121 14703 12155
rect 14645 12115 14703 12121
rect 15105 12155 15163 12161
rect 15105 12121 15117 12155
rect 15151 12152 15163 12155
rect 15454 12152 15482 12182
rect 16298 12180 16304 12192
rect 16356 12180 16362 12232
rect 17957 12223 18015 12229
rect 17957 12189 17969 12223
rect 18003 12220 18015 12223
rect 18046 12220 18052 12232
rect 18003 12192 18052 12220
rect 18003 12189 18015 12192
rect 17957 12183 18015 12189
rect 18046 12180 18052 12192
rect 18104 12180 18110 12232
rect 18138 12180 18144 12232
rect 18196 12220 18202 12232
rect 18417 12223 18475 12229
rect 18417 12220 18429 12223
rect 18196 12192 18429 12220
rect 18196 12180 18202 12192
rect 18417 12189 18429 12192
rect 18463 12189 18475 12223
rect 18417 12183 18475 12189
rect 18601 12223 18659 12229
rect 18601 12189 18613 12223
rect 18647 12189 18659 12223
rect 18601 12183 18659 12189
rect 15151 12124 15482 12152
rect 18325 12155 18383 12161
rect 15151 12121 15163 12124
rect 15105 12115 15163 12121
rect 18325 12121 18337 12155
rect 18371 12152 18383 12155
rect 18509 12155 18567 12161
rect 18509 12152 18521 12155
rect 18371 12124 18521 12152
rect 18371 12121 18383 12124
rect 18325 12115 18383 12121
rect 18509 12121 18521 12124
rect 18555 12121 18567 12155
rect 18509 12115 18567 12121
rect 15010 12084 15016 12096
rect 14476 12056 15016 12084
rect 15010 12044 15016 12056
rect 15068 12044 15074 12096
rect 15473 12087 15531 12093
rect 15473 12053 15485 12087
rect 15519 12084 15531 12087
rect 15562 12084 15568 12096
rect 15519 12056 15568 12084
rect 15519 12053 15531 12056
rect 15473 12047 15531 12053
rect 15562 12044 15568 12056
rect 15620 12044 15626 12096
rect 15654 12044 15660 12096
rect 15712 12044 15718 12096
rect 18138 12044 18144 12096
rect 18196 12084 18202 12096
rect 18616 12084 18644 12183
rect 18708 12152 18736 12260
rect 19150 12248 19156 12300
rect 19208 12288 19214 12300
rect 19245 12291 19303 12297
rect 19245 12288 19257 12291
rect 19208 12260 19257 12288
rect 19208 12248 19214 12260
rect 19245 12257 19257 12260
rect 19291 12257 19303 12291
rect 19245 12251 19303 12257
rect 18874 12180 18880 12232
rect 18932 12180 18938 12232
rect 19426 12210 19432 12232
rect 19352 12182 19432 12210
rect 19352 12152 19380 12182
rect 19426 12180 19432 12182
rect 19484 12180 19490 12232
rect 19534 12229 19656 12230
rect 19519 12223 19656 12229
rect 19519 12189 19531 12223
rect 19565 12222 19656 12223
rect 19565 12220 19840 12222
rect 19902 12220 19930 12396
rect 20254 12384 20260 12436
rect 20312 12384 20318 12436
rect 20714 12384 20720 12436
rect 20772 12384 20778 12436
rect 19565 12202 19930 12220
rect 19565 12189 19577 12202
rect 19628 12194 19930 12202
rect 19812 12192 19930 12194
rect 20272 12220 20300 12384
rect 23385 12359 23443 12365
rect 22066 12328 23244 12356
rect 21910 12248 21916 12300
rect 21968 12288 21974 12300
rect 22066 12288 22094 12328
rect 21968 12260 22094 12288
rect 21968 12248 21974 12260
rect 22186 12248 22192 12300
rect 22244 12248 22250 12300
rect 20625 12223 20683 12229
rect 20625 12220 20637 12223
rect 20272 12192 20637 12220
rect 19519 12183 19577 12189
rect 20625 12189 20637 12192
rect 20671 12189 20683 12223
rect 20625 12183 20683 12189
rect 20806 12180 20812 12232
rect 20864 12180 20870 12232
rect 21450 12180 21456 12232
rect 21508 12180 21514 12232
rect 21818 12180 21824 12232
rect 21876 12180 21882 12232
rect 22094 12180 22100 12232
rect 22152 12180 22158 12232
rect 23216 12229 23244 12328
rect 23385 12325 23397 12359
rect 23431 12356 23443 12359
rect 24854 12356 24860 12368
rect 23431 12328 24860 12356
rect 23431 12325 23443 12328
rect 23385 12319 23443 12325
rect 24854 12316 24860 12328
rect 24912 12316 24918 12368
rect 23201 12223 23259 12229
rect 23201 12189 23213 12223
rect 23247 12189 23259 12223
rect 23201 12183 23259 12189
rect 23474 12180 23480 12232
rect 23532 12220 23538 12232
rect 23661 12223 23719 12229
rect 23661 12220 23673 12223
rect 23532 12192 23673 12220
rect 23532 12180 23538 12192
rect 23661 12189 23673 12192
rect 23707 12189 23719 12223
rect 23661 12183 23719 12189
rect 18708 12124 19380 12152
rect 24026 12112 24032 12164
rect 24084 12112 24090 12164
rect 18196 12056 18644 12084
rect 18196 12044 18202 12056
rect 19150 12044 19156 12096
rect 19208 12084 19214 12096
rect 19426 12084 19432 12096
rect 19208 12056 19432 12084
rect 19208 12044 19214 12056
rect 19426 12044 19432 12056
rect 19484 12044 19490 12096
rect 1104 11994 24723 12016
rect 1104 11942 6814 11994
rect 6866 11942 6878 11994
rect 6930 11942 6942 11994
rect 6994 11942 7006 11994
rect 7058 11942 7070 11994
rect 7122 11942 12679 11994
rect 12731 11942 12743 11994
rect 12795 11942 12807 11994
rect 12859 11942 12871 11994
rect 12923 11942 12935 11994
rect 12987 11942 18544 11994
rect 18596 11942 18608 11994
rect 18660 11942 18672 11994
rect 18724 11942 18736 11994
rect 18788 11942 18800 11994
rect 18852 11942 24409 11994
rect 24461 11942 24473 11994
rect 24525 11942 24537 11994
rect 24589 11942 24601 11994
rect 24653 11942 24665 11994
rect 24717 11942 24723 11994
rect 1104 11920 24723 11942
rect 1854 11880 1860 11892
rect 1688 11852 1860 11880
rect 1688 11753 1716 11852
rect 1854 11840 1860 11852
rect 1912 11880 1918 11892
rect 1912 11852 3464 11880
rect 1912 11840 1918 11852
rect 3436 11812 3464 11852
rect 3510 11840 3516 11892
rect 3568 11880 3574 11892
rect 5626 11880 5632 11892
rect 3568 11852 5632 11880
rect 3568 11840 3574 11852
rect 5626 11840 5632 11852
rect 5684 11840 5690 11892
rect 6730 11880 6736 11892
rect 6380 11852 6736 11880
rect 3436 11784 3832 11812
rect 1673 11747 1731 11753
rect 1673 11713 1685 11747
rect 1719 11713 1731 11747
rect 1673 11707 1731 11713
rect 2406 11704 2412 11756
rect 2464 11704 2470 11756
rect 2498 11704 2504 11756
rect 2556 11753 2562 11756
rect 2556 11747 2584 11753
rect 2572 11713 2584 11747
rect 2556 11707 2584 11713
rect 2556 11704 2562 11707
rect 1486 11636 1492 11688
rect 1544 11676 1550 11688
rect 1854 11676 1860 11688
rect 1544 11648 1860 11676
rect 1544 11636 1550 11648
rect 1854 11636 1860 11648
rect 1912 11636 1918 11688
rect 2682 11636 2688 11688
rect 2740 11636 2746 11688
rect 3605 11679 3663 11685
rect 3605 11645 3617 11679
rect 3651 11676 3663 11679
rect 3694 11676 3700 11688
rect 3651 11648 3700 11676
rect 3651 11645 3663 11648
rect 3605 11639 3663 11645
rect 3694 11636 3700 11648
rect 3752 11636 3758 11688
rect 3804 11685 3832 11784
rect 4798 11704 4804 11756
rect 4856 11704 4862 11756
rect 6380 11753 6408 11852
rect 6730 11840 6736 11852
rect 6788 11880 6794 11892
rect 7098 11880 7104 11892
rect 6788 11852 7104 11880
rect 6788 11840 6794 11852
rect 7098 11840 7104 11852
rect 7156 11840 7162 11892
rect 7374 11840 7380 11892
rect 7432 11840 7438 11892
rect 7466 11840 7472 11892
rect 7524 11880 7530 11892
rect 9677 11883 9735 11889
rect 9677 11880 9689 11883
rect 7524 11852 9689 11880
rect 7524 11840 7530 11852
rect 9677 11849 9689 11852
rect 9723 11849 9735 11883
rect 9677 11843 9735 11849
rect 12084 11852 12296 11880
rect 6638 11783 6644 11824
rect 6623 11777 6644 11783
rect 6696 11812 6702 11824
rect 6822 11812 6828 11824
rect 6696 11784 6828 11812
rect 6365 11747 6423 11753
rect 6365 11713 6377 11747
rect 6411 11713 6423 11747
rect 6623 11743 6635 11777
rect 6696 11772 6702 11784
rect 6822 11772 6828 11784
rect 6880 11772 6886 11824
rect 6669 11746 6684 11772
rect 7837 11747 7895 11753
rect 6669 11743 6681 11746
rect 6623 11737 6681 11743
rect 6365 11707 6423 11713
rect 7837 11713 7849 11747
rect 7883 11744 7895 11747
rect 8202 11744 8208 11756
rect 7883 11716 8208 11744
rect 7883 11713 7895 11716
rect 7837 11707 7895 11713
rect 8202 11704 8208 11716
rect 8260 11704 8266 11756
rect 9030 11704 9036 11756
rect 9088 11704 9094 11756
rect 12084 11744 12112 11852
rect 12268 11812 12296 11852
rect 12434 11840 12440 11892
rect 12492 11880 12498 11892
rect 12710 11880 12716 11892
rect 12492 11852 12716 11880
rect 12492 11840 12498 11852
rect 12710 11840 12716 11852
rect 12768 11880 12774 11892
rect 12768 11852 13216 11880
rect 12768 11840 12774 11852
rect 13078 11812 13084 11824
rect 12268 11784 13084 11812
rect 13078 11772 13084 11784
rect 13136 11772 13142 11824
rect 13188 11812 13216 11852
rect 13262 11840 13268 11892
rect 13320 11880 13326 11892
rect 13449 11883 13507 11889
rect 13449 11880 13461 11883
rect 13320 11852 13461 11880
rect 13320 11840 13326 11852
rect 13449 11849 13461 11852
rect 13495 11849 13507 11883
rect 13449 11843 13507 11849
rect 14182 11840 14188 11892
rect 14240 11840 14246 11892
rect 14918 11840 14924 11892
rect 14976 11840 14982 11892
rect 15010 11840 15016 11892
rect 15068 11880 15074 11892
rect 15746 11880 15752 11892
rect 15068 11852 15752 11880
rect 15068 11840 15074 11852
rect 15746 11840 15752 11852
rect 15804 11840 15810 11892
rect 20625 11883 20683 11889
rect 17328 11852 19288 11880
rect 13906 11812 13912 11824
rect 13188 11784 13912 11812
rect 13906 11772 13912 11784
rect 13964 11772 13970 11824
rect 14200 11812 14228 11840
rect 14198 11784 14228 11812
rect 14198 11783 14226 11784
rect 14167 11777 14226 11783
rect 9600 11716 12112 11744
rect 9600 11688 9628 11716
rect 12618 11704 12624 11756
rect 12676 11744 12682 11756
rect 12711 11747 12769 11753
rect 12711 11744 12723 11747
rect 12676 11716 12723 11744
rect 12676 11704 12682 11716
rect 12711 11713 12723 11716
rect 12757 11744 12769 11747
rect 13538 11744 13544 11756
rect 12757 11716 13544 11744
rect 12757 11713 12769 11716
rect 12711 11707 12769 11713
rect 13538 11704 13544 11716
rect 13596 11704 13602 11756
rect 13814 11704 13820 11756
rect 13872 11744 13878 11756
rect 14167 11744 14179 11777
rect 13872 11743 14179 11744
rect 14213 11744 14226 11777
rect 16850 11744 16856 11756
rect 14213 11743 16856 11744
rect 13872 11716 16856 11743
rect 13872 11704 13878 11716
rect 16850 11704 16856 11716
rect 16908 11704 16914 11756
rect 17328 11753 17356 11852
rect 19260 11812 19288 11852
rect 20625 11849 20637 11883
rect 20671 11880 20683 11883
rect 20806 11880 20812 11892
rect 20671 11852 20812 11880
rect 20671 11849 20683 11852
rect 20625 11843 20683 11849
rect 20806 11840 20812 11852
rect 20864 11840 20870 11892
rect 22005 11883 22063 11889
rect 22005 11849 22017 11883
rect 22051 11880 22063 11883
rect 22094 11880 22100 11892
rect 22051 11852 22100 11880
rect 22051 11849 22063 11852
rect 22005 11843 22063 11849
rect 22094 11840 22100 11852
rect 22152 11840 22158 11892
rect 22278 11840 22284 11892
rect 22336 11880 22342 11892
rect 22646 11880 22652 11892
rect 22336 11852 22652 11880
rect 22336 11840 22342 11852
rect 22646 11840 22652 11852
rect 22704 11840 22710 11892
rect 24302 11812 24308 11824
rect 17420 11784 19196 11812
rect 19260 11784 24308 11812
rect 17420 11753 17448 11784
rect 17972 11756 18000 11784
rect 17313 11747 17371 11753
rect 17313 11713 17325 11747
rect 17359 11713 17371 11747
rect 17313 11707 17371 11713
rect 17405 11747 17463 11753
rect 17405 11713 17417 11747
rect 17451 11713 17463 11747
rect 17661 11747 17719 11753
rect 17661 11744 17673 11747
rect 17405 11707 17463 11713
rect 17512 11716 17673 11744
rect 3789 11679 3847 11685
rect 3789 11645 3801 11679
rect 3835 11676 3847 11679
rect 3835 11648 4384 11676
rect 3835 11645 3847 11648
rect 3789 11639 3847 11645
rect 2130 11568 2136 11620
rect 2188 11568 2194 11620
rect 4249 11611 4307 11617
rect 4249 11608 4261 11611
rect 3068 11580 4261 11608
rect 2774 11500 2780 11552
rect 2832 11540 2838 11552
rect 3068 11540 3096 11580
rect 4249 11577 4261 11580
rect 4295 11577 4307 11611
rect 4249 11571 4307 11577
rect 2832 11512 3096 11540
rect 2832 11500 2838 11512
rect 3326 11500 3332 11552
rect 3384 11500 3390 11552
rect 4356 11540 4384 11648
rect 4522 11636 4528 11688
rect 4580 11636 4586 11688
rect 4663 11679 4721 11685
rect 4663 11645 4675 11679
rect 4709 11676 4721 11679
rect 5718 11676 5724 11688
rect 4709 11648 5724 11676
rect 4709 11645 4721 11648
rect 4663 11639 4721 11645
rect 5718 11636 5724 11648
rect 5776 11636 5782 11688
rect 8021 11679 8079 11685
rect 8021 11676 8033 11679
rect 7944 11648 8033 11676
rect 7944 11552 7972 11648
rect 8021 11645 8033 11648
rect 8067 11645 8079 11679
rect 8757 11679 8815 11685
rect 8757 11676 8769 11679
rect 8021 11639 8079 11645
rect 8588 11648 8769 11676
rect 8478 11568 8484 11620
rect 8536 11568 8542 11620
rect 4614 11540 4620 11552
rect 4356 11512 4620 11540
rect 4614 11500 4620 11512
rect 4672 11540 4678 11552
rect 5166 11540 5172 11552
rect 4672 11512 5172 11540
rect 4672 11500 4678 11512
rect 5166 11500 5172 11512
rect 5224 11500 5230 11552
rect 5442 11500 5448 11552
rect 5500 11500 5506 11552
rect 7926 11500 7932 11552
rect 7984 11500 7990 11552
rect 8294 11500 8300 11552
rect 8352 11540 8358 11552
rect 8588 11540 8616 11648
rect 8757 11645 8769 11648
rect 8803 11645 8815 11679
rect 8757 11639 8815 11645
rect 8895 11679 8953 11685
rect 8895 11645 8907 11679
rect 8941 11676 8953 11679
rect 9582 11676 9588 11688
rect 8941 11648 9588 11676
rect 8941 11645 8953 11648
rect 8895 11639 8953 11645
rect 9582 11636 9588 11648
rect 9640 11636 9646 11688
rect 11514 11636 11520 11688
rect 11572 11676 11578 11688
rect 12437 11679 12495 11685
rect 12437 11676 12449 11679
rect 11572 11648 12449 11676
rect 11572 11636 11578 11648
rect 12437 11645 12449 11648
rect 12483 11645 12495 11679
rect 12437 11639 12495 11645
rect 13262 11636 13268 11688
rect 13320 11676 13326 11688
rect 13909 11679 13967 11685
rect 13909 11676 13921 11679
rect 13320 11648 13921 11676
rect 13320 11636 13326 11648
rect 13909 11645 13921 11648
rect 13955 11645 13967 11679
rect 17328 11676 17356 11707
rect 17512 11676 17540 11716
rect 17661 11713 17673 11716
rect 17707 11713 17719 11747
rect 17661 11707 17719 11713
rect 17954 11704 17960 11756
rect 18012 11704 18018 11756
rect 18138 11704 18144 11756
rect 18196 11744 18202 11756
rect 18196 11716 18736 11744
rect 18196 11704 18202 11716
rect 17328 11648 17540 11676
rect 18708 11676 18736 11716
rect 18782 11704 18788 11756
rect 18840 11744 18846 11756
rect 19168 11753 19196 11784
rect 24302 11772 24308 11784
rect 24360 11772 24366 11824
rect 19061 11747 19119 11753
rect 19061 11744 19073 11747
rect 18840 11716 19073 11744
rect 18840 11704 18846 11716
rect 19061 11713 19073 11716
rect 19107 11713 19119 11747
rect 19061 11707 19119 11713
rect 19153 11747 19211 11753
rect 19153 11713 19165 11747
rect 19199 11713 19211 11747
rect 19153 11707 19211 11713
rect 19420 11747 19478 11753
rect 19420 11713 19432 11747
rect 19466 11744 19478 11747
rect 19702 11744 19708 11756
rect 19466 11716 19708 11744
rect 19466 11713 19478 11716
rect 19420 11707 19478 11713
rect 19702 11704 19708 11716
rect 19760 11704 19766 11756
rect 20809 11747 20867 11753
rect 20809 11744 20821 11747
rect 20548 11716 20821 11744
rect 18708 11648 18920 11676
rect 13909 11639 13967 11645
rect 9416 11580 12572 11608
rect 9416 11540 9444 11580
rect 8352 11512 9444 11540
rect 8352 11500 8358 11512
rect 9490 11500 9496 11552
rect 9548 11540 9554 11552
rect 11974 11540 11980 11552
rect 9548 11512 11980 11540
rect 9548 11500 9554 11512
rect 11974 11500 11980 11512
rect 12032 11500 12038 11552
rect 12544 11540 12572 11580
rect 12894 11540 12900 11552
rect 12544 11512 12900 11540
rect 12894 11500 12900 11512
rect 12952 11500 12958 11552
rect 13924 11540 13952 11639
rect 14936 11580 17448 11608
rect 14936 11552 14964 11580
rect 14274 11540 14280 11552
rect 13924 11512 14280 11540
rect 14274 11500 14280 11512
rect 14332 11500 14338 11552
rect 14918 11500 14924 11552
rect 14976 11500 14982 11552
rect 17129 11543 17187 11549
rect 17129 11509 17141 11543
rect 17175 11540 17187 11543
rect 17310 11540 17316 11552
rect 17175 11512 17316 11540
rect 17175 11509 17187 11512
rect 17129 11503 17187 11509
rect 17310 11500 17316 11512
rect 17368 11500 17374 11552
rect 17420 11540 17448 11580
rect 18782 11568 18788 11620
rect 18840 11568 18846 11620
rect 18892 11617 18920 11648
rect 20548 11617 20576 11716
rect 20809 11713 20821 11716
rect 20855 11713 20867 11747
rect 20809 11707 20867 11713
rect 21450 11704 21456 11756
rect 21508 11744 21514 11756
rect 21821 11747 21879 11753
rect 21821 11744 21833 11747
rect 21508 11716 21833 11744
rect 21508 11704 21514 11716
rect 21821 11713 21833 11716
rect 21867 11713 21879 11747
rect 21821 11707 21879 11713
rect 22005 11745 22063 11751
rect 22005 11711 22017 11745
rect 22051 11711 22063 11745
rect 22005 11705 22063 11711
rect 22020 11676 22048 11705
rect 22370 11704 22376 11756
rect 22428 11704 22434 11756
rect 23075 11747 23133 11753
rect 23075 11744 23087 11747
rect 22572 11716 23087 11744
rect 22020 11648 22232 11676
rect 22204 11617 22232 11648
rect 18877 11611 18935 11617
rect 18877 11577 18889 11611
rect 18923 11577 18935 11611
rect 18877 11571 18935 11577
rect 20533 11611 20591 11617
rect 20533 11577 20545 11611
rect 20579 11577 20591 11611
rect 20533 11571 20591 11577
rect 22189 11611 22247 11617
rect 22189 11577 22201 11611
rect 22235 11577 22247 11611
rect 22189 11571 22247 11577
rect 21082 11540 21088 11552
rect 17420 11512 21088 11540
rect 21082 11500 21088 11512
rect 21140 11540 21146 11552
rect 22572 11540 22600 11716
rect 23075 11713 23087 11716
rect 23121 11713 23133 11747
rect 23075 11707 23133 11713
rect 22646 11636 22652 11688
rect 22704 11676 22710 11688
rect 22833 11679 22891 11685
rect 22833 11676 22845 11679
rect 22704 11648 22845 11676
rect 22704 11636 22710 11648
rect 22833 11645 22845 11648
rect 22879 11645 22891 11679
rect 22833 11639 22891 11645
rect 21140 11512 22600 11540
rect 21140 11500 21146 11512
rect 23842 11500 23848 11552
rect 23900 11500 23906 11552
rect 1104 11450 24564 11472
rect 1104 11398 3882 11450
rect 3934 11398 3946 11450
rect 3998 11398 4010 11450
rect 4062 11398 4074 11450
rect 4126 11398 4138 11450
rect 4190 11398 9747 11450
rect 9799 11398 9811 11450
rect 9863 11398 9875 11450
rect 9927 11398 9939 11450
rect 9991 11398 10003 11450
rect 10055 11398 15612 11450
rect 15664 11398 15676 11450
rect 15728 11398 15740 11450
rect 15792 11398 15804 11450
rect 15856 11398 15868 11450
rect 15920 11398 21477 11450
rect 21529 11398 21541 11450
rect 21593 11398 21605 11450
rect 21657 11398 21669 11450
rect 21721 11398 21733 11450
rect 21785 11398 24564 11450
rect 1104 11376 24564 11398
rect 1302 11296 1308 11348
rect 1360 11336 1366 11348
rect 1360 11308 2360 11336
rect 1360 11296 1366 11308
rect 2332 11268 2360 11308
rect 2682 11296 2688 11348
rect 2740 11296 2746 11348
rect 3329 11339 3387 11345
rect 3329 11305 3341 11339
rect 3375 11305 3387 11339
rect 3329 11299 3387 11305
rect 3344 11268 3372 11299
rect 3602 11296 3608 11348
rect 3660 11336 3666 11348
rect 4525 11339 4583 11345
rect 4525 11336 4537 11339
rect 3660 11308 4537 11336
rect 3660 11296 3666 11308
rect 4525 11305 4537 11308
rect 4571 11305 4583 11339
rect 4525 11299 4583 11305
rect 5534 11296 5540 11348
rect 5592 11336 5598 11348
rect 6917 11339 6975 11345
rect 6917 11336 6929 11339
rect 5592 11308 6929 11336
rect 5592 11296 5598 11308
rect 6917 11305 6929 11308
rect 6963 11305 6975 11339
rect 8294 11336 8300 11348
rect 6917 11299 6975 11305
rect 7024 11308 8300 11336
rect 2332 11240 3372 11268
rect 3528 11240 5856 11268
rect 2498 11160 2504 11212
rect 2556 11200 2562 11212
rect 3528 11200 3556 11240
rect 2556 11172 3556 11200
rect 2556 11160 2562 11172
rect 3602 11160 3608 11212
rect 3660 11200 3666 11212
rect 5442 11200 5448 11212
rect 3660 11172 4384 11200
rect 3660 11160 3666 11172
rect 1673 11135 1731 11141
rect 1673 11101 1685 11135
rect 1719 11101 1731 11135
rect 1673 11095 1731 11101
rect 1947 11135 2005 11141
rect 1947 11101 1959 11135
rect 1993 11132 2005 11135
rect 2314 11132 2320 11144
rect 1993 11104 2320 11132
rect 1993 11101 2005 11104
rect 1947 11095 2005 11101
rect 1688 11064 1716 11095
rect 2314 11092 2320 11104
rect 2372 11092 2378 11144
rect 3142 11092 3148 11144
rect 3200 11132 3206 11144
rect 3881 11135 3939 11141
rect 3881 11132 3893 11135
rect 3200 11104 3893 11132
rect 3200 11092 3206 11104
rect 3881 11101 3893 11104
rect 3927 11101 3939 11135
rect 3881 11095 3939 11101
rect 3237 11067 3295 11073
rect 1688 11036 1992 11064
rect 1964 11008 1992 11036
rect 3237 11033 3249 11067
rect 3283 11064 3295 11067
rect 4246 11064 4252 11076
rect 3283 11036 4252 11064
rect 3283 11033 3295 11036
rect 3237 11027 3295 11033
rect 4246 11024 4252 11036
rect 4304 11024 4310 11076
rect 4356 11064 4384 11172
rect 4448 11172 5448 11200
rect 4448 11141 4476 11172
rect 5442 11160 5448 11172
rect 5500 11160 5506 11212
rect 5718 11160 5724 11212
rect 5776 11160 5782 11212
rect 5828 11200 5856 11240
rect 5997 11203 6055 11209
rect 5997 11200 6009 11203
rect 5828 11172 6009 11200
rect 5997 11169 6009 11172
rect 6043 11169 6055 11203
rect 5997 11163 6055 11169
rect 6086 11160 6092 11212
rect 6144 11209 6150 11212
rect 6144 11203 6172 11209
rect 6160 11169 6172 11203
rect 6144 11163 6172 11169
rect 6273 11203 6331 11209
rect 6273 11169 6285 11203
rect 6319 11200 6331 11203
rect 6454 11200 6460 11212
rect 6319 11172 6460 11200
rect 6319 11169 6331 11172
rect 6273 11163 6331 11169
rect 6144 11160 6150 11163
rect 6454 11160 6460 11172
rect 6512 11160 6518 11212
rect 6638 11160 6644 11212
rect 6696 11200 6702 11212
rect 7024 11200 7052 11308
rect 8294 11296 8300 11308
rect 8352 11296 8358 11348
rect 8478 11296 8484 11348
rect 8536 11296 8542 11348
rect 9030 11296 9036 11348
rect 9088 11336 9094 11348
rect 9953 11339 10011 11345
rect 9953 11336 9965 11339
rect 9088 11308 9965 11336
rect 9088 11296 9094 11308
rect 9953 11305 9965 11308
rect 9999 11305 10011 11339
rect 9953 11299 10011 11305
rect 10686 11296 10692 11348
rect 10744 11336 10750 11348
rect 12253 11339 12311 11345
rect 12253 11336 12265 11339
rect 10744 11308 12265 11336
rect 10744 11296 10750 11308
rect 12253 11305 12265 11308
rect 12299 11305 12311 11339
rect 12253 11299 12311 11305
rect 12434 11296 12440 11348
rect 12492 11336 12498 11348
rect 14918 11336 14924 11348
rect 12492 11308 14924 11336
rect 12492 11296 12498 11308
rect 14918 11296 14924 11308
rect 14976 11296 14982 11348
rect 16298 11296 16304 11348
rect 16356 11296 16362 11348
rect 16850 11296 16856 11348
rect 16908 11336 16914 11348
rect 16908 11308 17264 11336
rect 16908 11296 16914 11308
rect 12066 11228 12072 11280
rect 12124 11268 12130 11280
rect 14550 11268 14556 11280
rect 12124 11240 14556 11268
rect 12124 11228 12130 11240
rect 14550 11228 14556 11240
rect 14608 11228 14614 11280
rect 14642 11228 14648 11280
rect 14700 11268 14706 11280
rect 16316 11268 16344 11296
rect 17236 11268 17264 11308
rect 18046 11296 18052 11348
rect 18104 11296 18110 11348
rect 18874 11296 18880 11348
rect 18932 11336 18938 11348
rect 19521 11339 19579 11345
rect 19521 11336 19533 11339
rect 18932 11308 19533 11336
rect 18932 11296 18938 11308
rect 19521 11305 19533 11308
rect 19567 11305 19579 11339
rect 19521 11299 19579 11305
rect 19904 11308 22131 11336
rect 19904 11268 19932 11308
rect 14700 11240 16436 11268
rect 17236 11240 19932 11268
rect 22103 11268 22131 11308
rect 22370 11296 22376 11348
rect 22428 11336 22434 11348
rect 22557 11339 22615 11345
rect 22557 11336 22569 11339
rect 22428 11308 22569 11336
rect 22428 11296 22434 11308
rect 22557 11305 22569 11308
rect 22603 11305 22615 11339
rect 22557 11299 22615 11305
rect 22103 11240 22600 11268
rect 14700 11228 14706 11240
rect 6696 11172 7052 11200
rect 6696 11160 6702 11172
rect 7098 11160 7104 11212
rect 7156 11200 7162 11212
rect 7469 11203 7527 11209
rect 7469 11200 7481 11203
rect 7156 11172 7481 11200
rect 7156 11160 7162 11172
rect 7469 11169 7481 11172
rect 7515 11169 7527 11203
rect 8941 11203 8999 11209
rect 8941 11200 8953 11203
rect 7469 11163 7527 11169
rect 8128 11172 8953 11200
rect 4433 11135 4491 11141
rect 4433 11101 4445 11135
rect 4479 11101 4491 11135
rect 4433 11095 4491 11101
rect 5077 11135 5135 11141
rect 5077 11101 5089 11135
rect 5123 11101 5135 11135
rect 5077 11095 5135 11101
rect 5092 11064 5120 11095
rect 5166 11092 5172 11144
rect 5224 11132 5230 11144
rect 5261 11135 5319 11141
rect 5261 11132 5273 11135
rect 5224 11104 5273 11132
rect 5224 11092 5230 11104
rect 5261 11101 5273 11104
rect 5307 11101 5319 11135
rect 5261 11095 5319 11101
rect 4356 11036 5120 11064
rect 7484 11064 7512 11163
rect 7743 11135 7801 11141
rect 7743 11101 7755 11135
rect 7789 11132 7801 11135
rect 7834 11132 7840 11144
rect 7789 11104 7840 11132
rect 7789 11101 7801 11104
rect 7743 11095 7801 11101
rect 7834 11092 7840 11104
rect 7892 11092 7898 11144
rect 8128 11132 8156 11172
rect 7944 11104 8156 11132
rect 7944 11064 7972 11104
rect 7484 11036 7972 11064
rect 8496 11064 8524 11172
rect 8941 11169 8953 11172
rect 8987 11169 8999 11203
rect 8941 11163 8999 11169
rect 10226 11160 10232 11212
rect 10284 11200 10290 11212
rect 10597 11203 10655 11209
rect 10597 11200 10609 11203
rect 10284 11172 10609 11200
rect 10284 11160 10290 11172
rect 10597 11169 10609 11172
rect 10643 11169 10655 11203
rect 10962 11200 10968 11212
rect 10597 11163 10655 11169
rect 10796 11172 10968 11200
rect 8570 11092 8576 11144
rect 8628 11132 8634 11144
rect 8754 11132 8760 11144
rect 8628 11104 8760 11132
rect 8628 11092 8634 11104
rect 8754 11092 8760 11104
rect 8812 11132 8818 11144
rect 9183 11135 9241 11141
rect 9183 11132 9195 11135
rect 8812 11104 9195 11132
rect 8812 11092 8818 11104
rect 9183 11101 9195 11104
rect 9229 11101 9241 11135
rect 9183 11095 9241 11101
rect 10134 11092 10140 11144
rect 10192 11132 10198 11144
rect 10413 11135 10471 11141
rect 10413 11132 10425 11135
rect 10192 11104 10425 11132
rect 10192 11092 10198 11104
rect 10413 11101 10425 11104
rect 10459 11132 10471 11135
rect 10796 11132 10824 11172
rect 10962 11160 10968 11172
rect 11020 11160 11026 11212
rect 11054 11160 11060 11212
rect 11112 11160 11118 11212
rect 11471 11203 11529 11209
rect 11471 11169 11483 11203
rect 11517 11200 11529 11203
rect 11517 11172 12204 11200
rect 11517 11169 11529 11172
rect 11471 11163 11529 11169
rect 10459 11104 10824 11132
rect 10459 11101 10471 11104
rect 10413 11095 10471 11101
rect 11330 11092 11336 11144
rect 11388 11092 11394 11144
rect 11606 11092 11612 11144
rect 11664 11092 11670 11144
rect 12176 11132 12204 11172
rect 14274 11160 14280 11212
rect 14332 11200 14338 11212
rect 15841 11203 15899 11209
rect 15841 11200 15853 11203
rect 14332 11172 15853 11200
rect 14332 11160 14338 11172
rect 15841 11169 15853 11172
rect 15887 11200 15899 11203
rect 15930 11200 15936 11212
rect 15887 11172 15936 11200
rect 15887 11169 15899 11172
rect 15841 11163 15899 11169
rect 15930 11160 15936 11172
rect 15988 11160 15994 11212
rect 16298 11160 16304 11212
rect 16356 11160 16362 11212
rect 16408 11200 16436 11240
rect 22572 11212 22600 11240
rect 16694 11203 16752 11209
rect 16694 11200 16706 11203
rect 16408 11172 16706 11200
rect 16694 11169 16706 11172
rect 16740 11169 16752 11203
rect 16694 11163 16752 11169
rect 17402 11160 17408 11212
rect 17460 11160 17466 11212
rect 19794 11200 19800 11212
rect 19628 11172 19800 11200
rect 12342 11132 12348 11144
rect 12176 11104 12348 11132
rect 12342 11092 12348 11104
rect 12400 11092 12406 11144
rect 12894 11092 12900 11144
rect 12952 11132 12958 11144
rect 15010 11132 15016 11144
rect 12952 11104 15016 11132
rect 12952 11092 12958 11104
rect 15010 11092 15016 11104
rect 15068 11092 15074 11144
rect 15657 11135 15715 11141
rect 15657 11101 15669 11135
rect 15703 11132 15715 11135
rect 15703 11104 15884 11132
rect 15703 11101 15715 11104
rect 15657 11095 15715 11101
rect 8496 11036 9674 11064
rect 1946 10956 1952 11008
rect 2004 10956 2010 11008
rect 3142 10956 3148 11008
rect 3200 10996 3206 11008
rect 3878 10996 3884 11008
rect 3200 10968 3884 10996
rect 3200 10956 3206 10968
rect 3878 10956 3884 10968
rect 3936 10956 3942 11008
rect 3970 10956 3976 11008
rect 4028 10956 4034 11008
rect 4338 10956 4344 11008
rect 4396 10996 4402 11008
rect 6086 10996 6092 11008
rect 4396 10968 6092 10996
rect 4396 10956 4402 10968
rect 6086 10956 6092 10968
rect 6144 10956 6150 11008
rect 9646 10996 9674 11036
rect 15856 11008 15884 11104
rect 16574 11092 16580 11144
rect 16632 11092 16638 11144
rect 16850 11092 16856 11144
rect 16908 11092 16914 11144
rect 17420 11132 17448 11160
rect 17957 11135 18015 11141
rect 17957 11132 17969 11135
rect 17420 11104 17969 11132
rect 17957 11101 17969 11104
rect 18003 11101 18015 11135
rect 17957 11095 18015 11101
rect 17402 11024 17408 11076
rect 17460 11064 17466 11076
rect 17497 11067 17555 11073
rect 17497 11064 17509 11067
rect 17460 11036 17509 11064
rect 17460 11024 17466 11036
rect 17497 11033 17509 11036
rect 17543 11033 17555 11067
rect 17497 11027 17555 11033
rect 18230 11024 18236 11076
rect 18288 11064 18294 11076
rect 18874 11064 18880 11076
rect 18288 11036 18880 11064
rect 18288 11024 18294 11036
rect 18874 11024 18880 11036
rect 18932 11024 18938 11076
rect 13262 10996 13268 11008
rect 9646 10968 13268 10996
rect 13262 10956 13268 10968
rect 13320 10956 13326 11008
rect 15838 10956 15844 11008
rect 15896 10956 15902 11008
rect 16942 10956 16948 11008
rect 17000 10996 17006 11008
rect 18046 10996 18052 11008
rect 17000 10968 18052 10996
rect 17000 10956 17006 10968
rect 18046 10956 18052 10968
rect 18104 10956 18110 11008
rect 19628 10996 19656 11172
rect 19794 11160 19800 11172
rect 19852 11160 19858 11212
rect 22554 11160 22560 11212
rect 22612 11160 22618 11212
rect 22738 11160 22744 11212
rect 22796 11160 22802 11212
rect 19702 11092 19708 11144
rect 19760 11092 19766 11144
rect 20070 11141 20076 11144
rect 20039 11135 20076 11141
rect 20039 11101 20051 11135
rect 20039 11095 20076 11101
rect 20070 11092 20076 11095
rect 20128 11092 20134 11144
rect 21177 11135 21235 11141
rect 21177 11101 21189 11135
rect 21223 11132 21235 11135
rect 21266 11132 21272 11144
rect 21223 11104 21272 11132
rect 21223 11101 21235 11104
rect 21177 11095 21235 11101
rect 21266 11092 21272 11104
rect 21324 11092 21330 11144
rect 22922 11092 22928 11144
rect 22980 11132 22986 11144
rect 23015 11135 23073 11141
rect 23015 11132 23027 11135
rect 22980 11104 23027 11132
rect 22980 11092 22986 11104
rect 23015 11101 23027 11104
rect 23061 11132 23073 11135
rect 23061 11104 23244 11132
rect 23061 11101 23073 11104
rect 23015 11095 23073 11101
rect 19720 11064 19748 11092
rect 23216 11076 23244 11104
rect 21444 11067 21502 11073
rect 19720 11036 21036 11064
rect 21008 11008 21036 11036
rect 21444 11033 21456 11067
rect 21490 11064 21502 11067
rect 22554 11064 22560 11076
rect 21490 11036 22560 11064
rect 21490 11033 21502 11036
rect 21444 11027 21502 11033
rect 22554 11024 22560 11036
rect 22612 11024 22618 11076
rect 23198 11024 23204 11076
rect 23256 11024 23262 11076
rect 20346 10996 20352 11008
rect 19628 10968 20352 10996
rect 20346 10956 20352 10968
rect 20404 10956 20410 11008
rect 20806 10956 20812 11008
rect 20864 10956 20870 11008
rect 20990 10956 20996 11008
rect 21048 10956 21054 11008
rect 22370 10956 22376 11008
rect 22428 10996 22434 11008
rect 23753 10999 23811 11005
rect 23753 10996 23765 10999
rect 22428 10968 23765 10996
rect 22428 10956 22434 10968
rect 23753 10965 23765 10968
rect 23799 10965 23811 10999
rect 23753 10959 23811 10965
rect 1104 10906 24723 10928
rect 1104 10854 6814 10906
rect 6866 10854 6878 10906
rect 6930 10854 6942 10906
rect 6994 10854 7006 10906
rect 7058 10854 7070 10906
rect 7122 10854 12679 10906
rect 12731 10854 12743 10906
rect 12795 10854 12807 10906
rect 12859 10854 12871 10906
rect 12923 10854 12935 10906
rect 12987 10854 18544 10906
rect 18596 10854 18608 10906
rect 18660 10854 18672 10906
rect 18724 10854 18736 10906
rect 18788 10854 18800 10906
rect 18852 10854 24409 10906
rect 24461 10854 24473 10906
rect 24525 10854 24537 10906
rect 24589 10854 24601 10906
rect 24653 10854 24665 10906
rect 24717 10854 24723 10906
rect 1104 10832 24723 10854
rect 658 10752 664 10804
rect 716 10792 722 10804
rect 1581 10795 1639 10801
rect 1581 10792 1593 10795
rect 716 10764 1593 10792
rect 716 10752 722 10764
rect 1581 10761 1593 10764
rect 1627 10761 1639 10795
rect 1581 10755 1639 10761
rect 2774 10752 2780 10804
rect 2832 10792 2838 10804
rect 2961 10795 3019 10801
rect 2961 10792 2973 10795
rect 2832 10764 2973 10792
rect 2832 10752 2838 10764
rect 2961 10761 2973 10764
rect 3007 10761 3019 10795
rect 4154 10792 4160 10804
rect 2961 10755 3019 10761
rect 3586 10764 4160 10792
rect 1964 10696 2360 10724
rect 1964 10665 1992 10696
rect 1489 10659 1547 10665
rect 1489 10625 1501 10659
rect 1535 10625 1547 10659
rect 1489 10619 1547 10625
rect 1949 10659 2007 10665
rect 1949 10625 1961 10659
rect 1995 10625 2007 10659
rect 2222 10656 2228 10668
rect 2183 10628 2228 10656
rect 1949 10619 2007 10625
rect 1504 10520 1532 10619
rect 2222 10616 2228 10628
rect 2280 10616 2286 10668
rect 2332 10656 2360 10696
rect 2406 10684 2412 10736
rect 2464 10724 2470 10736
rect 3586 10724 3614 10764
rect 4154 10752 4160 10764
rect 4212 10752 4218 10804
rect 4341 10795 4399 10801
rect 4341 10761 4353 10795
rect 4387 10792 4399 10795
rect 4798 10792 4804 10804
rect 4387 10764 4804 10792
rect 4387 10761 4399 10764
rect 4341 10755 4399 10761
rect 4798 10752 4804 10764
rect 4856 10752 4862 10804
rect 5718 10752 5724 10804
rect 5776 10752 5782 10804
rect 11054 10752 11060 10804
rect 11112 10752 11118 10804
rect 11606 10752 11612 10804
rect 11664 10792 11670 10804
rect 12529 10795 12587 10801
rect 12529 10792 12541 10795
rect 11664 10764 12541 10792
rect 11664 10752 11670 10764
rect 12529 10761 12541 10764
rect 12575 10761 12587 10795
rect 16209 10795 16267 10801
rect 12529 10755 12587 10761
rect 15120 10764 15608 10792
rect 2464 10696 3614 10724
rect 2464 10684 2470 10696
rect 3586 10695 3614 10696
rect 3586 10689 3645 10695
rect 3142 10656 3148 10668
rect 2332 10628 3148 10656
rect 3142 10616 3148 10628
rect 3200 10656 3206 10668
rect 3329 10659 3387 10665
rect 3329 10656 3341 10659
rect 3200 10628 3341 10656
rect 3200 10616 3206 10628
rect 3329 10625 3341 10628
rect 3375 10625 3387 10659
rect 3586 10658 3599 10689
rect 3587 10655 3599 10658
rect 3633 10655 3645 10689
rect 3878 10684 3884 10736
rect 3936 10724 3942 10736
rect 5258 10724 5264 10736
rect 3936 10696 5264 10724
rect 3936 10684 3942 10696
rect 4724 10665 4752 10696
rect 5258 10684 5264 10696
rect 5316 10724 5322 10736
rect 11514 10724 11520 10736
rect 5316 10684 5350 10724
rect 3587 10649 3645 10655
rect 4709 10659 4767 10665
rect 3329 10619 3387 10625
rect 4709 10625 4721 10659
rect 4755 10625 4767 10659
rect 4709 10619 4767 10625
rect 4890 10616 4896 10668
rect 4948 10656 4954 10668
rect 4983 10659 5041 10665
rect 4983 10656 4995 10659
rect 4948 10628 4995 10656
rect 4948 10616 4954 10628
rect 4983 10625 4995 10628
rect 5029 10625 5041 10659
rect 4983 10619 5041 10625
rect 5322 10588 5350 10684
rect 10060 10696 11520 10724
rect 7098 10616 7104 10668
rect 7156 10656 7162 10668
rect 7926 10656 7932 10668
rect 7156 10628 7932 10656
rect 7156 10616 7162 10628
rect 7926 10616 7932 10628
rect 7984 10616 7990 10668
rect 10060 10665 10088 10696
rect 10045 10659 10103 10665
rect 10045 10656 10057 10659
rect 9646 10628 10057 10656
rect 7374 10588 7380 10600
rect 5322 10560 7380 10588
rect 7374 10548 7380 10560
rect 7432 10588 7438 10600
rect 9646 10588 9674 10628
rect 10045 10625 10057 10628
rect 10091 10625 10103 10659
rect 10318 10656 10324 10668
rect 10279 10628 10324 10656
rect 10045 10619 10103 10625
rect 10318 10616 10324 10628
rect 10376 10656 10382 10668
rect 10962 10656 10968 10668
rect 10376 10628 10968 10656
rect 10376 10616 10382 10628
rect 10962 10616 10968 10628
rect 11020 10616 11026 10668
rect 7432 10560 9674 10588
rect 11164 10588 11192 10696
rect 11514 10684 11520 10696
rect 11572 10724 11578 10736
rect 13906 10724 13912 10736
rect 11572 10696 13912 10724
rect 11572 10684 11578 10696
rect 11238 10616 11244 10668
rect 11296 10656 11302 10668
rect 11759 10659 11817 10665
rect 11759 10656 11771 10659
rect 11296 10628 11771 10656
rect 11296 10616 11302 10628
rect 11759 10625 11771 10628
rect 11805 10656 11817 10659
rect 12158 10656 12164 10668
rect 11805 10628 12164 10656
rect 11805 10625 11817 10628
rect 11759 10619 11817 10625
rect 12158 10616 12164 10628
rect 12216 10616 12222 10668
rect 13464 10665 13492 10696
rect 13906 10684 13912 10696
rect 13964 10724 13970 10736
rect 15120 10724 15148 10764
rect 13964 10696 15148 10724
rect 13964 10684 13970 10696
rect 13449 10659 13507 10665
rect 13449 10625 13461 10659
rect 13495 10625 13507 10659
rect 13449 10619 13507 10625
rect 13723 10659 13781 10665
rect 13723 10625 13735 10659
rect 13769 10656 13781 10659
rect 13814 10656 13820 10668
rect 13769 10628 13820 10656
rect 13769 10625 13781 10628
rect 13723 10619 13781 10625
rect 13814 10616 13820 10628
rect 13872 10616 13878 10668
rect 11517 10591 11575 10597
rect 11517 10588 11529 10591
rect 11164 10560 11529 10588
rect 7432 10548 7438 10560
rect 11517 10557 11529 10560
rect 11563 10557 11575 10591
rect 15120 10588 15148 10696
rect 15194 10684 15200 10736
rect 15252 10724 15258 10736
rect 15580 10724 15608 10764
rect 16209 10761 16221 10795
rect 16255 10792 16267 10795
rect 16298 10792 16304 10804
rect 16255 10764 16304 10792
rect 16255 10761 16267 10764
rect 16209 10755 16267 10761
rect 16298 10752 16304 10764
rect 16356 10752 16362 10804
rect 16850 10752 16856 10804
rect 16908 10792 16914 10804
rect 17681 10795 17739 10801
rect 17681 10792 17693 10795
rect 16908 10764 17693 10792
rect 16908 10752 16914 10764
rect 17681 10761 17693 10764
rect 17727 10761 17739 10795
rect 17681 10755 17739 10761
rect 21818 10752 21824 10804
rect 21876 10792 21882 10804
rect 21913 10795 21971 10801
rect 21913 10792 21925 10795
rect 21876 10764 21925 10792
rect 21876 10752 21882 10764
rect 21913 10761 21925 10764
rect 21959 10761 21971 10795
rect 21913 10755 21971 10761
rect 23842 10752 23848 10804
rect 23900 10752 23906 10804
rect 18322 10724 18328 10736
rect 15252 10696 15482 10724
rect 15580 10696 18328 10724
rect 15252 10684 15258 10696
rect 15454 10665 15482 10696
rect 16684 10665 16712 10696
rect 18322 10684 18328 10696
rect 18380 10724 18386 10736
rect 22462 10724 22468 10736
rect 18380 10696 22468 10724
rect 18380 10684 18386 10696
rect 22462 10684 22468 10696
rect 22520 10684 22526 10736
rect 22738 10684 22744 10736
rect 22796 10684 22802 10736
rect 23106 10684 23112 10736
rect 23164 10684 23170 10736
rect 15439 10659 15497 10665
rect 15439 10625 15451 10659
rect 15485 10625 15497 10659
rect 15439 10619 15497 10625
rect 16669 10659 16727 10665
rect 16669 10625 16681 10659
rect 16715 10625 16727 10659
rect 16942 10656 16948 10668
rect 16903 10628 16948 10656
rect 16669 10619 16727 10625
rect 16942 10616 16948 10628
rect 17000 10616 17006 10668
rect 21821 10659 21879 10665
rect 21821 10625 21833 10659
rect 21867 10656 21879 10659
rect 22281 10659 22339 10665
rect 21867 10628 22140 10656
rect 21867 10625 21879 10628
rect 21821 10619 21879 10625
rect 15197 10591 15255 10597
rect 15197 10588 15209 10591
rect 15120 10560 15209 10588
rect 11517 10551 11575 10557
rect 15197 10557 15209 10560
rect 15243 10557 15255 10591
rect 15197 10551 15255 10557
rect 1504 10492 2084 10520
rect 2056 10452 2084 10492
rect 7006 10480 7012 10532
rect 7064 10520 7070 10532
rect 7466 10520 7472 10532
rect 7064 10492 7472 10520
rect 7064 10480 7070 10492
rect 7466 10480 7472 10492
rect 7524 10520 7530 10532
rect 7524 10492 8892 10520
rect 7524 10480 7530 10492
rect 8754 10452 8760 10464
rect 2056 10424 8760 10452
rect 8754 10412 8760 10424
rect 8812 10412 8818 10464
rect 8864 10452 8892 10492
rect 13262 10480 13268 10532
rect 13320 10520 13326 10532
rect 13446 10520 13452 10532
rect 13320 10492 13452 10520
rect 13320 10480 13326 10492
rect 13446 10480 13452 10492
rect 13504 10480 13510 10532
rect 14384 10492 14780 10520
rect 14384 10452 14412 10492
rect 14752 10464 14780 10492
rect 14918 10480 14924 10532
rect 14976 10480 14982 10532
rect 19426 10480 19432 10532
rect 19484 10520 19490 10532
rect 21818 10520 21824 10532
rect 19484 10492 21824 10520
rect 19484 10480 19490 10492
rect 21818 10480 21824 10492
rect 21876 10480 21882 10532
rect 22112 10529 22140 10628
rect 22281 10625 22293 10659
rect 22327 10656 22339 10659
rect 22554 10656 22560 10668
rect 22327 10628 22560 10656
rect 22327 10625 22339 10628
rect 22281 10619 22339 10625
rect 22554 10616 22560 10628
rect 22612 10616 22618 10668
rect 22649 10659 22707 10665
rect 22649 10625 22661 10659
rect 22695 10656 22707 10659
rect 22756 10656 22784 10684
rect 22695 10628 22784 10656
rect 22695 10625 22707 10628
rect 22649 10619 22707 10625
rect 22830 10616 22836 10668
rect 22888 10656 22894 10668
rect 22923 10659 22981 10665
rect 22923 10656 22935 10659
rect 22888 10628 22935 10656
rect 22888 10616 22894 10628
rect 22923 10625 22935 10628
rect 22969 10656 22981 10659
rect 23124 10656 23152 10684
rect 22969 10628 23152 10656
rect 23860 10656 23888 10752
rect 24213 10659 24271 10665
rect 24213 10656 24225 10659
rect 23860 10628 24225 10656
rect 22969 10625 22981 10628
rect 22923 10619 22981 10625
rect 24213 10625 24225 10628
rect 24259 10625 24271 10659
rect 24213 10619 24271 10625
rect 22097 10523 22155 10529
rect 22097 10489 22109 10523
rect 22143 10489 22155 10523
rect 22097 10483 22155 10489
rect 8864 10424 14412 10452
rect 14458 10412 14464 10464
rect 14516 10412 14522 10464
rect 14734 10412 14740 10464
rect 14792 10412 14798 10464
rect 14936 10452 14964 10480
rect 16942 10452 16948 10464
rect 14936 10424 16948 10452
rect 16942 10412 16948 10424
rect 17000 10412 17006 10464
rect 22646 10412 22652 10464
rect 22704 10452 22710 10464
rect 23661 10455 23719 10461
rect 23661 10452 23673 10455
rect 22704 10424 23673 10452
rect 22704 10412 22710 10424
rect 23661 10421 23673 10424
rect 23707 10421 23719 10455
rect 23661 10415 23719 10421
rect 24026 10412 24032 10464
rect 24084 10412 24090 10464
rect 1104 10362 24564 10384
rect 1104 10310 3882 10362
rect 3934 10310 3946 10362
rect 3998 10310 4010 10362
rect 4062 10310 4074 10362
rect 4126 10310 4138 10362
rect 4190 10310 9747 10362
rect 9799 10310 9811 10362
rect 9863 10310 9875 10362
rect 9927 10310 9939 10362
rect 9991 10310 10003 10362
rect 10055 10310 15612 10362
rect 15664 10310 15676 10362
rect 15728 10310 15740 10362
rect 15792 10310 15804 10362
rect 15856 10310 15868 10362
rect 15920 10310 21477 10362
rect 21529 10310 21541 10362
rect 21593 10310 21605 10362
rect 21657 10310 21669 10362
rect 21721 10310 21733 10362
rect 21785 10310 24564 10362
rect 1104 10288 24564 10310
rect 2130 10208 2136 10260
rect 2188 10248 2194 10260
rect 2409 10251 2467 10257
rect 2409 10248 2421 10251
rect 2188 10220 2421 10248
rect 2188 10208 2194 10220
rect 2409 10217 2421 10220
rect 2455 10217 2467 10251
rect 2409 10211 2467 10217
rect 2866 10208 2872 10260
rect 2924 10208 2930 10260
rect 2958 10208 2964 10260
rect 3016 10208 3022 10260
rect 3602 10208 3608 10260
rect 3660 10248 3666 10260
rect 5077 10251 5135 10257
rect 5077 10248 5089 10251
rect 3660 10220 5089 10248
rect 3660 10208 3666 10220
rect 5077 10217 5089 10220
rect 5123 10217 5135 10251
rect 5077 10211 5135 10217
rect 5629 10251 5687 10257
rect 5629 10217 5641 10251
rect 5675 10217 5687 10251
rect 8478 10248 8484 10260
rect 5629 10211 5687 10217
rect 7576 10220 8484 10248
rect 2884 10112 2912 10208
rect 3694 10140 3700 10192
rect 3752 10180 3758 10192
rect 5644 10180 5672 10211
rect 7576 10189 7604 10220
rect 8478 10208 8484 10220
rect 8536 10208 8542 10260
rect 8754 10208 8760 10260
rect 8812 10208 8818 10260
rect 9214 10208 9220 10260
rect 9272 10248 9278 10260
rect 11974 10248 11980 10260
rect 9272 10220 11980 10248
rect 9272 10208 9278 10220
rect 11974 10208 11980 10220
rect 12032 10208 12038 10260
rect 14458 10208 14464 10260
rect 14516 10248 14522 10260
rect 14516 10220 14688 10248
rect 14516 10208 14522 10220
rect 7561 10183 7619 10189
rect 3752 10152 5672 10180
rect 6472 10152 7512 10180
rect 3752 10140 3758 10152
rect 2332 10084 2912 10112
rect 4157 10115 4215 10121
rect 1397 10047 1455 10053
rect 1397 10013 1409 10047
rect 1443 10013 1455 10047
rect 1397 10007 1455 10013
rect 1671 10047 1729 10053
rect 1671 10013 1683 10047
rect 1717 10044 1729 10047
rect 2332 10044 2360 10084
rect 4157 10081 4169 10115
rect 4203 10112 4215 10115
rect 4338 10112 4344 10124
rect 4203 10084 4344 10112
rect 4203 10081 4215 10084
rect 4157 10075 4215 10081
rect 4338 10072 4344 10084
rect 4396 10072 4402 10124
rect 6472 10056 6500 10152
rect 6917 10115 6975 10121
rect 6917 10081 6929 10115
rect 6963 10112 6975 10115
rect 7006 10112 7012 10124
rect 6963 10084 7012 10112
rect 6963 10081 6975 10084
rect 6917 10075 6975 10081
rect 7006 10072 7012 10084
rect 7064 10072 7070 10124
rect 7098 10072 7104 10124
rect 7156 10072 7162 10124
rect 7484 10112 7512 10152
rect 7561 10149 7573 10183
rect 7607 10149 7619 10183
rect 7561 10143 7619 10149
rect 13449 10183 13507 10189
rect 13449 10149 13461 10183
rect 13495 10180 13507 10183
rect 14550 10180 14556 10192
rect 13495 10152 14556 10180
rect 13495 10149 13507 10152
rect 13449 10143 13507 10149
rect 14550 10140 14556 10152
rect 14608 10140 14614 10192
rect 7837 10115 7895 10121
rect 7837 10112 7849 10115
rect 7484 10084 7849 10112
rect 7837 10081 7849 10084
rect 7883 10081 7895 10115
rect 7837 10075 7895 10081
rect 8113 10115 8171 10121
rect 8113 10081 8125 10115
rect 8159 10112 8171 10115
rect 8294 10112 8300 10124
rect 8159 10084 8300 10112
rect 8159 10081 8171 10084
rect 8113 10075 8171 10081
rect 8294 10072 8300 10084
rect 8352 10072 8358 10124
rect 12434 10072 12440 10124
rect 12492 10072 12498 10124
rect 14274 10072 14280 10124
rect 14332 10072 14338 10124
rect 14660 10112 14688 10220
rect 14734 10208 14740 10260
rect 14792 10248 14798 10260
rect 22557 10251 22615 10257
rect 14792 10220 19334 10248
rect 14792 10208 14798 10220
rect 15746 10140 15752 10192
rect 15804 10180 15810 10192
rect 18693 10183 18751 10189
rect 18693 10180 18705 10183
rect 15804 10152 18705 10180
rect 15804 10140 15810 10152
rect 18693 10149 18705 10152
rect 18739 10149 18751 10183
rect 19306 10180 19334 10220
rect 22557 10217 22569 10251
rect 22603 10248 22615 10251
rect 24121 10251 24179 10257
rect 22603 10220 23118 10248
rect 22603 10217 22615 10220
rect 22557 10211 22615 10217
rect 20901 10183 20959 10189
rect 20901 10180 20913 10183
rect 19306 10152 20913 10180
rect 18693 10143 18751 10149
rect 20901 10149 20913 10152
rect 20947 10149 20959 10183
rect 20901 10143 20959 10149
rect 22281 10183 22339 10189
rect 22281 10149 22293 10183
rect 22327 10180 22339 10183
rect 22327 10152 23042 10180
rect 22327 10149 22339 10152
rect 22281 10143 22339 10149
rect 14737 10115 14795 10121
rect 14737 10112 14749 10115
rect 14660 10084 14749 10112
rect 14737 10081 14749 10084
rect 14783 10081 14795 10115
rect 14737 10075 14795 10081
rect 20806 10072 20812 10124
rect 20864 10072 20870 10124
rect 22370 10072 22376 10124
rect 22428 10112 22434 10124
rect 22428 10084 22508 10112
rect 22428 10072 22434 10084
rect 1717 10016 2360 10044
rect 1717 10013 1729 10016
rect 1671 10007 1729 10013
rect 1412 9976 1440 10007
rect 3234 10004 3240 10056
rect 3292 10044 3298 10056
rect 4433 10047 4491 10053
rect 4433 10044 4445 10047
rect 3292 10016 4445 10044
rect 3292 10004 3298 10016
rect 4433 10013 4445 10016
rect 4479 10013 4491 10047
rect 5537 10047 5595 10053
rect 4433 10007 4491 10013
rect 4908 10016 5488 10044
rect 1946 9976 1952 9988
rect 1412 9948 1952 9976
rect 1946 9936 1952 9948
rect 2004 9936 2010 9988
rect 2869 9979 2927 9985
rect 2869 9945 2881 9979
rect 2915 9945 2927 9979
rect 2869 9939 2927 9945
rect 2884 9908 2912 9939
rect 3786 9936 3792 9988
rect 3844 9976 3850 9988
rect 3881 9979 3939 9985
rect 3881 9976 3893 9979
rect 3844 9948 3893 9976
rect 3844 9936 3850 9948
rect 3881 9945 3893 9948
rect 3927 9945 3939 9979
rect 4908 9976 4936 10016
rect 3881 9939 3939 9945
rect 4080 9948 4936 9976
rect 4985 9979 5043 9985
rect 4080 9908 4108 9948
rect 4985 9945 4997 9979
rect 5031 9945 5043 9979
rect 5460 9976 5488 10016
rect 5537 10013 5549 10047
rect 5583 10044 5595 10047
rect 5626 10044 5632 10056
rect 5583 10016 5632 10044
rect 5583 10013 5595 10016
rect 5537 10007 5595 10013
rect 5626 10004 5632 10016
rect 5684 10004 5690 10056
rect 6454 10004 6460 10056
rect 6512 10004 6518 10056
rect 7282 10044 7288 10056
rect 7116 10016 7288 10044
rect 7116 9976 7144 10016
rect 7282 10004 7288 10016
rect 7340 10004 7346 10056
rect 8018 10053 8024 10056
rect 7975 10047 8024 10053
rect 7975 10013 7987 10047
rect 8021 10013 8024 10047
rect 7975 10007 8024 10013
rect 8018 10004 8024 10007
rect 8076 10004 8082 10056
rect 8754 10004 8760 10056
rect 8812 10044 8818 10056
rect 8941 10047 8999 10053
rect 8941 10044 8953 10047
rect 8812 10016 8953 10044
rect 8812 10004 8818 10016
rect 8941 10013 8953 10016
rect 8987 10013 8999 10047
rect 12618 10044 12624 10056
rect 9232 10023 12388 10044
rect 8941 10007 8999 10013
rect 9199 10017 12388 10023
rect 9199 9983 9211 10017
rect 9245 10016 12388 10017
rect 9245 9986 9260 10016
rect 9245 9983 9257 9986
rect 9199 9977 9257 9983
rect 10502 9976 10508 9988
rect 5460 9948 7144 9976
rect 9416 9948 10508 9976
rect 4985 9939 5043 9945
rect 2884 9880 4108 9908
rect 4154 9868 4160 9920
rect 4212 9908 4218 9920
rect 4525 9911 4583 9917
rect 4525 9908 4537 9911
rect 4212 9880 4537 9908
rect 4212 9868 4218 9880
rect 4525 9877 4537 9880
rect 4571 9877 4583 9911
rect 5000 9908 5028 9939
rect 9416 9908 9444 9948
rect 10502 9936 10508 9948
rect 10560 9936 10566 9988
rect 11882 9936 11888 9988
rect 11940 9976 11946 9988
rect 12066 9976 12072 9988
rect 11940 9948 12072 9976
rect 11940 9936 11946 9948
rect 12066 9936 12072 9948
rect 12124 9976 12130 9988
rect 12161 9979 12219 9985
rect 12161 9976 12173 9979
rect 12124 9948 12173 9976
rect 12124 9936 12130 9948
rect 12161 9945 12173 9948
rect 12207 9945 12219 9979
rect 12161 9939 12219 9945
rect 5000 9880 9444 9908
rect 4525 9871 4583 9877
rect 9490 9868 9496 9920
rect 9548 9908 9554 9920
rect 9953 9911 10011 9917
rect 9953 9908 9965 9911
rect 9548 9880 9965 9908
rect 9548 9868 9554 9880
rect 9953 9877 9965 9880
rect 9999 9877 10011 9911
rect 12360 9908 12388 10016
rect 12452 10016 12624 10044
rect 12452 9985 12480 10016
rect 12618 10004 12624 10016
rect 12676 10004 12682 10056
rect 12897 10047 12955 10053
rect 12897 10013 12909 10047
rect 12943 10044 12955 10047
rect 13354 10044 13360 10056
rect 12943 10016 13360 10044
rect 12943 10013 12955 10016
rect 12897 10007 12955 10013
rect 13354 10004 13360 10016
rect 13412 10004 13418 10056
rect 14093 10047 14151 10053
rect 14093 10013 14105 10047
rect 14139 10044 14151 10047
rect 14458 10044 14464 10056
rect 14139 10016 14464 10044
rect 14139 10013 14151 10016
rect 14093 10007 14151 10013
rect 14458 10004 14464 10016
rect 14516 10004 14522 10056
rect 15010 10004 15016 10056
rect 15068 10004 15074 10056
rect 15194 10053 15200 10056
rect 15151 10047 15200 10053
rect 15151 10013 15163 10047
rect 15197 10013 15200 10047
rect 15151 10007 15200 10013
rect 15194 10004 15200 10007
rect 15252 10004 15258 10056
rect 15286 10004 15292 10056
rect 15344 10004 15350 10056
rect 18049 10047 18107 10053
rect 18049 10013 18061 10047
rect 18095 10044 18107 10047
rect 18138 10044 18144 10056
rect 18095 10016 18144 10044
rect 18095 10013 18107 10016
rect 18049 10007 18107 10013
rect 18138 10004 18144 10016
rect 18196 10004 18202 10056
rect 18230 10004 18236 10056
rect 18288 10004 18294 10056
rect 18322 10004 18328 10056
rect 18380 10044 18386 10056
rect 18693 10047 18751 10053
rect 18693 10044 18705 10047
rect 18380 10016 18705 10044
rect 18380 10004 18386 10016
rect 18693 10013 18705 10016
rect 18739 10013 18751 10047
rect 18693 10007 18751 10013
rect 19797 10047 19855 10053
rect 19797 10013 19809 10047
rect 19843 10013 19855 10047
rect 19797 10007 19855 10013
rect 12437 9979 12495 9985
rect 12437 9945 12449 9979
rect 12483 9945 12495 9979
rect 12437 9939 12495 9945
rect 12526 9936 12532 9988
rect 12584 9936 12590 9988
rect 12636 9976 12664 10004
rect 13078 9976 13084 9988
rect 12636 9948 13084 9976
rect 13078 9936 13084 9948
rect 13136 9936 13142 9988
rect 14182 9976 14188 9988
rect 13188 9948 14188 9976
rect 13188 9908 13216 9948
rect 14182 9936 14188 9948
rect 14240 9936 14246 9988
rect 16482 9976 16488 9988
rect 15764 9948 16488 9976
rect 12360 9880 13216 9908
rect 9953 9871 10011 9877
rect 13262 9868 13268 9920
rect 13320 9917 13326 9920
rect 13320 9908 13327 9917
rect 13320 9880 13365 9908
rect 13320 9871 13327 9880
rect 13320 9868 13326 9871
rect 15010 9868 15016 9920
rect 15068 9908 15074 9920
rect 15764 9908 15792 9948
rect 16482 9936 16488 9948
rect 16540 9936 16546 9988
rect 19812 9920 19840 10007
rect 19978 10004 19984 10056
rect 20036 10004 20042 10056
rect 20898 10004 20904 10056
rect 20956 10004 20962 10056
rect 22480 10053 22508 10084
rect 22465 10047 22523 10053
rect 22465 10013 22477 10047
rect 22511 10013 22523 10047
rect 22465 10007 22523 10013
rect 22646 10004 22652 10056
rect 22704 10044 22710 10056
rect 22741 10047 22799 10053
rect 22741 10044 22753 10047
rect 22704 10016 22753 10044
rect 22704 10004 22710 10016
rect 22741 10013 22753 10016
rect 22787 10013 22799 10047
rect 22741 10007 22799 10013
rect 22833 10047 22891 10053
rect 22833 10013 22845 10047
rect 22879 10038 22891 10047
rect 23014 10038 23042 10152
rect 22879 10013 23042 10038
rect 22833 10010 23042 10013
rect 22833 10007 22891 10010
rect 21269 9979 21327 9985
rect 21269 9945 21281 9979
rect 21315 9976 21327 9979
rect 21542 9976 21548 9988
rect 21315 9948 21548 9976
rect 21315 9945 21327 9948
rect 21269 9939 21327 9945
rect 21542 9936 21548 9948
rect 21600 9936 21606 9988
rect 23090 9976 23118 10220
rect 24121 10217 24133 10251
rect 24167 10248 24179 10251
rect 24854 10248 24860 10260
rect 24167 10220 24860 10248
rect 24167 10217 24179 10220
rect 24121 10211 24179 10217
rect 24854 10208 24860 10220
rect 24912 10208 24918 10260
rect 23845 10047 23903 10053
rect 23845 10013 23857 10047
rect 23891 10044 23903 10047
rect 24026 10044 24032 10056
rect 23891 10016 24032 10044
rect 23891 10013 23903 10016
rect 23845 10007 23903 10013
rect 24026 10004 24032 10016
rect 24084 10004 24090 10056
rect 25130 10004 25136 10056
rect 25188 10004 25194 10056
rect 23293 9979 23351 9985
rect 23293 9976 23305 9979
rect 23090 9948 23305 9976
rect 23293 9945 23305 9948
rect 23339 9945 23351 9979
rect 23293 9939 23351 9945
rect 23661 9979 23719 9985
rect 23661 9945 23673 9979
rect 23707 9976 23719 9979
rect 24854 9976 24860 9988
rect 23707 9948 24860 9976
rect 23707 9945 23719 9948
rect 23661 9939 23719 9945
rect 24854 9936 24860 9948
rect 24912 9936 24918 9988
rect 15068 9880 15792 9908
rect 15068 9868 15074 9880
rect 15930 9868 15936 9920
rect 15988 9868 15994 9920
rect 17218 9868 17224 9920
rect 17276 9908 17282 9920
rect 18966 9908 18972 9920
rect 17276 9880 18972 9908
rect 17276 9868 17282 9880
rect 18966 9868 18972 9880
rect 19024 9868 19030 9920
rect 19794 9868 19800 9920
rect 19852 9868 19858 9920
rect 19981 9911 20039 9917
rect 19981 9877 19993 9911
rect 20027 9908 20039 9911
rect 20714 9908 20720 9920
rect 20027 9880 20720 9908
rect 20027 9877 20039 9880
rect 19981 9871 20039 9877
rect 20714 9868 20720 9880
rect 20772 9868 20778 9920
rect 23017 9911 23075 9917
rect 23017 9877 23029 9911
rect 23063 9908 23075 9911
rect 25148 9908 25176 10004
rect 23063 9880 25176 9908
rect 23063 9877 23075 9880
rect 23017 9871 23075 9877
rect 1104 9818 24723 9840
rect 1104 9766 6814 9818
rect 6866 9766 6878 9818
rect 6930 9766 6942 9818
rect 6994 9766 7006 9818
rect 7058 9766 7070 9818
rect 7122 9766 12679 9818
rect 12731 9766 12743 9818
rect 12795 9766 12807 9818
rect 12859 9766 12871 9818
rect 12923 9766 12935 9818
rect 12987 9766 18544 9818
rect 18596 9766 18608 9818
rect 18660 9766 18672 9818
rect 18724 9766 18736 9818
rect 18788 9766 18800 9818
rect 18852 9766 24409 9818
rect 24461 9766 24473 9818
rect 24525 9766 24537 9818
rect 24589 9766 24601 9818
rect 24653 9766 24665 9818
rect 24717 9766 24723 9818
rect 1104 9744 24723 9766
rect 1762 9664 1768 9716
rect 1820 9664 1826 9716
rect 2866 9664 2872 9716
rect 2924 9704 2930 9716
rect 3234 9704 3240 9716
rect 2924 9676 3240 9704
rect 2924 9664 2930 9676
rect 3234 9664 3240 9676
rect 3292 9704 3298 9716
rect 3510 9704 3516 9716
rect 3292 9676 3516 9704
rect 3292 9664 3298 9676
rect 3510 9664 3516 9676
rect 3568 9664 3574 9716
rect 4062 9664 4068 9716
rect 4120 9704 4126 9716
rect 5534 9704 5540 9716
rect 4120 9676 5540 9704
rect 4120 9664 4126 9676
rect 5534 9664 5540 9676
rect 5592 9664 5598 9716
rect 7374 9664 7380 9716
rect 7432 9664 7438 9716
rect 8018 9664 8024 9716
rect 8076 9704 8082 9716
rect 8202 9704 8208 9716
rect 8076 9676 8208 9704
rect 8076 9664 8082 9676
rect 8202 9664 8208 9676
rect 8260 9664 8266 9716
rect 8294 9664 8300 9716
rect 8352 9664 8358 9716
rect 10781 9707 10839 9713
rect 10781 9704 10793 9707
rect 8404 9676 10793 9704
rect 750 9596 756 9648
rect 808 9636 814 9648
rect 808 9608 2360 9636
rect 808 9596 814 9608
rect 1673 9571 1731 9577
rect 1673 9537 1685 9571
rect 1719 9568 1731 9571
rect 2130 9568 2136 9580
rect 1719 9540 2136 9568
rect 1719 9537 1731 9540
rect 1673 9531 1731 9537
rect 2130 9528 2136 9540
rect 2188 9528 2194 9580
rect 2332 9568 2360 9608
rect 5258 9596 5264 9648
rect 5316 9636 5322 9648
rect 6546 9636 6552 9648
rect 5316 9608 6552 9636
rect 5316 9596 5322 9608
rect 6546 9596 6552 9608
rect 6604 9596 6610 9648
rect 2593 9571 2651 9577
rect 2593 9568 2605 9571
rect 2332 9540 2605 9568
rect 2332 9512 2360 9540
rect 2593 9537 2605 9540
rect 2639 9537 2651 9571
rect 2593 9531 2651 9537
rect 3602 9528 3608 9580
rect 3660 9528 3666 9580
rect 4433 9571 4491 9577
rect 4433 9537 4445 9571
rect 4479 9568 4491 9571
rect 4522 9568 4528 9580
rect 4479 9540 4528 9568
rect 4479 9537 4491 9540
rect 4433 9531 4491 9537
rect 4522 9528 4528 9540
rect 4580 9528 4586 9580
rect 5167 9571 5225 9577
rect 5167 9537 5179 9571
rect 5213 9568 5225 9571
rect 7285 9571 7343 9577
rect 5213 9540 6868 9568
rect 5213 9537 5225 9540
rect 5167 9531 5225 9537
rect 2314 9460 2320 9512
rect 2372 9460 2378 9512
rect 2409 9503 2467 9509
rect 2409 9469 2421 9503
rect 2455 9469 2467 9503
rect 2409 9463 2467 9469
rect 2424 9432 2452 9463
rect 2774 9460 2780 9512
rect 2832 9500 2838 9512
rect 3510 9509 3516 9512
rect 3329 9503 3387 9509
rect 3329 9500 3341 9503
rect 2832 9472 3341 9500
rect 2832 9460 2838 9472
rect 3329 9469 3341 9472
rect 3375 9469 3387 9503
rect 3329 9463 3387 9469
rect 3467 9503 3516 9509
rect 3467 9469 3479 9503
rect 3513 9469 3516 9503
rect 3467 9463 3516 9469
rect 3510 9460 3516 9463
rect 3568 9500 3574 9512
rect 3568 9472 4474 9500
rect 3568 9460 3574 9472
rect 2866 9432 2872 9444
rect 2424 9404 2872 9432
rect 2866 9392 2872 9404
rect 2924 9392 2930 9444
rect 3050 9392 3056 9444
rect 3108 9392 3114 9444
rect 4249 9367 4307 9373
rect 4249 9333 4261 9367
rect 4295 9364 4307 9367
rect 4338 9364 4344 9376
rect 4295 9336 4344 9364
rect 4295 9333 4307 9336
rect 4249 9327 4307 9333
rect 4338 9324 4344 9336
rect 4396 9324 4402 9376
rect 4446 9364 4474 9472
rect 4890 9460 4896 9512
rect 4948 9460 4954 9512
rect 5626 9460 5632 9512
rect 5684 9500 5690 9512
rect 6730 9500 6736 9512
rect 5684 9472 6736 9500
rect 5684 9460 5690 9472
rect 6730 9460 6736 9472
rect 6788 9460 6794 9512
rect 4709 9435 4767 9441
rect 4709 9401 4721 9435
rect 4755 9432 4767 9435
rect 4798 9432 4804 9444
rect 4755 9404 4804 9432
rect 4755 9401 4767 9404
rect 4709 9395 4767 9401
rect 4798 9392 4804 9404
rect 4856 9392 4862 9444
rect 6178 9432 6184 9444
rect 5552 9404 6184 9432
rect 5552 9364 5580 9404
rect 6178 9392 6184 9404
rect 6236 9392 6242 9444
rect 4446 9336 5580 9364
rect 5902 9324 5908 9376
rect 5960 9324 5966 9376
rect 6840 9364 6868 9540
rect 7285 9537 7297 9571
rect 7331 9568 7343 9571
rect 7392 9568 7420 9664
rect 8220 9636 8248 9664
rect 8404 9636 8432 9676
rect 10781 9673 10793 9676
rect 10827 9673 10839 9707
rect 10781 9667 10839 9673
rect 12526 9664 12532 9716
rect 12584 9704 12590 9716
rect 13357 9707 13415 9713
rect 13357 9704 13369 9707
rect 12584 9676 13369 9704
rect 12584 9664 12590 9676
rect 13357 9673 13369 9676
rect 13403 9673 13415 9707
rect 13357 9667 13415 9673
rect 13998 9664 14004 9716
rect 14056 9704 14062 9716
rect 15010 9704 15016 9716
rect 14056 9676 15016 9704
rect 14056 9664 14062 9676
rect 15010 9664 15016 9676
rect 15068 9664 15074 9716
rect 15105 9707 15163 9713
rect 15105 9673 15117 9707
rect 15151 9704 15163 9707
rect 15286 9704 15292 9716
rect 15151 9676 15292 9704
rect 15151 9673 15163 9676
rect 15105 9667 15163 9673
rect 15286 9664 15292 9676
rect 15344 9664 15350 9716
rect 17862 9664 17868 9716
rect 17920 9704 17926 9716
rect 20622 9704 20628 9716
rect 17920 9676 20628 9704
rect 17920 9664 17926 9676
rect 20622 9664 20628 9676
rect 20680 9664 20686 9716
rect 20806 9664 20812 9716
rect 20864 9664 20870 9716
rect 20898 9664 20904 9716
rect 20956 9704 20962 9716
rect 21269 9707 21327 9713
rect 21269 9704 21281 9707
rect 20956 9676 21281 9704
rect 20956 9664 20962 9676
rect 21269 9673 21281 9676
rect 21315 9673 21327 9707
rect 21269 9667 21327 9673
rect 21542 9664 21548 9716
rect 21600 9664 21606 9716
rect 21818 9664 21824 9716
rect 21876 9704 21882 9716
rect 23934 9704 23940 9716
rect 21876 9676 23940 9704
rect 21876 9664 21882 9676
rect 23934 9664 23940 9676
rect 23992 9664 23998 9716
rect 8220 9608 8432 9636
rect 9214 9596 9220 9648
rect 9272 9636 9278 9648
rect 9398 9636 9404 9648
rect 9272 9608 9404 9636
rect 9272 9596 9278 9608
rect 9398 9596 9404 9608
rect 9456 9636 9462 9648
rect 9493 9639 9551 9645
rect 9493 9636 9505 9639
rect 9456 9608 9505 9636
rect 9456 9596 9462 9608
rect 9493 9605 9505 9608
rect 9539 9605 9551 9639
rect 9493 9599 9551 9605
rect 9861 9639 9919 9645
rect 9861 9605 9873 9639
rect 9907 9636 9919 9639
rect 10318 9636 10324 9648
rect 9907 9608 10324 9636
rect 9907 9605 9919 9608
rect 9861 9599 9919 9605
rect 10318 9596 10324 9608
rect 10376 9596 10382 9648
rect 10594 9596 10600 9648
rect 10652 9596 10658 9648
rect 14550 9636 14556 9648
rect 12820 9608 14556 9636
rect 7558 9568 7564 9580
rect 7331 9540 7420 9568
rect 7519 9540 7564 9568
rect 7331 9537 7343 9540
rect 7285 9531 7343 9537
rect 7558 9528 7564 9540
rect 7616 9528 7622 9580
rect 9769 9571 9827 9577
rect 9769 9537 9781 9571
rect 9815 9568 9827 9571
rect 10134 9568 10140 9580
rect 9815 9540 10140 9568
rect 9815 9537 9827 9540
rect 9769 9531 9827 9537
rect 10134 9528 10140 9540
rect 10192 9528 10198 9580
rect 10226 9528 10232 9580
rect 10284 9528 10290 9580
rect 12619 9571 12677 9577
rect 12619 9537 12631 9571
rect 12665 9568 12677 9571
rect 12820 9568 12848 9608
rect 14550 9596 14556 9608
rect 14608 9636 14614 9648
rect 16022 9636 16028 9648
rect 14608 9608 16028 9636
rect 14608 9596 14614 9608
rect 16022 9596 16028 9608
rect 16080 9596 16086 9648
rect 16482 9596 16488 9648
rect 16540 9596 16546 9648
rect 18046 9596 18052 9648
rect 18104 9636 18110 9648
rect 18104 9608 18828 9636
rect 18104 9596 18110 9608
rect 18800 9602 18828 9608
rect 18859 9602 18917 9607
rect 18800 9601 18917 9602
rect 12665 9540 12848 9568
rect 12665 9537 12677 9540
rect 12619 9531 12677 9537
rect 13906 9528 13912 9580
rect 13964 9568 13970 9580
rect 14093 9571 14151 9577
rect 14093 9568 14105 9571
rect 13964 9540 14105 9568
rect 13964 9528 13970 9540
rect 14093 9537 14105 9540
rect 14139 9537 14151 9571
rect 14093 9531 14151 9537
rect 14366 9528 14372 9580
rect 14424 9568 14430 9580
rect 15010 9568 15016 9580
rect 14424 9540 15016 9568
rect 14424 9528 14430 9540
rect 15010 9528 15016 9540
rect 15068 9528 15074 9580
rect 9496 9512 9548 9518
rect 11422 9460 11428 9512
rect 11480 9500 11486 9512
rect 12345 9503 12403 9509
rect 12345 9500 12357 9503
rect 11480 9472 12357 9500
rect 11480 9460 11486 9472
rect 12345 9469 12357 9472
rect 12391 9469 12403 9503
rect 12345 9463 12403 9469
rect 15102 9460 15108 9512
rect 15160 9500 15166 9512
rect 15378 9500 15384 9512
rect 15160 9472 15384 9500
rect 15160 9460 15166 9472
rect 15378 9460 15384 9472
rect 15436 9460 15442 9512
rect 15838 9460 15844 9512
rect 15896 9500 15902 9512
rect 16022 9500 16028 9512
rect 15896 9472 16028 9500
rect 15896 9460 15902 9472
rect 16022 9460 16028 9472
rect 16080 9460 16086 9512
rect 9496 9454 9548 9460
rect 16500 9376 16528 9596
rect 17310 9528 17316 9580
rect 17368 9528 17374 9580
rect 17678 9528 17684 9580
rect 17736 9568 17742 9580
rect 17954 9568 17960 9580
rect 17736 9540 17960 9568
rect 17736 9528 17742 9540
rect 17954 9528 17960 9540
rect 18012 9528 18018 9580
rect 18800 9574 18871 9601
rect 18859 9567 18871 9574
rect 18905 9567 18917 9601
rect 19150 9596 19156 9648
rect 19208 9636 19214 9648
rect 20824 9636 20852 9664
rect 19208 9608 19334 9636
rect 20824 9608 21496 9636
rect 19208 9596 19214 9608
rect 18859 9561 18917 9567
rect 19306 9568 19334 9608
rect 19426 9568 19432 9580
rect 19306 9540 19432 9568
rect 19426 9528 19432 9540
rect 19484 9528 19490 9580
rect 19610 9528 19616 9580
rect 19668 9568 19674 9580
rect 20349 9571 20407 9577
rect 20349 9568 20361 9571
rect 19668 9540 20361 9568
rect 19668 9528 19674 9540
rect 20349 9537 20361 9540
rect 20395 9537 20407 9571
rect 20349 9531 20407 9537
rect 20714 9528 20720 9580
rect 20772 9568 20778 9580
rect 20809 9571 20867 9577
rect 20809 9568 20821 9571
rect 20772 9540 20821 9568
rect 20772 9528 20778 9540
rect 20809 9537 20821 9540
rect 20855 9537 20867 9571
rect 20809 9531 20867 9537
rect 21174 9528 21180 9580
rect 21232 9528 21238 9580
rect 21468 9577 21496 9608
rect 21453 9571 21511 9577
rect 21453 9537 21465 9571
rect 21499 9537 21511 9571
rect 21453 9531 21511 9537
rect 21637 9571 21695 9577
rect 21637 9537 21649 9571
rect 21683 9568 21695 9571
rect 21683 9540 21864 9568
rect 21683 9537 21695 9540
rect 21637 9531 21695 9537
rect 16850 9460 16856 9512
rect 16908 9500 16914 9512
rect 17037 9503 17095 9509
rect 17037 9500 17049 9503
rect 16908 9472 17049 9500
rect 16908 9460 16914 9472
rect 17037 9469 17049 9472
rect 17083 9469 17095 9503
rect 18598 9500 18604 9512
rect 17037 9463 17095 9469
rect 17880 9472 18604 9500
rect 7650 9364 7656 9376
rect 6840 9336 7656 9364
rect 7650 9324 7656 9336
rect 7708 9324 7714 9376
rect 10686 9324 10692 9376
rect 10744 9364 10750 9376
rect 14918 9364 14924 9376
rect 10744 9336 14924 9364
rect 10744 9324 10750 9336
rect 14918 9324 14924 9336
rect 14976 9324 14982 9376
rect 16482 9324 16488 9376
rect 16540 9324 16546 9376
rect 17052 9364 17080 9463
rect 17402 9364 17408 9376
rect 17052 9336 17408 9364
rect 17402 9324 17408 9336
rect 17460 9364 17466 9376
rect 17880 9364 17908 9472
rect 18598 9460 18604 9472
rect 18656 9460 18662 9512
rect 19794 9500 19800 9512
rect 19628 9472 19800 9500
rect 19628 9441 19656 9472
rect 19794 9460 19800 9472
rect 19852 9500 19858 9512
rect 20073 9503 20131 9509
rect 20073 9500 20085 9503
rect 19852 9472 20085 9500
rect 19852 9460 19858 9472
rect 20073 9469 20085 9472
rect 20119 9469 20131 9503
rect 20073 9463 20131 9469
rect 20254 9460 20260 9512
rect 20312 9500 20318 9512
rect 20312 9472 20944 9500
rect 20312 9460 20318 9472
rect 19613 9435 19671 9441
rect 19613 9401 19625 9435
rect 19659 9401 19671 9435
rect 19613 9395 19671 9401
rect 20809 9435 20867 9441
rect 20809 9401 20821 9435
rect 20855 9401 20867 9435
rect 20809 9395 20867 9401
rect 17460 9336 17908 9364
rect 18049 9367 18107 9373
rect 17460 9324 17466 9336
rect 18049 9333 18061 9367
rect 18095 9364 18107 9367
rect 18138 9364 18144 9376
rect 18095 9336 18144 9364
rect 18095 9333 18107 9336
rect 18049 9327 18107 9333
rect 18138 9324 18144 9336
rect 18196 9324 18202 9376
rect 18506 9324 18512 9376
rect 18564 9364 18570 9376
rect 20824 9364 20852 9395
rect 18564 9336 20852 9364
rect 20916 9364 20944 9472
rect 21836 9441 21864 9540
rect 22002 9528 22008 9580
rect 22060 9528 22066 9580
rect 23075 9571 23133 9577
rect 23075 9568 23087 9571
rect 22572 9540 23087 9568
rect 21821 9435 21879 9441
rect 21821 9401 21833 9435
rect 21867 9401 21879 9435
rect 21821 9395 21879 9401
rect 22572 9364 22600 9540
rect 23075 9537 23087 9540
rect 23121 9537 23133 9571
rect 23075 9531 23133 9537
rect 22738 9460 22744 9512
rect 22796 9500 22802 9512
rect 22833 9503 22891 9509
rect 22833 9500 22845 9503
rect 22796 9472 22845 9500
rect 22796 9460 22802 9472
rect 22833 9469 22845 9472
rect 22879 9469 22891 9503
rect 22833 9463 22891 9469
rect 20916 9336 22600 9364
rect 18564 9324 18570 9336
rect 23842 9324 23848 9376
rect 23900 9324 23906 9376
rect 1104 9274 24564 9296
rect 1104 9222 3882 9274
rect 3934 9222 3946 9274
rect 3998 9222 4010 9274
rect 4062 9222 4074 9274
rect 4126 9222 4138 9274
rect 4190 9222 9747 9274
rect 9799 9222 9811 9274
rect 9863 9222 9875 9274
rect 9927 9222 9939 9274
rect 9991 9222 10003 9274
rect 10055 9222 15612 9274
rect 15664 9222 15676 9274
rect 15728 9222 15740 9274
rect 15792 9222 15804 9274
rect 15856 9222 15868 9274
rect 15920 9222 21477 9274
rect 21529 9222 21541 9274
rect 21593 9222 21605 9274
rect 21657 9222 21669 9274
rect 21721 9222 21733 9274
rect 21785 9222 24564 9274
rect 1104 9200 24564 9222
rect 2869 9163 2927 9169
rect 2869 9129 2881 9163
rect 2915 9160 2927 9163
rect 3050 9160 3056 9172
rect 2915 9132 3056 9160
rect 2915 9129 2927 9132
rect 2869 9123 2927 9129
rect 3050 9120 3056 9132
rect 3108 9120 3114 9172
rect 3786 9120 3792 9172
rect 3844 9160 3850 9172
rect 3844 9132 5856 9160
rect 3844 9120 3850 9132
rect 4890 9052 4896 9104
rect 4948 9092 4954 9104
rect 5718 9092 5724 9104
rect 4948 9064 5724 9092
rect 4948 9052 4954 9064
rect 5718 9052 5724 9064
rect 5776 9052 5782 9104
rect 5626 8984 5632 9036
rect 5684 8984 5690 9036
rect 5828 9024 5856 9132
rect 5902 9120 5908 9172
rect 5960 9120 5966 9172
rect 6086 9120 6092 9172
rect 6144 9160 6150 9172
rect 6144 9132 8432 9160
rect 6144 9120 6150 9132
rect 5920 9092 5948 9120
rect 6181 9095 6239 9101
rect 6181 9092 6193 9095
rect 5920 9064 6193 9092
rect 6181 9061 6193 9064
rect 6227 9061 6239 9095
rect 8404 9092 8432 9132
rect 8478 9120 8484 9172
rect 8536 9120 8542 9172
rect 10042 9160 10048 9172
rect 9646 9132 10048 9160
rect 9646 9092 9674 9132
rect 10042 9120 10048 9132
rect 10100 9120 10106 9172
rect 10318 9120 10324 9172
rect 10376 9160 10382 9172
rect 10597 9163 10655 9169
rect 10597 9160 10609 9163
rect 10376 9132 10609 9160
rect 10376 9120 10382 9132
rect 10597 9129 10609 9132
rect 10643 9129 10655 9163
rect 10597 9123 10655 9129
rect 11532 9132 12112 9160
rect 8404 9064 9674 9092
rect 6181 9055 6239 9061
rect 8496 9036 8524 9064
rect 10502 9052 10508 9104
rect 10560 9092 10566 9104
rect 11532 9092 11560 9132
rect 10560 9064 11560 9092
rect 12084 9092 12112 9132
rect 12434 9120 12440 9172
rect 12492 9120 12498 9172
rect 14936 9132 17540 9160
rect 14936 9092 14964 9132
rect 12084 9064 14964 9092
rect 10560 9052 10566 9064
rect 15102 9052 15108 9104
rect 15160 9092 15166 9104
rect 16206 9092 16212 9104
rect 15160 9064 16212 9092
rect 15160 9052 15166 9064
rect 7377 9027 7435 9033
rect 7377 9024 7389 9027
rect 5828 8996 7389 9024
rect 7377 8993 7389 8996
rect 7423 8993 7435 9027
rect 7377 8987 7435 8993
rect 8478 8984 8484 9036
rect 8536 8984 8542 9036
rect 11422 8984 11428 9036
rect 11480 8984 11486 9036
rect 15856 9033 15884 9064
rect 16206 9052 16212 9064
rect 16264 9052 16270 9104
rect 17512 9101 17540 9132
rect 17586 9120 17592 9172
rect 17644 9160 17650 9172
rect 20254 9160 20260 9172
rect 17644 9132 20260 9160
rect 17644 9120 17650 9132
rect 20254 9120 20260 9132
rect 20312 9120 20318 9172
rect 20530 9120 20536 9172
rect 20588 9160 20594 9172
rect 20588 9132 21680 9160
rect 20588 9120 20594 9132
rect 17497 9095 17555 9101
rect 17497 9061 17509 9095
rect 17543 9061 17555 9095
rect 17497 9055 17555 9061
rect 18598 9052 18604 9104
rect 18656 9092 18662 9104
rect 19150 9092 19156 9104
rect 18656 9064 19156 9092
rect 18656 9052 18662 9064
rect 19150 9052 19156 9064
rect 19208 9052 19214 9104
rect 21652 9092 21680 9132
rect 22002 9120 22008 9172
rect 22060 9160 22066 9172
rect 22097 9163 22155 9169
rect 22097 9160 22109 9163
rect 22060 9132 22109 9160
rect 22060 9120 22066 9132
rect 22097 9129 22109 9132
rect 22143 9129 22155 9163
rect 22097 9123 22155 9129
rect 23842 9120 23848 9172
rect 23900 9120 23906 9172
rect 24118 9120 24124 9172
rect 24176 9120 24182 9172
rect 22738 9092 22744 9104
rect 21652 9064 22744 9092
rect 22738 9052 22744 9064
rect 22796 9052 22802 9104
rect 15841 9027 15899 9033
rect 15841 8993 15853 9027
rect 15887 8993 15899 9027
rect 15841 8987 15899 8993
rect 16298 8984 16304 9036
rect 16356 8984 16362 9036
rect 16390 8984 16396 9036
rect 16448 9024 16454 9036
rect 16758 9033 16764 9036
rect 16577 9027 16635 9033
rect 16577 9024 16589 9027
rect 16448 8996 16589 9024
rect 16448 8984 16454 8996
rect 16577 8993 16589 8996
rect 16623 8993 16635 9027
rect 16577 8987 16635 8993
rect 16715 9027 16764 9033
rect 16715 8993 16727 9027
rect 16761 8993 16764 9027
rect 16715 8987 16764 8993
rect 16758 8984 16764 8987
rect 16816 9024 16822 9036
rect 16816 8996 17540 9024
rect 16816 8984 16822 8996
rect 1854 8916 1860 8968
rect 1912 8916 1918 8968
rect 2131 8959 2189 8965
rect 2131 8925 2143 8959
rect 2177 8956 2189 8959
rect 2222 8956 2228 8968
rect 2177 8928 2228 8956
rect 2177 8925 2189 8928
rect 2131 8919 2189 8925
rect 2222 8916 2228 8928
rect 2280 8916 2286 8968
rect 3326 8916 3332 8968
rect 3384 8956 3390 8968
rect 4062 8956 4068 8968
rect 3384 8928 4068 8956
rect 3384 8916 3390 8928
rect 4062 8916 4068 8928
rect 4120 8916 4126 8968
rect 4157 8959 4215 8965
rect 4157 8925 4169 8959
rect 4203 8956 4215 8959
rect 4430 8956 4436 8968
rect 4203 8928 4292 8956
rect 4391 8928 4436 8956
rect 4203 8925 4215 8928
rect 4157 8919 4215 8925
rect 3050 8848 3056 8900
rect 3108 8888 3114 8900
rect 3510 8888 3516 8900
rect 3108 8860 3516 8888
rect 3108 8848 3114 8860
rect 3510 8848 3516 8860
rect 3568 8848 3574 8900
rect 4264 8832 4292 8928
rect 4430 8916 4436 8928
rect 4488 8916 4494 8968
rect 5537 8959 5595 8965
rect 5537 8925 5549 8959
rect 5583 8956 5595 8959
rect 5644 8956 5672 8984
rect 17512 8968 17540 8996
rect 22094 8984 22100 9036
rect 22152 9024 22158 9036
rect 23109 9027 23167 9033
rect 22152 8996 22600 9024
rect 22152 8984 22158 8996
rect 5583 8928 5672 8956
rect 5721 8959 5779 8965
rect 5583 8925 5595 8928
rect 5537 8919 5595 8925
rect 5721 8925 5733 8959
rect 5767 8956 5779 8959
rect 5902 8956 5908 8968
rect 5767 8928 5908 8956
rect 5767 8925 5779 8928
rect 5721 8919 5779 8925
rect 5902 8916 5908 8928
rect 5960 8916 5966 8968
rect 6454 8916 6460 8968
rect 6512 8916 6518 8968
rect 6546 8916 6552 8968
rect 6604 8965 6610 8968
rect 6604 8959 6632 8965
rect 6620 8925 6632 8959
rect 6604 8919 6632 8925
rect 6604 8916 6610 8919
rect 6730 8916 6736 8968
rect 6788 8916 6794 8968
rect 7469 8959 7527 8965
rect 7469 8956 7481 8959
rect 7392 8928 7481 8956
rect 7392 8900 7420 8928
rect 7469 8925 7481 8928
rect 7515 8925 7527 8959
rect 7469 8919 7527 8925
rect 7650 8916 7656 8968
rect 7708 8956 7714 8968
rect 7743 8959 7801 8965
rect 7743 8956 7755 8959
rect 7708 8928 7755 8956
rect 7708 8916 7714 8928
rect 7743 8925 7755 8928
rect 7789 8925 7801 8959
rect 7743 8919 7801 8925
rect 8754 8916 8760 8968
rect 8812 8956 8818 8968
rect 9585 8959 9643 8965
rect 9585 8956 9597 8959
rect 8812 8928 9597 8956
rect 8812 8916 8818 8928
rect 9585 8925 9597 8928
rect 9631 8925 9643 8959
rect 9585 8919 9643 8925
rect 9859 8959 9917 8965
rect 9859 8925 9871 8959
rect 9905 8956 9917 8959
rect 11699 8959 11757 8965
rect 9905 8928 11652 8956
rect 9905 8925 9917 8928
rect 9859 8919 9917 8925
rect 4540 8860 5764 8888
rect 4540 8832 4568 8860
rect 2038 8780 2044 8832
rect 2096 8820 2102 8832
rect 2774 8820 2780 8832
rect 2096 8792 2780 8820
rect 2096 8780 2102 8792
rect 2774 8780 2780 8792
rect 2832 8780 2838 8832
rect 4246 8780 4252 8832
rect 4304 8780 4310 8832
rect 4522 8780 4528 8832
rect 4580 8780 4586 8832
rect 5074 8780 5080 8832
rect 5132 8820 5138 8832
rect 5169 8823 5227 8829
rect 5169 8820 5181 8823
rect 5132 8792 5181 8820
rect 5132 8780 5138 8792
rect 5169 8789 5181 8792
rect 5215 8789 5227 8823
rect 5736 8820 5764 8860
rect 7374 8848 7380 8900
rect 7432 8848 7438 8900
rect 11164 8832 11192 8928
rect 11624 8888 11652 8928
rect 11699 8925 11711 8959
rect 11745 8956 11757 8959
rect 12342 8956 12348 8968
rect 11745 8928 12348 8956
rect 11745 8925 11757 8928
rect 11699 8919 11757 8925
rect 12342 8916 12348 8928
rect 12400 8956 12406 8968
rect 14826 8956 14832 8968
rect 12400 8928 14832 8956
rect 12400 8916 12406 8928
rect 14826 8916 14832 8928
rect 14884 8916 14890 8968
rect 14918 8916 14924 8968
rect 14976 8956 14982 8968
rect 15657 8959 15715 8965
rect 15657 8956 15669 8959
rect 14976 8928 15669 8956
rect 14976 8916 14982 8928
rect 15657 8925 15669 8928
rect 15703 8925 15715 8959
rect 15657 8919 15715 8925
rect 16850 8916 16856 8968
rect 16908 8916 16914 8968
rect 17494 8916 17500 8968
rect 17552 8916 17558 8968
rect 17589 8959 17647 8965
rect 17589 8925 17601 8959
rect 17635 8956 17647 8959
rect 17678 8956 17684 8968
rect 17635 8928 17684 8956
rect 17635 8925 17647 8928
rect 17589 8919 17647 8925
rect 17678 8916 17684 8928
rect 17736 8956 17742 8968
rect 19245 8959 19303 8965
rect 19245 8956 19257 8959
rect 17736 8928 19257 8956
rect 17736 8916 17742 8928
rect 19245 8925 19257 8928
rect 19291 8925 19303 8959
rect 19245 8919 19303 8925
rect 20717 8959 20775 8965
rect 20717 8925 20729 8959
rect 20763 8956 20775 8959
rect 21266 8956 21272 8968
rect 20763 8928 21272 8956
rect 20763 8925 20775 8928
rect 20717 8919 20775 8925
rect 21266 8916 21272 8928
rect 21324 8956 21330 8968
rect 22186 8956 22192 8968
rect 21324 8928 22192 8956
rect 21324 8916 21330 8928
rect 22186 8916 22192 8928
rect 22244 8916 22250 8968
rect 22278 8916 22284 8968
rect 22336 8916 22342 8968
rect 22572 8965 22600 8996
rect 23109 8993 23121 9027
rect 23155 8993 23167 9027
rect 23109 8987 23167 8993
rect 22557 8959 22615 8965
rect 22557 8925 22569 8959
rect 22603 8925 22615 8959
rect 22557 8919 22615 8925
rect 23014 8916 23020 8968
rect 23072 8916 23078 8968
rect 15194 8888 15200 8900
rect 11624 8860 15200 8888
rect 15194 8848 15200 8860
rect 15252 8848 15258 8900
rect 17856 8891 17914 8897
rect 17856 8857 17868 8891
rect 17902 8888 17914 8891
rect 19334 8888 19340 8900
rect 17902 8860 19340 8888
rect 17902 8857 17914 8860
rect 17856 8851 17914 8857
rect 19334 8848 19340 8860
rect 19392 8848 19398 8900
rect 19512 8891 19570 8897
rect 19512 8857 19524 8891
rect 19558 8857 19570 8891
rect 19512 8851 19570 8857
rect 10318 8820 10324 8832
rect 5736 8792 10324 8820
rect 5169 8783 5227 8789
rect 10318 8780 10324 8792
rect 10376 8780 10382 8832
rect 11146 8780 11152 8832
rect 11204 8780 11210 8832
rect 14458 8780 14464 8832
rect 14516 8820 14522 8832
rect 16390 8820 16396 8832
rect 14516 8792 16396 8820
rect 14516 8780 14522 8792
rect 16390 8780 16396 8792
rect 16448 8780 16454 8832
rect 18969 8823 19027 8829
rect 18969 8789 18981 8823
rect 19015 8820 19027 8823
rect 19150 8820 19156 8832
rect 19015 8792 19156 8820
rect 19015 8789 19027 8792
rect 18969 8783 19027 8789
rect 19150 8780 19156 8792
rect 19208 8780 19214 8832
rect 19527 8820 19555 8851
rect 19702 8848 19708 8900
rect 19760 8888 19766 8900
rect 20990 8897 20996 8900
rect 20984 8888 20996 8897
rect 19760 8860 20760 8888
rect 20951 8860 20996 8888
rect 19760 8848 19766 8860
rect 19886 8820 19892 8832
rect 19527 8792 19892 8820
rect 19886 8780 19892 8792
rect 19944 8780 19950 8832
rect 20622 8780 20628 8832
rect 20680 8780 20686 8832
rect 20732 8820 20760 8860
rect 20984 8851 20996 8860
rect 20990 8848 20996 8851
rect 21048 8848 21054 8900
rect 23124 8888 23152 8987
rect 23566 8916 23572 8968
rect 23624 8916 23630 8968
rect 23860 8965 23888 9120
rect 23845 8959 23903 8965
rect 23845 8925 23857 8959
rect 23891 8925 23903 8959
rect 23845 8919 23903 8925
rect 23937 8959 23995 8965
rect 23937 8925 23949 8959
rect 23983 8925 23995 8959
rect 23937 8919 23995 8925
rect 23952 8888 23980 8919
rect 22066 8860 23152 8888
rect 23676 8860 23980 8888
rect 22066 8820 22094 8860
rect 20732 8792 22094 8820
rect 23382 8780 23388 8832
rect 23440 8780 23446 8832
rect 23676 8829 23704 8860
rect 23661 8823 23719 8829
rect 23661 8789 23673 8823
rect 23707 8789 23719 8823
rect 23661 8783 23719 8789
rect 1104 8730 24723 8752
rect 1104 8678 6814 8730
rect 6866 8678 6878 8730
rect 6930 8678 6942 8730
rect 6994 8678 7006 8730
rect 7058 8678 7070 8730
rect 7122 8678 12679 8730
rect 12731 8678 12743 8730
rect 12795 8678 12807 8730
rect 12859 8678 12871 8730
rect 12923 8678 12935 8730
rect 12987 8678 18544 8730
rect 18596 8678 18608 8730
rect 18660 8678 18672 8730
rect 18724 8678 18736 8730
rect 18788 8678 18800 8730
rect 18852 8678 24409 8730
rect 24461 8678 24473 8730
rect 24525 8678 24537 8730
rect 24589 8678 24601 8730
rect 24653 8678 24665 8730
rect 24717 8678 24723 8730
rect 1104 8656 24723 8678
rect 2314 8576 2320 8628
rect 2372 8616 2378 8628
rect 5721 8619 5779 8625
rect 5721 8616 5733 8619
rect 2372 8588 5733 8616
rect 2372 8576 2378 8588
rect 5721 8585 5733 8588
rect 5767 8585 5779 8619
rect 5721 8579 5779 8585
rect 6730 8576 6736 8628
rect 6788 8616 6794 8628
rect 7377 8619 7435 8625
rect 7377 8616 7389 8619
rect 6788 8588 7389 8616
rect 6788 8576 6794 8588
rect 7377 8585 7389 8588
rect 7423 8585 7435 8619
rect 7377 8579 7435 8585
rect 7650 8576 7656 8628
rect 7708 8616 7714 8628
rect 11238 8616 11244 8628
rect 7708 8588 11244 8616
rect 7708 8576 7714 8588
rect 11238 8576 11244 8588
rect 11296 8576 11302 8628
rect 11330 8576 11336 8628
rect 11388 8616 11394 8628
rect 13262 8616 13268 8628
rect 11388 8588 13268 8616
rect 11388 8576 11394 8588
rect 13262 8576 13268 8588
rect 13320 8616 13326 8628
rect 16758 8616 16764 8628
rect 13320 8588 16764 8616
rect 13320 8576 13326 8588
rect 16758 8576 16764 8588
rect 16816 8576 16822 8628
rect 16850 8576 16856 8628
rect 16908 8616 16914 8628
rect 17681 8619 17739 8625
rect 17681 8616 17693 8619
rect 16908 8588 17693 8616
rect 16908 8576 16914 8588
rect 17681 8585 17693 8588
rect 17727 8585 17739 8619
rect 17681 8579 17739 8585
rect 18141 8619 18199 8625
rect 18141 8585 18153 8619
rect 18187 8616 18199 8619
rect 18230 8616 18236 8628
rect 18187 8588 18236 8616
rect 18187 8585 18199 8588
rect 18141 8579 18199 8585
rect 18230 8576 18236 8588
rect 18288 8576 18294 8628
rect 18322 8576 18328 8628
rect 18380 8616 18386 8628
rect 18417 8619 18475 8625
rect 18417 8616 18429 8619
rect 18380 8588 18429 8616
rect 18380 8576 18386 8588
rect 18417 8585 18429 8588
rect 18463 8585 18475 8619
rect 18417 8579 18475 8585
rect 19610 8576 19616 8628
rect 19668 8576 19674 8628
rect 19702 8576 19708 8628
rect 19760 8576 19766 8628
rect 19978 8576 19984 8628
rect 20036 8616 20042 8628
rect 20165 8619 20223 8625
rect 20165 8616 20177 8619
rect 20036 8588 20177 8616
rect 20036 8576 20042 8588
rect 20165 8585 20177 8588
rect 20211 8585 20223 8619
rect 20165 8579 20223 8585
rect 20622 8576 20628 8628
rect 20680 8576 20686 8628
rect 20809 8619 20867 8625
rect 20809 8585 20821 8619
rect 20855 8616 20867 8619
rect 21174 8616 21180 8628
rect 20855 8588 21180 8616
rect 20855 8585 20867 8588
rect 20809 8579 20867 8585
rect 21174 8576 21180 8588
rect 21232 8576 21238 8628
rect 23750 8576 23756 8628
rect 23808 8576 23814 8628
rect 24029 8619 24087 8625
rect 24029 8585 24041 8619
rect 24075 8585 24087 8619
rect 24029 8579 24087 8585
rect 3234 8508 3240 8560
rect 3292 8548 3298 8560
rect 3292 8520 4108 8548
rect 3292 8508 3298 8520
rect 1670 8440 1676 8492
rect 1728 8440 1734 8492
rect 2409 8483 2467 8489
rect 2409 8449 2421 8483
rect 2455 8449 2467 8483
rect 2409 8443 2467 8449
rect 1302 8372 1308 8424
rect 1360 8372 1366 8424
rect 1486 8372 1492 8424
rect 1544 8372 1550 8424
rect 2038 8372 2044 8424
rect 2096 8412 2102 8424
rect 2424 8412 2452 8443
rect 2682 8440 2688 8492
rect 2740 8440 2746 8492
rect 3694 8440 3700 8492
rect 3752 8480 3758 8492
rect 4080 8489 4108 8520
rect 6623 8513 6681 8519
rect 3881 8483 3939 8489
rect 3881 8480 3893 8483
rect 3752 8452 3893 8480
rect 3752 8440 3758 8452
rect 3881 8449 3893 8452
rect 3927 8449 3939 8483
rect 3881 8443 3939 8449
rect 4065 8483 4123 8489
rect 4065 8449 4077 8483
rect 4111 8449 4123 8483
rect 4065 8443 4123 8449
rect 5074 8440 5080 8492
rect 5132 8440 5138 8492
rect 5994 8440 6000 8492
rect 6052 8440 6058 8492
rect 6623 8479 6635 8513
rect 6669 8510 6681 8513
rect 6669 8482 6776 8510
rect 10042 8508 10048 8560
rect 10100 8548 10106 8560
rect 19720 8548 19748 8576
rect 10100 8520 19748 8548
rect 10100 8508 10106 8520
rect 6669 8479 6681 8482
rect 6623 8473 6681 8479
rect 6748 8480 6776 8482
rect 7558 8480 7564 8492
rect 6748 8452 7564 8480
rect 7558 8440 7564 8452
rect 7616 8440 7622 8492
rect 8295 8483 8353 8489
rect 8295 8449 8307 8483
rect 8341 8480 8353 8483
rect 8386 8480 8392 8492
rect 8341 8452 8392 8480
rect 8341 8449 8353 8452
rect 8295 8443 8353 8449
rect 8386 8440 8392 8452
rect 8444 8480 8450 8492
rect 8846 8480 8852 8492
rect 8444 8452 8852 8480
rect 8444 8440 8450 8452
rect 8846 8440 8852 8452
rect 8904 8440 8910 8492
rect 10594 8440 10600 8492
rect 10652 8480 10658 8492
rect 10962 8480 10968 8492
rect 10652 8452 10968 8480
rect 10652 8440 10658 8452
rect 10962 8440 10968 8452
rect 11020 8480 11026 8492
rect 15470 8480 15476 8492
rect 11020 8452 15476 8480
rect 11020 8440 11026 8452
rect 15470 8440 15476 8452
rect 15528 8440 15534 8492
rect 16943 8483 17001 8489
rect 16943 8449 16955 8483
rect 16989 8480 17001 8483
rect 17310 8480 17316 8492
rect 16989 8452 17316 8480
rect 16989 8449 17001 8452
rect 16943 8443 17001 8449
rect 17310 8440 17316 8452
rect 17368 8440 17374 8492
rect 18049 8483 18107 8489
rect 18049 8449 18061 8483
rect 18095 8449 18107 8483
rect 18049 8443 18107 8449
rect 2096 8384 2452 8412
rect 2547 8415 2605 8421
rect 2096 8372 2102 8384
rect 2547 8381 2559 8415
rect 2593 8412 2605 8415
rect 3050 8412 3056 8424
rect 2593 8384 3056 8412
rect 2593 8381 2605 8384
rect 2547 8375 2605 8381
rect 3050 8372 3056 8384
rect 3108 8412 3114 8424
rect 3786 8412 3792 8424
rect 3108 8384 3792 8412
rect 3108 8372 3114 8384
rect 3786 8372 3792 8384
rect 3844 8372 3850 8424
rect 4614 8372 4620 8424
rect 4672 8412 4678 8424
rect 4801 8415 4859 8421
rect 4801 8412 4813 8415
rect 4672 8384 4813 8412
rect 4672 8372 4678 8384
rect 4801 8381 4813 8384
rect 4847 8381 4859 8415
rect 4801 8375 4859 8381
rect 4890 8372 4896 8424
rect 4948 8421 4954 8424
rect 4948 8415 4997 8421
rect 4948 8381 4951 8415
rect 4985 8412 4997 8415
rect 6012 8412 6040 8440
rect 4985 8384 6040 8412
rect 4985 8381 4997 8384
rect 4948 8375 4997 8381
rect 4948 8372 4954 8375
rect 6178 8372 6184 8424
rect 6236 8412 6242 8424
rect 6365 8415 6423 8421
rect 6365 8412 6377 8415
rect 6236 8384 6377 8412
rect 6236 8372 6242 8384
rect 6365 8381 6377 8384
rect 6411 8381 6423 8415
rect 6365 8375 6423 8381
rect 7374 8372 7380 8424
rect 7432 8412 7438 8424
rect 8021 8415 8079 8421
rect 8021 8412 8033 8415
rect 7432 8384 8033 8412
rect 7432 8372 7438 8384
rect 8021 8381 8033 8384
rect 8067 8381 8079 8415
rect 8021 8375 8079 8381
rect 14734 8372 14740 8424
rect 14792 8412 14798 8424
rect 15197 8415 15255 8421
rect 15197 8412 15209 8415
rect 14792 8384 15209 8412
rect 14792 8372 14798 8384
rect 15197 8381 15209 8384
rect 15243 8381 15255 8415
rect 16669 8415 16727 8421
rect 16669 8412 16681 8415
rect 15197 8375 15255 8381
rect 15856 8384 16681 8412
rect 1320 8344 1348 8372
rect 2056 8344 2084 8372
rect 1320 8316 2084 8344
rect 2130 8304 2136 8356
rect 2188 8304 2194 8356
rect 3878 8344 3884 8356
rect 3804 8316 3884 8344
rect 2038 8236 2044 8288
rect 2096 8276 2102 8288
rect 3329 8279 3387 8285
rect 3329 8276 3341 8279
rect 2096 8248 3341 8276
rect 2096 8236 2102 8248
rect 3329 8245 3341 8248
rect 3375 8245 3387 8279
rect 3329 8239 3387 8245
rect 3605 8279 3663 8285
rect 3605 8245 3617 8279
rect 3651 8276 3663 8279
rect 3804 8276 3832 8316
rect 3878 8304 3884 8316
rect 3936 8304 3942 8356
rect 4522 8304 4528 8356
rect 4580 8304 4586 8356
rect 5718 8304 5724 8356
rect 5776 8344 5782 8356
rect 6196 8344 6224 8372
rect 11054 8344 11060 8356
rect 5776 8316 6224 8344
rect 7024 8316 8156 8344
rect 5776 8304 5782 8316
rect 3651 8248 3832 8276
rect 3651 8245 3663 8248
rect 3605 8239 3663 8245
rect 4062 8236 4068 8288
rect 4120 8276 4126 8288
rect 4982 8276 4988 8288
rect 4120 8248 4988 8276
rect 4120 8236 4126 8248
rect 4982 8236 4988 8248
rect 5040 8236 5046 8288
rect 5902 8236 5908 8288
rect 5960 8276 5966 8288
rect 7024 8276 7052 8316
rect 5960 8248 7052 8276
rect 5960 8236 5966 8248
rect 7650 8236 7656 8288
rect 7708 8276 7714 8288
rect 7834 8276 7840 8288
rect 7708 8248 7840 8276
rect 7708 8236 7714 8248
rect 7834 8236 7840 8248
rect 7892 8236 7898 8288
rect 8128 8276 8156 8316
rect 8680 8316 11060 8344
rect 8680 8276 8708 8316
rect 11054 8304 11060 8316
rect 11112 8304 11118 8356
rect 8128 8248 8708 8276
rect 8938 8236 8944 8288
rect 8996 8276 9002 8288
rect 9033 8279 9091 8285
rect 9033 8276 9045 8279
rect 8996 8248 9045 8276
rect 8996 8236 9002 8248
rect 9033 8245 9045 8248
rect 9079 8245 9091 8279
rect 15212 8276 15240 8375
rect 15856 8276 15884 8384
rect 16669 8381 16681 8384
rect 16715 8381 16727 8415
rect 16669 8375 16727 8381
rect 15212 8248 15884 8276
rect 16209 8279 16267 8285
rect 9033 8239 9091 8245
rect 16209 8245 16221 8279
rect 16255 8276 16267 8279
rect 16298 8276 16304 8288
rect 16255 8248 16304 8276
rect 16255 8245 16267 8248
rect 16209 8239 16267 8245
rect 16298 8236 16304 8248
rect 16356 8236 16362 8288
rect 16684 8276 16712 8375
rect 18064 8344 18092 8443
rect 18138 8440 18144 8492
rect 18196 8480 18202 8492
rect 18325 8483 18383 8489
rect 18325 8480 18337 8483
rect 18196 8452 18337 8480
rect 18196 8440 18202 8452
rect 18325 8449 18337 8452
rect 18371 8449 18383 8483
rect 18325 8443 18383 8449
rect 18509 8483 18567 8489
rect 18509 8449 18521 8483
rect 18555 8449 18567 8483
rect 18509 8443 18567 8449
rect 18785 8483 18843 8489
rect 18785 8449 18797 8483
rect 18831 8480 18843 8483
rect 19061 8483 19119 8489
rect 18831 8452 19012 8480
rect 18831 8449 18843 8452
rect 18785 8443 18843 8449
rect 18524 8412 18552 8443
rect 18984 8412 19012 8452
rect 19061 8449 19073 8483
rect 19107 8480 19119 8483
rect 19150 8480 19156 8492
rect 19107 8452 19156 8480
rect 19107 8449 19119 8452
rect 19061 8443 19119 8449
rect 19150 8440 19156 8452
rect 19208 8440 19214 8492
rect 19521 8483 19579 8489
rect 19521 8449 19533 8483
rect 19567 8480 19579 8483
rect 19567 8452 19840 8480
rect 19567 8449 19579 8452
rect 19521 8443 19579 8449
rect 19334 8412 19340 8424
rect 18524 8384 18920 8412
rect 18984 8384 19340 8412
rect 18892 8353 18920 8384
rect 19334 8372 19340 8384
rect 19392 8372 19398 8424
rect 18601 8347 18659 8353
rect 18601 8344 18613 8347
rect 18064 8316 18613 8344
rect 18601 8313 18613 8316
rect 18647 8313 18659 8347
rect 18601 8307 18659 8313
rect 18877 8347 18935 8353
rect 18877 8313 18889 8347
rect 18923 8313 18935 8347
rect 18877 8307 18935 8313
rect 17862 8276 17868 8288
rect 16684 8248 17868 8276
rect 17862 8236 17868 8248
rect 17920 8236 17926 8288
rect 19352 8276 19380 8372
rect 19812 8353 19840 8452
rect 19886 8440 19892 8492
rect 19944 8480 19950 8492
rect 19981 8483 20039 8489
rect 19981 8480 19993 8483
rect 19944 8452 19993 8480
rect 19944 8440 19950 8452
rect 19981 8449 19993 8452
rect 20027 8449 20039 8483
rect 19981 8443 20039 8449
rect 20349 8483 20407 8489
rect 20349 8449 20361 8483
rect 20395 8480 20407 8483
rect 20640 8480 20668 8576
rect 22548 8551 22606 8557
rect 22548 8517 22560 8551
rect 22594 8548 22606 8551
rect 23198 8548 23204 8560
rect 22594 8520 23204 8548
rect 22594 8517 22606 8520
rect 22548 8511 22606 8517
rect 23198 8508 23204 8520
rect 23256 8548 23262 8560
rect 24044 8548 24072 8579
rect 23256 8520 24072 8548
rect 23256 8508 23262 8520
rect 20395 8452 20668 8480
rect 20395 8449 20407 8452
rect 20349 8443 20407 8449
rect 19996 8412 20024 8443
rect 20990 8440 20996 8492
rect 21048 8480 21054 8492
rect 21048 8452 21864 8480
rect 21048 8440 21054 8452
rect 20714 8412 20720 8424
rect 19996 8384 20720 8412
rect 20714 8372 20720 8384
rect 20772 8372 20778 8424
rect 21836 8356 21864 8452
rect 22002 8440 22008 8492
rect 22060 8440 22066 8492
rect 22370 8440 22376 8492
rect 22428 8440 22434 8492
rect 23937 8483 23995 8489
rect 23937 8480 23949 8483
rect 23676 8452 23949 8480
rect 22094 8372 22100 8424
rect 22152 8372 22158 8424
rect 22186 8372 22192 8424
rect 22244 8412 22250 8424
rect 22281 8415 22339 8421
rect 22281 8412 22293 8415
rect 22244 8384 22293 8412
rect 22244 8372 22250 8384
rect 22281 8381 22293 8384
rect 22327 8412 22339 8415
rect 22388 8412 22416 8440
rect 22327 8384 22416 8412
rect 22327 8381 22339 8384
rect 22281 8375 22339 8381
rect 19797 8347 19855 8353
rect 19797 8313 19809 8347
rect 19843 8313 19855 8347
rect 19797 8307 19855 8313
rect 21818 8304 21824 8356
rect 21876 8304 21882 8356
rect 23676 8353 23704 8452
rect 23937 8449 23949 8452
rect 23983 8449 23995 8483
rect 23937 8443 23995 8449
rect 24210 8440 24216 8492
rect 24268 8440 24274 8492
rect 23661 8347 23719 8353
rect 23661 8313 23673 8347
rect 23707 8313 23719 8347
rect 23661 8307 23719 8313
rect 19352 8248 24624 8276
rect 1104 8186 24564 8208
rect 1104 8134 3882 8186
rect 3934 8134 3946 8186
rect 3998 8134 4010 8186
rect 4062 8134 4074 8186
rect 4126 8134 4138 8186
rect 4190 8134 9747 8186
rect 9799 8134 9811 8186
rect 9863 8134 9875 8186
rect 9927 8134 9939 8186
rect 9991 8134 10003 8186
rect 10055 8134 15612 8186
rect 15664 8134 15676 8186
rect 15728 8134 15740 8186
rect 15792 8134 15804 8186
rect 15856 8134 15868 8186
rect 15920 8134 21477 8186
rect 21529 8134 21541 8186
rect 21593 8134 21605 8186
rect 21657 8134 21669 8186
rect 21721 8134 21733 8186
rect 21785 8134 24564 8186
rect 1104 8112 24564 8134
rect 1854 8032 1860 8084
rect 1912 8032 1918 8084
rect 1946 8032 1952 8084
rect 2004 8032 2010 8084
rect 3329 8075 3387 8081
rect 2332 8044 3004 8072
rect 1872 8004 1900 8032
rect 2332 8004 2360 8044
rect 1872 7976 2360 8004
rect 2332 7945 2360 7976
rect 2317 7939 2375 7945
rect 2317 7905 2329 7939
rect 2363 7905 2375 7939
rect 2976 7936 3004 8044
rect 3329 8041 3341 8075
rect 3375 8072 3387 8075
rect 3602 8072 3608 8084
rect 3375 8044 3608 8072
rect 3375 8041 3387 8044
rect 3329 8035 3387 8041
rect 3602 8032 3608 8044
rect 3660 8032 3666 8084
rect 4246 8072 4252 8084
rect 3804 8044 4252 8072
rect 3602 7936 3608 7948
rect 2976 7908 3608 7936
rect 2317 7899 2375 7905
rect 3602 7896 3608 7908
rect 3660 7896 3666 7948
rect 3804 7945 3832 8044
rect 4246 8032 4252 8044
rect 4304 8032 4310 8084
rect 4522 8032 4528 8084
rect 4580 8072 4586 8084
rect 4801 8075 4859 8081
rect 4801 8072 4813 8075
rect 4580 8044 4813 8072
rect 4580 8032 4586 8044
rect 4801 8041 4813 8044
rect 4847 8041 4859 8075
rect 4801 8035 4859 8041
rect 5534 8032 5540 8084
rect 5592 8072 5598 8084
rect 5905 8075 5963 8081
rect 5905 8072 5917 8075
rect 5592 8044 5917 8072
rect 5592 8032 5598 8044
rect 5905 8041 5917 8044
rect 5951 8041 5963 8075
rect 7374 8072 7380 8084
rect 5905 8035 5963 8041
rect 7300 8044 7380 8072
rect 3789 7939 3847 7945
rect 3789 7905 3801 7939
rect 3835 7905 3847 7939
rect 3789 7899 3847 7905
rect 2498 7828 2504 7880
rect 2556 7868 2562 7880
rect 2591 7871 2649 7877
rect 2591 7868 2603 7871
rect 2556 7840 2603 7868
rect 2556 7828 2562 7840
rect 2591 7837 2603 7840
rect 2637 7837 2649 7871
rect 4062 7868 4068 7880
rect 4023 7840 4068 7868
rect 2591 7831 2649 7837
rect 4062 7828 4068 7840
rect 4120 7828 4126 7880
rect 5166 7828 5172 7880
rect 5224 7868 5230 7880
rect 5813 7871 5871 7877
rect 5813 7868 5825 7871
rect 5224 7840 5825 7868
rect 5224 7828 5230 7840
rect 5813 7837 5825 7840
rect 5859 7837 5871 7871
rect 5813 7831 5871 7837
rect 6086 7828 6092 7880
rect 6144 7868 6150 7880
rect 7300 7877 7328 8044
rect 7374 8032 7380 8044
rect 7432 8032 7438 8084
rect 8662 8032 8668 8084
rect 8720 8072 8726 8084
rect 8720 8044 11008 8072
rect 8720 8032 8726 8044
rect 10980 7948 11008 8044
rect 11330 8032 11336 8084
rect 11388 8072 11394 8084
rect 12158 8072 12164 8084
rect 11388 8044 12164 8072
rect 11388 8032 11394 8044
rect 12158 8032 12164 8044
rect 12216 8032 12222 8084
rect 13817 8075 13875 8081
rect 13817 8041 13829 8075
rect 13863 8072 13875 8075
rect 13998 8072 14004 8084
rect 13863 8044 14004 8072
rect 13863 8041 13875 8044
rect 13817 8035 13875 8041
rect 13998 8032 14004 8044
rect 14056 8032 14062 8084
rect 22186 8032 22192 8084
rect 22244 8072 22250 8084
rect 22833 8075 22891 8081
rect 22833 8072 22845 8075
rect 22244 8044 22845 8072
rect 22244 8032 22250 8044
rect 22833 8041 22845 8044
rect 22879 8041 22891 8075
rect 22833 8035 22891 8041
rect 23014 8032 23020 8084
rect 23072 8072 23078 8084
rect 23201 8075 23259 8081
rect 23201 8072 23213 8075
rect 23072 8044 23213 8072
rect 23072 8032 23078 8044
rect 23201 8041 23213 8044
rect 23247 8041 23259 8075
rect 23201 8035 23259 8041
rect 23750 8032 23756 8084
rect 23808 8032 23814 8084
rect 24213 8075 24271 8081
rect 24213 8041 24225 8075
rect 24259 8072 24271 8075
rect 24596 8072 24624 8248
rect 24259 8044 24624 8072
rect 24259 8041 24271 8044
rect 24213 8035 24271 8041
rect 22278 7964 22284 8016
rect 22336 8004 22342 8016
rect 22465 8007 22523 8013
rect 22465 8004 22477 8007
rect 22336 7976 22477 8004
rect 22336 7964 22342 7976
rect 22465 7973 22477 7976
rect 22511 7973 22523 8007
rect 22465 7967 22523 7973
rect 13544 7948 13596 7954
rect 9858 7896 9864 7948
rect 9916 7936 9922 7948
rect 9916 7908 10732 7936
rect 9916 7896 9922 7908
rect 7285 7871 7343 7877
rect 7285 7868 7297 7871
rect 6144 7840 7297 7868
rect 6144 7828 6150 7840
rect 7285 7837 7297 7840
rect 7331 7837 7343 7871
rect 7285 7831 7343 7837
rect 7559 7871 7617 7877
rect 7559 7837 7571 7871
rect 7605 7868 7617 7871
rect 7650 7868 7656 7880
rect 7605 7840 7656 7868
rect 7605 7837 7617 7840
rect 7559 7831 7617 7837
rect 7650 7828 7656 7840
rect 7708 7828 7714 7880
rect 8754 7828 8760 7880
rect 8812 7868 8818 7880
rect 9125 7871 9183 7877
rect 9125 7868 9137 7871
rect 8812 7840 9137 7868
rect 8812 7828 8818 7840
rect 9125 7837 9137 7840
rect 9171 7837 9183 7871
rect 9125 7831 9183 7837
rect 9399 7871 9457 7877
rect 9399 7837 9411 7871
rect 9445 7868 9457 7871
rect 10594 7868 10600 7880
rect 9445 7840 10600 7868
rect 9445 7837 9457 7840
rect 9399 7831 9457 7837
rect 1857 7803 1915 7809
rect 1857 7769 1869 7803
rect 1903 7800 1915 7803
rect 4338 7800 4344 7812
rect 1903 7772 4344 7800
rect 1903 7769 1915 7772
rect 1857 7763 1915 7769
rect 4338 7760 4344 7772
rect 4396 7760 4402 7812
rect 4430 7760 4436 7812
rect 4488 7800 4494 7812
rect 5261 7803 5319 7809
rect 5261 7800 5273 7803
rect 4488 7772 5273 7800
rect 4488 7760 4494 7772
rect 5261 7769 5273 7772
rect 5307 7769 5319 7803
rect 9508 7800 9536 7840
rect 10594 7828 10600 7840
rect 10652 7828 10658 7880
rect 10704 7868 10732 7908
rect 10962 7896 10968 7948
rect 11020 7896 11026 7948
rect 22480 7936 22508 7967
rect 22554 7964 22560 8016
rect 22612 8004 22618 8016
rect 23569 8007 23627 8013
rect 23569 8004 23581 8007
rect 22612 7976 23581 8004
rect 22612 7964 22618 7976
rect 23569 7973 23581 7976
rect 23615 7973 23627 8007
rect 23569 7967 23627 7973
rect 23768 7936 23796 8032
rect 25590 7936 25596 7948
rect 22480 7908 23152 7936
rect 13544 7890 13596 7896
rect 11207 7871 11265 7877
rect 11207 7868 11219 7871
rect 10704 7840 11219 7868
rect 11207 7837 11219 7840
rect 11253 7837 11265 7871
rect 12897 7871 12955 7877
rect 11207 7831 11265 7837
rect 11716 7840 12434 7868
rect 5261 7763 5319 7769
rect 6748 7772 9536 7800
rect 6748 7744 6776 7772
rect 10318 7760 10324 7812
rect 10376 7800 10382 7812
rect 11716 7800 11744 7840
rect 10376 7772 11744 7800
rect 10376 7760 10382 7772
rect 11790 7760 11796 7812
rect 11848 7800 11854 7812
rect 12406 7800 12434 7840
rect 12897 7837 12909 7871
rect 12943 7868 12955 7871
rect 12943 7840 13492 7868
rect 12943 7837 12955 7840
rect 12897 7831 12955 7837
rect 12805 7803 12863 7809
rect 11848 7772 12112 7800
rect 12406 7772 12756 7800
rect 11848 7760 11854 7772
rect 12084 7744 12112 7772
rect 4062 7692 4068 7744
rect 4120 7732 4126 7744
rect 5353 7735 5411 7741
rect 5353 7732 5365 7735
rect 4120 7704 5365 7732
rect 4120 7692 4126 7704
rect 5353 7701 5365 7704
rect 5399 7701 5411 7735
rect 5353 7695 5411 7701
rect 6730 7692 6736 7744
rect 6788 7692 6794 7744
rect 8294 7692 8300 7744
rect 8352 7692 8358 7744
rect 8662 7692 8668 7744
rect 8720 7732 8726 7744
rect 9306 7732 9312 7744
rect 8720 7704 9312 7732
rect 8720 7692 8726 7704
rect 9306 7692 9312 7704
rect 9364 7692 9370 7744
rect 9398 7692 9404 7744
rect 9456 7732 9462 7744
rect 9674 7732 9680 7744
rect 9456 7704 9680 7732
rect 9456 7692 9462 7704
rect 9674 7692 9680 7704
rect 9732 7692 9738 7744
rect 10042 7692 10048 7744
rect 10100 7732 10106 7744
rect 10137 7735 10195 7741
rect 10137 7732 10149 7735
rect 10100 7704 10149 7732
rect 10100 7692 10106 7704
rect 10137 7701 10149 7704
rect 10183 7701 10195 7735
rect 10137 7695 10195 7701
rect 11882 7692 11888 7744
rect 11940 7732 11946 7744
rect 11977 7735 12035 7741
rect 11977 7732 11989 7735
rect 11940 7704 11989 7732
rect 11940 7692 11946 7704
rect 11977 7701 11989 7704
rect 12023 7701 12035 7735
rect 11977 7695 12035 7701
rect 12066 7692 12072 7744
rect 12124 7732 12130 7744
rect 12526 7732 12532 7744
rect 12124 7704 12532 7732
rect 12124 7692 12130 7704
rect 12526 7692 12532 7704
rect 12584 7692 12590 7744
rect 12728 7732 12756 7772
rect 12805 7769 12817 7803
rect 12851 7800 12863 7803
rect 13078 7800 13084 7812
rect 12851 7772 13084 7800
rect 12851 7769 12863 7772
rect 12805 7763 12863 7769
rect 13078 7760 13084 7772
rect 13136 7760 13142 7812
rect 13265 7803 13323 7809
rect 13265 7769 13277 7803
rect 13311 7800 13323 7803
rect 13354 7800 13360 7812
rect 13311 7772 13360 7800
rect 13311 7769 13323 7772
rect 13265 7763 13323 7769
rect 13354 7760 13360 7772
rect 13412 7760 13418 7812
rect 13464 7800 13492 7840
rect 13906 7828 13912 7880
rect 13964 7868 13970 7880
rect 14734 7868 14740 7880
rect 13964 7840 14740 7868
rect 13964 7828 13970 7840
rect 14734 7828 14740 7840
rect 14792 7868 14798 7880
rect 14829 7871 14887 7877
rect 14829 7868 14841 7871
rect 14792 7840 14841 7868
rect 14792 7828 14798 7840
rect 14829 7837 14841 7840
rect 14875 7837 14887 7871
rect 15102 7868 15108 7880
rect 15063 7840 15108 7868
rect 14829 7831 14887 7837
rect 15102 7828 15108 7840
rect 15160 7828 15166 7880
rect 15194 7828 15200 7880
rect 15252 7868 15258 7880
rect 16114 7868 16120 7880
rect 15252 7840 16120 7868
rect 15252 7828 15258 7840
rect 16114 7828 16120 7840
rect 16172 7828 16178 7880
rect 19426 7828 19432 7880
rect 19484 7868 19490 7880
rect 23124 7877 23152 7908
rect 23308 7908 23796 7936
rect 25424 7908 25596 7936
rect 21453 7871 21511 7877
rect 21453 7868 21465 7871
rect 19484 7840 21465 7868
rect 19484 7828 19490 7840
rect 21453 7837 21465 7840
rect 21499 7837 21511 7871
rect 21695 7871 21753 7877
rect 21695 7868 21707 7871
rect 21453 7831 21511 7837
rect 21560 7840 21707 7868
rect 13464 7772 13584 7800
rect 13446 7732 13452 7744
rect 12728 7704 13452 7732
rect 13446 7692 13452 7704
rect 13504 7692 13510 7744
rect 13556 7732 13584 7772
rect 13630 7760 13636 7812
rect 13688 7760 13694 7812
rect 21358 7760 21364 7812
rect 21416 7800 21422 7812
rect 21560 7800 21588 7840
rect 21695 7837 21707 7840
rect 21741 7837 21753 7871
rect 21695 7831 21753 7837
rect 23017 7871 23075 7877
rect 23017 7837 23029 7871
rect 23063 7837 23075 7871
rect 23017 7831 23075 7837
rect 23109 7871 23167 7877
rect 23109 7837 23121 7871
rect 23155 7837 23167 7871
rect 23109 7831 23167 7837
rect 21416 7772 21588 7800
rect 23032 7800 23060 7831
rect 23198 7828 23204 7880
rect 23256 7828 23262 7880
rect 23308 7877 23336 7908
rect 23293 7871 23351 7877
rect 23293 7837 23305 7871
rect 23339 7837 23351 7871
rect 23293 7831 23351 7837
rect 23382 7828 23388 7880
rect 23440 7828 23446 7880
rect 23845 7871 23903 7877
rect 23845 7837 23857 7871
rect 23891 7868 23903 7871
rect 23934 7868 23940 7880
rect 23891 7840 23940 7868
rect 23891 7837 23903 7840
rect 23845 7831 23903 7837
rect 23934 7828 23940 7840
rect 23992 7828 23998 7880
rect 24026 7828 24032 7880
rect 24084 7828 24090 7880
rect 23216 7800 23244 7828
rect 23032 7772 23244 7800
rect 21416 7760 21422 7772
rect 25424 7744 25452 7908
rect 25590 7896 25596 7908
rect 25648 7896 25654 7948
rect 14182 7732 14188 7744
rect 13556 7704 14188 7732
rect 14182 7692 14188 7704
rect 14240 7692 14246 7744
rect 15654 7692 15660 7744
rect 15712 7732 15718 7744
rect 15841 7735 15899 7741
rect 15841 7732 15853 7735
rect 15712 7704 15853 7732
rect 15712 7692 15718 7704
rect 15841 7701 15853 7704
rect 15887 7701 15899 7735
rect 15841 7695 15899 7701
rect 16850 7692 16856 7744
rect 16908 7732 16914 7744
rect 17310 7732 17316 7744
rect 16908 7704 17316 7732
rect 16908 7692 16914 7704
rect 17310 7692 17316 7704
rect 17368 7692 17374 7744
rect 23658 7692 23664 7744
rect 23716 7692 23722 7744
rect 25406 7692 25412 7744
rect 25464 7692 25470 7744
rect 1104 7642 24723 7664
rect 1104 7590 6814 7642
rect 6866 7590 6878 7642
rect 6930 7590 6942 7642
rect 6994 7590 7006 7642
rect 7058 7590 7070 7642
rect 7122 7590 12679 7642
rect 12731 7590 12743 7642
rect 12795 7590 12807 7642
rect 12859 7590 12871 7642
rect 12923 7590 12935 7642
rect 12987 7590 18544 7642
rect 18596 7590 18608 7642
rect 18660 7590 18672 7642
rect 18724 7590 18736 7642
rect 18788 7590 18800 7642
rect 18852 7590 24409 7642
rect 24461 7590 24473 7642
rect 24525 7590 24537 7642
rect 24589 7590 24601 7642
rect 24653 7590 24665 7642
rect 24717 7590 24723 7642
rect 1104 7568 24723 7590
rect 1762 7488 1768 7540
rect 1820 7488 1826 7540
rect 2501 7531 2559 7537
rect 2501 7497 2513 7531
rect 2547 7528 2559 7531
rect 2682 7528 2688 7540
rect 2547 7500 2688 7528
rect 2547 7497 2559 7500
rect 2501 7491 2559 7497
rect 2682 7488 2688 7500
rect 2740 7488 2746 7540
rect 3068 7500 3832 7528
rect 1780 7460 1808 7488
rect 1504 7432 1808 7460
rect 1394 7352 1400 7404
rect 1452 7392 1458 7404
rect 1504 7401 1532 7432
rect 1489 7395 1547 7401
rect 1489 7392 1501 7395
rect 1452 7364 1501 7392
rect 1452 7352 1458 7364
rect 1489 7361 1501 7364
rect 1535 7361 1547 7395
rect 1489 7355 1547 7361
rect 1763 7395 1821 7401
rect 1763 7361 1775 7395
rect 1809 7392 1821 7395
rect 1809 7364 2774 7392
rect 1809 7361 1821 7364
rect 1763 7355 1821 7361
rect 2746 7188 2774 7364
rect 3068 7324 3096 7500
rect 3142 7420 3148 7472
rect 3200 7420 3206 7472
rect 3160 7392 3188 7420
rect 3403 7405 3461 7411
rect 3403 7402 3415 7405
rect 3344 7392 3415 7402
rect 3160 7374 3415 7392
rect 3160 7364 3372 7374
rect 3403 7371 3415 7374
rect 3449 7371 3461 7405
rect 3403 7365 3461 7371
rect 3510 7352 3516 7404
rect 3568 7392 3574 7404
rect 3804 7392 3832 7500
rect 4062 7488 4068 7540
rect 4120 7528 4126 7540
rect 5813 7531 5871 7537
rect 5813 7528 5825 7531
rect 4120 7500 5825 7528
rect 4120 7488 4126 7500
rect 5813 7497 5825 7500
rect 5859 7497 5871 7531
rect 5813 7491 5871 7497
rect 7374 7488 7380 7540
rect 7432 7528 7438 7540
rect 7432 7500 13366 7528
rect 7432 7488 7438 7500
rect 4154 7420 4160 7472
rect 4212 7460 4218 7472
rect 4522 7460 4528 7472
rect 4212 7432 4528 7460
rect 4212 7420 4218 7432
rect 4522 7420 4528 7432
rect 4580 7420 4586 7472
rect 4617 7463 4675 7469
rect 4617 7429 4629 7463
rect 4663 7460 4675 7463
rect 7466 7460 7472 7472
rect 4663 7432 7472 7460
rect 4663 7429 4675 7432
rect 4617 7423 4675 7429
rect 7466 7420 7472 7432
rect 7524 7420 7530 7472
rect 9582 7420 9588 7472
rect 9640 7420 9646 7472
rect 9674 7420 9680 7472
rect 9732 7460 9738 7472
rect 9861 7463 9919 7469
rect 9861 7460 9873 7463
rect 9732 7432 9873 7460
rect 9732 7420 9738 7432
rect 9861 7429 9873 7432
rect 9907 7429 9919 7463
rect 9861 7423 9919 7429
rect 10060 7432 10732 7460
rect 4246 7392 4252 7404
rect 3568 7364 3765 7392
rect 3804 7364 4252 7392
rect 3568 7352 3574 7364
rect 3145 7327 3203 7333
rect 3145 7324 3157 7327
rect 3068 7296 3157 7324
rect 3145 7293 3157 7296
rect 3191 7293 3203 7327
rect 3737 7324 3765 7364
rect 4246 7352 4252 7364
rect 4304 7352 4310 7404
rect 4982 7352 4988 7404
rect 5040 7352 5046 7404
rect 5169 7395 5227 7401
rect 5169 7361 5181 7395
rect 5215 7392 5227 7395
rect 5442 7392 5448 7404
rect 5215 7364 5448 7392
rect 5215 7361 5227 7364
rect 5169 7355 5227 7361
rect 5442 7352 5448 7364
rect 5500 7352 5506 7404
rect 5721 7395 5779 7401
rect 5721 7361 5733 7395
rect 5767 7361 5779 7395
rect 5721 7355 5779 7361
rect 5000 7324 5028 7352
rect 5736 7324 5764 7355
rect 6362 7352 6368 7404
rect 6420 7352 6426 7404
rect 7558 7352 7564 7404
rect 7616 7392 7622 7404
rect 7745 7395 7803 7401
rect 7745 7392 7757 7395
rect 7616 7364 7757 7392
rect 7616 7352 7622 7364
rect 7745 7361 7757 7364
rect 7791 7361 7803 7395
rect 7745 7355 7803 7361
rect 8662 7352 8668 7404
rect 8720 7352 8726 7404
rect 8938 7352 8944 7404
rect 8996 7352 9002 7404
rect 9600 7392 9628 7420
rect 10060 7392 10088 7432
rect 9600 7364 10088 7392
rect 3737 7296 4844 7324
rect 5000 7296 5764 7324
rect 3145 7287 3203 7293
rect 4062 7216 4068 7268
rect 4120 7216 4126 7268
rect 4080 7188 4108 7216
rect 2746 7160 4108 7188
rect 4157 7191 4215 7197
rect 4157 7157 4169 7191
rect 4203 7188 4215 7191
rect 4338 7188 4344 7200
rect 4203 7160 4344 7188
rect 4203 7157 4215 7160
rect 4157 7151 4215 7157
rect 4338 7148 4344 7160
rect 4396 7148 4402 7200
rect 4706 7148 4712 7200
rect 4764 7148 4770 7200
rect 4816 7188 4844 7296
rect 6380 7256 6408 7352
rect 7926 7284 7932 7336
rect 7984 7284 7990 7336
rect 8294 7284 8300 7336
rect 8352 7324 8358 7336
rect 8389 7327 8447 7333
rect 8389 7324 8401 7327
rect 8352 7296 8401 7324
rect 8352 7284 8358 7296
rect 8389 7293 8401 7296
rect 8435 7293 8447 7327
rect 8389 7287 8447 7293
rect 8803 7327 8861 7333
rect 8803 7293 8815 7327
rect 8849 7324 8861 7327
rect 9600 7324 9628 7364
rect 10134 7352 10140 7404
rect 10192 7352 10198 7404
rect 10226 7352 10232 7404
rect 10284 7352 10290 7404
rect 10318 7352 10324 7404
rect 10376 7392 10382 7404
rect 10597 7395 10655 7401
rect 10597 7392 10609 7395
rect 10376 7364 10609 7392
rect 10376 7352 10382 7364
rect 10597 7361 10609 7364
rect 10643 7361 10655 7395
rect 10704 7392 10732 7432
rect 10778 7420 10784 7472
rect 10836 7460 10842 7472
rect 10965 7463 11023 7469
rect 10965 7460 10977 7463
rect 10836 7432 10977 7460
rect 10836 7420 10842 7432
rect 10965 7429 10977 7432
rect 11011 7429 11023 7463
rect 10965 7423 11023 7429
rect 11701 7463 11759 7469
rect 11701 7429 11713 7463
rect 11747 7460 11759 7463
rect 11790 7460 11796 7472
rect 11747 7432 11796 7460
rect 11747 7429 11759 7432
rect 11701 7423 11759 7429
rect 11790 7420 11796 7432
rect 11848 7420 11854 7472
rect 12066 7420 12072 7472
rect 12124 7420 12130 7472
rect 12158 7420 12164 7472
rect 12216 7460 12222 7472
rect 12342 7460 12348 7472
rect 12216 7432 12348 7460
rect 12216 7420 12222 7432
rect 12342 7420 12348 7432
rect 12400 7420 12406 7472
rect 12434 7420 12440 7472
rect 12492 7420 12498 7472
rect 12805 7463 12863 7469
rect 12805 7429 12817 7463
rect 12851 7460 12863 7463
rect 12986 7460 12992 7472
rect 12851 7432 12992 7460
rect 12851 7429 12863 7432
rect 12805 7423 12863 7429
rect 12986 7420 12992 7432
rect 13044 7460 13050 7472
rect 13044 7432 13216 7460
rect 13044 7420 13050 7432
rect 11977 7395 12035 7401
rect 10704 7364 11192 7392
rect 10597 7355 10655 7361
rect 8849 7296 9628 7324
rect 8849 7293 8861 7296
rect 8803 7287 8861 7293
rect 10042 7284 10048 7336
rect 10100 7284 10106 7336
rect 11164 7265 11192 7364
rect 11977 7361 11989 7395
rect 12023 7392 12035 7395
rect 13078 7392 13084 7404
rect 12023 7364 13084 7392
rect 12023 7361 12035 7364
rect 11977 7355 12035 7361
rect 13078 7352 13084 7364
rect 13136 7352 13142 7404
rect 11882 7284 11888 7336
rect 11940 7284 11946 7336
rect 11149 7259 11207 7265
rect 6380 7228 7696 7256
rect 5261 7191 5319 7197
rect 5261 7188 5273 7191
rect 4816 7160 5273 7188
rect 5261 7157 5273 7160
rect 5307 7157 5319 7191
rect 5261 7151 5319 7157
rect 6270 7148 6276 7200
rect 6328 7188 6334 7200
rect 7558 7188 7564 7200
rect 6328 7160 7564 7188
rect 6328 7148 6334 7160
rect 7558 7148 7564 7160
rect 7616 7148 7622 7200
rect 7668 7188 7696 7228
rect 11149 7225 11161 7259
rect 11195 7225 11207 7259
rect 13188 7256 13216 7432
rect 13338 7392 13366 7500
rect 13446 7488 13452 7540
rect 13504 7528 13510 7540
rect 16301 7531 16359 7537
rect 16301 7528 16313 7531
rect 13504 7500 16313 7528
rect 13504 7488 13510 7500
rect 16301 7497 16313 7500
rect 16347 7497 16359 7531
rect 16301 7491 16359 7497
rect 16574 7488 16580 7540
rect 16632 7528 16638 7540
rect 17770 7528 17776 7540
rect 16632 7500 17776 7528
rect 16632 7488 16638 7500
rect 17770 7488 17776 7500
rect 17828 7488 17834 7540
rect 20622 7488 20628 7540
rect 20680 7528 20686 7540
rect 21174 7528 21180 7540
rect 20680 7500 21180 7528
rect 20680 7488 20686 7500
rect 21174 7488 21180 7500
rect 21232 7528 21238 7540
rect 23937 7531 23995 7537
rect 23937 7528 23949 7531
rect 21232 7500 23949 7528
rect 21232 7488 21238 7500
rect 23937 7497 23949 7500
rect 23983 7497 23995 7531
rect 23937 7491 23995 7497
rect 24026 7488 24032 7540
rect 24084 7528 24090 7540
rect 24213 7531 24271 7537
rect 24213 7528 24225 7531
rect 24084 7500 24225 7528
rect 24084 7488 24090 7500
rect 24213 7497 24225 7500
rect 24259 7497 24271 7531
rect 24213 7491 24271 7497
rect 16390 7420 16396 7472
rect 16448 7460 16454 7472
rect 16448 7432 19932 7460
rect 16448 7420 16454 7432
rect 13338 7364 13768 7392
rect 13630 7256 13636 7268
rect 13188 7228 13636 7256
rect 11149 7219 11207 7225
rect 13630 7216 13636 7228
rect 13688 7216 13694 7268
rect 9585 7191 9643 7197
rect 9585 7188 9597 7191
rect 7668 7160 9597 7188
rect 9585 7157 9597 7160
rect 9631 7157 9643 7191
rect 9585 7151 9643 7157
rect 12989 7191 13047 7197
rect 12989 7157 13001 7191
rect 13035 7188 13047 7191
rect 13262 7188 13268 7200
rect 13035 7160 13268 7188
rect 13035 7157 13047 7160
rect 12989 7151 13047 7157
rect 13262 7148 13268 7160
rect 13320 7148 13326 7200
rect 13740 7188 13768 7364
rect 14274 7352 14280 7404
rect 14332 7392 14338 7404
rect 14645 7395 14703 7401
rect 14645 7392 14657 7395
rect 14332 7364 14657 7392
rect 14332 7352 14338 7364
rect 14645 7361 14657 7364
rect 14691 7361 14703 7395
rect 14645 7355 14703 7361
rect 15654 7352 15660 7404
rect 15712 7352 15718 7404
rect 16482 7352 16488 7404
rect 16540 7352 16546 7404
rect 16942 7352 16948 7404
rect 17000 7392 17006 7404
rect 17405 7395 17463 7401
rect 17405 7392 17417 7395
rect 17000 7364 17417 7392
rect 17000 7352 17006 7364
rect 17405 7361 17417 7364
rect 17451 7361 17463 7395
rect 17405 7355 17463 7361
rect 17957 7395 18015 7401
rect 17957 7361 17969 7395
rect 18003 7392 18015 7395
rect 18138 7392 18144 7404
rect 18003 7364 18144 7392
rect 18003 7361 18015 7364
rect 17957 7355 18015 7361
rect 18138 7352 18144 7364
rect 18196 7352 18202 7404
rect 19426 7352 19432 7404
rect 19484 7392 19490 7404
rect 19797 7395 19855 7401
rect 19797 7392 19809 7395
rect 19484 7364 19809 7392
rect 19484 7352 19490 7364
rect 19797 7361 19809 7364
rect 19843 7361 19855 7395
rect 19904 7392 19932 7432
rect 20346 7420 20352 7472
rect 20404 7460 20410 7472
rect 22094 7460 22100 7472
rect 20404 7432 22100 7460
rect 20404 7420 20410 7432
rect 22094 7420 22100 7432
rect 22152 7420 22158 7472
rect 23293 7404 23351 7405
rect 20070 7392 20076 7404
rect 19904 7364 20076 7392
rect 19797 7355 19855 7361
rect 20070 7352 20076 7364
rect 20128 7352 20134 7404
rect 20162 7352 20168 7404
rect 20220 7392 20226 7404
rect 23014 7392 23020 7404
rect 20220 7364 23020 7392
rect 20220 7352 20226 7364
rect 23014 7352 23020 7364
rect 23072 7352 23078 7404
rect 23290 7352 23296 7404
rect 23348 7396 23354 7404
rect 23348 7368 23389 7396
rect 23661 7395 23719 7401
rect 23348 7352 23354 7368
rect 23661 7361 23673 7395
rect 23707 7361 23719 7395
rect 23661 7355 23719 7361
rect 23753 7395 23811 7401
rect 23753 7361 23765 7395
rect 23799 7392 23811 7395
rect 23842 7392 23848 7404
rect 23799 7364 23848 7392
rect 23799 7361 23811 7364
rect 23753 7355 23811 7361
rect 14461 7327 14519 7333
rect 14461 7293 14473 7327
rect 14507 7324 14519 7327
rect 14826 7324 14832 7336
rect 14507 7296 14832 7324
rect 14507 7293 14519 7296
rect 14461 7287 14519 7293
rect 14826 7284 14832 7296
rect 14884 7284 14890 7336
rect 15010 7284 15016 7336
rect 15068 7324 15074 7336
rect 15381 7327 15439 7333
rect 15381 7324 15393 7327
rect 15068 7296 15393 7324
rect 15068 7284 15074 7296
rect 15381 7293 15393 7296
rect 15427 7293 15439 7327
rect 15381 7287 15439 7293
rect 15519 7327 15577 7333
rect 15519 7293 15531 7327
rect 15565 7324 15577 7327
rect 16022 7324 16028 7336
rect 15565 7296 16028 7324
rect 15565 7293 15577 7296
rect 15519 7287 15577 7293
rect 16022 7284 16028 7296
rect 16080 7324 16086 7336
rect 16500 7324 16528 7352
rect 16080 7296 16528 7324
rect 16080 7284 16086 7296
rect 17218 7284 17224 7336
rect 17276 7284 17282 7336
rect 20806 7284 20812 7336
rect 20864 7324 20870 7336
rect 21358 7324 21364 7336
rect 20864 7296 21364 7324
rect 20864 7284 20870 7296
rect 21358 7284 21364 7296
rect 21416 7284 21422 7336
rect 23676 7324 23704 7355
rect 23842 7352 23848 7364
rect 23900 7352 23906 7404
rect 24026 7352 24032 7404
rect 24084 7352 24090 7404
rect 25038 7352 25044 7404
rect 25096 7392 25102 7404
rect 25096 7364 25176 7392
rect 25096 7352 25102 7364
rect 24854 7324 24860 7336
rect 23676 7296 24860 7324
rect 24854 7284 24860 7296
rect 24912 7284 24918 7336
rect 15105 7259 15163 7265
rect 15105 7225 15117 7259
rect 15151 7256 15163 7259
rect 15194 7256 15200 7268
rect 15151 7228 15200 7256
rect 15151 7225 15163 7228
rect 15105 7219 15163 7225
rect 15194 7216 15200 7228
rect 15252 7216 15258 7268
rect 16206 7216 16212 7268
rect 16264 7256 16270 7268
rect 17865 7259 17923 7265
rect 17865 7256 17877 7259
rect 16264 7228 17877 7256
rect 16264 7216 16270 7228
rect 17865 7225 17877 7228
rect 17911 7225 17923 7259
rect 23477 7259 23535 7265
rect 23477 7256 23489 7259
rect 17865 7219 17923 7225
rect 20456 7228 23489 7256
rect 17126 7188 17132 7200
rect 13740 7160 17132 7188
rect 17126 7148 17132 7160
rect 17184 7148 17190 7200
rect 19886 7148 19892 7200
rect 19944 7188 19950 7200
rect 20456 7188 20484 7228
rect 23477 7225 23489 7228
rect 23523 7225 23535 7259
rect 23477 7219 23535 7225
rect 25148 7200 25176 7364
rect 19944 7160 20484 7188
rect 19944 7148 19950 7160
rect 20806 7148 20812 7200
rect 20864 7148 20870 7200
rect 23109 7191 23167 7197
rect 23109 7157 23121 7191
rect 23155 7188 23167 7191
rect 23566 7188 23572 7200
rect 23155 7160 23572 7188
rect 23155 7157 23167 7160
rect 23109 7151 23167 7157
rect 23566 7148 23572 7160
rect 23624 7148 23630 7200
rect 25130 7148 25136 7200
rect 25188 7148 25194 7200
rect 1104 7098 24564 7120
rect 1104 7046 3882 7098
rect 3934 7046 3946 7098
rect 3998 7046 4010 7098
rect 4062 7046 4074 7098
rect 4126 7046 4138 7098
rect 4190 7046 9747 7098
rect 9799 7046 9811 7098
rect 9863 7046 9875 7098
rect 9927 7046 9939 7098
rect 9991 7046 10003 7098
rect 10055 7046 15612 7098
rect 15664 7046 15676 7098
rect 15728 7046 15740 7098
rect 15792 7046 15804 7098
rect 15856 7046 15868 7098
rect 15920 7046 21477 7098
rect 21529 7046 21541 7098
rect 21593 7046 21605 7098
rect 21657 7046 21669 7098
rect 21721 7046 21733 7098
rect 21785 7046 24564 7098
rect 1104 7024 24564 7046
rect 1578 6944 1584 6996
rect 1636 6944 1642 6996
rect 1670 6944 1676 6996
rect 1728 6984 1734 6996
rect 7374 6984 7380 6996
rect 1728 6956 7380 6984
rect 1728 6944 1734 6956
rect 7374 6944 7380 6956
rect 7432 6944 7438 6996
rect 7466 6944 7472 6996
rect 7524 6944 7530 6996
rect 10226 6944 10232 6996
rect 10284 6984 10290 6996
rect 10873 6987 10931 6993
rect 10873 6984 10885 6987
rect 10284 6956 10885 6984
rect 10284 6944 10290 6956
rect 10873 6953 10885 6956
rect 10919 6953 10931 6987
rect 10873 6947 10931 6953
rect 12066 6944 12072 6996
rect 12124 6984 12130 6996
rect 12253 6987 12311 6993
rect 12253 6984 12265 6987
rect 12124 6956 12265 6984
rect 12124 6944 12130 6956
rect 12253 6953 12265 6956
rect 12299 6953 12311 6987
rect 12253 6947 12311 6953
rect 12434 6944 12440 6996
rect 12492 6984 12498 6996
rect 13354 6984 13360 6996
rect 12492 6956 13360 6984
rect 12492 6944 12498 6956
rect 13354 6944 13360 6956
rect 13412 6944 13418 6996
rect 13538 6944 13544 6996
rect 13596 6984 13602 6996
rect 13633 6987 13691 6993
rect 13633 6984 13645 6987
rect 13596 6956 13645 6984
rect 13596 6944 13602 6956
rect 13633 6953 13645 6956
rect 13679 6953 13691 6987
rect 13633 6947 13691 6953
rect 13740 6956 14872 6984
rect 7282 6876 7288 6928
rect 7340 6916 7346 6928
rect 9490 6916 9496 6928
rect 7340 6888 9496 6916
rect 7340 6876 7346 6888
rect 9490 6876 9496 6888
rect 9548 6876 9554 6928
rect 5626 6808 5632 6860
rect 5684 6808 5690 6860
rect 5813 6851 5871 6857
rect 5813 6817 5825 6851
rect 5859 6848 5871 6851
rect 5902 6848 5908 6860
rect 5859 6820 5908 6848
rect 5859 6817 5871 6820
rect 5813 6811 5871 6817
rect 5902 6808 5908 6820
rect 5960 6808 5966 6860
rect 6270 6808 6276 6860
rect 6328 6808 6334 6860
rect 6638 6808 6644 6860
rect 6696 6857 6702 6860
rect 6696 6851 6724 6857
rect 6712 6817 6724 6851
rect 6696 6811 6724 6817
rect 6825 6851 6883 6857
rect 6825 6817 6837 6851
rect 6871 6848 6883 6851
rect 7374 6848 7380 6860
rect 6871 6820 7380 6848
rect 6871 6817 6883 6820
rect 6825 6811 6883 6817
rect 6696 6808 6702 6811
rect 7374 6808 7380 6820
rect 7432 6808 7438 6860
rect 7926 6808 7932 6860
rect 7984 6848 7990 6860
rect 9766 6848 9772 6860
rect 7984 6820 9772 6848
rect 7984 6808 7990 6820
rect 9766 6808 9772 6820
rect 9824 6808 9830 6860
rect 11054 6808 11060 6860
rect 11112 6848 11118 6860
rect 11241 6851 11299 6857
rect 11241 6848 11253 6851
rect 11112 6820 11253 6848
rect 11112 6808 11118 6820
rect 11241 6817 11253 6820
rect 11287 6817 11299 6851
rect 11241 6811 11299 6817
rect 2590 6789 2596 6792
rect 2317 6783 2375 6789
rect 2317 6749 2329 6783
rect 2363 6749 2375 6783
rect 2317 6743 2375 6749
rect 2559 6783 2596 6789
rect 2559 6749 2571 6783
rect 2559 6743 2596 6749
rect 1486 6672 1492 6724
rect 1544 6672 1550 6724
rect 2332 6712 2360 6743
rect 2590 6740 2596 6743
rect 2648 6740 2654 6792
rect 4246 6740 4252 6792
rect 4304 6740 4310 6792
rect 4523 6783 4581 6789
rect 4523 6749 4535 6783
rect 4569 6780 4581 6783
rect 5534 6780 5540 6792
rect 4569 6752 5540 6780
rect 4569 6749 4581 6752
rect 4523 6743 4581 6749
rect 5534 6740 5540 6752
rect 5592 6740 5598 6792
rect 6546 6740 6552 6792
rect 6604 6740 6610 6792
rect 9306 6740 9312 6792
rect 9364 6780 9370 6792
rect 9861 6783 9919 6789
rect 9861 6780 9873 6783
rect 9364 6752 9873 6780
rect 9364 6740 9370 6752
rect 9861 6749 9873 6752
rect 9907 6749 9919 6783
rect 9861 6743 9919 6749
rect 10042 6740 10048 6792
rect 10100 6780 10106 6792
rect 10135 6783 10193 6789
rect 10135 6780 10147 6783
rect 10100 6752 10147 6780
rect 10100 6740 10106 6752
rect 10135 6749 10147 6752
rect 10181 6780 10193 6783
rect 10181 6752 10548 6780
rect 10181 6749 10193 6752
rect 10135 6743 10193 6749
rect 4264 6712 4292 6740
rect 2332 6684 4292 6712
rect 9214 6672 9220 6724
rect 9272 6712 9278 6724
rect 10226 6712 10232 6724
rect 9272 6684 10232 6712
rect 9272 6672 9278 6684
rect 10226 6672 10232 6684
rect 10284 6672 10290 6724
rect 10520 6712 10548 6752
rect 10594 6740 10600 6792
rect 10652 6780 10658 6792
rect 10652 6759 11542 6780
rect 10652 6753 11557 6759
rect 10652 6752 11511 6753
rect 10652 6740 10658 6752
rect 11330 6712 11336 6724
rect 10520 6684 11336 6712
rect 11330 6672 11336 6684
rect 11388 6672 11394 6724
rect 11499 6719 11511 6752
rect 11545 6719 11557 6753
rect 12066 6740 12072 6792
rect 12124 6740 12130 6792
rect 12342 6740 12348 6792
rect 12400 6780 12406 6792
rect 12621 6783 12679 6789
rect 12621 6780 12633 6783
rect 12400 6752 12633 6780
rect 12400 6740 12406 6752
rect 12621 6749 12633 6752
rect 12667 6749 12679 6783
rect 12621 6743 12679 6749
rect 12802 6740 12808 6792
rect 12860 6780 12866 6792
rect 12895 6783 12953 6789
rect 12895 6780 12907 6783
rect 12860 6752 12907 6780
rect 12860 6740 12866 6752
rect 12895 6749 12907 6752
rect 12941 6780 12953 6783
rect 13740 6780 13768 6956
rect 14844 6916 14872 6956
rect 15194 6944 15200 6996
rect 15252 6944 15258 6996
rect 16390 6944 16396 6996
rect 16448 6944 16454 6996
rect 16485 6987 16543 6993
rect 16485 6953 16497 6987
rect 16531 6984 16543 6987
rect 16942 6984 16948 6996
rect 16531 6956 16948 6984
rect 16531 6953 16543 6956
rect 16485 6947 16543 6953
rect 16942 6944 16948 6956
rect 17000 6944 17006 6996
rect 17126 6944 17132 6996
rect 17184 6984 17190 6996
rect 17184 6956 21496 6984
rect 17184 6944 17190 6956
rect 16408 6916 16436 6944
rect 14844 6888 16436 6916
rect 18230 6876 18236 6928
rect 18288 6916 18294 6928
rect 21468 6925 21496 6956
rect 23014 6944 23020 6996
rect 23072 6984 23078 6996
rect 23072 6956 23796 6984
rect 23072 6944 23078 6956
rect 18417 6919 18475 6925
rect 18417 6916 18429 6919
rect 18288 6888 18429 6916
rect 18288 6876 18294 6888
rect 18417 6885 18429 6888
rect 18463 6885 18475 6919
rect 18417 6879 18475 6885
rect 21453 6919 21511 6925
rect 21453 6885 21465 6919
rect 21499 6885 21511 6919
rect 21453 6879 21511 6885
rect 21818 6876 21824 6928
rect 21876 6916 21882 6928
rect 23768 6925 23796 6956
rect 23753 6919 23811 6925
rect 21876 6888 22048 6916
rect 21876 6876 21882 6888
rect 14185 6851 14243 6857
rect 14185 6848 14197 6851
rect 12941 6752 13768 6780
rect 14016 6820 14197 6848
rect 12941 6749 12953 6752
rect 12895 6743 12953 6749
rect 11499 6713 11557 6719
rect 12084 6712 12112 6740
rect 13906 6712 13912 6724
rect 12084 6684 13912 6712
rect 13906 6672 13912 6684
rect 13964 6712 13970 6724
rect 14016 6712 14044 6820
rect 14185 6817 14197 6820
rect 14231 6817 14243 6851
rect 20714 6848 20720 6860
rect 14185 6811 14243 6817
rect 18064 6820 20720 6848
rect 14090 6740 14096 6792
rect 14148 6780 14154 6792
rect 16393 6783 16451 6789
rect 14148 6753 14504 6780
rect 14148 6752 14455 6753
rect 14148 6740 14154 6752
rect 14443 6719 14455 6752
rect 14489 6722 14504 6753
rect 16393 6749 16405 6783
rect 16439 6780 16451 6783
rect 16853 6783 16911 6789
rect 16439 6752 16712 6780
rect 16439 6749 16451 6752
rect 16393 6743 16451 6749
rect 14489 6719 14501 6722
rect 14443 6713 14501 6719
rect 13964 6684 14044 6712
rect 13964 6672 13970 6684
rect 14642 6672 14648 6724
rect 14700 6672 14706 6724
rect 2222 6604 2228 6656
rect 2280 6644 2286 6656
rect 3234 6644 3240 6656
rect 2280 6616 3240 6644
rect 2280 6604 2286 6616
rect 3234 6604 3240 6616
rect 3292 6604 3298 6656
rect 3326 6604 3332 6656
rect 3384 6604 3390 6656
rect 5261 6647 5319 6653
rect 5261 6613 5273 6647
rect 5307 6644 5319 6647
rect 5626 6644 5632 6656
rect 5307 6616 5632 6644
rect 5307 6613 5319 6616
rect 5261 6607 5319 6613
rect 5626 6604 5632 6616
rect 5684 6604 5690 6656
rect 5718 6604 5724 6656
rect 5776 6644 5782 6656
rect 14660 6644 14688 6672
rect 16684 6653 16712 6752
rect 16853 6749 16865 6783
rect 16899 6749 16911 6783
rect 16853 6743 16911 6749
rect 16945 6783 17003 6789
rect 16945 6749 16957 6783
rect 16991 6780 17003 6783
rect 17770 6780 17776 6792
rect 16991 6752 17776 6780
rect 16991 6749 17003 6752
rect 16945 6743 17003 6749
rect 16868 6712 16896 6743
rect 17770 6740 17776 6752
rect 17828 6740 17834 6792
rect 17212 6715 17270 6721
rect 17212 6712 17224 6715
rect 16868 6684 17224 6712
rect 17212 6681 17224 6684
rect 17258 6712 17270 6715
rect 18064 6712 18092 6820
rect 20714 6808 20720 6820
rect 20772 6808 20778 6860
rect 20806 6808 20812 6860
rect 20864 6848 20870 6860
rect 21913 6851 21971 6857
rect 21913 6848 21925 6851
rect 20864 6820 21128 6848
rect 20864 6808 20870 6820
rect 18601 6783 18659 6789
rect 18601 6749 18613 6783
rect 18647 6749 18659 6783
rect 18601 6743 18659 6749
rect 18616 6712 18644 6743
rect 19242 6740 19248 6792
rect 19300 6740 19306 6792
rect 20533 6783 20591 6789
rect 20533 6749 20545 6783
rect 20579 6780 20591 6783
rect 20622 6780 20628 6792
rect 20579 6752 20628 6780
rect 20579 6749 20591 6752
rect 20533 6743 20591 6749
rect 20622 6740 20628 6752
rect 20680 6740 20686 6792
rect 20990 6740 20996 6792
rect 21048 6740 21054 6792
rect 17258 6684 18092 6712
rect 18340 6684 18644 6712
rect 21100 6712 21128 6820
rect 21560 6820 21925 6848
rect 21560 6789 21588 6820
rect 21913 6817 21925 6820
rect 21959 6817 21971 6851
rect 22020 6848 22048 6888
rect 23753 6885 23765 6919
rect 23799 6885 23811 6919
rect 23753 6879 23811 6885
rect 22020 6820 22784 6848
rect 21913 6811 21971 6817
rect 21545 6783 21603 6789
rect 21545 6749 21557 6783
rect 21591 6749 21603 6783
rect 21545 6743 21603 6749
rect 21821 6783 21879 6789
rect 21821 6749 21833 6783
rect 21867 6749 21879 6783
rect 21821 6743 21879 6749
rect 22005 6783 22063 6789
rect 22005 6749 22017 6783
rect 22051 6749 22063 6783
rect 22005 6743 22063 6749
rect 21836 6712 21864 6743
rect 21100 6684 21864 6712
rect 17258 6681 17270 6684
rect 17212 6675 17270 6681
rect 18340 6653 18368 6684
rect 5776 6616 14688 6644
rect 16669 6647 16727 6653
rect 5776 6604 5782 6616
rect 16669 6613 16681 6647
rect 16715 6613 16727 6647
rect 16669 6607 16727 6613
rect 18325 6647 18383 6653
rect 18325 6613 18337 6647
rect 18371 6613 18383 6647
rect 18325 6607 18383 6613
rect 19337 6647 19395 6653
rect 19337 6613 19349 6647
rect 19383 6644 19395 6647
rect 19610 6644 19616 6656
rect 19383 6616 19616 6644
rect 19383 6613 19395 6616
rect 19337 6607 19395 6613
rect 19610 6604 19616 6616
rect 19668 6604 19674 6656
rect 20349 6647 20407 6653
rect 20349 6613 20361 6647
rect 20395 6644 20407 6647
rect 20622 6644 20628 6656
rect 20395 6616 20628 6644
rect 20395 6613 20407 6616
rect 20349 6607 20407 6613
rect 20622 6604 20628 6616
rect 20680 6604 20686 6656
rect 22020 6644 22048 6743
rect 22278 6740 22284 6792
rect 22336 6740 22342 6792
rect 22554 6740 22560 6792
rect 22612 6740 22618 6792
rect 22756 6653 22784 6820
rect 23106 6740 23112 6792
rect 23164 6740 23170 6792
rect 23474 6740 23480 6792
rect 23532 6740 23538 6792
rect 23842 6740 23848 6792
rect 23900 6740 23906 6792
rect 22097 6647 22155 6653
rect 22097 6644 22109 6647
rect 22020 6616 22109 6644
rect 22097 6613 22109 6616
rect 22143 6613 22155 6647
rect 22097 6607 22155 6613
rect 22741 6647 22799 6653
rect 22741 6613 22753 6647
rect 22787 6613 22799 6647
rect 22741 6607 22799 6613
rect 1104 6554 24723 6576
rect 1104 6502 6814 6554
rect 6866 6502 6878 6554
rect 6930 6502 6942 6554
rect 6994 6502 7006 6554
rect 7058 6502 7070 6554
rect 7122 6502 12679 6554
rect 12731 6502 12743 6554
rect 12795 6502 12807 6554
rect 12859 6502 12871 6554
rect 12923 6502 12935 6554
rect 12987 6502 18544 6554
rect 18596 6502 18608 6554
rect 18660 6502 18672 6554
rect 18724 6502 18736 6554
rect 18788 6502 18800 6554
rect 18852 6502 24409 6554
rect 24461 6502 24473 6554
rect 24525 6502 24537 6554
rect 24589 6502 24601 6554
rect 24653 6502 24665 6554
rect 24717 6502 24723 6554
rect 1104 6480 24723 6502
rect 2130 6400 2136 6452
rect 2188 6440 2194 6452
rect 2409 6443 2467 6449
rect 2409 6440 2421 6443
rect 2188 6412 2421 6440
rect 2188 6400 2194 6412
rect 2409 6409 2421 6412
rect 2455 6409 2467 6443
rect 2774 6440 2780 6452
rect 2409 6403 2467 6409
rect 2746 6400 2780 6440
rect 2832 6400 2838 6452
rect 3234 6440 3240 6452
rect 2976 6412 3240 6440
rect 1671 6307 1729 6313
rect 1671 6273 1683 6307
rect 1717 6304 1729 6307
rect 2746 6304 2774 6400
rect 2976 6313 3004 6412
rect 3234 6400 3240 6412
rect 3292 6440 3298 6452
rect 5718 6440 5724 6452
rect 3292 6412 5724 6440
rect 3292 6400 3298 6412
rect 5718 6400 5724 6412
rect 5776 6400 5782 6452
rect 5905 6443 5963 6449
rect 5905 6409 5917 6443
rect 5951 6440 5963 6443
rect 6270 6440 6276 6452
rect 5951 6412 6276 6440
rect 5951 6409 5963 6412
rect 5905 6403 5963 6409
rect 6270 6400 6276 6412
rect 6328 6400 6334 6452
rect 10042 6440 10048 6452
rect 6840 6412 10048 6440
rect 5534 6332 5540 6384
rect 5592 6372 5598 6384
rect 6840 6372 6868 6412
rect 10042 6400 10048 6412
rect 10100 6400 10106 6452
rect 10612 6412 14136 6440
rect 9674 6372 9680 6384
rect 5592 6344 6868 6372
rect 6932 6344 9680 6372
rect 5592 6332 5598 6344
rect 6932 6343 6960 6344
rect 6899 6337 6960 6343
rect 1717 6276 2774 6304
rect 2961 6307 3019 6313
rect 1717 6273 1729 6276
rect 1671 6267 1729 6273
rect 2961 6273 2973 6307
rect 3007 6273 3019 6307
rect 2961 6267 3019 6273
rect 3786 6264 3792 6316
rect 3844 6313 3850 6316
rect 3844 6307 3872 6313
rect 3860 6273 3872 6307
rect 3844 6267 3872 6273
rect 5167 6307 5225 6313
rect 5167 6273 5179 6307
rect 5213 6304 5225 6307
rect 6899 6304 6911 6337
rect 5213 6303 6911 6304
rect 6945 6303 6960 6337
rect 9674 6332 9680 6344
rect 9732 6332 9738 6384
rect 9766 6332 9772 6384
rect 9824 6372 9830 6384
rect 10612 6372 10640 6412
rect 12342 6372 12348 6384
rect 9824 6344 10640 6372
rect 12268 6344 12348 6372
rect 9824 6332 9830 6344
rect 5213 6276 6960 6303
rect 5213 6273 5225 6276
rect 5167 6267 5225 6273
rect 3844 6264 3850 6267
rect 7466 6264 7472 6316
rect 7524 6304 7530 6316
rect 8295 6307 8353 6313
rect 8295 6304 8307 6307
rect 7524 6276 8307 6304
rect 7524 6264 7530 6276
rect 8295 6273 8307 6276
rect 8341 6304 8353 6307
rect 9122 6304 9128 6316
rect 8341 6276 9128 6304
rect 8341 6273 8353 6276
rect 8295 6267 8353 6273
rect 9122 6264 9128 6276
rect 9180 6264 9186 6316
rect 9306 6264 9312 6316
rect 9364 6304 9370 6316
rect 11422 6304 11428 6316
rect 9364 6276 11428 6304
rect 9364 6264 9370 6276
rect 11422 6264 11428 6276
rect 11480 6304 11486 6316
rect 12268 6304 12296 6344
rect 12342 6332 12348 6344
rect 12400 6372 12406 6384
rect 12400 6344 13216 6372
rect 12400 6332 12406 6344
rect 11480 6276 12296 6304
rect 11480 6264 11486 6276
rect 1394 6196 1400 6248
rect 1452 6196 1458 6248
rect 2777 6239 2835 6245
rect 2777 6205 2789 6239
rect 2823 6236 2835 6239
rect 2823 6208 3280 6236
rect 2823 6205 2835 6208
rect 2777 6199 2835 6205
rect 3252 6180 3280 6208
rect 3326 6196 3332 6248
rect 3384 6236 3390 6248
rect 3421 6239 3479 6245
rect 3421 6236 3433 6239
rect 3384 6208 3433 6236
rect 3384 6196 3390 6208
rect 3421 6205 3433 6208
rect 3467 6205 3479 6239
rect 3697 6239 3755 6245
rect 3697 6236 3709 6239
rect 3421 6199 3479 6205
rect 3528 6208 3709 6236
rect 3234 6128 3240 6180
rect 3292 6128 3298 6180
rect 1302 6060 1308 6112
rect 1360 6100 1366 6112
rect 2406 6100 2412 6112
rect 1360 6072 2412 6100
rect 1360 6060 1366 6072
rect 2406 6060 2412 6072
rect 2464 6100 2470 6112
rect 3528 6100 3556 6208
rect 3697 6205 3709 6208
rect 3743 6205 3755 6239
rect 3697 6199 3755 6205
rect 3973 6239 4031 6245
rect 3973 6205 3985 6239
rect 4019 6236 4031 6239
rect 4338 6236 4344 6248
rect 4019 6208 4344 6236
rect 4019 6205 4031 6208
rect 3973 6199 4031 6205
rect 4338 6196 4344 6208
rect 4396 6196 4402 6248
rect 4893 6239 4951 6245
rect 4893 6205 4905 6239
rect 4939 6205 4951 6239
rect 4893 6199 4951 6205
rect 4908 6168 4936 6199
rect 6178 6196 6184 6248
rect 6236 6236 6242 6248
rect 6641 6239 6699 6245
rect 6641 6236 6653 6239
rect 6236 6208 6653 6236
rect 6236 6196 6242 6208
rect 6641 6205 6653 6208
rect 6687 6205 6699 6239
rect 6641 6199 6699 6205
rect 8021 6239 8079 6245
rect 8021 6205 8033 6239
rect 8067 6205 8079 6239
rect 8021 6199 8079 6205
rect 4356 6140 4936 6168
rect 4356 6112 4384 6140
rect 2464 6072 3556 6100
rect 2464 6060 2470 6072
rect 4338 6060 4344 6112
rect 4396 6060 4402 6112
rect 4614 6060 4620 6112
rect 4672 6060 4678 6112
rect 4908 6100 4936 6140
rect 6362 6128 6368 6180
rect 6420 6128 6426 6180
rect 6380 6100 6408 6128
rect 4908 6072 6408 6100
rect 6656 6100 6684 6199
rect 8036 6168 8064 6199
rect 8938 6196 8944 6248
rect 8996 6236 9002 6248
rect 10594 6236 10600 6248
rect 8996 6208 10600 6236
rect 8996 6196 9002 6208
rect 10594 6196 10600 6208
rect 10652 6196 10658 6248
rect 13188 6245 13216 6344
rect 13722 6332 13728 6384
rect 13780 6332 13786 6384
rect 14108 6372 14136 6412
rect 14182 6400 14188 6452
rect 14240 6400 14246 6452
rect 17218 6400 17224 6452
rect 17276 6440 17282 6452
rect 17681 6443 17739 6449
rect 17681 6440 17693 6443
rect 17276 6412 17693 6440
rect 17276 6400 17282 6412
rect 17681 6409 17693 6412
rect 17727 6409 17739 6443
rect 17681 6403 17739 6409
rect 14108 6344 17632 6372
rect 13354 6264 13360 6316
rect 13412 6304 13418 6316
rect 13447 6307 13505 6313
rect 13447 6304 13459 6307
rect 13412 6276 13459 6304
rect 13412 6264 13418 6276
rect 13447 6273 13459 6276
rect 13493 6304 13505 6307
rect 13740 6304 13768 6332
rect 13493 6276 13860 6304
rect 13493 6273 13505 6276
rect 13447 6267 13505 6273
rect 13173 6239 13231 6245
rect 13173 6205 13185 6239
rect 13219 6205 13231 6239
rect 13832 6236 13860 6276
rect 15470 6264 15476 6316
rect 15528 6304 15534 6316
rect 16911 6307 16969 6313
rect 16911 6304 16923 6307
rect 15528 6276 16923 6304
rect 15528 6264 15534 6276
rect 16911 6273 16923 6276
rect 16957 6273 16969 6307
rect 16911 6267 16969 6273
rect 16298 6236 16304 6248
rect 13832 6208 16304 6236
rect 13173 6199 13231 6205
rect 12066 6168 12072 6180
rect 7300 6140 8064 6168
rect 7300 6100 7328 6140
rect 6656 6072 7328 6100
rect 7650 6060 7656 6112
rect 7708 6060 7714 6112
rect 8036 6100 8064 6140
rect 8680 6140 12072 6168
rect 8680 6100 8708 6140
rect 12066 6128 12072 6140
rect 12124 6128 12130 6180
rect 8036 6072 8708 6100
rect 8846 6060 8852 6112
rect 8904 6100 8910 6112
rect 9033 6103 9091 6109
rect 9033 6100 9045 6103
rect 8904 6072 9045 6100
rect 8904 6060 8910 6072
rect 9033 6069 9045 6072
rect 9079 6069 9091 6103
rect 9033 6063 9091 6069
rect 9122 6060 9128 6112
rect 9180 6100 9186 6112
rect 11606 6100 11612 6112
rect 9180 6072 11612 6100
rect 9180 6060 9186 6072
rect 11606 6060 11612 6072
rect 11664 6060 11670 6112
rect 13188 6100 13216 6199
rect 16298 6196 16304 6208
rect 16356 6196 16362 6248
rect 16666 6196 16672 6248
rect 16724 6196 16730 6248
rect 15470 6128 15476 6180
rect 15528 6168 15534 6180
rect 16022 6168 16028 6180
rect 15528 6140 16028 6168
rect 15528 6128 15534 6140
rect 16022 6128 16028 6140
rect 16080 6128 16086 6180
rect 16206 6128 16212 6180
rect 16264 6168 16270 6180
rect 17604 6168 17632 6344
rect 17696 6304 17724 6403
rect 18138 6400 18144 6452
rect 18196 6400 18202 6452
rect 18230 6400 18236 6452
rect 18288 6400 18294 6452
rect 18325 6443 18383 6449
rect 18325 6409 18337 6443
rect 18371 6440 18383 6443
rect 19242 6440 19248 6452
rect 18371 6412 19248 6440
rect 18371 6409 18383 6412
rect 18325 6403 18383 6409
rect 19242 6400 19248 6412
rect 19300 6400 19306 6452
rect 19334 6400 19340 6452
rect 19392 6440 19398 6452
rect 19978 6440 19984 6452
rect 19392 6412 19984 6440
rect 19392 6400 19398 6412
rect 19978 6400 19984 6412
rect 20036 6400 20042 6452
rect 20349 6443 20407 6449
rect 20349 6409 20361 6443
rect 20395 6409 20407 6443
rect 20349 6403 20407 6409
rect 18248 6313 18276 6400
rect 18868 6375 18926 6381
rect 18868 6372 18880 6375
rect 18524 6344 18880 6372
rect 18524 6313 18552 6344
rect 18868 6341 18880 6344
rect 18914 6372 18926 6375
rect 19886 6372 19892 6384
rect 18914 6344 19892 6372
rect 18914 6341 18926 6344
rect 18868 6335 18926 6341
rect 19886 6332 19892 6344
rect 19944 6332 19950 6384
rect 18049 6307 18107 6313
rect 18049 6304 18061 6307
rect 17696 6276 18061 6304
rect 18049 6273 18061 6276
rect 18095 6273 18107 6307
rect 18049 6267 18107 6273
rect 18233 6307 18291 6313
rect 18233 6273 18245 6307
rect 18279 6273 18291 6307
rect 18233 6267 18291 6273
rect 18509 6307 18567 6313
rect 18509 6273 18521 6307
rect 18555 6273 18567 6307
rect 18509 6267 18567 6273
rect 19426 6264 19432 6316
rect 19484 6304 19490 6316
rect 20073 6307 20131 6313
rect 20073 6304 20085 6307
rect 19484 6276 20085 6304
rect 19484 6264 19490 6276
rect 20073 6273 20085 6276
rect 20119 6273 20131 6307
rect 20073 6267 20131 6273
rect 20257 6307 20315 6313
rect 20257 6273 20269 6307
rect 20303 6304 20315 6307
rect 20364 6304 20392 6403
rect 20622 6400 20628 6452
rect 20680 6400 20686 6452
rect 20990 6400 20996 6452
rect 21048 6400 21054 6452
rect 21082 6400 21088 6452
rect 21140 6440 21146 6452
rect 21821 6443 21879 6449
rect 21821 6440 21833 6443
rect 21140 6412 21833 6440
rect 21140 6400 21146 6412
rect 21821 6409 21833 6412
rect 21867 6409 21879 6443
rect 23014 6440 23020 6452
rect 21821 6403 21879 6409
rect 22066 6412 23020 6440
rect 20303 6276 20392 6304
rect 20533 6307 20591 6313
rect 20303 6273 20315 6276
rect 20257 6267 20315 6273
rect 20533 6273 20545 6307
rect 20579 6273 20591 6307
rect 20640 6304 20668 6400
rect 22066 6372 22094 6412
rect 23014 6400 23020 6412
rect 23072 6400 23078 6452
rect 23106 6400 23112 6452
rect 23164 6400 23170 6452
rect 23474 6400 23480 6452
rect 23532 6440 23538 6452
rect 23569 6443 23627 6449
rect 23569 6440 23581 6443
rect 23532 6412 23581 6440
rect 23532 6400 23538 6412
rect 23569 6409 23581 6412
rect 23615 6409 23627 6443
rect 23569 6403 23627 6409
rect 23658 6400 23664 6452
rect 23716 6400 23722 6452
rect 23842 6400 23848 6452
rect 23900 6400 23906 6452
rect 24213 6443 24271 6449
rect 24213 6409 24225 6443
rect 24259 6440 24271 6443
rect 24302 6440 24308 6452
rect 24259 6412 24308 6440
rect 24259 6409 24271 6412
rect 24213 6403 24271 6409
rect 24302 6400 24308 6412
rect 24360 6400 24366 6452
rect 21100 6344 22094 6372
rect 20901 6307 20959 6313
rect 20901 6304 20913 6307
rect 20640 6276 20913 6304
rect 20533 6267 20591 6273
rect 20901 6273 20913 6276
rect 20947 6273 20959 6307
rect 20901 6267 20959 6273
rect 17770 6196 17776 6248
rect 17828 6236 17834 6248
rect 18598 6236 18604 6248
rect 17828 6208 18604 6236
rect 17828 6196 17834 6208
rect 18598 6196 18604 6208
rect 18656 6196 18662 6248
rect 20548 6236 20576 6267
rect 19996 6208 20576 6236
rect 18506 6168 18512 6180
rect 16264 6140 16528 6168
rect 17604 6140 18512 6168
rect 16264 6128 16270 6140
rect 16390 6100 16396 6112
rect 13188 6072 16396 6100
rect 16390 6060 16396 6072
rect 16448 6060 16454 6112
rect 16500 6100 16528 6140
rect 18506 6128 18512 6140
rect 18564 6128 18570 6180
rect 19996 6177 20024 6208
rect 19981 6171 20039 6177
rect 19981 6137 19993 6171
rect 20027 6137 20039 6171
rect 21100 6168 21128 6344
rect 21177 6307 21235 6313
rect 21177 6273 21189 6307
rect 21223 6304 21235 6307
rect 21266 6304 21272 6316
rect 21223 6276 21272 6304
rect 21223 6273 21235 6276
rect 21177 6267 21235 6273
rect 21266 6264 21272 6276
rect 21324 6264 21330 6316
rect 21358 6264 21364 6316
rect 21416 6264 21422 6316
rect 21453 6307 21511 6313
rect 21453 6273 21465 6307
rect 21499 6273 21511 6307
rect 21453 6267 21511 6273
rect 21468 6236 21496 6267
rect 21818 6264 21824 6316
rect 21876 6304 21882 6316
rect 22005 6307 22063 6313
rect 22005 6304 22017 6307
rect 21876 6276 22017 6304
rect 21876 6264 21882 6276
rect 22005 6273 22017 6276
rect 22051 6273 22063 6307
rect 22005 6267 22063 6273
rect 22094 6264 22100 6316
rect 22152 6264 22158 6316
rect 22371 6307 22429 6313
rect 22371 6273 22383 6307
rect 22417 6304 22429 6307
rect 22830 6304 22836 6316
rect 22417 6276 22836 6304
rect 22417 6273 22429 6276
rect 22371 6267 22429 6273
rect 22830 6264 22836 6276
rect 22888 6264 22894 6316
rect 19981 6131 20039 6137
rect 20548 6140 21128 6168
rect 21192 6208 21496 6236
rect 23124 6236 23152 6400
rect 23676 6372 23704 6400
rect 23676 6344 23980 6372
rect 23477 6307 23535 6313
rect 23477 6273 23489 6307
rect 23523 6304 23535 6307
rect 23566 6304 23572 6316
rect 23523 6276 23572 6304
rect 23523 6273 23535 6276
rect 23477 6267 23535 6273
rect 23566 6264 23572 6276
rect 23624 6264 23630 6316
rect 23952 6313 23980 6344
rect 23753 6307 23811 6313
rect 23753 6273 23765 6307
rect 23799 6273 23811 6307
rect 23753 6267 23811 6273
rect 23937 6307 23995 6313
rect 23937 6273 23949 6307
rect 23983 6273 23995 6307
rect 23937 6267 23995 6273
rect 23768 6236 23796 6267
rect 24026 6264 24032 6316
rect 24084 6264 24090 6316
rect 23124 6208 23796 6236
rect 20548 6112 20576 6140
rect 19518 6100 19524 6112
rect 16500 6072 19524 6100
rect 19518 6060 19524 6072
rect 19576 6060 19582 6112
rect 20162 6060 20168 6112
rect 20220 6060 20226 6112
rect 20530 6060 20536 6112
rect 20588 6060 20594 6112
rect 20714 6060 20720 6112
rect 20772 6100 20778 6112
rect 21192 6100 21220 6208
rect 21269 6171 21327 6177
rect 21269 6137 21281 6171
rect 21315 6168 21327 6171
rect 21315 6140 22094 6168
rect 21315 6137 21327 6140
rect 21269 6131 21327 6137
rect 20772 6072 21220 6100
rect 20772 6060 20778 6072
rect 21542 6060 21548 6112
rect 21600 6100 21606 6112
rect 21637 6103 21695 6109
rect 21637 6100 21649 6103
rect 21600 6072 21649 6100
rect 21600 6060 21606 6072
rect 21637 6069 21649 6072
rect 21683 6069 21695 6103
rect 22066 6100 22094 6140
rect 22370 6100 22376 6112
rect 22066 6072 22376 6100
rect 21637 6063 21695 6069
rect 22370 6060 22376 6072
rect 22428 6060 22434 6112
rect 22554 6060 22560 6112
rect 22612 6100 22618 6112
rect 23106 6100 23112 6112
rect 22612 6072 23112 6100
rect 22612 6060 22618 6072
rect 23106 6060 23112 6072
rect 23164 6060 23170 6112
rect 1104 6010 24564 6032
rect 1104 5958 3882 6010
rect 3934 5958 3946 6010
rect 3998 5958 4010 6010
rect 4062 5958 4074 6010
rect 4126 5958 4138 6010
rect 4190 5958 9747 6010
rect 9799 5958 9811 6010
rect 9863 5958 9875 6010
rect 9927 5958 9939 6010
rect 9991 5958 10003 6010
rect 10055 5958 15612 6010
rect 15664 5958 15676 6010
rect 15728 5958 15740 6010
rect 15792 5958 15804 6010
rect 15856 5958 15868 6010
rect 15920 5958 21477 6010
rect 21529 5958 21541 6010
rect 21593 5958 21605 6010
rect 21657 5958 21669 6010
rect 21721 5958 21733 6010
rect 21785 5958 24564 6010
rect 1104 5936 24564 5958
rect 3329 5899 3387 5905
rect 3329 5865 3341 5899
rect 3375 5896 3387 5899
rect 4430 5896 4436 5908
rect 3375 5868 4436 5896
rect 3375 5865 3387 5868
rect 3329 5859 3387 5865
rect 4430 5856 4436 5868
rect 4488 5856 4494 5908
rect 4890 5856 4896 5908
rect 4948 5856 4954 5908
rect 6454 5896 6460 5908
rect 5184 5868 6460 5896
rect 1670 5720 1676 5772
rect 1728 5720 1734 5772
rect 2130 5720 2136 5772
rect 2188 5720 2194 5772
rect 2406 5720 2412 5772
rect 2464 5720 2470 5772
rect 2547 5763 2605 5769
rect 2547 5729 2559 5763
rect 2593 5760 2605 5763
rect 3786 5760 3792 5772
rect 2593 5732 3792 5760
rect 2593 5729 2605 5732
rect 2547 5723 2605 5729
rect 3786 5720 3792 5732
rect 3844 5720 3850 5772
rect 4617 5763 4675 5769
rect 4617 5729 4629 5763
rect 4663 5760 4675 5763
rect 4908 5760 4936 5856
rect 4663 5732 4936 5760
rect 4663 5729 4675 5732
rect 4617 5723 4675 5729
rect 5074 5720 5080 5772
rect 5132 5720 5138 5772
rect 5184 5760 5212 5868
rect 6454 5856 6460 5868
rect 6512 5896 6518 5908
rect 6512 5868 7052 5896
rect 6512 5856 6518 5868
rect 7024 5828 7052 5868
rect 7374 5856 7380 5908
rect 7432 5856 7438 5908
rect 7650 5856 7656 5908
rect 7708 5896 7714 5908
rect 8294 5896 8300 5908
rect 7708 5868 8300 5896
rect 7708 5856 7714 5868
rect 8294 5856 8300 5868
rect 8352 5856 8358 5908
rect 8754 5856 8760 5908
rect 8812 5896 8818 5908
rect 9306 5896 9312 5908
rect 8812 5868 9312 5896
rect 8812 5856 8818 5868
rect 9306 5856 9312 5868
rect 9364 5856 9370 5908
rect 11054 5896 11060 5908
rect 9968 5868 11060 5896
rect 7024 5800 8708 5828
rect 8680 5772 8708 5800
rect 5470 5763 5528 5769
rect 5470 5760 5482 5763
rect 5184 5732 5482 5760
rect 5470 5729 5482 5732
rect 5516 5729 5528 5763
rect 5470 5723 5528 5729
rect 5626 5720 5632 5772
rect 5684 5720 5690 5772
rect 7466 5720 7472 5772
rect 7524 5720 7530 5772
rect 8662 5720 8668 5772
rect 8720 5720 8726 5772
rect 1489 5695 1547 5701
rect 1489 5661 1501 5695
rect 1535 5661 1547 5695
rect 1489 5655 1547 5661
rect 1504 5556 1532 5655
rect 2682 5652 2688 5704
rect 2740 5652 2746 5704
rect 3418 5652 3424 5704
rect 3476 5652 3482 5704
rect 4062 5652 4068 5704
rect 4120 5652 4126 5704
rect 4433 5695 4491 5701
rect 4433 5661 4445 5695
rect 4479 5692 4491 5695
rect 4522 5692 4528 5704
rect 4479 5664 4528 5692
rect 4479 5661 4491 5664
rect 4433 5655 4491 5661
rect 4522 5652 4528 5664
rect 4580 5652 4586 5704
rect 5350 5652 5356 5704
rect 5408 5652 5414 5704
rect 6362 5652 6368 5704
rect 6420 5652 6426 5704
rect 6639 5695 6697 5701
rect 6639 5661 6651 5695
rect 6685 5692 6697 5695
rect 7484 5692 7512 5720
rect 6685 5664 7512 5692
rect 6685 5661 6697 5664
rect 6639 5655 6697 5661
rect 9306 5652 9312 5704
rect 9364 5692 9370 5704
rect 9968 5701 9996 5868
rect 11054 5856 11060 5868
rect 11112 5856 11118 5908
rect 11606 5856 11612 5908
rect 11664 5896 11670 5908
rect 22094 5896 22100 5908
rect 11664 5868 22100 5896
rect 11664 5856 11670 5868
rect 22094 5856 22100 5868
rect 22152 5856 22158 5908
rect 22189 5899 22247 5905
rect 22189 5865 22201 5899
rect 22235 5896 22247 5899
rect 22278 5896 22284 5908
rect 22235 5868 22284 5896
rect 22235 5865 22247 5868
rect 22189 5859 22247 5865
rect 22278 5856 22284 5868
rect 22336 5856 22342 5908
rect 23934 5856 23940 5908
rect 23992 5896 23998 5908
rect 24213 5899 24271 5905
rect 24213 5896 24225 5899
rect 23992 5868 24225 5896
rect 23992 5856 23998 5868
rect 24213 5865 24225 5868
rect 24259 5865 24271 5899
rect 24213 5859 24271 5865
rect 13906 5788 13912 5840
rect 13964 5828 13970 5840
rect 14734 5828 14740 5840
rect 13964 5800 14740 5828
rect 13964 5788 13970 5800
rect 14734 5788 14740 5800
rect 14792 5788 14798 5840
rect 15028 5800 15240 5828
rect 15028 5772 15056 5800
rect 13814 5720 13820 5772
rect 13872 5760 13878 5772
rect 14274 5760 14280 5772
rect 13872 5732 14280 5760
rect 13872 5720 13878 5732
rect 14274 5720 14280 5732
rect 14332 5760 14338 5772
rect 14645 5763 14703 5769
rect 14645 5760 14657 5763
rect 14332 5732 14657 5760
rect 14332 5720 14338 5732
rect 14645 5729 14657 5732
rect 14691 5729 14703 5763
rect 14645 5723 14703 5729
rect 15010 5720 15016 5772
rect 15068 5720 15074 5772
rect 15102 5720 15108 5772
rect 15160 5720 15166 5772
rect 15212 5760 15240 5800
rect 18506 5788 18512 5840
rect 18564 5828 18570 5840
rect 20073 5831 20131 5837
rect 20073 5828 20085 5831
rect 18564 5800 20085 5828
rect 18564 5788 18570 5800
rect 20073 5797 20085 5800
rect 20119 5797 20131 5831
rect 20073 5791 20131 5797
rect 22462 5788 22468 5840
rect 22520 5788 22526 5840
rect 22557 5831 22615 5837
rect 22557 5797 22569 5831
rect 22603 5828 22615 5831
rect 22646 5828 22652 5840
rect 22603 5800 22652 5828
rect 22603 5797 22615 5800
rect 22557 5791 22615 5797
rect 22646 5788 22652 5800
rect 22704 5788 22710 5840
rect 15381 5763 15439 5769
rect 15381 5760 15393 5763
rect 15212 5732 15393 5760
rect 15381 5729 15393 5732
rect 15427 5729 15439 5763
rect 15381 5723 15439 5729
rect 15470 5720 15476 5772
rect 15528 5769 15534 5772
rect 15528 5763 15556 5769
rect 15544 5729 15556 5763
rect 15528 5723 15556 5729
rect 15657 5763 15715 5769
rect 15657 5729 15669 5763
rect 15703 5760 15715 5763
rect 16022 5760 16028 5772
rect 15703 5732 16028 5760
rect 15703 5729 15715 5732
rect 15657 5723 15715 5729
rect 15528 5720 15534 5723
rect 16022 5720 16028 5732
rect 16080 5720 16086 5772
rect 16666 5720 16672 5772
rect 16724 5760 16730 5772
rect 17402 5760 17408 5772
rect 16724 5732 17408 5760
rect 16724 5720 16730 5732
rect 17402 5720 17408 5732
rect 17460 5760 17466 5772
rect 17770 5760 17776 5772
rect 17460 5732 17776 5760
rect 17460 5720 17466 5732
rect 17770 5720 17776 5732
rect 17828 5720 17834 5772
rect 18598 5720 18604 5772
rect 18656 5760 18662 5772
rect 20809 5763 20867 5769
rect 20809 5760 20821 5763
rect 18656 5732 20821 5760
rect 18656 5720 18662 5732
rect 20456 5704 20484 5732
rect 20809 5729 20821 5732
rect 20855 5729 20867 5763
rect 22186 5760 22192 5772
rect 20809 5723 20867 5729
rect 21836 5732 22192 5760
rect 9953 5695 10011 5701
rect 9953 5692 9965 5695
rect 9364 5664 9965 5692
rect 9364 5652 9370 5664
rect 9953 5661 9965 5664
rect 9999 5661 10011 5695
rect 9953 5655 10011 5661
rect 10227 5695 10285 5701
rect 10227 5661 10239 5695
rect 10273 5692 10285 5695
rect 11698 5692 11704 5704
rect 10273 5664 11704 5692
rect 10273 5661 10285 5664
rect 10227 5655 10285 5661
rect 11698 5652 11704 5664
rect 11756 5652 11762 5704
rect 14461 5695 14519 5701
rect 14461 5661 14473 5695
rect 14507 5692 14519 5695
rect 14826 5692 14832 5704
rect 14507 5664 14832 5692
rect 14507 5661 14519 5664
rect 14461 5655 14519 5661
rect 14826 5652 14832 5664
rect 14884 5652 14890 5704
rect 16298 5652 16304 5704
rect 16356 5692 16362 5704
rect 18015 5695 18073 5701
rect 18015 5692 18027 5695
rect 16356 5664 18027 5692
rect 16356 5652 16362 5664
rect 18015 5661 18027 5664
rect 18061 5661 18073 5695
rect 18015 5655 18073 5661
rect 19242 5652 19248 5704
rect 19300 5652 19306 5704
rect 19426 5652 19432 5704
rect 19484 5652 19490 5704
rect 19610 5652 19616 5704
rect 19668 5652 19674 5704
rect 20162 5652 20168 5704
rect 20220 5652 20226 5704
rect 20438 5652 20444 5704
rect 20496 5652 20502 5704
rect 20530 5652 20536 5704
rect 20588 5652 20594 5704
rect 20717 5695 20775 5701
rect 20717 5661 20729 5695
rect 20763 5661 20775 5695
rect 20824 5692 20852 5723
rect 21836 5692 21864 5732
rect 22186 5720 22192 5732
rect 22244 5760 22250 5772
rect 22833 5763 22891 5769
rect 22833 5760 22845 5763
rect 22244 5732 22845 5760
rect 22244 5720 22250 5732
rect 22833 5729 22845 5732
rect 22879 5729 22891 5763
rect 22833 5723 22891 5729
rect 20824 5664 21864 5692
rect 20717 5655 20775 5661
rect 4080 5624 4108 5652
rect 3528 5596 4108 5624
rect 8036 5596 12434 5624
rect 3528 5556 3556 5596
rect 8036 5568 8064 5596
rect 1504 5528 3556 5556
rect 3605 5559 3663 5565
rect 3605 5525 3617 5559
rect 3651 5556 3663 5559
rect 4982 5556 4988 5568
rect 3651 5528 4988 5556
rect 3651 5525 3663 5528
rect 3605 5519 3663 5525
rect 4982 5516 4988 5528
rect 5040 5516 5046 5568
rect 6270 5516 6276 5568
rect 6328 5516 6334 5568
rect 8018 5516 8024 5568
rect 8076 5516 8082 5568
rect 8570 5516 8576 5568
rect 8628 5556 8634 5568
rect 9398 5556 9404 5568
rect 8628 5528 9404 5556
rect 8628 5516 8634 5528
rect 9398 5516 9404 5528
rect 9456 5516 9462 5568
rect 10134 5516 10140 5568
rect 10192 5556 10198 5568
rect 10965 5559 11023 5565
rect 10965 5556 10977 5559
rect 10192 5528 10977 5556
rect 10192 5516 10198 5528
rect 10965 5525 10977 5528
rect 11011 5525 11023 5559
rect 12406 5556 12434 5596
rect 17678 5584 17684 5636
rect 17736 5624 17742 5636
rect 19260 5624 19288 5652
rect 17736 5596 19288 5624
rect 17736 5584 17742 5596
rect 16301 5559 16359 5565
rect 16301 5556 16313 5559
rect 12406 5528 16313 5556
rect 10965 5519 11023 5525
rect 16301 5525 16313 5528
rect 16347 5525 16359 5559
rect 16301 5519 16359 5525
rect 17770 5516 17776 5568
rect 17828 5556 17834 5568
rect 18046 5556 18052 5568
rect 17828 5528 18052 5556
rect 17828 5516 17834 5528
rect 18046 5516 18052 5528
rect 18104 5516 18110 5568
rect 18785 5559 18843 5565
rect 18785 5525 18797 5559
rect 18831 5556 18843 5559
rect 19444 5556 19472 5652
rect 19518 5584 19524 5636
rect 19576 5624 19582 5636
rect 20732 5624 20760 5655
rect 22278 5652 22284 5704
rect 22336 5652 22342 5704
rect 22738 5652 22744 5704
rect 22796 5652 22802 5704
rect 19576 5596 20760 5624
rect 21076 5627 21134 5633
rect 19576 5584 19582 5596
rect 21076 5593 21088 5627
rect 21122 5624 21134 5627
rect 21174 5624 21180 5636
rect 21122 5596 21180 5624
rect 21122 5593 21134 5596
rect 21076 5587 21134 5593
rect 21174 5584 21180 5596
rect 21232 5584 21238 5636
rect 23100 5627 23158 5633
rect 23100 5593 23112 5627
rect 23146 5624 23158 5627
rect 23290 5624 23296 5636
rect 23146 5596 23296 5624
rect 23146 5593 23158 5596
rect 23100 5587 23158 5593
rect 23290 5584 23296 5596
rect 23348 5624 23354 5636
rect 23658 5624 23664 5636
rect 23348 5596 23664 5624
rect 23348 5584 23354 5596
rect 23658 5584 23664 5596
rect 23716 5584 23722 5636
rect 18831 5528 19472 5556
rect 18831 5525 18843 5528
rect 18785 5519 18843 5525
rect 19978 5516 19984 5568
rect 20036 5556 20042 5568
rect 20530 5556 20536 5568
rect 20036 5528 20536 5556
rect 20036 5516 20042 5528
rect 20530 5516 20536 5528
rect 20588 5516 20594 5568
rect 20717 5559 20775 5565
rect 20717 5525 20729 5559
rect 20763 5556 20775 5559
rect 23474 5556 23480 5568
rect 20763 5528 23480 5556
rect 20763 5525 20775 5528
rect 20717 5519 20775 5525
rect 23474 5516 23480 5528
rect 23532 5516 23538 5568
rect 1104 5466 24723 5488
rect 1104 5414 6814 5466
rect 6866 5414 6878 5466
rect 6930 5414 6942 5466
rect 6994 5414 7006 5466
rect 7058 5414 7070 5466
rect 7122 5414 12679 5466
rect 12731 5414 12743 5466
rect 12795 5414 12807 5466
rect 12859 5414 12871 5466
rect 12923 5414 12935 5466
rect 12987 5414 18544 5466
rect 18596 5414 18608 5466
rect 18660 5414 18672 5466
rect 18724 5414 18736 5466
rect 18788 5414 18800 5466
rect 18852 5414 24409 5466
rect 24461 5414 24473 5466
rect 24525 5414 24537 5466
rect 24589 5414 24601 5466
rect 24653 5414 24665 5466
rect 24717 5414 24723 5466
rect 1104 5392 24723 5414
rect 2409 5355 2467 5361
rect 2409 5321 2421 5355
rect 2455 5352 2467 5355
rect 2682 5352 2688 5364
rect 2455 5324 2688 5352
rect 2455 5321 2467 5324
rect 2409 5315 2467 5321
rect 2682 5312 2688 5324
rect 2740 5312 2746 5364
rect 3234 5312 3240 5364
rect 3292 5312 3298 5364
rect 3510 5312 3516 5364
rect 3568 5352 3574 5364
rect 3789 5355 3847 5361
rect 3789 5352 3801 5355
rect 3568 5324 3801 5352
rect 3568 5312 3574 5324
rect 3789 5321 3801 5324
rect 3835 5321 3847 5355
rect 3789 5315 3847 5321
rect 5074 5312 5080 5364
rect 5132 5352 5138 5364
rect 5169 5355 5227 5361
rect 5169 5352 5181 5355
rect 5132 5324 5181 5352
rect 5132 5312 5138 5324
rect 5169 5321 5181 5324
rect 5215 5321 5227 5355
rect 5169 5315 5227 5321
rect 6546 5312 6552 5364
rect 6604 5352 6610 5364
rect 8570 5352 8576 5364
rect 6604 5324 8576 5352
rect 6604 5312 6610 5324
rect 8570 5312 8576 5324
rect 8628 5312 8634 5364
rect 9122 5312 9128 5364
rect 9180 5352 9186 5364
rect 9674 5352 9680 5364
rect 9180 5324 9680 5352
rect 9180 5312 9186 5324
rect 9674 5312 9680 5324
rect 9732 5352 9738 5364
rect 9769 5355 9827 5361
rect 9769 5352 9781 5355
rect 9732 5324 9781 5352
rect 9732 5312 9738 5324
rect 9769 5321 9781 5324
rect 9815 5321 9827 5355
rect 9769 5315 9827 5321
rect 10318 5312 10324 5364
rect 10376 5352 10382 5364
rect 10376 5324 10548 5352
rect 10376 5312 10382 5324
rect 1670 5255 1676 5296
rect 1655 5249 1676 5255
rect 1394 5176 1400 5228
rect 1452 5176 1458 5228
rect 1655 5215 1667 5249
rect 1728 5244 1734 5296
rect 3145 5287 3203 5293
rect 3145 5253 3157 5287
rect 3191 5284 3203 5287
rect 6270 5284 6276 5296
rect 3191 5256 6276 5284
rect 3191 5253 3203 5256
rect 3145 5247 3203 5253
rect 6270 5244 6276 5256
rect 6328 5244 6334 5296
rect 9398 5244 9404 5296
rect 9456 5284 9462 5296
rect 10520 5293 10548 5324
rect 15194 5312 15200 5364
rect 15252 5352 15258 5364
rect 15749 5355 15807 5361
rect 15749 5352 15761 5355
rect 15252 5324 15761 5352
rect 15252 5312 15258 5324
rect 15749 5321 15761 5324
rect 15795 5321 15807 5355
rect 19334 5352 19340 5364
rect 15749 5315 15807 5321
rect 19306 5312 19340 5352
rect 19392 5312 19398 5364
rect 20441 5355 20499 5361
rect 20441 5321 20453 5355
rect 20487 5321 20499 5355
rect 20441 5315 20499 5321
rect 10505 5287 10563 5293
rect 9456 5256 10364 5284
rect 9456 5244 9462 5256
rect 1701 5218 1716 5244
rect 2777 5219 2835 5225
rect 1701 5215 1713 5218
rect 1655 5209 1713 5215
rect 2777 5185 2789 5219
rect 2823 5185 2835 5219
rect 2777 5179 2835 5185
rect 3697 5219 3755 5225
rect 3697 5185 3709 5219
rect 3743 5185 3755 5219
rect 3697 5179 3755 5185
rect 1210 4972 1216 5024
rect 1268 5012 1274 5024
rect 2792 5012 2820 5179
rect 3712 5080 3740 5179
rect 4154 5176 4160 5228
rect 4212 5176 4218 5228
rect 4431 5219 4489 5225
rect 4431 5185 4443 5219
rect 4477 5216 4489 5219
rect 6730 5216 6736 5228
rect 4477 5188 6736 5216
rect 4477 5185 4489 5188
rect 4431 5179 4489 5185
rect 6730 5176 6736 5188
rect 6788 5176 6794 5228
rect 7653 5219 7711 5225
rect 7653 5185 7665 5219
rect 7699 5216 7711 5219
rect 7699 5188 7972 5216
rect 7699 5185 7711 5188
rect 7653 5179 7711 5185
rect 5902 5108 5908 5160
rect 5960 5148 5966 5160
rect 7837 5151 7895 5157
rect 7837 5148 7849 5151
rect 5960 5120 7849 5148
rect 5960 5108 5966 5120
rect 7837 5117 7849 5120
rect 7883 5117 7895 5151
rect 7944 5148 7972 5188
rect 8570 5176 8576 5228
rect 8628 5176 8634 5228
rect 8846 5176 8852 5228
rect 8904 5176 8910 5228
rect 9490 5176 9496 5228
rect 9548 5176 9554 5228
rect 9674 5176 9680 5228
rect 9732 5216 9738 5228
rect 9950 5216 9956 5228
rect 9732 5188 9956 5216
rect 9732 5176 9738 5188
rect 9950 5176 9956 5188
rect 10008 5216 10014 5228
rect 10045 5219 10103 5225
rect 10045 5216 10057 5219
rect 10008 5188 10057 5216
rect 10008 5176 10014 5188
rect 10045 5185 10057 5188
rect 10091 5185 10103 5219
rect 10045 5179 10103 5185
rect 10134 5176 10140 5228
rect 10192 5176 10198 5228
rect 10336 5216 10364 5256
rect 10505 5253 10517 5287
rect 10551 5253 10563 5287
rect 10505 5247 10563 5253
rect 10778 5244 10784 5296
rect 10836 5284 10842 5296
rect 10873 5287 10931 5293
rect 10873 5284 10885 5287
rect 10836 5256 10885 5284
rect 10836 5244 10842 5256
rect 10873 5253 10885 5256
rect 10919 5253 10931 5287
rect 10873 5247 10931 5253
rect 15102 5244 15108 5296
rect 15160 5284 15166 5296
rect 19306 5284 19334 5312
rect 15160 5256 19334 5284
rect 20456 5284 20484 5315
rect 20898 5312 20904 5364
rect 20956 5352 20962 5364
rect 21085 5355 21143 5361
rect 21085 5352 21097 5355
rect 20956 5324 21097 5352
rect 20956 5312 20962 5324
rect 21085 5321 21097 5324
rect 21131 5321 21143 5355
rect 21085 5315 21143 5321
rect 21637 5355 21695 5361
rect 21637 5321 21649 5355
rect 21683 5352 21695 5355
rect 21683 5324 22692 5352
rect 21683 5321 21695 5324
rect 21637 5315 21695 5321
rect 20456 5256 21864 5284
rect 15160 5244 15166 5256
rect 10336 5188 10916 5216
rect 8202 5148 8208 5160
rect 7944 5120 8208 5148
rect 7837 5111 7895 5117
rect 8202 5108 8208 5120
rect 8260 5108 8266 5160
rect 8294 5108 8300 5160
rect 8352 5108 8358 5160
rect 8662 5108 8668 5160
rect 8720 5157 8726 5160
rect 8720 5151 8769 5157
rect 8720 5117 8723 5151
rect 8757 5117 8769 5151
rect 8720 5111 8769 5117
rect 8720 5108 8726 5111
rect 10226 5108 10232 5160
rect 10284 5108 10290 5160
rect 3712 5052 4292 5080
rect 1268 4984 2820 5012
rect 2961 5015 3019 5021
rect 1268 4972 1274 4984
rect 2961 4981 2973 5015
rect 3007 5012 3019 5015
rect 3510 5012 3516 5024
rect 3007 4984 3516 5012
rect 3007 4981 3019 4984
rect 2961 4975 3019 4981
rect 3510 4972 3516 4984
rect 3568 4972 3574 5024
rect 4264 5012 4292 5052
rect 5534 5040 5540 5092
rect 5592 5080 5598 5092
rect 10888 5080 10916 5188
rect 12526 5176 12532 5228
rect 12584 5216 12590 5228
rect 12805 5219 12863 5225
rect 12805 5216 12817 5219
rect 12584 5188 12817 5216
rect 12584 5176 12590 5188
rect 12805 5185 12817 5188
rect 12851 5185 12863 5219
rect 12805 5179 12863 5185
rect 13998 5176 14004 5228
rect 14056 5176 14062 5228
rect 14642 5176 14648 5228
rect 14700 5176 14706 5228
rect 14734 5176 14740 5228
rect 14792 5176 14798 5228
rect 14918 5176 14924 5228
rect 14976 5216 14982 5228
rect 15011 5219 15069 5225
rect 15011 5216 15023 5219
rect 14976 5188 15023 5216
rect 14976 5176 14982 5188
rect 15011 5185 15023 5188
rect 15057 5216 15069 5219
rect 19242 5216 19248 5228
rect 15057 5188 19248 5216
rect 15057 5185 15069 5188
rect 15011 5179 15069 5185
rect 19242 5176 19248 5188
rect 19300 5176 19306 5228
rect 19337 5219 19395 5225
rect 19337 5185 19349 5219
rect 19383 5185 19395 5219
rect 19337 5179 19395 5185
rect 19424 5220 19482 5225
rect 19518 5220 19524 5238
rect 19424 5219 19524 5220
rect 19424 5185 19436 5219
rect 19470 5192 19524 5219
rect 19470 5185 19482 5192
rect 19518 5186 19524 5192
rect 19576 5186 19582 5238
rect 19671 5229 19729 5235
rect 19671 5195 19683 5229
rect 19717 5226 19729 5229
rect 19717 5216 19748 5226
rect 19794 5216 19800 5228
rect 19717 5195 19800 5216
rect 19671 5189 19800 5195
rect 19720 5188 19800 5189
rect 19424 5179 19482 5185
rect 12434 5108 12440 5160
rect 12492 5148 12498 5160
rect 12989 5151 13047 5157
rect 12989 5148 13001 5151
rect 12492 5120 13001 5148
rect 12492 5108 12498 5120
rect 12989 5117 13001 5120
rect 13035 5148 13047 5151
rect 13078 5148 13084 5160
rect 13035 5120 13084 5148
rect 13035 5117 13047 5120
rect 12989 5111 13047 5117
rect 13078 5108 13084 5120
rect 13136 5108 13142 5160
rect 13722 5108 13728 5160
rect 13780 5108 13786 5160
rect 13863 5151 13921 5157
rect 13863 5117 13875 5151
rect 13909 5148 13921 5151
rect 14660 5148 14688 5176
rect 19352 5148 19380 5179
rect 19794 5176 19800 5188
rect 19852 5176 19858 5228
rect 20898 5176 20904 5228
rect 20956 5176 20962 5228
rect 20990 5176 20996 5228
rect 21048 5216 21054 5228
rect 21468 5225 21496 5256
rect 21836 5225 21864 5256
rect 21361 5219 21419 5225
rect 21361 5216 21373 5219
rect 21048 5188 21373 5216
rect 21048 5176 21054 5188
rect 21361 5185 21373 5188
rect 21407 5185 21419 5219
rect 21361 5179 21419 5185
rect 21453 5219 21511 5225
rect 21453 5185 21465 5219
rect 21499 5185 21511 5219
rect 21453 5179 21511 5185
rect 21637 5219 21695 5225
rect 21637 5185 21649 5219
rect 21683 5185 21695 5219
rect 21637 5179 21695 5185
rect 21821 5219 21879 5225
rect 21821 5185 21833 5219
rect 21867 5185 21879 5219
rect 21821 5179 21879 5185
rect 13909 5120 14688 5148
rect 19306 5120 19380 5148
rect 13909 5117 13921 5120
rect 13863 5111 13921 5117
rect 12618 5080 12624 5092
rect 5592 5052 8432 5080
rect 10888 5052 12624 5080
rect 5592 5040 5598 5052
rect 8018 5012 8024 5024
rect 4264 4984 8024 5012
rect 8018 4972 8024 4984
rect 8076 4972 8082 5024
rect 8404 5012 8432 5052
rect 12618 5040 12624 5052
rect 12676 5040 12682 5092
rect 13446 5040 13452 5092
rect 13504 5040 13510 5092
rect 9398 5012 9404 5024
rect 8404 4984 9404 5012
rect 9398 4972 9404 4984
rect 9456 4972 9462 5024
rect 10962 4972 10968 5024
rect 11020 5012 11026 5024
rect 11057 5015 11115 5021
rect 11057 5012 11069 5015
rect 11020 4984 11069 5012
rect 11020 4972 11026 4984
rect 11057 4981 11069 4984
rect 11103 4981 11115 5015
rect 11057 4975 11115 4981
rect 11790 4972 11796 5024
rect 11848 5012 11854 5024
rect 14645 5015 14703 5021
rect 14645 5012 14657 5015
rect 11848 4984 14657 5012
rect 11848 4972 11854 4984
rect 14645 4981 14657 4984
rect 14691 4981 14703 5015
rect 14645 4975 14703 4981
rect 19150 4972 19156 5024
rect 19208 4972 19214 5024
rect 19306 5012 19334 5120
rect 20162 5108 20168 5160
rect 20220 5148 20226 5160
rect 21652 5148 21680 5179
rect 21910 5176 21916 5228
rect 21968 5216 21974 5228
rect 22664 5225 22692 5324
rect 23845 5287 23903 5293
rect 23845 5253 23857 5287
rect 23891 5284 23903 5287
rect 24118 5284 24124 5296
rect 23891 5256 24124 5284
rect 23891 5253 23903 5256
rect 23845 5247 23903 5253
rect 24118 5244 24124 5256
rect 24176 5244 24182 5296
rect 22189 5219 22247 5225
rect 22189 5216 22201 5219
rect 21968 5188 22201 5216
rect 21968 5176 21974 5188
rect 22189 5185 22201 5188
rect 22235 5185 22247 5219
rect 22189 5179 22247 5185
rect 22649 5219 22707 5225
rect 22649 5185 22661 5219
rect 22695 5185 22707 5219
rect 22649 5179 22707 5185
rect 23014 5176 23020 5228
rect 23072 5176 23078 5228
rect 20220 5120 21680 5148
rect 20220 5108 20226 5120
rect 20254 5040 20260 5092
rect 20312 5080 20318 5092
rect 21358 5080 21364 5092
rect 20312 5052 21364 5080
rect 20312 5040 20318 5052
rect 21358 5040 21364 5052
rect 21416 5040 21422 5092
rect 22094 5040 22100 5092
rect 22152 5080 22158 5092
rect 22649 5083 22707 5089
rect 22649 5080 22661 5083
rect 22152 5052 22661 5080
rect 22152 5040 22158 5052
rect 22649 5049 22661 5052
rect 22695 5049 22707 5083
rect 22649 5043 22707 5049
rect 20346 5012 20352 5024
rect 19306 4984 20352 5012
rect 20346 4972 20352 4984
rect 20404 4972 20410 5024
rect 21174 4972 21180 5024
rect 21232 4972 21238 5024
rect 22002 4972 22008 5024
rect 22060 5012 22066 5024
rect 23382 5012 23388 5024
rect 22060 4984 23388 5012
rect 22060 4972 22066 4984
rect 23382 4972 23388 4984
rect 23440 4972 23446 5024
rect 1104 4922 24564 4944
rect 1104 4870 3882 4922
rect 3934 4870 3946 4922
rect 3998 4870 4010 4922
rect 4062 4870 4074 4922
rect 4126 4870 4138 4922
rect 4190 4870 9747 4922
rect 9799 4870 9811 4922
rect 9863 4870 9875 4922
rect 9927 4870 9939 4922
rect 9991 4870 10003 4922
rect 10055 4870 15612 4922
rect 15664 4870 15676 4922
rect 15728 4870 15740 4922
rect 15792 4870 15804 4922
rect 15856 4870 15868 4922
rect 15920 4870 21477 4922
rect 21529 4870 21541 4922
rect 21593 4870 21605 4922
rect 21657 4870 21669 4922
rect 21721 4870 21733 4922
rect 21785 4870 24564 4922
rect 1104 4848 24564 4870
rect 1302 4768 1308 4820
rect 1360 4808 1366 4820
rect 3237 4811 3295 4817
rect 3237 4808 3249 4811
rect 1360 4780 3249 4808
rect 1360 4768 1366 4780
rect 3237 4777 3249 4780
rect 3283 4777 3295 4811
rect 3237 4771 3295 4777
rect 3694 4768 3700 4820
rect 3752 4808 3758 4820
rect 4525 4811 4583 4817
rect 4525 4808 4537 4811
rect 3752 4780 4537 4808
rect 3752 4768 3758 4780
rect 4525 4777 4537 4780
rect 4571 4777 4583 4811
rect 4525 4771 4583 4777
rect 5074 4768 5080 4820
rect 5132 4768 5138 4820
rect 5534 4768 5540 4820
rect 5592 4768 5598 4820
rect 6362 4808 6368 4820
rect 5920 4780 6368 4808
rect 2130 4700 2136 4752
rect 2188 4740 2194 4752
rect 2409 4743 2467 4749
rect 2409 4740 2421 4743
rect 2188 4712 2421 4740
rect 2188 4700 2194 4712
rect 2409 4709 2421 4712
rect 2455 4709 2467 4743
rect 2409 4703 2467 4709
rect 2590 4700 2596 4752
rect 2648 4740 2654 4752
rect 4065 4743 4123 4749
rect 4065 4740 4077 4743
rect 2648 4712 4077 4740
rect 2648 4700 2654 4712
rect 4065 4709 4077 4712
rect 4111 4709 4123 4743
rect 4065 4703 4123 4709
rect 4430 4700 4436 4752
rect 4488 4740 4494 4752
rect 4488 4712 5764 4740
rect 4488 4700 4494 4712
rect 1394 4632 1400 4684
rect 1452 4632 1458 4684
rect 3142 4632 3148 4684
rect 3200 4672 3206 4684
rect 3200 4644 5304 4672
rect 3200 4632 3206 4644
rect 1670 4604 1676 4616
rect 1631 4576 1676 4604
rect 1670 4564 1676 4576
rect 1728 4564 1734 4616
rect 2590 4564 2596 4616
rect 2648 4604 2654 4616
rect 2777 4607 2835 4613
rect 2777 4604 2789 4607
rect 2648 4576 2789 4604
rect 2648 4564 2654 4576
rect 2777 4573 2789 4576
rect 2823 4573 2835 4607
rect 2777 4567 2835 4573
rect 3881 4607 3939 4613
rect 3881 4573 3893 4607
rect 3927 4604 3939 4607
rect 4614 4604 4620 4616
rect 3927 4576 4620 4604
rect 3927 4573 3939 4576
rect 3881 4567 3939 4573
rect 4614 4564 4620 4576
rect 4672 4564 4678 4616
rect 4893 4607 4951 4613
rect 4893 4573 4905 4607
rect 4939 4604 4951 4607
rect 5074 4604 5080 4616
rect 4939 4576 5080 4604
rect 4939 4573 4951 4576
rect 4893 4567 4951 4573
rect 5074 4564 5080 4576
rect 5132 4564 5138 4616
rect 5276 4613 5304 4644
rect 5736 4613 5764 4712
rect 5920 4681 5948 4780
rect 6362 4768 6368 4780
rect 6420 4808 6426 4820
rect 6420 4780 6592 4808
rect 6420 4768 6426 4780
rect 6564 4740 6592 4780
rect 7098 4768 7104 4820
rect 7156 4808 7162 4820
rect 10137 4811 10195 4817
rect 7156 4780 10088 4808
rect 7156 4768 7162 4780
rect 6564 4712 7328 4740
rect 5905 4675 5963 4681
rect 5905 4641 5917 4675
rect 5951 4641 5963 4675
rect 5905 4635 5963 4641
rect 7300 4616 7328 4712
rect 8294 4700 8300 4752
rect 8352 4700 8358 4752
rect 8662 4700 8668 4752
rect 8720 4740 8726 4752
rect 10060 4740 10088 4780
rect 10137 4777 10149 4811
rect 10183 4808 10195 4811
rect 10226 4808 10232 4820
rect 10183 4780 10232 4808
rect 10183 4777 10195 4780
rect 10137 4771 10195 4777
rect 10226 4768 10232 4780
rect 10284 4768 10290 4820
rect 12618 4768 12624 4820
rect 12676 4808 12682 4820
rect 15194 4808 15200 4820
rect 12676 4780 15200 4808
rect 12676 4768 12682 4780
rect 15194 4768 15200 4780
rect 15252 4768 15258 4820
rect 15749 4811 15807 4817
rect 15749 4777 15761 4811
rect 15795 4808 15807 4811
rect 16022 4808 16028 4820
rect 15795 4780 16028 4808
rect 15795 4777 15807 4780
rect 15749 4771 15807 4777
rect 16022 4768 16028 4780
rect 16080 4768 16086 4820
rect 19150 4768 19156 4820
rect 19208 4768 19214 4820
rect 19337 4811 19395 4817
rect 19337 4777 19349 4811
rect 19383 4808 19395 4811
rect 20162 4808 20168 4820
rect 19383 4780 20168 4808
rect 19383 4777 19395 4780
rect 19337 4771 19395 4777
rect 20162 4768 20168 4780
rect 20220 4768 20226 4820
rect 20257 4811 20315 4817
rect 20257 4777 20269 4811
rect 20303 4808 20315 4811
rect 21910 4808 21916 4820
rect 20303 4780 21916 4808
rect 20303 4777 20315 4780
rect 20257 4771 20315 4777
rect 21910 4768 21916 4780
rect 21968 4768 21974 4820
rect 24121 4811 24179 4817
rect 24121 4777 24133 4811
rect 24167 4808 24179 4811
rect 25498 4808 25504 4820
rect 24167 4780 25504 4808
rect 24167 4777 24179 4780
rect 24121 4771 24179 4777
rect 25498 4768 25504 4780
rect 25556 4768 25562 4820
rect 11238 4740 11244 4752
rect 8720 4712 9076 4740
rect 10060 4712 11244 4740
rect 8720 4700 8726 4712
rect 5261 4607 5319 4613
rect 5261 4573 5273 4607
rect 5307 4573 5319 4607
rect 5261 4567 5319 4573
rect 5721 4607 5779 4613
rect 5721 4573 5733 4607
rect 5767 4573 5779 4607
rect 5721 4567 5779 4573
rect 6179 4607 6237 4613
rect 6179 4573 6191 4607
rect 6225 4604 6237 4607
rect 7098 4604 7104 4616
rect 6225 4576 7104 4604
rect 6225 4573 6237 4576
rect 6179 4567 6237 4573
rect 7098 4564 7104 4576
rect 7156 4564 7162 4616
rect 7282 4564 7288 4616
rect 7340 4564 7346 4616
rect 7559 4607 7617 4613
rect 7559 4573 7571 4607
rect 7605 4604 7617 4607
rect 8018 4604 8024 4616
rect 7605 4576 8024 4604
rect 7605 4573 7617 4576
rect 7559 4567 7617 4573
rect 8018 4564 8024 4576
rect 8076 4564 8082 4616
rect 3145 4539 3203 4545
rect 3145 4505 3157 4539
rect 3191 4536 3203 4539
rect 4433 4539 4491 4545
rect 3191 4508 4384 4536
rect 3191 4505 3203 4508
rect 3145 4499 3203 4505
rect 842 4428 848 4480
rect 900 4468 906 4480
rect 2961 4471 3019 4477
rect 2961 4468 2973 4471
rect 900 4440 2973 4468
rect 900 4428 906 4440
rect 2961 4437 2973 4440
rect 3007 4437 3019 4471
rect 2961 4431 3019 4437
rect 3694 4428 3700 4480
rect 3752 4468 3758 4480
rect 4246 4468 4252 4480
rect 3752 4440 4252 4468
rect 3752 4428 3758 4440
rect 4246 4428 4252 4440
rect 4304 4428 4310 4480
rect 4356 4468 4384 4508
rect 4433 4505 4445 4539
rect 4479 4536 4491 4539
rect 4798 4536 4804 4548
rect 4479 4508 4804 4536
rect 4479 4505 4491 4508
rect 4433 4499 4491 4505
rect 4798 4496 4804 4508
rect 4856 4496 4862 4548
rect 8938 4536 8944 4548
rect 5000 4508 8944 4536
rect 5000 4468 5028 4508
rect 8938 4496 8944 4508
rect 8996 4496 9002 4548
rect 9048 4536 9076 4712
rect 11238 4700 11244 4712
rect 11296 4700 11302 4752
rect 11882 4632 11888 4684
rect 11940 4632 11946 4684
rect 14734 4632 14740 4684
rect 14792 4632 14798 4684
rect 18966 4672 18972 4684
rect 18800 4644 18972 4672
rect 9125 4607 9183 4613
rect 9125 4573 9137 4607
rect 9171 4604 9183 4607
rect 9306 4604 9312 4616
rect 9171 4576 9312 4604
rect 9171 4573 9183 4576
rect 9125 4567 9183 4573
rect 9306 4564 9312 4576
rect 9364 4564 9370 4616
rect 9399 4607 9457 4613
rect 9399 4573 9411 4607
rect 9445 4604 9457 4607
rect 11422 4604 11428 4616
rect 9445 4576 11428 4604
rect 9445 4573 9457 4576
rect 9399 4567 9457 4573
rect 11422 4564 11428 4576
rect 11480 4564 11486 4616
rect 11606 4564 11612 4616
rect 11664 4564 11670 4616
rect 11701 4607 11759 4613
rect 11701 4573 11713 4607
rect 11747 4604 11759 4607
rect 12526 4604 12532 4616
rect 11747 4576 12532 4604
rect 11747 4573 11759 4576
rect 11701 4567 11759 4573
rect 12526 4564 12532 4576
rect 12584 4564 12590 4616
rect 15011 4607 15069 4613
rect 15011 4573 15023 4607
rect 15057 4604 15069 4607
rect 15102 4604 15108 4616
rect 15057 4576 15108 4604
rect 15057 4573 15069 4576
rect 15011 4567 15069 4573
rect 15102 4564 15108 4576
rect 15160 4564 15166 4616
rect 17221 4607 17279 4613
rect 17221 4573 17233 4607
rect 17267 4573 17279 4607
rect 17221 4567 17279 4573
rect 17495 4607 17553 4613
rect 17495 4573 17507 4607
rect 17541 4604 17553 4607
rect 17586 4604 17592 4616
rect 17541 4576 17592 4604
rect 17541 4573 17553 4576
rect 17495 4567 17553 4573
rect 10962 4536 10968 4548
rect 9048 4508 10968 4536
rect 10962 4496 10968 4508
rect 11020 4496 11026 4548
rect 11054 4496 11060 4548
rect 11112 4536 11118 4548
rect 12069 4539 12127 4545
rect 12069 4536 12081 4539
rect 11112 4508 12081 4536
rect 11112 4496 11118 4508
rect 12069 4505 12081 4508
rect 12115 4505 12127 4539
rect 17236 4536 17264 4567
rect 17586 4564 17592 4576
rect 17644 4564 17650 4616
rect 18230 4564 18236 4616
rect 18288 4564 18294 4616
rect 18800 4613 18828 4644
rect 18966 4632 18972 4644
rect 19024 4632 19030 4684
rect 19168 4672 19196 4768
rect 19613 4743 19671 4749
rect 19613 4709 19625 4743
rect 19659 4740 19671 4743
rect 19659 4712 20300 4740
rect 19659 4709 19671 4712
rect 19613 4703 19671 4709
rect 20272 4684 20300 4712
rect 19168 4644 20208 4672
rect 18785 4607 18843 4613
rect 18785 4573 18797 4607
rect 18831 4573 18843 4607
rect 18785 4567 18843 4573
rect 18877 4607 18935 4613
rect 18877 4573 18889 4607
rect 18923 4604 18935 4607
rect 19521 4607 19579 4613
rect 18923 4576 19472 4604
rect 18923 4573 18935 4576
rect 18877 4567 18935 4573
rect 18248 4536 18276 4564
rect 17236 4508 18276 4536
rect 12069 4499 12127 4505
rect 4356 4440 5028 4468
rect 5442 4428 5448 4480
rect 5500 4428 5506 4480
rect 6917 4471 6975 4477
rect 6917 4437 6929 4471
rect 6963 4468 6975 4471
rect 7374 4468 7380 4480
rect 6963 4440 7380 4468
rect 6963 4437 6975 4440
rect 6917 4431 6975 4437
rect 7374 4428 7380 4440
rect 7432 4428 7438 4480
rect 7466 4428 7472 4480
rect 7524 4468 7530 4480
rect 10778 4468 10784 4480
rect 7524 4440 10784 4468
rect 7524 4428 7530 4440
rect 10778 4428 10784 4440
rect 10836 4428 10842 4480
rect 11330 4428 11336 4480
rect 11388 4428 11394 4480
rect 11422 4428 11428 4480
rect 11480 4468 11486 4480
rect 12437 4471 12495 4477
rect 12437 4468 12449 4471
rect 11480 4440 12449 4468
rect 11480 4428 11486 4440
rect 12437 4437 12449 4440
rect 12483 4437 12495 4471
rect 12437 4431 12495 4437
rect 17770 4428 17776 4480
rect 17828 4468 17834 4480
rect 18233 4471 18291 4477
rect 18233 4468 18245 4471
rect 17828 4440 18245 4468
rect 17828 4428 17834 4440
rect 18233 4437 18245 4440
rect 18279 4437 18291 4471
rect 18233 4431 18291 4437
rect 18414 4428 18420 4480
rect 18472 4468 18478 4480
rect 18601 4471 18659 4477
rect 18601 4468 18613 4471
rect 18472 4440 18613 4468
rect 18472 4428 18478 4440
rect 18601 4437 18613 4440
rect 18647 4437 18659 4471
rect 18601 4431 18659 4437
rect 18969 4471 19027 4477
rect 18969 4437 18981 4471
rect 19015 4468 19027 4471
rect 19334 4468 19340 4480
rect 19015 4440 19340 4468
rect 19015 4437 19027 4440
rect 18969 4431 19027 4437
rect 19334 4428 19340 4440
rect 19392 4428 19398 4480
rect 19444 4468 19472 4576
rect 19521 4573 19533 4607
rect 19567 4573 19579 4607
rect 19521 4567 19579 4573
rect 19536 4536 19564 4567
rect 19794 4564 19800 4616
rect 19852 4564 19858 4616
rect 20070 4564 20076 4616
rect 20128 4564 20134 4616
rect 20180 4613 20208 4644
rect 20254 4632 20260 4684
rect 20312 4632 20318 4684
rect 20346 4632 20352 4684
rect 20404 4672 20410 4684
rect 20404 4644 20576 4672
rect 20404 4632 20410 4644
rect 20165 4607 20223 4613
rect 20165 4573 20177 4607
rect 20211 4573 20223 4607
rect 20165 4567 20223 4573
rect 20438 4564 20444 4616
rect 20496 4564 20502 4616
rect 20548 4536 20576 4644
rect 22186 4632 22192 4684
rect 22244 4632 22250 4684
rect 23201 4675 23259 4681
rect 23201 4672 23213 4675
rect 22296 4644 23213 4672
rect 21910 4564 21916 4616
rect 21968 4564 21974 4616
rect 22094 4564 22100 4616
rect 22152 4604 22158 4616
rect 22296 4604 22324 4644
rect 23201 4641 23213 4644
rect 23247 4641 23259 4675
rect 23201 4635 23259 4641
rect 22152 4576 22324 4604
rect 22152 4564 22158 4576
rect 22646 4564 22652 4616
rect 22704 4564 22710 4616
rect 22830 4564 22836 4616
rect 22888 4564 22894 4616
rect 20708 4539 20766 4545
rect 20708 4536 20720 4539
rect 19536 4508 20392 4536
rect 20548 4508 20720 4536
rect 19794 4468 19800 4480
rect 19444 4440 19800 4468
rect 19794 4428 19800 4440
rect 19852 4428 19858 4480
rect 19889 4471 19947 4477
rect 19889 4437 19901 4471
rect 19935 4468 19947 4471
rect 20254 4468 20260 4480
rect 19935 4440 20260 4468
rect 19935 4437 19947 4440
rect 19889 4431 19947 4437
rect 20254 4428 20260 4440
rect 20312 4428 20318 4480
rect 20364 4468 20392 4508
rect 20708 4505 20720 4508
rect 20754 4536 20766 4539
rect 22664 4536 22692 4564
rect 20754 4508 22692 4536
rect 24029 4539 24087 4545
rect 20754 4505 20766 4508
rect 20708 4499 20766 4505
rect 24029 4505 24041 4539
rect 24075 4536 24087 4539
rect 25498 4536 25504 4548
rect 24075 4508 25504 4536
rect 24075 4505 24087 4508
rect 24029 4499 24087 4505
rect 25498 4496 25504 4508
rect 25556 4496 25562 4548
rect 21821 4471 21879 4477
rect 21821 4468 21833 4471
rect 20364 4440 21833 4468
rect 21821 4437 21833 4440
rect 21867 4437 21879 4471
rect 21821 4431 21879 4437
rect 1104 4378 24723 4400
rect 1104 4326 6814 4378
rect 6866 4326 6878 4378
rect 6930 4326 6942 4378
rect 6994 4326 7006 4378
rect 7058 4326 7070 4378
rect 7122 4326 12679 4378
rect 12731 4326 12743 4378
rect 12795 4326 12807 4378
rect 12859 4326 12871 4378
rect 12923 4326 12935 4378
rect 12987 4326 18544 4378
rect 18596 4326 18608 4378
rect 18660 4326 18672 4378
rect 18724 4326 18736 4378
rect 18788 4326 18800 4378
rect 18852 4326 24409 4378
rect 24461 4326 24473 4378
rect 24525 4326 24537 4378
rect 24589 4326 24601 4378
rect 24653 4326 24665 4378
rect 24717 4326 24723 4378
rect 1104 4304 24723 4326
rect 2222 4224 2228 4276
rect 2280 4264 2286 4276
rect 3694 4264 3700 4276
rect 2280 4236 3700 4264
rect 2280 4224 2286 4236
rect 3694 4224 3700 4236
rect 3752 4224 3758 4276
rect 4338 4224 4344 4276
rect 4396 4264 4402 4276
rect 4890 4264 4896 4276
rect 4396 4236 4896 4264
rect 4396 4224 4402 4236
rect 4890 4224 4896 4236
rect 4948 4224 4954 4276
rect 5074 4224 5080 4276
rect 5132 4264 5138 4276
rect 5132 4236 8800 4264
rect 5132 4224 5138 4236
rect 1857 4199 1915 4205
rect 1857 4165 1869 4199
rect 1903 4196 1915 4199
rect 1946 4196 1952 4208
rect 1903 4168 1952 4196
rect 1903 4165 1915 4168
rect 1857 4159 1915 4165
rect 1946 4156 1952 4168
rect 2004 4156 2010 4208
rect 2038 4156 2044 4208
rect 2096 4196 2102 4208
rect 2409 4199 2467 4205
rect 2409 4196 2421 4199
rect 2096 4168 2421 4196
rect 2096 4156 2102 4168
rect 2409 4165 2421 4168
rect 2455 4165 2467 4199
rect 6270 4196 6276 4208
rect 2409 4159 2467 4165
rect 4632 4168 6276 4196
rect 1394 4088 1400 4140
rect 1452 4088 1458 4140
rect 2498 4088 2504 4140
rect 2556 4088 2562 4140
rect 2682 4088 2688 4140
rect 2740 4088 2746 4140
rect 3602 4088 3608 4140
rect 3660 4088 3666 4140
rect 4632 4137 4660 4168
rect 6270 4156 6276 4168
rect 6328 4156 6334 4208
rect 8772 4196 8800 4236
rect 8938 4224 8944 4276
rect 8996 4224 9002 4276
rect 11422 4264 11428 4276
rect 9646 4236 11428 4264
rect 9646 4196 9674 4236
rect 11422 4224 11428 4236
rect 11480 4224 11486 4276
rect 12526 4224 12532 4276
rect 12584 4224 12590 4276
rect 13998 4224 14004 4276
rect 14056 4264 14062 4276
rect 14093 4267 14151 4273
rect 14093 4264 14105 4267
rect 14056 4236 14105 4264
rect 14056 4224 14062 4236
rect 14093 4233 14105 4236
rect 14139 4233 14151 4267
rect 14093 4227 14151 4233
rect 14550 4224 14556 4276
rect 14608 4224 14614 4276
rect 18230 4224 18236 4276
rect 18288 4264 18294 4276
rect 18690 4264 18696 4276
rect 18288 4236 18696 4264
rect 18288 4224 18294 4236
rect 18690 4224 18696 4236
rect 18748 4264 18754 4276
rect 19518 4264 19524 4276
rect 18748 4236 19524 4264
rect 18748 4224 18754 4236
rect 19518 4224 19524 4236
rect 19576 4264 19582 4276
rect 23566 4264 23572 4276
rect 19576 4236 21128 4264
rect 19576 4224 19582 4236
rect 8772 4168 9674 4196
rect 10137 4199 10195 4205
rect 10137 4165 10149 4199
rect 10183 4196 10195 4199
rect 10502 4196 10508 4208
rect 10183 4168 10508 4196
rect 10183 4165 10195 4168
rect 10137 4159 10195 4165
rect 10502 4156 10508 4168
rect 10560 4156 10566 4208
rect 11146 4156 11152 4208
rect 11204 4156 11210 4208
rect 11238 4156 11244 4208
rect 11296 4196 11302 4208
rect 14182 4196 14188 4208
rect 11296 4168 14188 4196
rect 11296 4156 11302 4168
rect 14182 4156 14188 4168
rect 14240 4156 14246 4208
rect 4617 4131 4675 4137
rect 4617 4097 4629 4131
rect 4663 4097 4675 4131
rect 4617 4091 4675 4097
rect 4891 4131 4949 4137
rect 4891 4097 4903 4131
rect 4937 4128 4949 4131
rect 5350 4128 5356 4140
rect 4937 4100 5356 4128
rect 4937 4097 4949 4100
rect 4891 4091 4949 4097
rect 5350 4088 5356 4100
rect 5408 4088 5414 4140
rect 5626 4088 5632 4140
rect 5684 4128 5690 4140
rect 6181 4131 6239 4137
rect 6181 4128 6193 4131
rect 5684 4100 6193 4128
rect 5684 4088 5690 4100
rect 6181 4097 6193 4100
rect 6227 4097 6239 4131
rect 6181 4091 6239 4097
rect 6638 4088 6644 4140
rect 6696 4128 6702 4140
rect 7285 4131 7343 4137
rect 7285 4128 7297 4131
rect 6696 4100 7297 4128
rect 6696 4088 6702 4100
rect 7285 4097 7297 4100
rect 7331 4128 7343 4131
rect 7466 4128 7472 4140
rect 7331 4100 7472 4128
rect 7331 4097 7343 4100
rect 7285 4091 7343 4097
rect 7466 4088 7472 4100
rect 7524 4088 7530 4140
rect 8294 4088 8300 4140
rect 8352 4088 8358 4140
rect 8938 4088 8944 4140
rect 8996 4128 9002 4140
rect 10042 4128 10048 4140
rect 8996 4100 10048 4128
rect 8996 4088 9002 4100
rect 10042 4088 10048 4100
rect 10100 4128 10106 4140
rect 10686 4128 10692 4140
rect 10100 4100 10692 4128
rect 10100 4088 10106 4100
rect 10686 4088 10692 4100
rect 10744 4088 10750 4140
rect 11164 4128 11192 4156
rect 11759 4131 11817 4137
rect 11759 4128 11771 4131
rect 11164 4100 11771 4128
rect 11759 4097 11771 4100
rect 11805 4097 11817 4131
rect 11759 4091 11817 4097
rect 13262 4088 13268 4140
rect 13320 4128 13326 4140
rect 13355 4131 13413 4137
rect 13355 4128 13367 4131
rect 13320 4100 13367 4128
rect 13320 4088 13326 4100
rect 13355 4097 13367 4100
rect 13401 4128 13413 4131
rect 14568 4128 14596 4224
rect 17126 4156 17132 4208
rect 17184 4196 17190 4208
rect 19426 4196 19432 4208
rect 17184 4168 19432 4196
rect 17184 4156 17190 4168
rect 19426 4156 19432 4168
rect 19484 4156 19490 4208
rect 13401 4100 14596 4128
rect 17681 4131 17739 4137
rect 13401 4097 13413 4100
rect 13355 4091 13413 4097
rect 17681 4097 17693 4131
rect 17727 4128 17739 4131
rect 17770 4128 17776 4140
rect 17727 4100 17776 4128
rect 17727 4097 17739 4100
rect 17681 4091 17739 4097
rect 17770 4088 17776 4100
rect 17828 4088 17834 4140
rect 17862 4088 17868 4140
rect 17920 4088 17926 4140
rect 18230 4088 18236 4140
rect 18288 4088 18294 4140
rect 18509 4131 18567 4137
rect 18509 4097 18521 4131
rect 18555 4128 18567 4131
rect 18690 4128 18696 4140
rect 18555 4100 18696 4128
rect 18555 4097 18567 4100
rect 18509 4091 18567 4097
rect 18690 4088 18696 4100
rect 18748 4088 18754 4140
rect 18783 4131 18841 4137
rect 18783 4097 18795 4131
rect 18829 4128 18841 4131
rect 19242 4128 19248 4140
rect 18829 4100 19248 4128
rect 18829 4097 18841 4100
rect 18783 4091 18841 4097
rect 19242 4088 19248 4100
rect 19300 4088 19306 4140
rect 20088 4128 20116 4236
rect 20165 4199 20223 4205
rect 20165 4165 20177 4199
rect 20211 4196 20223 4199
rect 20530 4196 20536 4208
rect 20211 4168 20536 4196
rect 20211 4165 20223 4168
rect 20165 4159 20223 4165
rect 20530 4156 20536 4168
rect 20588 4156 20594 4208
rect 20254 4128 20260 4140
rect 20088 4100 20260 4128
rect 20254 4088 20260 4100
rect 20312 4088 20318 4140
rect 20346 4088 20352 4140
rect 20404 4128 20410 4140
rect 20809 4131 20867 4137
rect 20809 4128 20821 4131
rect 20404 4100 20821 4128
rect 20404 4088 20410 4100
rect 20809 4097 20821 4100
rect 20855 4097 20867 4131
rect 21100 4128 21128 4236
rect 21468 4236 23572 4264
rect 21468 4205 21496 4236
rect 23566 4224 23572 4236
rect 23624 4224 23630 4276
rect 21453 4199 21511 4205
rect 21453 4165 21465 4199
rect 21499 4165 21511 4199
rect 21453 4159 21511 4165
rect 21634 4156 21640 4208
rect 21692 4156 21698 4208
rect 21910 4156 21916 4208
rect 21968 4196 21974 4208
rect 21968 4168 23060 4196
rect 21968 4156 21974 4168
rect 21100 4100 21864 4128
rect 20809 4091 20867 4097
rect 2516 4060 2544 4088
rect 2593 4063 2651 4069
rect 2593 4060 2605 4063
rect 2516 4032 2605 4060
rect 2593 4029 2605 4032
rect 2639 4029 2651 4063
rect 2593 4023 2651 4029
rect 2869 4063 2927 4069
rect 2869 4029 2881 4063
rect 2915 4060 2927 4063
rect 3722 4063 3780 4069
rect 3722 4060 3734 4063
rect 2915 4032 3280 4060
rect 2915 4029 2927 4032
rect 2869 4023 2927 4029
rect 3252 4004 3280 4032
rect 3436 4032 3734 4060
rect 2133 3995 2191 4001
rect 2133 3961 2145 3995
rect 2179 3992 2191 3995
rect 2958 3992 2964 4004
rect 2179 3964 2964 3992
rect 2179 3961 2191 3964
rect 2133 3955 2191 3961
rect 2958 3952 2964 3964
rect 3016 3952 3022 4004
rect 3234 3952 3240 4004
rect 3292 3952 3298 4004
rect 3326 3952 3332 4004
rect 3384 3952 3390 4004
rect 1581 3927 1639 3933
rect 1581 3893 1593 3927
rect 1627 3924 1639 3927
rect 1946 3924 1952 3936
rect 1627 3896 1952 3924
rect 1627 3893 1639 3896
rect 1581 3887 1639 3893
rect 1946 3884 1952 3896
rect 2004 3884 2010 3936
rect 3436 3924 3464 4032
rect 3722 4029 3734 4032
rect 3768 4029 3780 4063
rect 3722 4023 3780 4029
rect 3878 4020 3884 4072
rect 3936 4020 3942 4072
rect 7101 4063 7159 4069
rect 7101 4029 7113 4063
rect 7147 4029 7159 4063
rect 7101 4023 7159 4029
rect 7116 3992 7144 4023
rect 7374 4020 7380 4072
rect 7432 4060 7438 4072
rect 7745 4063 7803 4069
rect 7745 4060 7757 4063
rect 7432 4032 7757 4060
rect 7432 4020 7438 4032
rect 7745 4029 7757 4032
rect 7791 4029 7803 4063
rect 7745 4023 7803 4029
rect 8018 4020 8024 4072
rect 8076 4020 8082 4072
rect 8159 4063 8217 4069
rect 8159 4029 8171 4063
rect 8205 4060 8217 4063
rect 8478 4060 8484 4072
rect 8205 4032 8484 4060
rect 8205 4029 8217 4032
rect 8159 4023 8217 4029
rect 8478 4020 8484 4032
rect 8536 4020 8542 4072
rect 11054 4060 11060 4072
rect 8680 4032 11060 4060
rect 7834 3992 7840 4004
rect 7116 3964 7840 3992
rect 7834 3952 7840 3964
rect 7892 3952 7898 4004
rect 4246 3924 4252 3936
rect 3436 3896 4252 3924
rect 4246 3884 4252 3896
rect 4304 3884 4310 3936
rect 4522 3884 4528 3936
rect 4580 3884 4586 3936
rect 4982 3884 4988 3936
rect 5040 3924 5046 3936
rect 5629 3927 5687 3933
rect 5629 3924 5641 3927
rect 5040 3896 5641 3924
rect 5040 3884 5046 3896
rect 5629 3893 5641 3896
rect 5675 3893 5687 3927
rect 5629 3887 5687 3893
rect 5997 3927 6055 3933
rect 5997 3893 6009 3927
rect 6043 3924 6055 3927
rect 8680 3924 8708 4032
rect 11054 4020 11060 4032
rect 11112 4020 11118 4072
rect 11514 4020 11520 4072
rect 11572 4020 11578 4072
rect 13081 4063 13139 4069
rect 13081 4029 13093 4063
rect 13127 4029 13139 4063
rect 21726 4060 21732 4072
rect 13081 4023 13139 4029
rect 19168 4032 21732 4060
rect 9306 3952 9312 4004
rect 9364 3992 9370 4004
rect 11532 3992 11560 4020
rect 9364 3964 11560 3992
rect 9364 3952 9370 3964
rect 6043 3896 8708 3924
rect 6043 3893 6055 3896
rect 5997 3887 6055 3893
rect 10594 3884 10600 3936
rect 10652 3884 10658 3936
rect 11146 3884 11152 3936
rect 11204 3924 11210 3936
rect 12434 3924 12440 3936
rect 11204 3896 12440 3924
rect 11204 3884 11210 3896
rect 12434 3884 12440 3896
rect 12492 3884 12498 3936
rect 12986 3884 12992 3936
rect 13044 3924 13050 3936
rect 13096 3924 13124 4023
rect 14826 3952 14832 4004
rect 14884 3992 14890 4004
rect 17865 3995 17923 4001
rect 17865 3992 17877 3995
rect 14884 3964 17877 3992
rect 14884 3952 14890 3964
rect 17865 3961 17877 3964
rect 17911 3961 17923 3995
rect 17865 3955 17923 3961
rect 18046 3952 18052 4004
rect 18104 3992 18110 4004
rect 18506 3992 18512 4004
rect 18104 3964 18512 3992
rect 18104 3952 18110 3964
rect 18506 3952 18512 3964
rect 18564 3952 18570 4004
rect 13906 3924 13912 3936
rect 13044 3896 13912 3924
rect 13044 3884 13050 3896
rect 13906 3884 13912 3896
rect 13964 3924 13970 3936
rect 14642 3924 14648 3936
rect 13964 3896 14648 3924
rect 13964 3884 13970 3896
rect 14642 3884 14648 3896
rect 14700 3884 14706 3936
rect 18966 3884 18972 3936
rect 19024 3924 19030 3936
rect 19168 3924 19196 4032
rect 21726 4020 21732 4032
rect 21784 4020 21790 4072
rect 21836 4060 21864 4100
rect 22002 4088 22008 4140
rect 22060 4088 22066 4140
rect 22371 4131 22429 4137
rect 22371 4097 22383 4131
rect 22417 4128 22429 4131
rect 22922 4128 22928 4140
rect 22417 4100 22928 4128
rect 22417 4097 22429 4100
rect 22371 4091 22429 4097
rect 22922 4088 22928 4100
rect 22980 4088 22986 4140
rect 22094 4060 22100 4072
rect 21836 4032 22100 4060
rect 22094 4020 22100 4032
rect 22152 4020 22158 4072
rect 23032 4060 23060 4168
rect 24026 4156 24032 4208
rect 24084 4156 24090 4208
rect 23290 4088 23296 4140
rect 23348 4128 23354 4140
rect 23569 4131 23627 4137
rect 23569 4128 23581 4131
rect 23348 4100 23581 4128
rect 23348 4088 23354 4100
rect 23569 4097 23581 4100
rect 23615 4097 23627 4131
rect 23569 4091 23627 4097
rect 23750 4088 23756 4140
rect 23808 4088 23814 4140
rect 24213 4131 24271 4137
rect 24213 4097 24225 4131
rect 24259 4128 24271 4131
rect 24946 4128 24952 4140
rect 24259 4100 24952 4128
rect 24259 4097 24271 4100
rect 24213 4091 24271 4097
rect 24946 4088 24952 4100
rect 25004 4088 25010 4140
rect 23032 4032 23980 4060
rect 21082 3952 21088 4004
rect 21140 3992 21146 4004
rect 21266 3992 21272 4004
rect 21140 3964 21272 3992
rect 21140 3952 21146 3964
rect 21266 3952 21272 3964
rect 21324 3952 21330 4004
rect 21542 3952 21548 4004
rect 21600 3952 21606 4004
rect 22922 3952 22928 4004
rect 22980 3992 22986 4004
rect 23658 3992 23664 4004
rect 22980 3964 23664 3992
rect 22980 3952 22986 3964
rect 23658 3952 23664 3964
rect 23716 3952 23722 4004
rect 19024 3896 19196 3924
rect 19024 3884 19030 3896
rect 19242 3884 19248 3936
rect 19300 3924 19306 3936
rect 19521 3927 19579 3933
rect 19521 3924 19533 3927
rect 19300 3896 19533 3924
rect 19300 3884 19306 3896
rect 19521 3893 19533 3896
rect 19567 3893 19579 3927
rect 19521 3887 19579 3893
rect 19702 3884 19708 3936
rect 19760 3924 19766 3936
rect 20257 3927 20315 3933
rect 20257 3924 20269 3927
rect 19760 3896 20269 3924
rect 19760 3884 19766 3896
rect 20257 3893 20269 3896
rect 20303 3893 20315 3927
rect 20257 3887 20315 3893
rect 20530 3884 20536 3936
rect 20588 3924 20594 3936
rect 20901 3927 20959 3933
rect 20901 3924 20913 3927
rect 20588 3896 20913 3924
rect 20588 3884 20594 3896
rect 20901 3893 20913 3896
rect 20947 3893 20959 3927
rect 21560 3924 21588 3952
rect 23952 3936 23980 4032
rect 21821 3927 21879 3933
rect 21821 3924 21833 3927
rect 21560 3896 21833 3924
rect 20901 3887 20959 3893
rect 21821 3893 21833 3896
rect 21867 3893 21879 3927
rect 21821 3887 21879 3893
rect 23106 3884 23112 3936
rect 23164 3884 23170 3936
rect 23934 3884 23940 3936
rect 23992 3884 23998 3936
rect 1104 3834 24564 3856
rect 1104 3782 3882 3834
rect 3934 3782 3946 3834
rect 3998 3782 4010 3834
rect 4062 3782 4074 3834
rect 4126 3782 4138 3834
rect 4190 3782 9747 3834
rect 9799 3782 9811 3834
rect 9863 3782 9875 3834
rect 9927 3782 9939 3834
rect 9991 3782 10003 3834
rect 10055 3782 15612 3834
rect 15664 3782 15676 3834
rect 15728 3782 15740 3834
rect 15792 3782 15804 3834
rect 15856 3782 15868 3834
rect 15920 3782 21477 3834
rect 21529 3782 21541 3834
rect 21593 3782 21605 3834
rect 21657 3782 21669 3834
rect 21721 3782 21733 3834
rect 21785 3782 24564 3834
rect 1104 3760 24564 3782
rect 1578 3680 1584 3732
rect 1636 3680 1642 3732
rect 2777 3723 2835 3729
rect 2777 3689 2789 3723
rect 2823 3720 2835 3723
rect 3326 3720 3332 3732
rect 2823 3692 3332 3720
rect 2823 3689 2835 3692
rect 2777 3683 2835 3689
rect 3326 3680 3332 3692
rect 3384 3680 3390 3732
rect 4338 3680 4344 3732
rect 4396 3680 4402 3732
rect 4890 3720 4896 3732
rect 4448 3692 4896 3720
rect 3050 3612 3056 3664
rect 3108 3652 3114 3664
rect 3421 3655 3479 3661
rect 3421 3652 3433 3655
rect 3108 3624 3433 3652
rect 3108 3612 3114 3624
rect 3421 3621 3433 3624
rect 3467 3621 3479 3655
rect 4356 3652 4384 3680
rect 4448 3661 4476 3692
rect 4890 3680 4896 3692
rect 4948 3680 4954 3732
rect 5074 3680 5080 3732
rect 5132 3720 5138 3732
rect 5132 3692 5396 3720
rect 5132 3680 5138 3692
rect 3421 3615 3479 3621
rect 3988 3624 4384 3652
rect 4433 3655 4491 3661
rect 1486 3544 1492 3596
rect 1544 3584 1550 3596
rect 1765 3587 1823 3593
rect 1765 3584 1777 3587
rect 1544 3556 1777 3584
rect 1544 3544 1550 3556
rect 1765 3553 1777 3556
rect 1811 3553 1823 3587
rect 1765 3547 1823 3553
rect 3786 3544 3792 3596
rect 3844 3544 3850 3596
rect 658 3476 664 3528
rect 716 3516 722 3528
rect 1397 3519 1455 3525
rect 1397 3516 1409 3519
rect 716 3488 1409 3516
rect 716 3476 722 3488
rect 1397 3485 1409 3488
rect 1443 3485 1455 3519
rect 1397 3479 1455 3485
rect 2039 3519 2097 3525
rect 2039 3485 2051 3519
rect 2085 3516 2097 3519
rect 2958 3516 2964 3528
rect 2085 3488 2964 3516
rect 2085 3485 2097 3488
rect 2039 3479 2097 3485
rect 2958 3476 2964 3488
rect 3016 3476 3022 3528
rect 3418 3516 3424 3528
rect 3068 3488 3424 3516
rect 2314 3340 2320 3392
rect 2372 3380 2378 3392
rect 3068 3380 3096 3488
rect 3418 3476 3424 3488
rect 3476 3476 3482 3528
rect 3988 3525 4016 3624
rect 4433 3621 4445 3655
rect 4479 3621 4491 3655
rect 4433 3615 4491 3621
rect 4338 3544 4344 3596
rect 4396 3584 4402 3596
rect 5368 3584 5396 3692
rect 5718 3680 5724 3732
rect 5776 3720 5782 3732
rect 5776 3692 7328 3720
rect 5776 3680 5782 3692
rect 5736 3593 5764 3680
rect 7300 3652 7328 3692
rect 7558 3680 7564 3732
rect 7616 3680 7622 3732
rect 7834 3680 7840 3732
rect 7892 3720 7898 3732
rect 9122 3720 9128 3732
rect 7892 3692 9128 3720
rect 7892 3680 7898 3692
rect 9122 3680 9128 3692
rect 9180 3680 9186 3732
rect 11882 3680 11888 3732
rect 11940 3680 11946 3732
rect 12986 3720 12992 3732
rect 12544 3692 12992 3720
rect 5828 3624 6500 3652
rect 7300 3624 8248 3652
rect 5721 3587 5779 3593
rect 4396 3556 4752 3584
rect 4396 3544 4402 3556
rect 4724 3525 4752 3556
rect 4914 3556 5672 3584
rect 3973 3519 4031 3525
rect 3973 3485 3985 3519
rect 4019 3485 4031 3519
rect 3973 3479 4031 3485
rect 4709 3519 4767 3525
rect 4709 3485 4721 3519
rect 4755 3485 4767 3519
rect 4709 3479 4767 3485
rect 4826 3519 4884 3525
rect 4826 3485 4838 3519
rect 4872 3516 4884 3519
rect 4914 3516 4942 3556
rect 4872 3488 4942 3516
rect 4872 3485 4884 3488
rect 4826 3479 4884 3485
rect 4982 3476 4988 3528
rect 5040 3476 5046 3528
rect 5644 3516 5672 3556
rect 5721 3553 5733 3587
rect 5767 3553 5779 3587
rect 5721 3547 5779 3553
rect 5828 3516 5856 3624
rect 6472 3596 6500 3624
rect 8220 3596 8248 3624
rect 8944 3596 8996 3602
rect 5902 3544 5908 3596
rect 5960 3544 5966 3596
rect 6362 3544 6368 3596
rect 6420 3544 6426 3596
rect 6454 3544 6460 3596
rect 6512 3584 6518 3596
rect 6822 3593 6828 3596
rect 6641 3587 6699 3593
rect 6641 3584 6653 3587
rect 6512 3556 6653 3584
rect 6512 3544 6518 3556
rect 6641 3553 6653 3556
rect 6687 3553 6699 3587
rect 6641 3547 6699 3553
rect 6779 3587 6828 3593
rect 6779 3553 6791 3587
rect 6825 3553 6828 3587
rect 6779 3547 6828 3553
rect 6822 3544 6828 3547
rect 6880 3544 6886 3596
rect 7282 3584 7288 3596
rect 6932 3556 7288 3584
rect 6932 3525 6960 3556
rect 7282 3544 7288 3556
rect 7340 3544 7346 3596
rect 8202 3544 8208 3596
rect 8260 3544 8266 3596
rect 12544 3593 12572 3692
rect 12986 3680 12992 3692
rect 13044 3680 13050 3732
rect 13446 3680 13452 3732
rect 13504 3720 13510 3732
rect 13541 3723 13599 3729
rect 13541 3720 13553 3723
rect 13504 3692 13553 3720
rect 13504 3680 13510 3692
rect 13541 3689 13553 3692
rect 13587 3689 13599 3723
rect 17678 3720 17684 3732
rect 13541 3683 13599 3689
rect 17144 3692 17684 3720
rect 12529 3587 12587 3593
rect 12529 3553 12541 3587
rect 12575 3553 12587 3587
rect 12529 3547 12587 3553
rect 8944 3538 8996 3544
rect 5644 3488 5856 3516
rect 6917 3519 6975 3525
rect 6917 3485 6929 3519
rect 6963 3485 6975 3519
rect 6917 3479 6975 3485
rect 7837 3519 7895 3525
rect 7837 3485 7849 3519
rect 7883 3485 7895 3519
rect 7837 3479 7895 3485
rect 3237 3451 3295 3457
rect 3237 3417 3249 3451
rect 3283 3448 3295 3451
rect 7852 3448 7880 3479
rect 7926 3476 7932 3528
rect 7984 3516 7990 3528
rect 8113 3519 8171 3525
rect 8113 3516 8125 3519
rect 7984 3488 8125 3516
rect 7984 3476 7990 3488
rect 8113 3485 8125 3488
rect 8159 3485 8171 3519
rect 8113 3479 8171 3485
rect 8757 3519 8815 3525
rect 8757 3485 8769 3519
rect 8803 3485 8815 3519
rect 8757 3479 8815 3485
rect 9401 3519 9459 3525
rect 9401 3485 9413 3519
rect 9447 3516 9459 3519
rect 9582 3516 9588 3528
rect 9447 3488 9588 3516
rect 9447 3485 9459 3488
rect 9401 3479 9459 3485
rect 3283 3420 4016 3448
rect 3283 3417 3295 3420
rect 3237 3411 3295 3417
rect 2372 3352 3096 3380
rect 3988 3380 4016 3420
rect 7392 3420 7880 3448
rect 8772 3448 8800 3479
rect 9582 3476 9588 3488
rect 9640 3476 9646 3528
rect 10778 3476 10784 3528
rect 10836 3476 10842 3528
rect 10873 3519 10931 3525
rect 10873 3485 10885 3519
rect 10919 3485 10931 3519
rect 10873 3479 10931 3485
rect 11147 3519 11205 3525
rect 11147 3485 11159 3519
rect 11193 3516 11205 3519
rect 11238 3516 11244 3528
rect 11193 3488 11244 3516
rect 11193 3485 11205 3488
rect 11147 3479 11205 3485
rect 8772 3420 9444 3448
rect 5629 3383 5687 3389
rect 5629 3380 5641 3383
rect 3988 3352 5641 3380
rect 2372 3340 2378 3352
rect 5629 3349 5641 3352
rect 5675 3349 5687 3383
rect 5629 3343 5687 3349
rect 6546 3340 6552 3392
rect 6604 3380 6610 3392
rect 7392 3380 7420 3420
rect 6604 3352 7420 3380
rect 6604 3340 6610 3352
rect 7650 3340 7656 3392
rect 7708 3340 7714 3392
rect 7926 3340 7932 3392
rect 7984 3340 7990 3392
rect 8570 3340 8576 3392
rect 8628 3340 8634 3392
rect 9122 3340 9128 3392
rect 9180 3340 9186 3392
rect 9416 3380 9444 3420
rect 9490 3408 9496 3460
rect 9548 3408 9554 3460
rect 9861 3451 9919 3457
rect 9861 3417 9873 3451
rect 9907 3417 9919 3451
rect 9861 3411 9919 3417
rect 10229 3451 10287 3457
rect 10229 3417 10241 3451
rect 10275 3448 10287 3451
rect 10796 3448 10824 3476
rect 10275 3420 10824 3448
rect 10888 3448 10916 3479
rect 11238 3476 11244 3488
rect 11296 3476 11302 3528
rect 11514 3476 11520 3528
rect 11572 3476 11578 3528
rect 12158 3476 12164 3528
rect 12216 3516 12222 3528
rect 17144 3525 17172 3692
rect 17678 3680 17684 3692
rect 17736 3680 17742 3732
rect 17773 3723 17831 3729
rect 17773 3689 17785 3723
rect 17819 3720 17831 3723
rect 17862 3720 17868 3732
rect 17819 3692 17868 3720
rect 17819 3689 17831 3692
rect 17773 3683 17831 3689
rect 17862 3680 17868 3692
rect 17920 3680 17926 3732
rect 18230 3680 18236 3732
rect 18288 3680 18294 3732
rect 19334 3680 19340 3732
rect 19392 3680 19398 3732
rect 19426 3680 19432 3732
rect 19484 3720 19490 3732
rect 19705 3723 19763 3729
rect 19705 3720 19717 3723
rect 19484 3692 19717 3720
rect 19484 3680 19490 3692
rect 19705 3689 19717 3692
rect 19751 3689 19763 3723
rect 19705 3683 19763 3689
rect 20254 3680 20260 3732
rect 20312 3720 20318 3732
rect 20312 3692 20760 3720
rect 20312 3680 20318 3692
rect 17497 3655 17555 3661
rect 17497 3621 17509 3655
rect 17543 3652 17555 3655
rect 18248 3652 18276 3680
rect 17543 3624 18276 3652
rect 19352 3652 19380 3680
rect 19352 3624 20576 3652
rect 17543 3621 17555 3624
rect 17497 3615 17555 3621
rect 17218 3544 17224 3596
rect 17276 3544 17282 3596
rect 17770 3584 17776 3596
rect 17420 3556 17776 3584
rect 17420 3525 17448 3556
rect 17770 3544 17776 3556
rect 17828 3544 17834 3596
rect 17880 3556 19840 3584
rect 12771 3519 12829 3525
rect 12771 3516 12783 3519
rect 12216 3488 12783 3516
rect 12216 3476 12222 3488
rect 12771 3485 12783 3488
rect 12817 3485 12829 3519
rect 12771 3479 12829 3485
rect 17129 3519 17187 3525
rect 17129 3485 17141 3519
rect 17175 3485 17187 3519
rect 17129 3479 17187 3485
rect 17405 3519 17463 3525
rect 17405 3485 17417 3519
rect 17451 3485 17463 3519
rect 17405 3479 17463 3485
rect 17586 3476 17592 3528
rect 17644 3476 17650 3528
rect 17678 3476 17684 3528
rect 17736 3476 17742 3528
rect 11532 3448 11560 3476
rect 10888 3420 11560 3448
rect 10275 3417 10287 3420
rect 10229 3411 10287 3417
rect 9582 3380 9588 3392
rect 9416 3352 9588 3380
rect 9582 3340 9588 3352
rect 9640 3340 9646 3392
rect 9876 3380 9904 3411
rect 16942 3408 16948 3460
rect 17000 3448 17006 3460
rect 17880 3448 17908 3556
rect 18414 3476 18420 3528
rect 18472 3516 18478 3528
rect 18601 3519 18659 3525
rect 18601 3516 18613 3519
rect 18472 3488 18613 3516
rect 18472 3476 18478 3488
rect 18601 3485 18613 3488
rect 18647 3485 18659 3519
rect 18601 3479 18659 3485
rect 19242 3476 19248 3528
rect 19300 3476 19306 3528
rect 19426 3476 19432 3528
rect 19484 3476 19490 3528
rect 19812 3525 19840 3556
rect 20346 3544 20352 3596
rect 20404 3544 20410 3596
rect 19797 3519 19855 3525
rect 19797 3485 19809 3519
rect 19843 3485 19855 3519
rect 19797 3479 19855 3485
rect 19978 3476 19984 3528
rect 20036 3476 20042 3528
rect 17000 3420 17908 3448
rect 18049 3451 18107 3457
rect 17000 3408 17006 3420
rect 18049 3417 18061 3451
rect 18095 3448 18107 3451
rect 19334 3448 19340 3460
rect 18095 3420 19340 3448
rect 18095 3417 18107 3420
rect 18049 3411 18107 3417
rect 19334 3408 19340 3420
rect 19392 3408 19398 3460
rect 20364 3448 20392 3544
rect 19444 3420 20392 3448
rect 10318 3380 10324 3392
rect 9876 3352 10324 3380
rect 10318 3340 10324 3352
rect 10376 3340 10382 3392
rect 10410 3340 10416 3392
rect 10468 3340 10474 3392
rect 18138 3340 18144 3392
rect 18196 3340 18202 3392
rect 18230 3340 18236 3392
rect 18288 3380 18294 3392
rect 18693 3383 18751 3389
rect 18693 3380 18705 3383
rect 18288 3352 18705 3380
rect 18288 3340 18294 3352
rect 18693 3349 18705 3352
rect 18739 3349 18751 3383
rect 18693 3343 18751 3349
rect 19150 3340 19156 3392
rect 19208 3380 19214 3392
rect 19444 3380 19472 3420
rect 19208 3352 19472 3380
rect 19208 3340 19214 3352
rect 19518 3340 19524 3392
rect 19576 3380 19582 3392
rect 20073 3383 20131 3389
rect 20073 3380 20085 3383
rect 19576 3352 20085 3380
rect 19576 3340 19582 3352
rect 20073 3349 20085 3352
rect 20119 3349 20131 3383
rect 20073 3343 20131 3349
rect 20346 3340 20352 3392
rect 20404 3380 20410 3392
rect 20441 3383 20499 3389
rect 20441 3380 20453 3383
rect 20404 3352 20453 3380
rect 20404 3340 20410 3352
rect 20441 3349 20453 3352
rect 20487 3349 20499 3383
rect 20548 3380 20576 3624
rect 20732 3593 20760 3692
rect 21729 3655 21787 3661
rect 21729 3621 21741 3655
rect 21775 3621 21787 3655
rect 21729 3615 21787 3621
rect 20717 3587 20775 3593
rect 20717 3553 20729 3587
rect 20763 3553 20775 3587
rect 20717 3547 20775 3553
rect 20625 3519 20683 3525
rect 20625 3485 20637 3519
rect 20671 3485 20683 3519
rect 20625 3479 20683 3485
rect 20640 3448 20668 3479
rect 20898 3476 20904 3528
rect 20956 3516 20962 3528
rect 20991 3519 21049 3525
rect 20991 3516 21003 3519
rect 20956 3488 21003 3516
rect 20956 3476 20962 3488
rect 20991 3485 21003 3488
rect 21037 3485 21049 3519
rect 20991 3479 21049 3485
rect 21082 3476 21088 3528
rect 21140 3516 21146 3528
rect 21744 3516 21772 3615
rect 22278 3612 22284 3664
rect 22336 3612 22342 3664
rect 23658 3652 23664 3664
rect 23032 3624 23664 3652
rect 21818 3544 21824 3596
rect 21876 3584 21882 3596
rect 23032 3584 23060 3624
rect 23658 3612 23664 3624
rect 23716 3612 23722 3664
rect 23842 3612 23848 3664
rect 23900 3612 23906 3664
rect 21876 3556 23060 3584
rect 21876 3544 21882 3556
rect 23106 3544 23112 3596
rect 23164 3544 23170 3596
rect 22097 3519 22155 3525
rect 22097 3516 22109 3519
rect 21140 3488 22109 3516
rect 21140 3476 21146 3488
rect 22097 3485 22109 3488
rect 22143 3485 22155 3519
rect 22097 3479 22155 3485
rect 22186 3476 22192 3528
rect 22244 3516 22250 3528
rect 22281 3519 22339 3525
rect 22281 3516 22293 3519
rect 22244 3488 22293 3516
rect 22244 3476 22250 3488
rect 22281 3485 22293 3488
rect 22327 3485 22339 3519
rect 22281 3479 22339 3485
rect 22462 3476 22468 3528
rect 22520 3516 22526 3528
rect 22649 3519 22707 3525
rect 22649 3516 22661 3519
rect 22520 3488 22661 3516
rect 22520 3476 22526 3488
rect 22649 3485 22661 3488
rect 22695 3485 22707 3519
rect 22649 3479 22707 3485
rect 23293 3519 23351 3525
rect 23293 3485 23305 3519
rect 23339 3485 23351 3519
rect 23293 3479 23351 3485
rect 21818 3448 21824 3460
rect 20640 3420 21824 3448
rect 21818 3408 21824 3420
rect 21876 3408 21882 3460
rect 22738 3408 22744 3460
rect 22796 3448 22802 3460
rect 23106 3448 23112 3460
rect 22796 3420 23112 3448
rect 22796 3408 22802 3420
rect 23106 3408 23112 3420
rect 23164 3408 23170 3460
rect 23308 3380 23336 3479
rect 23474 3476 23480 3528
rect 23532 3516 23538 3528
rect 23753 3519 23811 3525
rect 23753 3516 23765 3519
rect 23532 3488 23765 3516
rect 23532 3476 23538 3488
rect 23753 3485 23765 3488
rect 23799 3485 23811 3519
rect 23753 3479 23811 3485
rect 23842 3408 23848 3460
rect 23900 3448 23906 3460
rect 25222 3448 25228 3460
rect 23900 3420 25228 3448
rect 23900 3408 23906 3420
rect 25222 3408 25228 3420
rect 25280 3408 25286 3460
rect 20548 3352 23336 3380
rect 20441 3343 20499 3349
rect 1104 3290 24723 3312
rect 1104 3238 6814 3290
rect 6866 3238 6878 3290
rect 6930 3238 6942 3290
rect 6994 3238 7006 3290
rect 7058 3238 7070 3290
rect 7122 3238 12679 3290
rect 12731 3238 12743 3290
rect 12795 3238 12807 3290
rect 12859 3238 12871 3290
rect 12923 3238 12935 3290
rect 12987 3238 18544 3290
rect 18596 3238 18608 3290
rect 18660 3238 18672 3290
rect 18724 3238 18736 3290
rect 18788 3238 18800 3290
rect 18852 3238 24409 3290
rect 24461 3238 24473 3290
rect 24525 3238 24537 3290
rect 24589 3238 24601 3290
rect 24653 3238 24665 3290
rect 24717 3238 24723 3290
rect 1104 3216 24723 3238
rect 1765 3179 1823 3185
rect 1765 3145 1777 3179
rect 1811 3176 1823 3179
rect 1854 3176 1860 3188
rect 1811 3148 1860 3176
rect 1811 3145 1823 3148
rect 1765 3139 1823 3145
rect 1854 3136 1860 3148
rect 1912 3136 1918 3188
rect 4522 3176 4528 3188
rect 2746 3148 4528 3176
rect 1673 3111 1731 3117
rect 1673 3077 1685 3111
rect 1719 3108 1731 3111
rect 2746 3108 2774 3148
rect 4522 3136 4528 3148
rect 4580 3136 4586 3188
rect 4617 3179 4675 3185
rect 4617 3145 4629 3179
rect 4663 3176 4675 3179
rect 5166 3176 5172 3188
rect 4663 3148 5172 3176
rect 4663 3145 4675 3148
rect 4617 3139 4675 3145
rect 5166 3136 5172 3148
rect 5224 3136 5230 3188
rect 5905 3179 5963 3185
rect 5905 3145 5917 3179
rect 5951 3176 5963 3179
rect 6362 3176 6368 3188
rect 5951 3148 6368 3176
rect 5951 3145 5963 3148
rect 5905 3139 5963 3145
rect 6362 3136 6368 3148
rect 6420 3136 6426 3188
rect 6549 3179 6607 3185
rect 6549 3145 6561 3179
rect 6595 3176 6607 3179
rect 6638 3176 6644 3188
rect 6595 3148 6644 3176
rect 6595 3145 6607 3148
rect 6549 3139 6607 3145
rect 6638 3136 6644 3148
rect 6696 3136 6702 3188
rect 7190 3136 7196 3188
rect 7248 3136 7254 3188
rect 8573 3179 8631 3185
rect 8573 3145 8585 3179
rect 8619 3176 8631 3179
rect 8938 3176 8944 3188
rect 8619 3148 8944 3176
rect 8619 3145 8631 3148
rect 8573 3139 8631 3145
rect 8938 3136 8944 3148
rect 8996 3136 9002 3188
rect 9490 3136 9496 3188
rect 9548 3176 9554 3188
rect 9953 3179 10011 3185
rect 9953 3176 9965 3179
rect 9548 3148 9965 3176
rect 9548 3136 9554 3148
rect 9953 3145 9965 3148
rect 9999 3145 10011 3179
rect 12158 3176 12164 3188
rect 9953 3139 10011 3145
rect 11882 3148 12164 3176
rect 1719 3080 2774 3108
rect 1719 3077 1731 3080
rect 1673 3071 1731 3077
rect 4982 3068 4988 3120
rect 5040 3068 5046 3120
rect 6270 3108 6276 3120
rect 5552 3080 6276 3108
rect 5151 3073 5209 3079
rect 2222 3000 2228 3052
rect 2280 3000 2286 3052
rect 2593 3043 2651 3049
rect 2593 3009 2605 3043
rect 2639 3040 2651 3043
rect 2866 3040 2872 3052
rect 2639 3012 2872 3040
rect 2639 3009 2651 3012
rect 2593 3003 2651 3009
rect 2866 3000 2872 3012
rect 2924 3000 2930 3052
rect 3970 3000 3976 3052
rect 4028 3000 4034 3052
rect 5000 3040 5028 3068
rect 4538 3012 5028 3040
rect 5151 3039 5163 3073
rect 5197 3070 5209 3073
rect 5197 3052 5210 3070
rect 5224 3040 5230 3052
rect 5552 3040 5580 3080
rect 6270 3068 6276 3080
rect 6328 3068 6334 3120
rect 7208 3108 7236 3136
rect 7208 3080 9352 3108
rect 5151 3033 5172 3039
rect 2682 2932 2688 2984
rect 2740 2972 2746 2984
rect 2777 2975 2835 2981
rect 2777 2972 2789 2975
rect 2740 2944 2789 2972
rect 2740 2932 2746 2944
rect 2777 2941 2789 2944
rect 2823 2941 2835 2975
rect 2777 2935 2835 2941
rect 2961 2975 3019 2981
rect 2961 2941 2973 2975
rect 3007 2941 3019 2975
rect 2961 2935 3019 2941
rect 2976 2904 3004 2935
rect 3510 2932 3516 2984
rect 3568 2972 3574 2984
rect 3697 2975 3755 2981
rect 3697 2972 3709 2975
rect 3568 2944 3709 2972
rect 3568 2932 3574 2944
rect 3697 2941 3709 2944
rect 3743 2941 3755 2975
rect 3697 2935 3755 2941
rect 3835 2975 3893 2981
rect 3835 2941 3847 2975
rect 3881 2972 3893 2975
rect 4338 2972 4344 2984
rect 3881 2944 4344 2972
rect 3881 2941 3893 2944
rect 3835 2935 3893 2941
rect 4338 2932 4344 2944
rect 4396 2972 4402 2984
rect 4538 2972 4566 3012
rect 5166 3000 5172 3033
rect 5224 3012 5580 3040
rect 5224 3000 5230 3012
rect 5626 3000 5632 3052
rect 5684 3040 5690 3052
rect 6457 3043 6515 3049
rect 6457 3040 6469 3043
rect 5684 3012 6469 3040
rect 5684 3000 5690 3012
rect 6457 3009 6469 3012
rect 6503 3009 6515 3043
rect 6457 3003 6515 3009
rect 6917 3043 6975 3049
rect 6917 3009 6929 3043
rect 6963 3009 6975 3043
rect 6917 3003 6975 3009
rect 4396 2944 4566 2972
rect 4893 2975 4951 2981
rect 4396 2932 4402 2944
rect 4893 2941 4905 2975
rect 4939 2941 4951 2975
rect 6932 2972 6960 3003
rect 7190 3000 7196 3052
rect 7248 3000 7254 3052
rect 7466 3000 7472 3052
rect 7524 3000 7530 3052
rect 7742 3000 7748 3052
rect 7800 3040 7806 3052
rect 7835 3043 7893 3049
rect 7835 3040 7847 3043
rect 7800 3012 7847 3040
rect 7800 3000 7806 3012
rect 7835 3009 7847 3012
rect 7881 3040 7893 3043
rect 7881 3012 8294 3040
rect 7881 3009 7893 3012
rect 7835 3003 7893 3009
rect 7374 2972 7380 2984
rect 6932 2944 7380 2972
rect 4893 2935 4951 2941
rect 3234 2904 3240 2916
rect 2976 2876 3240 2904
rect 3234 2864 3240 2876
rect 3292 2864 3298 2916
rect 3418 2864 3424 2916
rect 3476 2864 3482 2916
rect 3510 2796 3516 2848
rect 3568 2836 3574 2848
rect 4430 2836 4436 2848
rect 3568 2808 4436 2836
rect 3568 2796 3574 2808
rect 4430 2796 4436 2808
rect 4488 2796 4494 2848
rect 4908 2836 4936 2935
rect 7374 2932 7380 2944
rect 7432 2932 7438 2984
rect 7561 2975 7619 2981
rect 7561 2941 7573 2975
rect 7607 2941 7619 2975
rect 7561 2935 7619 2941
rect 6454 2864 6460 2916
rect 6512 2904 6518 2916
rect 6512 2876 7328 2904
rect 6512 2864 6518 2876
rect 5902 2836 5908 2848
rect 4908 2808 5908 2836
rect 5902 2796 5908 2808
rect 5960 2796 5966 2848
rect 6730 2796 6736 2848
rect 6788 2796 6794 2848
rect 7006 2796 7012 2848
rect 7064 2796 7070 2848
rect 7300 2845 7328 2876
rect 7285 2839 7343 2845
rect 7285 2805 7297 2839
rect 7331 2805 7343 2839
rect 7576 2836 7604 2935
rect 8266 2904 8294 3012
rect 8846 3000 8852 3052
rect 8904 3040 8910 3052
rect 9215 3043 9273 3049
rect 9215 3040 9227 3043
rect 8904 3012 9227 3040
rect 8904 3000 8910 3012
rect 9215 3009 9227 3012
rect 9261 3009 9273 3043
rect 9324 3040 9352 3080
rect 9398 3068 9404 3120
rect 9456 3108 9462 3120
rect 10686 3108 10692 3120
rect 9456 3080 10692 3108
rect 9456 3068 9462 3080
rect 10686 3068 10692 3080
rect 10744 3068 10750 3120
rect 10870 3068 10876 3120
rect 10928 3068 10934 3120
rect 11882 3059 11910 3148
rect 12158 3136 12164 3148
rect 12216 3136 12222 3188
rect 16942 3136 16948 3188
rect 17000 3136 17006 3188
rect 17313 3179 17371 3185
rect 17313 3145 17325 3179
rect 17359 3176 17371 3179
rect 17678 3176 17684 3188
rect 17359 3148 17684 3176
rect 17359 3145 17371 3148
rect 17313 3139 17371 3145
rect 17678 3136 17684 3148
rect 17736 3136 17742 3188
rect 19242 3176 19248 3188
rect 18248 3148 19248 3176
rect 16482 3068 16488 3120
rect 16540 3068 16546 3120
rect 18248 3108 18276 3148
rect 19242 3136 19248 3148
rect 19300 3136 19306 3188
rect 19334 3136 19340 3188
rect 19392 3176 19398 3188
rect 21453 3179 21511 3185
rect 21453 3176 21465 3179
rect 19392 3148 21465 3176
rect 19392 3136 19398 3148
rect 21453 3145 21465 3148
rect 21499 3145 21511 3179
rect 21453 3139 21511 3145
rect 22646 3136 22652 3188
rect 22704 3176 22710 3188
rect 23106 3176 23112 3188
rect 22704 3148 23112 3176
rect 22704 3136 22710 3148
rect 23106 3136 23112 3148
rect 23164 3136 23170 3188
rect 24946 3136 24952 3188
rect 25004 3176 25010 3188
rect 25590 3176 25596 3188
rect 25004 3148 25596 3176
rect 25004 3136 25010 3148
rect 25590 3136 25596 3148
rect 25648 3136 25654 3188
rect 18782 3108 18788 3120
rect 16776 3080 18276 3108
rect 18340 3080 18788 3108
rect 11882 3053 11941 3059
rect 10410 3040 10416 3052
rect 9324 3012 10416 3040
rect 9215 3003 9273 3009
rect 10410 3000 10416 3012
rect 10468 3000 10474 3052
rect 11514 3000 11520 3052
rect 11572 3040 11578 3052
rect 11609 3043 11667 3049
rect 11609 3040 11621 3043
rect 11572 3012 11621 3040
rect 11572 3000 11578 3012
rect 11609 3009 11621 3012
rect 11655 3009 11667 3043
rect 11882 3022 11895 3053
rect 11883 3019 11895 3022
rect 11929 3019 11941 3053
rect 16776 3049 16804 3080
rect 11883 3013 11941 3019
rect 16761 3043 16819 3049
rect 11609 3003 11667 3009
rect 16761 3009 16773 3043
rect 16807 3009 16819 3043
rect 16761 3003 16819 3009
rect 16945 3043 17003 3049
rect 16945 3009 16957 3043
rect 16991 3040 17003 3043
rect 17126 3040 17132 3052
rect 16991 3012 17132 3040
rect 16991 3009 17003 3012
rect 16945 3003 17003 3009
rect 17126 3000 17132 3012
rect 17184 3000 17190 3052
rect 17221 3043 17279 3049
rect 17221 3009 17233 3043
rect 17267 3040 17279 3043
rect 17402 3040 17408 3052
rect 17267 3012 17408 3040
rect 17267 3009 17279 3012
rect 17221 3003 17279 3009
rect 17402 3000 17408 3012
rect 17460 3000 17466 3052
rect 17494 3000 17500 3052
rect 17552 3000 17558 3052
rect 17586 3000 17592 3052
rect 17644 3000 17650 3052
rect 18340 3049 18368 3080
rect 18782 3068 18788 3080
rect 18840 3068 18846 3120
rect 19058 3068 19064 3120
rect 19116 3068 19122 3120
rect 19610 3068 19616 3120
rect 19668 3068 19674 3120
rect 21910 3068 21916 3120
rect 21968 3108 21974 3120
rect 22986 3111 23044 3117
rect 22986 3108 22998 3111
rect 21968 3080 22998 3108
rect 21968 3068 21974 3080
rect 22986 3077 22998 3080
rect 23032 3077 23044 3111
rect 22986 3071 23044 3077
rect 17681 3043 17739 3049
rect 17681 3009 17693 3043
rect 17727 3009 17739 3043
rect 17681 3003 17739 3009
rect 18325 3043 18383 3049
rect 18325 3009 18337 3043
rect 18371 3009 18383 3043
rect 18325 3003 18383 3009
rect 18509 3043 18567 3049
rect 18509 3009 18521 3043
rect 18555 3040 18567 3043
rect 18966 3040 18972 3052
rect 18555 3012 18972 3040
rect 18555 3009 18567 3012
rect 18509 3003 18567 3009
rect 8754 2932 8760 2984
rect 8812 2972 8818 2984
rect 8941 2975 8999 2981
rect 8941 2972 8953 2975
rect 8812 2944 8953 2972
rect 8812 2932 8818 2944
rect 8941 2941 8953 2944
rect 8987 2941 8999 2975
rect 8941 2935 8999 2941
rect 12526 2932 12532 2984
rect 12584 2972 12590 2984
rect 13446 2972 13452 2984
rect 12584 2944 13452 2972
rect 12584 2932 12590 2944
rect 13446 2932 13452 2944
rect 13504 2972 13510 2984
rect 14458 2972 14464 2984
rect 13504 2944 14464 2972
rect 13504 2932 13510 2944
rect 14458 2932 14464 2944
rect 14516 2932 14522 2984
rect 8662 2904 8668 2916
rect 8266 2876 8668 2904
rect 8662 2864 8668 2876
rect 8720 2864 8726 2916
rect 8772 2836 8800 2932
rect 17218 2864 17224 2916
rect 17276 2904 17282 2916
rect 17512 2904 17540 3000
rect 17276 2876 17540 2904
rect 17604 2904 17632 3000
rect 17696 2972 17724 3003
rect 18966 3000 18972 3012
rect 19024 3000 19030 3052
rect 20254 3000 20260 3052
rect 20312 3000 20318 3052
rect 20346 3000 20352 3052
rect 20404 3000 20410 3052
rect 21634 3000 21640 3052
rect 21692 3000 21698 3052
rect 22094 3000 22100 3052
rect 22152 3000 22158 3052
rect 22278 3000 22284 3052
rect 22336 3040 22342 3052
rect 22741 3043 22799 3049
rect 22741 3040 22753 3043
rect 22336 3012 22753 3040
rect 22336 3000 22342 3012
rect 22741 3009 22753 3012
rect 22787 3009 22799 3043
rect 22741 3003 22799 3009
rect 22848 3012 25268 3040
rect 18414 2972 18420 2984
rect 17696 2944 18420 2972
rect 18414 2932 18420 2944
rect 18472 2932 18478 2984
rect 20901 2975 20959 2981
rect 18616 2944 18828 2972
rect 18616 2904 18644 2944
rect 17604 2876 18644 2904
rect 17276 2864 17282 2876
rect 18690 2864 18696 2916
rect 18748 2864 18754 2916
rect 18800 2904 18828 2944
rect 20901 2941 20913 2975
rect 20947 2941 20959 2975
rect 20901 2935 20959 2941
rect 21821 2975 21879 2981
rect 21821 2941 21833 2975
rect 21867 2972 21879 2975
rect 22848 2972 22876 3012
rect 25240 2984 25268 3012
rect 21867 2944 22876 2972
rect 21867 2941 21879 2944
rect 21821 2935 21879 2941
rect 20073 2907 20131 2913
rect 20073 2904 20085 2907
rect 18800 2876 20085 2904
rect 20073 2873 20085 2876
rect 20119 2873 20131 2907
rect 20073 2867 20131 2873
rect 7576 2808 8800 2836
rect 7285 2799 7343 2805
rect 10962 2796 10968 2848
rect 11020 2796 11026 2848
rect 12342 2796 12348 2848
rect 12400 2836 12406 2848
rect 12621 2839 12679 2845
rect 12621 2836 12633 2839
rect 12400 2808 12633 2836
rect 12400 2796 12406 2808
rect 12621 2805 12633 2808
rect 12667 2805 12679 2839
rect 12621 2799 12679 2805
rect 17037 2839 17095 2845
rect 17037 2805 17049 2839
rect 17083 2836 17095 2839
rect 17402 2836 17408 2848
rect 17083 2808 17408 2836
rect 17083 2805 17095 2808
rect 17037 2799 17095 2805
rect 17402 2796 17408 2808
rect 17460 2796 17466 2848
rect 17494 2796 17500 2848
rect 17552 2836 17558 2848
rect 17773 2839 17831 2845
rect 17773 2836 17785 2839
rect 17552 2808 17785 2836
rect 17552 2796 17558 2808
rect 17773 2805 17785 2808
rect 17819 2805 17831 2839
rect 17773 2799 17831 2805
rect 18141 2839 18199 2845
rect 18141 2805 18153 2839
rect 18187 2836 18199 2839
rect 19058 2836 19064 2848
rect 18187 2808 19064 2836
rect 18187 2805 18199 2808
rect 18141 2799 18199 2805
rect 19058 2796 19064 2808
rect 19116 2796 19122 2848
rect 19150 2796 19156 2848
rect 19208 2796 19214 2848
rect 19242 2796 19248 2848
rect 19300 2836 19306 2848
rect 19705 2839 19763 2845
rect 19705 2836 19717 2839
rect 19300 2808 19717 2836
rect 19300 2796 19306 2808
rect 19705 2805 19717 2808
rect 19751 2805 19763 2839
rect 19705 2799 19763 2805
rect 19794 2796 19800 2848
rect 19852 2836 19858 2848
rect 20916 2836 20944 2935
rect 23934 2932 23940 2984
rect 23992 2972 23998 2984
rect 24854 2972 24860 2984
rect 23992 2944 24860 2972
rect 23992 2932 23998 2944
rect 24854 2932 24860 2944
rect 24912 2932 24918 2984
rect 25222 2932 25228 2984
rect 25280 2932 25286 2984
rect 21266 2864 21272 2916
rect 21324 2904 21330 2916
rect 21324 2876 22094 2904
rect 21324 2864 21330 2876
rect 19852 2808 20944 2836
rect 22066 2836 22094 2876
rect 22186 2864 22192 2916
rect 22244 2904 22250 2916
rect 22738 2904 22744 2916
rect 22244 2876 22744 2904
rect 22244 2864 22250 2876
rect 22738 2864 22744 2876
rect 22796 2864 22802 2916
rect 23014 2836 23020 2848
rect 22066 2808 23020 2836
rect 19852 2796 19858 2808
rect 23014 2796 23020 2808
rect 23072 2796 23078 2848
rect 23474 2796 23480 2848
rect 23532 2836 23538 2848
rect 24121 2839 24179 2845
rect 24121 2836 24133 2839
rect 23532 2808 24133 2836
rect 23532 2796 23538 2808
rect 24121 2805 24133 2808
rect 24167 2805 24179 2839
rect 24121 2799 24179 2805
rect 1104 2746 24564 2768
rect 1104 2694 3882 2746
rect 3934 2694 3946 2746
rect 3998 2694 4010 2746
rect 4062 2694 4074 2746
rect 4126 2694 4138 2746
rect 4190 2694 9747 2746
rect 9799 2694 9811 2746
rect 9863 2694 9875 2746
rect 9927 2694 9939 2746
rect 9991 2694 10003 2746
rect 10055 2694 15612 2746
rect 15664 2694 15676 2746
rect 15728 2694 15740 2746
rect 15792 2694 15804 2746
rect 15856 2694 15868 2746
rect 15920 2694 21477 2746
rect 21529 2694 21541 2746
rect 21593 2694 21605 2746
rect 21657 2694 21669 2746
rect 21721 2694 21733 2746
rect 21785 2694 24564 2746
rect 1104 2672 24564 2694
rect 1762 2592 1768 2644
rect 1820 2592 1826 2644
rect 2682 2632 2688 2644
rect 2332 2604 2688 2632
rect 1486 2456 1492 2508
rect 1544 2496 1550 2508
rect 2332 2505 2360 2604
rect 2682 2592 2688 2604
rect 2740 2632 2746 2644
rect 2740 2604 3832 2632
rect 2740 2592 2746 2604
rect 3329 2567 3387 2573
rect 3329 2533 3341 2567
rect 3375 2564 3387 2567
rect 3694 2564 3700 2576
rect 3375 2536 3700 2564
rect 3375 2533 3387 2536
rect 3329 2527 3387 2533
rect 3694 2524 3700 2536
rect 3752 2524 3758 2576
rect 3804 2505 3832 2604
rect 5350 2592 5356 2644
rect 5408 2592 5414 2644
rect 5442 2592 5448 2644
rect 5500 2632 5506 2644
rect 6917 2635 6975 2641
rect 5500 2604 6592 2632
rect 5500 2592 5506 2604
rect 4614 2524 4620 2576
rect 4672 2564 4678 2576
rect 5813 2567 5871 2573
rect 5813 2564 5825 2567
rect 4672 2536 5825 2564
rect 4672 2524 4678 2536
rect 5813 2533 5825 2536
rect 5859 2533 5871 2567
rect 6564 2564 6592 2604
rect 6917 2601 6929 2635
rect 6963 2632 6975 2635
rect 7282 2632 7288 2644
rect 6963 2604 7288 2632
rect 6963 2601 6975 2604
rect 6917 2595 6975 2601
rect 7282 2592 7288 2604
rect 7340 2592 7346 2644
rect 9858 2632 9864 2644
rect 7392 2604 9864 2632
rect 7392 2564 7420 2604
rect 9858 2592 9864 2604
rect 9916 2592 9922 2644
rect 13446 2592 13452 2644
rect 13504 2592 13510 2644
rect 15841 2635 15899 2641
rect 15841 2601 15853 2635
rect 15887 2632 15899 2635
rect 16206 2632 16212 2644
rect 15887 2604 16212 2632
rect 15887 2601 15899 2604
rect 15841 2595 15899 2601
rect 16206 2592 16212 2604
rect 16264 2592 16270 2644
rect 17678 2632 17684 2644
rect 17328 2604 17684 2632
rect 6564 2536 7420 2564
rect 5813 2527 5871 2533
rect 7742 2524 7748 2576
rect 7800 2564 7806 2576
rect 8941 2567 8999 2573
rect 8941 2564 8953 2567
rect 7800 2536 8953 2564
rect 7800 2524 7806 2536
rect 8941 2533 8953 2536
rect 8987 2533 8999 2567
rect 8941 2527 8999 2533
rect 9122 2524 9128 2576
rect 9180 2524 9186 2576
rect 17328 2564 17356 2604
rect 17678 2592 17684 2604
rect 17736 2592 17742 2644
rect 17954 2592 17960 2644
rect 18012 2632 18018 2644
rect 18322 2632 18328 2644
rect 18012 2604 18328 2632
rect 18012 2592 18018 2604
rect 18322 2592 18328 2604
rect 18380 2592 18386 2644
rect 18506 2592 18512 2644
rect 18564 2632 18570 2644
rect 20254 2632 20260 2644
rect 18564 2604 19196 2632
rect 18564 2592 18570 2604
rect 19168 2576 19196 2604
rect 19352 2604 20260 2632
rect 16040 2536 17356 2564
rect 18693 2567 18751 2573
rect 2317 2499 2375 2505
rect 2317 2496 2329 2499
rect 1544 2468 2329 2496
rect 1544 2456 1550 2468
rect 2317 2465 2329 2468
rect 2363 2465 2375 2499
rect 2317 2459 2375 2465
rect 3789 2499 3847 2505
rect 3789 2465 3801 2499
rect 3835 2465 3847 2499
rect 3789 2459 3847 2465
rect 5902 2456 5908 2508
rect 5960 2456 5966 2508
rect 7561 2499 7619 2505
rect 7561 2465 7573 2499
rect 7607 2496 7619 2499
rect 9140 2496 9168 2524
rect 7607 2468 9168 2496
rect 10968 2508 11020 2514
rect 7607 2465 7619 2468
rect 7561 2459 7619 2465
rect 10968 2450 11020 2456
rect 11072 2468 11894 2496
rect 1673 2431 1731 2437
rect 1673 2397 1685 2431
rect 1719 2428 1731 2431
rect 2130 2428 2136 2440
rect 1719 2400 2136 2428
rect 1719 2397 1731 2400
rect 1673 2391 1731 2397
rect 2130 2388 2136 2400
rect 2188 2388 2194 2440
rect 2591 2431 2649 2437
rect 2591 2397 2603 2431
rect 2637 2397 2649 2431
rect 5166 2428 5172 2440
rect 4078 2407 5172 2428
rect 2591 2391 2649 2397
rect 4047 2401 5172 2407
rect 2406 2320 2412 2372
rect 2464 2360 2470 2372
rect 2606 2360 2634 2391
rect 4047 2367 4059 2401
rect 4093 2400 5172 2401
rect 4093 2370 4106 2400
rect 5166 2388 5172 2400
rect 5224 2388 5230 2440
rect 5629 2431 5687 2437
rect 5629 2397 5641 2431
rect 5675 2397 5687 2431
rect 6178 2428 6184 2440
rect 6139 2400 6184 2428
rect 5629 2391 5687 2397
rect 4093 2367 4105 2370
rect 4047 2361 4105 2367
rect 5261 2363 5319 2369
rect 2464 2332 2634 2360
rect 2464 2320 2470 2332
rect 5261 2329 5273 2363
rect 5307 2360 5319 2363
rect 5442 2360 5448 2372
rect 5307 2332 5448 2360
rect 5307 2329 5319 2332
rect 5261 2323 5319 2329
rect 5442 2320 5448 2332
rect 5500 2320 5506 2372
rect 5644 2360 5672 2391
rect 6178 2388 6184 2400
rect 6236 2388 6242 2440
rect 7650 2428 7656 2440
rect 6288 2400 7656 2428
rect 6288 2360 6316 2400
rect 7650 2388 7656 2400
rect 7708 2388 7714 2440
rect 8294 2388 8300 2440
rect 8352 2428 8358 2440
rect 8389 2431 8447 2437
rect 8389 2428 8401 2431
rect 8352 2400 8401 2428
rect 8352 2388 8358 2400
rect 8389 2397 8401 2400
rect 8435 2397 8447 2431
rect 8389 2391 8447 2397
rect 8662 2388 8668 2440
rect 8720 2388 8726 2440
rect 9122 2388 9128 2440
rect 9180 2388 9186 2440
rect 9398 2388 9404 2440
rect 9456 2388 9462 2440
rect 9677 2431 9735 2437
rect 9677 2397 9689 2431
rect 9723 2397 9735 2431
rect 9677 2391 9735 2397
rect 5644 2332 6316 2360
rect 6362 2320 6368 2372
rect 6420 2360 6426 2372
rect 7377 2363 7435 2369
rect 7377 2360 7389 2363
rect 6420 2332 7389 2360
rect 6420 2320 6426 2332
rect 7377 2329 7389 2332
rect 7423 2329 7435 2363
rect 7377 2323 7435 2329
rect 7745 2363 7803 2369
rect 7745 2329 7757 2363
rect 7791 2360 7803 2363
rect 7791 2332 8248 2360
rect 7791 2329 7803 2332
rect 7745 2323 7803 2329
rect 3418 2252 3424 2304
rect 3476 2292 3482 2304
rect 4801 2295 4859 2301
rect 4801 2292 4813 2295
rect 3476 2264 4813 2292
rect 3476 2252 3482 2264
rect 4801 2261 4813 2264
rect 4847 2261 4859 2295
rect 4801 2255 4859 2261
rect 5994 2252 6000 2304
rect 6052 2292 6058 2304
rect 7006 2292 7012 2304
rect 6052 2264 7012 2292
rect 6052 2252 6058 2264
rect 7006 2252 7012 2264
rect 7064 2252 7070 2304
rect 7466 2252 7472 2304
rect 7524 2292 7530 2304
rect 8220 2301 8248 2332
rect 8754 2320 8760 2372
rect 8812 2360 8818 2372
rect 9692 2360 9720 2391
rect 9858 2388 9864 2440
rect 9916 2428 9922 2440
rect 9916 2400 10640 2428
rect 9916 2388 9922 2400
rect 8812 2332 9720 2360
rect 8812 2320 8818 2332
rect 10226 2320 10232 2372
rect 10284 2320 10290 2372
rect 10321 2363 10379 2369
rect 10321 2329 10333 2363
rect 10367 2360 10379 2363
rect 10502 2360 10508 2372
rect 10367 2332 10508 2360
rect 10367 2329 10379 2332
rect 10321 2323 10379 2329
rect 10502 2320 10508 2332
rect 10560 2320 10566 2372
rect 10612 2360 10640 2400
rect 10686 2388 10692 2440
rect 10744 2388 10750 2440
rect 11072 2418 11100 2468
rect 11866 2428 11894 2468
rect 12342 2456 12348 2508
rect 12400 2456 12406 2508
rect 13906 2456 13912 2508
rect 13964 2456 13970 2508
rect 13817 2431 13875 2437
rect 10888 2390 11100 2418
rect 11348 2400 11836 2428
rect 11866 2400 13308 2428
rect 10888 2360 10916 2390
rect 11348 2360 11376 2400
rect 11808 2372 11836 2400
rect 10612 2332 10916 2360
rect 10980 2332 11376 2360
rect 7837 2295 7895 2301
rect 7837 2292 7849 2295
rect 7524 2264 7849 2292
rect 7524 2252 7530 2264
rect 7837 2261 7849 2264
rect 7883 2261 7895 2295
rect 7837 2255 7895 2261
rect 8205 2295 8263 2301
rect 8205 2261 8217 2295
rect 8251 2261 8263 2295
rect 8205 2255 8263 2261
rect 8478 2252 8484 2304
rect 8536 2252 8542 2304
rect 9214 2252 9220 2304
rect 9272 2252 9278 2304
rect 9306 2252 9312 2304
rect 9364 2292 9370 2304
rect 9493 2295 9551 2301
rect 9493 2292 9505 2295
rect 9364 2264 9505 2292
rect 9364 2252 9370 2264
rect 9493 2261 9505 2264
rect 9539 2261 9551 2295
rect 9493 2255 9551 2261
rect 9953 2295 10011 2301
rect 9953 2261 9965 2295
rect 9999 2292 10011 2295
rect 10980 2292 11008 2332
rect 11790 2320 11796 2372
rect 11848 2320 11854 2372
rect 11974 2320 11980 2372
rect 12032 2360 12038 2372
rect 12161 2363 12219 2369
rect 12161 2360 12173 2363
rect 12032 2332 12173 2360
rect 12032 2320 12038 2332
rect 12161 2329 12173 2332
rect 12207 2329 12219 2363
rect 12161 2323 12219 2329
rect 12433 2363 12491 2369
rect 12433 2329 12445 2363
rect 12479 2329 12491 2363
rect 12433 2323 12491 2329
rect 9999 2264 11008 2292
rect 9999 2261 10011 2264
rect 9953 2255 10011 2261
rect 11054 2252 11060 2304
rect 11112 2252 11118 2304
rect 11238 2252 11244 2304
rect 11296 2252 11302 2304
rect 11701 2295 11759 2301
rect 11701 2261 11713 2295
rect 11747 2292 11759 2295
rect 12452 2292 12480 2323
rect 12526 2320 12532 2372
rect 12584 2320 12590 2372
rect 12897 2363 12955 2369
rect 12897 2329 12909 2363
rect 12943 2360 12955 2363
rect 13078 2360 13084 2372
rect 12943 2332 13084 2360
rect 12943 2329 12955 2332
rect 12897 2323 12955 2329
rect 13078 2320 13084 2332
rect 13136 2320 13142 2372
rect 13170 2320 13176 2372
rect 13228 2320 13234 2372
rect 13280 2369 13308 2400
rect 13817 2397 13829 2431
rect 13863 2428 13875 2431
rect 13924 2428 13952 2456
rect 16040 2437 16068 2536
rect 18693 2533 18705 2567
rect 18739 2533 18751 2567
rect 18693 2527 18751 2533
rect 17034 2496 17040 2508
rect 16592 2468 17040 2496
rect 13863 2400 13952 2428
rect 16025 2431 16083 2437
rect 13863 2397 13875 2400
rect 13817 2391 13875 2397
rect 16025 2397 16037 2431
rect 16071 2397 16083 2431
rect 16025 2391 16083 2397
rect 16301 2431 16359 2437
rect 16301 2397 16313 2431
rect 16347 2428 16359 2431
rect 16482 2428 16488 2440
rect 16347 2400 16488 2428
rect 16347 2397 16359 2400
rect 16301 2391 16359 2397
rect 16482 2388 16488 2400
rect 16540 2388 16546 2440
rect 16592 2437 16620 2468
rect 17034 2456 17040 2468
rect 17092 2456 17098 2508
rect 18708 2496 18736 2527
rect 19150 2524 19156 2576
rect 19208 2524 19214 2576
rect 19352 2564 19380 2604
rect 20254 2592 20260 2604
rect 20312 2592 20318 2644
rect 20438 2592 20444 2644
rect 20496 2632 20502 2644
rect 21542 2632 21548 2644
rect 20496 2604 21548 2632
rect 20496 2592 20502 2604
rect 21542 2592 21548 2604
rect 21600 2632 21606 2644
rect 22278 2632 22284 2644
rect 21600 2604 22284 2632
rect 21600 2592 21606 2604
rect 22278 2592 22284 2604
rect 22336 2592 22342 2644
rect 23845 2635 23903 2641
rect 23845 2601 23857 2635
rect 23891 2632 23903 2635
rect 25314 2632 25320 2644
rect 23891 2604 25320 2632
rect 23891 2601 23903 2604
rect 23845 2595 23903 2601
rect 25314 2592 25320 2604
rect 25372 2592 25378 2644
rect 19260 2536 19380 2564
rect 19444 2536 20484 2564
rect 19260 2496 19288 2536
rect 19444 2496 19472 2536
rect 18708 2468 19288 2496
rect 19352 2468 19472 2496
rect 16577 2431 16635 2437
rect 16577 2397 16589 2431
rect 16623 2397 16635 2431
rect 16577 2391 16635 2397
rect 16850 2388 16856 2440
rect 16908 2388 16914 2440
rect 17126 2388 17132 2440
rect 17184 2388 17190 2440
rect 17313 2431 17371 2437
rect 17313 2397 17325 2431
rect 17359 2428 17371 2431
rect 18785 2431 18843 2437
rect 17359 2400 18368 2428
rect 17359 2397 17371 2400
rect 17313 2391 17371 2397
rect 13265 2363 13323 2369
rect 13265 2329 13277 2363
rect 13311 2329 13323 2363
rect 13265 2323 13323 2329
rect 15746 2320 15752 2372
rect 15804 2320 15810 2372
rect 16408 2332 17172 2360
rect 13188 2292 13216 2320
rect 11747 2264 13216 2292
rect 11747 2261 11759 2264
rect 11701 2255 11759 2261
rect 13354 2252 13360 2304
rect 13412 2292 13418 2304
rect 13633 2295 13691 2301
rect 13633 2292 13645 2295
rect 13412 2264 13645 2292
rect 13412 2252 13418 2264
rect 13633 2261 13645 2264
rect 13679 2261 13691 2295
rect 13633 2255 13691 2261
rect 16114 2252 16120 2304
rect 16172 2252 16178 2304
rect 16408 2301 16436 2332
rect 16393 2295 16451 2301
rect 16393 2261 16405 2295
rect 16439 2261 16451 2295
rect 16393 2255 16451 2261
rect 16666 2252 16672 2304
rect 16724 2252 16730 2304
rect 16942 2252 16948 2304
rect 17000 2252 17006 2304
rect 17144 2292 17172 2332
rect 17218 2320 17224 2372
rect 17276 2360 17282 2372
rect 17558 2363 17616 2369
rect 17558 2360 17570 2363
rect 17276 2332 17570 2360
rect 17276 2320 17282 2332
rect 17558 2329 17570 2332
rect 17604 2329 17616 2363
rect 18340 2360 18368 2400
rect 18785 2397 18797 2431
rect 18831 2428 18843 2431
rect 19352 2428 19380 2468
rect 19886 2456 19892 2508
rect 19944 2456 19950 2508
rect 20456 2496 20484 2536
rect 20622 2524 20628 2576
rect 20680 2564 20686 2576
rect 21913 2567 21971 2573
rect 21913 2564 21925 2567
rect 20680 2536 21925 2564
rect 20680 2524 20686 2536
rect 21913 2533 21925 2536
rect 21959 2533 21971 2567
rect 21913 2527 21971 2533
rect 22094 2524 22100 2576
rect 22152 2564 22158 2576
rect 24029 2567 24087 2573
rect 24029 2564 24041 2567
rect 22152 2536 24041 2564
rect 22152 2524 22158 2536
rect 24029 2533 24041 2536
rect 24075 2533 24087 2567
rect 24029 2527 24087 2533
rect 23014 2496 23020 2508
rect 20456 2468 23020 2496
rect 23014 2456 23020 2468
rect 23072 2456 23078 2508
rect 23293 2499 23351 2505
rect 23293 2465 23305 2499
rect 23339 2496 23351 2499
rect 23382 2496 23388 2508
rect 23339 2468 23388 2496
rect 23339 2465 23351 2468
rect 23293 2459 23351 2465
rect 23382 2456 23388 2468
rect 23440 2456 23446 2508
rect 18831 2400 19380 2428
rect 19429 2431 19487 2437
rect 18831 2397 18843 2400
rect 18785 2391 18843 2397
rect 19429 2397 19441 2431
rect 19475 2428 19487 2431
rect 19610 2428 19616 2440
rect 19475 2400 19616 2428
rect 19475 2397 19487 2400
rect 19429 2391 19487 2397
rect 19610 2388 19616 2400
rect 19668 2388 19674 2440
rect 19705 2431 19763 2437
rect 19705 2397 19717 2431
rect 19751 2428 19763 2431
rect 20806 2428 20812 2440
rect 19751 2400 20812 2428
rect 19751 2397 19763 2400
rect 19705 2391 19763 2397
rect 20806 2388 20812 2400
rect 20864 2388 20870 2440
rect 21818 2388 21824 2440
rect 21876 2428 21882 2440
rect 22557 2431 22615 2437
rect 22557 2428 22569 2431
rect 21876 2400 22569 2428
rect 21876 2388 21882 2400
rect 22557 2397 22569 2400
rect 22603 2397 22615 2431
rect 24213 2431 24271 2437
rect 24213 2428 24225 2431
rect 22557 2391 22615 2397
rect 22664 2400 24225 2428
rect 19334 2360 19340 2372
rect 18340 2332 19340 2360
rect 17558 2323 17616 2329
rect 19334 2320 19340 2332
rect 19392 2320 19398 2372
rect 20622 2320 20628 2372
rect 20680 2320 20686 2372
rect 20714 2320 20720 2372
rect 20772 2360 20778 2372
rect 21358 2360 21364 2372
rect 20772 2332 21364 2360
rect 20772 2320 20778 2332
rect 21358 2320 21364 2332
rect 21416 2360 21422 2372
rect 22664 2360 22692 2400
rect 24213 2397 24225 2400
rect 24259 2397 24271 2431
rect 24213 2391 24271 2397
rect 21416 2332 22692 2360
rect 23753 2363 23811 2369
rect 21416 2320 21422 2332
rect 23753 2329 23765 2363
rect 23799 2360 23811 2363
rect 24118 2360 24124 2372
rect 23799 2332 24124 2360
rect 23799 2329 23811 2332
rect 23753 2323 23811 2329
rect 24118 2320 24124 2332
rect 24176 2320 24182 2372
rect 17954 2292 17960 2304
rect 17144 2264 17960 2292
rect 17954 2252 17960 2264
rect 18012 2252 18018 2304
rect 18598 2252 18604 2304
rect 18656 2292 18662 2304
rect 18969 2295 19027 2301
rect 18969 2292 18981 2295
rect 18656 2264 18981 2292
rect 18656 2252 18662 2264
rect 18969 2261 18981 2264
rect 19015 2261 19027 2295
rect 18969 2255 19027 2261
rect 19150 2252 19156 2304
rect 19208 2292 19214 2304
rect 19245 2295 19303 2301
rect 19245 2292 19257 2295
rect 19208 2264 19257 2292
rect 19208 2252 19214 2264
rect 19245 2261 19257 2264
rect 19291 2261 19303 2295
rect 19245 2255 19303 2261
rect 1104 2202 24723 2224
rect 1104 2150 6814 2202
rect 6866 2150 6878 2202
rect 6930 2150 6942 2202
rect 6994 2150 7006 2202
rect 7058 2150 7070 2202
rect 7122 2150 12679 2202
rect 12731 2150 12743 2202
rect 12795 2150 12807 2202
rect 12859 2150 12871 2202
rect 12923 2150 12935 2202
rect 12987 2150 18544 2202
rect 18596 2150 18608 2202
rect 18660 2150 18672 2202
rect 18724 2150 18736 2202
rect 18788 2150 18800 2202
rect 18852 2150 24409 2202
rect 24461 2150 24473 2202
rect 24525 2150 24537 2202
rect 24589 2150 24601 2202
rect 24653 2150 24665 2202
rect 24717 2150 24723 2202
rect 1104 2128 24723 2150
rect 25406 2116 25412 2168
rect 25464 2116 25470 2168
rect 3786 2048 3792 2100
rect 3844 2088 3850 2100
rect 3881 2091 3939 2097
rect 3881 2088 3893 2091
rect 3844 2060 3893 2088
rect 3844 2048 3850 2060
rect 3881 2057 3893 2060
rect 3927 2057 3939 2091
rect 3881 2051 3939 2057
rect 4890 2048 4896 2100
rect 4948 2088 4954 2100
rect 5261 2091 5319 2097
rect 5261 2088 5273 2091
rect 4948 2060 5273 2088
rect 4948 2048 4954 2060
rect 5261 2057 5273 2060
rect 5307 2057 5319 2091
rect 5261 2051 5319 2057
rect 6086 2048 6092 2100
rect 6144 2048 6150 2100
rect 6638 2088 6644 2100
rect 6194 2060 6644 2088
rect 1489 2023 1547 2029
rect 1489 1989 1501 2023
rect 1535 2020 1547 2023
rect 1670 2020 1676 2032
rect 1535 1992 1676 2020
rect 1535 1989 1547 1992
rect 1489 1983 1547 1989
rect 1670 1980 1676 1992
rect 1728 1980 1734 2032
rect 1857 2023 1915 2029
rect 1857 1989 1869 2023
rect 1903 2020 1915 2023
rect 2774 2020 2780 2032
rect 1903 1992 2780 2020
rect 1903 1989 1915 1992
rect 1857 1983 1915 1989
rect 2774 1980 2780 1992
rect 2832 1980 2838 2032
rect 6194 2020 6222 2060
rect 6638 2048 6644 2060
rect 6696 2048 6702 2100
rect 6917 2091 6975 2097
rect 6917 2057 6929 2091
rect 6963 2088 6975 2091
rect 7282 2088 7288 2100
rect 6963 2060 7288 2088
rect 6963 2057 6975 2060
rect 6917 2051 6975 2057
rect 7282 2048 7288 2060
rect 7340 2048 7346 2100
rect 7650 2048 7656 2100
rect 7708 2048 7714 2100
rect 7742 2048 7748 2100
rect 7800 2048 7806 2100
rect 8021 2091 8079 2097
rect 8021 2057 8033 2091
rect 8067 2088 8079 2091
rect 8110 2088 8116 2100
rect 8067 2060 8116 2088
rect 8067 2057 8079 2060
rect 8021 2051 8079 2057
rect 8110 2048 8116 2060
rect 8168 2048 8174 2100
rect 8757 2091 8815 2097
rect 8757 2057 8769 2091
rect 8803 2088 8815 2091
rect 8846 2088 8852 2100
rect 8803 2060 8852 2088
rect 8803 2057 8815 2060
rect 8757 2051 8815 2057
rect 8846 2048 8852 2060
rect 8904 2048 8910 2100
rect 9214 2048 9220 2100
rect 9272 2048 9278 2100
rect 9508 2060 10732 2088
rect 2884 1992 4292 2020
rect 2225 1955 2283 1961
rect 2225 1921 2237 1955
rect 2271 1921 2283 1955
rect 2225 1915 2283 1921
rect 934 1844 940 1896
rect 992 1884 998 1896
rect 2240 1884 2268 1915
rect 2682 1912 2688 1964
rect 2740 1952 2746 1964
rect 2884 1961 2912 1992
rect 2869 1955 2927 1961
rect 2869 1952 2881 1955
rect 2740 1924 2881 1952
rect 2740 1912 2746 1924
rect 2869 1921 2881 1924
rect 2915 1921 2927 1955
rect 2869 1915 2927 1921
rect 3143 1955 3201 1961
rect 3143 1921 3155 1955
rect 3189 1952 3201 1955
rect 3970 1952 3976 1964
rect 3189 1924 3976 1952
rect 3189 1921 3201 1924
rect 3143 1915 3201 1921
rect 3970 1912 3976 1924
rect 4028 1912 4034 1964
rect 4264 1961 4292 1992
rect 4538 1992 6222 2020
rect 4538 1961 4566 1992
rect 6454 1980 6460 2032
rect 6512 1980 6518 2032
rect 6730 1980 6736 2032
rect 6788 1980 6794 2032
rect 6825 2023 6883 2029
rect 6825 1989 6837 2023
rect 6871 1989 6883 2023
rect 6825 1983 6883 1989
rect 7561 2023 7619 2029
rect 7561 1989 7573 2023
rect 7607 2020 7619 2023
rect 7760 2020 7788 2048
rect 7607 1992 7788 2020
rect 7929 2023 7987 2029
rect 7607 1989 7619 1992
rect 7561 1983 7619 1989
rect 7929 1989 7941 2023
rect 7975 2020 7987 2023
rect 9232 2020 9260 2048
rect 7975 1992 9260 2020
rect 7975 1989 7987 1992
rect 7929 1983 7987 1989
rect 4249 1955 4307 1961
rect 4249 1921 4261 1955
rect 4295 1921 4307 1955
rect 4249 1915 4307 1921
rect 4523 1955 4581 1961
rect 4523 1921 4535 1955
rect 4569 1921 4581 1955
rect 4523 1915 4581 1921
rect 5350 1912 5356 1964
rect 5408 1952 5414 1964
rect 5813 1955 5871 1961
rect 5813 1952 5825 1955
rect 5408 1924 5825 1952
rect 5408 1912 5414 1924
rect 5813 1921 5825 1924
rect 5859 1921 5871 1955
rect 5813 1915 5871 1921
rect 5997 1955 6055 1961
rect 5997 1921 6009 1955
rect 6043 1952 6055 1955
rect 6748 1952 6776 1980
rect 6043 1924 6776 1952
rect 6043 1921 6055 1924
rect 5997 1915 6055 1921
rect 992 1856 2268 1884
rect 992 1844 998 1856
rect 2501 1819 2559 1825
rect 2501 1785 2513 1819
rect 2547 1785 2559 1819
rect 2501 1779 2559 1785
rect 5629 1819 5687 1825
rect 5629 1785 5641 1819
rect 5675 1816 5687 1819
rect 6840 1816 6868 1983
rect 7193 1955 7251 1961
rect 7193 1921 7205 1955
rect 7239 1921 7251 1955
rect 7193 1915 7251 1921
rect 7377 1955 7435 1961
rect 7377 1921 7389 1955
rect 7423 1952 7435 1955
rect 8018 1952 8024 1964
rect 7423 1924 8024 1952
rect 7423 1921 7435 1924
rect 7377 1915 7435 1921
rect 7208 1884 7236 1915
rect 8018 1912 8024 1924
rect 8076 1912 8082 1964
rect 8205 1955 8263 1961
rect 8205 1921 8217 1955
rect 8251 1952 8263 1955
rect 8386 1952 8392 1964
rect 8251 1924 8392 1952
rect 8251 1921 8263 1924
rect 8205 1915 8263 1921
rect 8386 1912 8392 1924
rect 8444 1912 8450 1964
rect 8478 1912 8484 1964
rect 8536 1912 8542 1964
rect 8665 1955 8723 1961
rect 8665 1921 8677 1955
rect 8711 1952 8723 1955
rect 9508 1952 9536 2060
rect 10042 1980 10048 2032
rect 10100 2020 10106 2032
rect 10704 2020 10732 2060
rect 10778 2048 10784 2100
rect 10836 2088 10842 2100
rect 11057 2091 11115 2097
rect 11057 2088 11069 2091
rect 10836 2060 11069 2088
rect 10836 2048 10842 2060
rect 11057 2057 11069 2060
rect 11103 2057 11115 2091
rect 11057 2051 11115 2057
rect 11330 2048 11336 2100
rect 11388 2088 11394 2100
rect 11388 2060 11744 2088
rect 11388 2048 11394 2060
rect 11606 2020 11612 2032
rect 10100 1992 10178 2020
rect 10704 1992 11612 2020
rect 10100 1980 10106 1992
rect 10150 1962 10178 1992
rect 11606 1980 11612 1992
rect 11664 1980 11670 2032
rect 10287 1965 10345 1971
rect 10287 1962 10299 1965
rect 8711 1924 9536 1952
rect 9585 1955 9643 1961
rect 8711 1921 8723 1924
rect 8665 1915 8723 1921
rect 9585 1921 9597 1955
rect 9631 1921 9643 1955
rect 10150 1934 10299 1962
rect 10287 1931 10299 1934
rect 10333 1931 10345 1965
rect 10287 1925 10345 1931
rect 9585 1915 9643 1921
rect 8496 1884 8524 1912
rect 7208 1856 8524 1884
rect 9217 1887 9275 1893
rect 9217 1853 9229 1887
rect 9263 1884 9275 1887
rect 9490 1884 9496 1896
rect 9263 1856 9496 1884
rect 9263 1853 9275 1856
rect 9217 1847 9275 1853
rect 9490 1844 9496 1856
rect 9548 1884 9554 1896
rect 9600 1884 9628 1915
rect 11514 1912 11520 1964
rect 11572 1912 11578 1964
rect 11716 1961 11744 2060
rect 12526 2048 12532 2100
rect 12584 2088 12590 2100
rect 13357 2091 13415 2097
rect 13357 2088 13369 2091
rect 12584 2060 13369 2088
rect 12584 2048 12590 2060
rect 13357 2057 13369 2060
rect 13403 2057 13415 2091
rect 13357 2051 13415 2057
rect 14458 2048 14464 2100
rect 14516 2048 14522 2100
rect 16666 2048 16672 2100
rect 16724 2048 16730 2100
rect 16942 2048 16948 2100
rect 17000 2088 17006 2100
rect 17000 2060 18920 2088
rect 17000 2048 17006 2060
rect 11882 1980 11888 2032
rect 11940 1980 11946 2032
rect 13262 2020 13268 2032
rect 12802 1992 13268 2020
rect 12603 1985 12661 1991
rect 12603 1982 12615 1985
rect 11701 1955 11759 1961
rect 11701 1921 11713 1955
rect 11747 1921 11759 1955
rect 11701 1915 11759 1921
rect 12250 1912 12256 1964
rect 12308 1952 12314 1964
rect 12544 1954 12615 1982
rect 12544 1952 12572 1954
rect 12308 1924 12572 1952
rect 12603 1951 12615 1954
rect 12649 1982 12661 1985
rect 12802 1982 12830 1992
rect 12649 1954 12830 1982
rect 13262 1980 13268 1992
rect 13320 1980 13326 2032
rect 13909 1955 13967 1961
rect 12649 1951 12661 1954
rect 12603 1945 12661 1951
rect 12308 1912 12314 1924
rect 13909 1921 13921 1955
rect 13955 1921 13967 1955
rect 14476 1952 14504 2048
rect 15378 1980 15384 2032
rect 15436 2020 15442 2032
rect 15473 2023 15531 2029
rect 15473 2020 15485 2023
rect 15436 1992 15485 2020
rect 15436 1980 15442 1992
rect 15473 1989 15485 1992
rect 15519 1989 15531 2023
rect 16684 2020 16712 2048
rect 16761 2023 16819 2029
rect 16761 2020 16773 2023
rect 16684 1992 16773 2020
rect 15473 1983 15531 1989
rect 16761 1989 16773 1992
rect 16807 1989 16819 2023
rect 16761 1983 16819 1989
rect 17126 1980 17132 2032
rect 17184 2020 17190 2032
rect 17313 2023 17371 2029
rect 17313 2020 17325 2023
rect 17184 1992 17325 2020
rect 17184 1980 17190 1992
rect 17313 1989 17325 1992
rect 17359 1989 17371 2023
rect 17313 1983 17371 1989
rect 17402 1980 17408 2032
rect 17460 2020 17466 2032
rect 17865 2023 17923 2029
rect 17865 2020 17877 2023
rect 17460 1992 17877 2020
rect 17460 1980 17466 1992
rect 17865 1989 17877 1992
rect 17911 1989 17923 2023
rect 17865 1983 17923 1989
rect 17954 1980 17960 2032
rect 18012 2020 18018 2032
rect 18417 2023 18475 2029
rect 18417 2020 18429 2023
rect 18012 1992 18429 2020
rect 18012 1980 18018 1992
rect 18417 1989 18429 1992
rect 18463 1989 18475 2023
rect 18417 1983 18475 1989
rect 14829 1955 14887 1961
rect 14829 1952 14841 1955
rect 14476 1924 14841 1952
rect 13909 1915 13967 1921
rect 14829 1921 14841 1924
rect 14875 1921 14887 1955
rect 14829 1915 14887 1921
rect 9548 1856 9628 1884
rect 9548 1844 9554 1856
rect 10042 1844 10048 1896
rect 10100 1844 10106 1896
rect 11532 1884 11560 1912
rect 12345 1887 12403 1893
rect 12345 1884 12357 1887
rect 11532 1856 12357 1884
rect 12345 1853 12357 1856
rect 12391 1853 12403 1887
rect 12345 1847 12403 1853
rect 7926 1816 7932 1828
rect 5675 1788 6776 1816
rect 6840 1788 7932 1816
rect 5675 1785 5687 1788
rect 5629 1779 5687 1785
rect 2516 1748 2544 1779
rect 3602 1748 3608 1760
rect 2516 1720 3608 1748
rect 3602 1708 3608 1720
rect 3660 1708 3666 1760
rect 4982 1708 4988 1760
rect 5040 1748 5046 1760
rect 6549 1751 6607 1757
rect 6549 1748 6561 1751
rect 5040 1720 6561 1748
rect 5040 1708 5046 1720
rect 6549 1717 6561 1720
rect 6595 1717 6607 1751
rect 6748 1748 6776 1788
rect 7926 1776 7932 1788
rect 7984 1776 7990 1828
rect 8386 1776 8392 1828
rect 8444 1776 8450 1828
rect 8478 1776 8484 1828
rect 8536 1816 8542 1828
rect 9674 1816 9680 1828
rect 8536 1788 9680 1816
rect 8536 1776 8542 1788
rect 9674 1776 9680 1788
rect 9732 1776 9738 1828
rect 9950 1816 9956 1828
rect 9784 1788 9956 1816
rect 9784 1748 9812 1788
rect 9950 1776 9956 1788
rect 10008 1776 10014 1828
rect 10778 1776 10784 1828
rect 10836 1816 10842 1828
rect 13924 1816 13952 1915
rect 16022 1912 16028 1964
rect 16080 1912 16086 1964
rect 16298 1912 16304 1964
rect 16356 1952 16362 1964
rect 18892 1961 18920 2060
rect 19058 2048 19064 2100
rect 19116 2048 19122 2100
rect 19886 2088 19892 2100
rect 19168 2060 19892 2088
rect 18785 1955 18843 1961
rect 18785 1952 18797 1955
rect 16356 1924 18797 1952
rect 16356 1912 16362 1924
rect 18785 1921 18797 1924
rect 18831 1921 18843 1955
rect 18785 1915 18843 1921
rect 18877 1955 18935 1961
rect 18877 1921 18889 1955
rect 18923 1921 18935 1955
rect 18877 1915 18935 1921
rect 18141 1887 18199 1893
rect 18141 1853 18153 1887
rect 18187 1884 18199 1887
rect 18230 1884 18236 1896
rect 18187 1856 18236 1884
rect 18187 1853 18199 1856
rect 18141 1847 18199 1853
rect 18230 1844 18236 1856
rect 18288 1844 18294 1896
rect 18322 1844 18328 1896
rect 18380 1884 18386 1896
rect 19168 1884 19196 2060
rect 19886 2048 19892 2060
rect 19944 2048 19950 2100
rect 20070 2048 20076 2100
rect 20128 2088 20134 2100
rect 20625 2091 20683 2097
rect 20625 2088 20637 2091
rect 20128 2060 20637 2088
rect 20128 2048 20134 2060
rect 20625 2057 20637 2060
rect 20671 2057 20683 2091
rect 23201 2091 23259 2097
rect 23201 2088 23213 2091
rect 20625 2051 20683 2057
rect 20732 2060 23213 2088
rect 19978 2020 19984 2032
rect 19444 1992 19984 2020
rect 19245 1955 19303 1961
rect 19245 1921 19257 1955
rect 19291 1952 19303 1955
rect 19334 1952 19340 1964
rect 19291 1924 19340 1952
rect 19291 1921 19303 1924
rect 19245 1915 19303 1921
rect 19334 1912 19340 1924
rect 19392 1952 19398 1964
rect 19444 1952 19472 1992
rect 19978 1980 19984 1992
rect 20036 1980 20042 2032
rect 20162 1980 20168 2032
rect 20220 2020 20226 2032
rect 20732 2020 20760 2060
rect 23201 2057 23213 2060
rect 23247 2057 23259 2091
rect 23201 2051 23259 2057
rect 23658 2048 23664 2100
rect 23716 2088 23722 2100
rect 24029 2091 24087 2097
rect 24029 2088 24041 2091
rect 23716 2060 24041 2088
rect 23716 2048 23722 2060
rect 24029 2057 24041 2060
rect 24075 2057 24087 2091
rect 24029 2051 24087 2057
rect 20220 1992 20760 2020
rect 20220 1980 20226 1992
rect 20898 1980 20904 2032
rect 20956 2020 20962 2032
rect 22066 2023 22124 2029
rect 22066 2020 22078 2023
rect 20956 1992 22078 2020
rect 20956 1980 20962 1992
rect 22066 1989 22078 1992
rect 22112 1989 22124 2023
rect 25424 2020 25452 2116
rect 22066 1983 22124 1989
rect 22204 1992 25452 2020
rect 19392 1924 19472 1952
rect 19512 1955 19570 1961
rect 19392 1912 19398 1924
rect 19512 1921 19524 1955
rect 19558 1952 19570 1955
rect 21821 1955 21879 1961
rect 21821 1952 21833 1955
rect 19558 1924 20392 1952
rect 19558 1921 19570 1924
rect 19512 1915 19570 1921
rect 18380 1856 19196 1884
rect 20364 1884 20392 1924
rect 21560 1924 21833 1952
rect 21560 1896 21588 1924
rect 21821 1921 21833 1924
rect 21867 1921 21879 1955
rect 22204 1952 22232 1992
rect 21821 1915 21879 1921
rect 21928 1924 22232 1952
rect 20714 1884 20720 1896
rect 20364 1856 20720 1884
rect 18380 1844 18386 1856
rect 20714 1844 20720 1856
rect 20772 1844 20778 1896
rect 20809 1887 20867 1893
rect 20809 1853 20821 1887
rect 20855 1853 20867 1887
rect 20809 1847 20867 1853
rect 10836 1788 12434 1816
rect 10836 1776 10842 1788
rect 6748 1720 9812 1748
rect 9861 1751 9919 1757
rect 6549 1711 6607 1717
rect 9861 1717 9873 1751
rect 9907 1748 9919 1751
rect 10502 1748 10508 1760
rect 9907 1720 10508 1748
rect 9907 1717 9919 1720
rect 9861 1711 9919 1717
rect 10502 1708 10508 1720
rect 10560 1708 10566 1760
rect 11517 1751 11575 1757
rect 11517 1717 11529 1751
rect 11563 1748 11575 1751
rect 11790 1748 11796 1760
rect 11563 1720 11796 1748
rect 11563 1717 11575 1720
rect 11517 1711 11575 1717
rect 11790 1708 11796 1720
rect 11848 1708 11854 1760
rect 11974 1708 11980 1760
rect 12032 1708 12038 1760
rect 12406 1748 12434 1788
rect 13188 1788 13952 1816
rect 13188 1748 13216 1788
rect 16666 1776 16672 1828
rect 16724 1816 16730 1828
rect 19058 1816 19064 1828
rect 16724 1788 19064 1816
rect 16724 1776 16730 1788
rect 19058 1776 19064 1788
rect 19116 1776 19122 1828
rect 12406 1720 13216 1748
rect 13722 1708 13728 1760
rect 13780 1708 13786 1760
rect 14182 1708 14188 1760
rect 14240 1748 14246 1760
rect 15013 1751 15071 1757
rect 15013 1748 15025 1751
rect 14240 1720 15025 1748
rect 14240 1708 14246 1720
rect 15013 1717 15025 1720
rect 15059 1717 15071 1751
rect 15013 1711 15071 1717
rect 15286 1708 15292 1760
rect 15344 1748 15350 1760
rect 15565 1751 15623 1757
rect 15565 1748 15577 1751
rect 15344 1720 15577 1748
rect 15344 1708 15350 1720
rect 15565 1717 15577 1720
rect 15611 1717 15623 1751
rect 15565 1711 15623 1717
rect 15930 1708 15936 1760
rect 15988 1748 15994 1760
rect 16117 1751 16175 1757
rect 16117 1748 16129 1751
rect 15988 1720 16129 1748
rect 15988 1708 15994 1720
rect 16117 1717 16129 1720
rect 16163 1717 16175 1751
rect 16117 1711 16175 1717
rect 16390 1708 16396 1760
rect 16448 1748 16454 1760
rect 16853 1751 16911 1757
rect 16853 1748 16865 1751
rect 16448 1720 16865 1748
rect 16448 1708 16454 1720
rect 16853 1717 16865 1720
rect 16899 1717 16911 1751
rect 16853 1711 16911 1717
rect 16942 1708 16948 1760
rect 17000 1748 17006 1760
rect 17405 1751 17463 1757
rect 17405 1748 17417 1751
rect 17000 1720 17417 1748
rect 17000 1708 17006 1720
rect 17405 1717 17417 1720
rect 17451 1717 17463 1751
rect 17405 1711 17463 1717
rect 17678 1708 17684 1760
rect 17736 1748 17742 1760
rect 20162 1748 20168 1760
rect 17736 1720 20168 1748
rect 17736 1708 17742 1720
rect 20162 1708 20168 1720
rect 20220 1708 20226 1760
rect 20824 1748 20852 1847
rect 21082 1844 21088 1896
rect 21140 1844 21146 1896
rect 21542 1844 21548 1896
rect 21600 1844 21606 1896
rect 21928 1884 21956 1924
rect 23750 1912 23756 1964
rect 23808 1952 23814 1964
rect 24213 1955 24271 1961
rect 24213 1952 24225 1955
rect 23808 1924 24225 1952
rect 23808 1912 23814 1924
rect 24213 1921 24225 1924
rect 24259 1921 24271 1955
rect 24213 1915 24271 1921
rect 21836 1856 21956 1884
rect 20898 1776 20904 1828
rect 20956 1816 20962 1828
rect 21836 1816 21864 1856
rect 20956 1788 21864 1816
rect 20956 1776 20962 1788
rect 24670 1748 24676 1760
rect 20824 1720 24676 1748
rect 24670 1708 24676 1720
rect 24728 1708 24734 1760
rect 1104 1658 24564 1680
rect 1104 1606 3882 1658
rect 3934 1606 3946 1658
rect 3998 1606 4010 1658
rect 4062 1606 4074 1658
rect 4126 1606 4138 1658
rect 4190 1606 9747 1658
rect 9799 1606 9811 1658
rect 9863 1606 9875 1658
rect 9927 1606 9939 1658
rect 9991 1606 10003 1658
rect 10055 1606 15612 1658
rect 15664 1606 15676 1658
rect 15728 1606 15740 1658
rect 15792 1606 15804 1658
rect 15856 1606 15868 1658
rect 15920 1606 21477 1658
rect 21529 1606 21541 1658
rect 21593 1606 21605 1658
rect 21657 1606 21669 1658
rect 21721 1606 21733 1658
rect 21785 1606 24564 1658
rect 1104 1584 24564 1606
rect 14 1504 20 1556
rect 72 1544 78 1556
rect 6086 1544 6092 1556
rect 72 1516 6092 1544
rect 72 1504 78 1516
rect 6086 1504 6092 1516
rect 6144 1504 6150 1556
rect 8478 1504 8484 1556
rect 8536 1504 8542 1556
rect 8665 1547 8723 1553
rect 8665 1513 8677 1547
rect 8711 1544 8723 1547
rect 9309 1547 9367 1553
rect 8711 1516 9260 1544
rect 8711 1513 8723 1516
rect 8665 1507 8723 1513
rect 1118 1436 1124 1488
rect 1176 1476 1182 1488
rect 4982 1476 4988 1488
rect 1176 1448 4988 1476
rect 1176 1436 1182 1448
rect 4982 1436 4988 1448
rect 5040 1436 5046 1488
rect 6181 1479 6239 1485
rect 6181 1445 6193 1479
rect 6227 1476 6239 1479
rect 6270 1476 6276 1488
rect 6227 1448 6276 1476
rect 6227 1445 6239 1448
rect 6181 1439 6239 1445
rect 6270 1436 6276 1448
rect 6328 1436 6334 1488
rect 3252 1380 3464 1408
rect 566 1300 572 1352
rect 624 1340 630 1352
rect 1489 1343 1547 1349
rect 1489 1340 1501 1343
rect 624 1312 1501 1340
rect 624 1300 630 1312
rect 1489 1309 1501 1312
rect 1535 1309 1547 1343
rect 1489 1303 1547 1309
rect 2225 1343 2283 1349
rect 2225 1309 2237 1343
rect 2271 1309 2283 1343
rect 2225 1303 2283 1309
rect 2593 1343 2651 1349
rect 2593 1309 2605 1343
rect 2639 1340 2651 1343
rect 3252 1340 3280 1380
rect 2639 1312 3280 1340
rect 2639 1309 2651 1312
rect 2593 1303 2651 1309
rect 1026 1232 1032 1284
rect 1084 1232 1090 1284
rect 1946 1232 1952 1284
rect 2004 1232 2010 1284
rect 2240 1272 2268 1303
rect 3326 1300 3332 1352
rect 3384 1300 3390 1352
rect 3436 1340 3464 1380
rect 3602 1368 3608 1420
rect 3660 1408 3666 1420
rect 8496 1408 8524 1504
rect 9232 1476 9260 1516
rect 9309 1513 9321 1547
rect 9355 1544 9367 1547
rect 9490 1544 9496 1556
rect 9355 1516 9496 1544
rect 9355 1513 9367 1516
rect 9309 1507 9367 1513
rect 9490 1504 9496 1516
rect 9548 1504 9554 1556
rect 10597 1547 10655 1553
rect 9692 1516 10548 1544
rect 9692 1476 9720 1516
rect 9232 1448 9720 1476
rect 10520 1476 10548 1516
rect 10597 1513 10609 1547
rect 10643 1544 10655 1547
rect 10962 1544 10968 1556
rect 10643 1516 10968 1544
rect 10643 1513 10655 1516
rect 10597 1507 10655 1513
rect 10962 1504 10968 1516
rect 11020 1504 11026 1556
rect 11238 1504 11244 1556
rect 11296 1504 11302 1556
rect 11606 1504 11612 1556
rect 11664 1544 11670 1556
rect 13722 1544 13728 1556
rect 11664 1516 13728 1544
rect 11664 1504 11670 1516
rect 13722 1504 13728 1516
rect 13780 1504 13786 1556
rect 14458 1504 14464 1556
rect 14516 1544 14522 1556
rect 15381 1547 15439 1553
rect 15381 1544 15393 1547
rect 14516 1516 15393 1544
rect 14516 1504 14522 1516
rect 15381 1513 15393 1516
rect 15427 1513 15439 1547
rect 15381 1507 15439 1513
rect 15933 1547 15991 1553
rect 15933 1513 15945 1547
rect 15979 1513 15991 1547
rect 15933 1507 15991 1513
rect 11146 1476 11152 1488
rect 10520 1448 11152 1476
rect 11146 1436 11152 1448
rect 11204 1436 11210 1488
rect 13630 1436 13636 1488
rect 13688 1476 13694 1488
rect 14737 1479 14795 1485
rect 14737 1476 14749 1479
rect 13688 1448 14749 1476
rect 13688 1436 13694 1448
rect 14737 1445 14749 1448
rect 14783 1445 14795 1479
rect 14737 1439 14795 1445
rect 14918 1436 14924 1488
rect 14976 1476 14982 1488
rect 15948 1476 15976 1507
rect 16022 1504 16028 1556
rect 16080 1544 16086 1556
rect 16301 1547 16359 1553
rect 16301 1544 16313 1547
rect 16080 1516 16313 1544
rect 16080 1504 16086 1516
rect 16301 1513 16313 1516
rect 16347 1513 16359 1547
rect 16301 1507 16359 1513
rect 16482 1504 16488 1556
rect 16540 1544 16546 1556
rect 20898 1544 20904 1556
rect 16540 1516 20904 1544
rect 16540 1504 16546 1516
rect 20898 1504 20904 1516
rect 20956 1504 20962 1556
rect 23106 1504 23112 1556
rect 23164 1504 23170 1556
rect 23845 1547 23903 1553
rect 23845 1513 23857 1547
rect 23891 1544 23903 1547
rect 25130 1544 25136 1556
rect 23891 1516 25136 1544
rect 23891 1513 23903 1516
rect 23845 1507 23903 1513
rect 25130 1504 25136 1516
rect 25188 1504 25194 1556
rect 14976 1448 15976 1476
rect 17497 1479 17555 1485
rect 14976 1436 14982 1448
rect 17497 1445 17509 1479
rect 17543 1445 17555 1479
rect 17497 1439 17555 1445
rect 3660 1380 8524 1408
rect 9585 1411 9643 1417
rect 3660 1368 3666 1380
rect 9585 1377 9597 1411
rect 9631 1377 9643 1411
rect 9585 1371 9643 1377
rect 3694 1340 3700 1352
rect 3436 1312 3700 1340
rect 3694 1300 3700 1312
rect 3752 1300 3758 1352
rect 3786 1300 3792 1352
rect 3844 1300 3850 1352
rect 3970 1300 3976 1352
rect 4028 1340 4034 1352
rect 4157 1343 4215 1349
rect 4157 1340 4169 1343
rect 4028 1312 4169 1340
rect 4028 1300 4034 1312
rect 4157 1309 4169 1312
rect 4203 1309 4215 1343
rect 4157 1303 4215 1309
rect 4430 1300 4436 1352
rect 4488 1300 4494 1352
rect 5810 1300 5816 1352
rect 5868 1300 5874 1352
rect 5994 1300 6000 1352
rect 6052 1300 6058 1352
rect 6086 1300 6092 1352
rect 6144 1340 6150 1352
rect 6365 1343 6423 1349
rect 6365 1340 6377 1343
rect 6144 1312 6377 1340
rect 6144 1300 6150 1312
rect 6365 1309 6377 1312
rect 6411 1309 6423 1343
rect 6365 1303 6423 1309
rect 6638 1300 6644 1352
rect 6696 1300 6702 1352
rect 7285 1343 7343 1349
rect 7285 1309 7297 1343
rect 7331 1309 7343 1343
rect 7285 1303 7343 1309
rect 7561 1343 7619 1349
rect 7561 1309 7573 1343
rect 7607 1309 7619 1343
rect 7561 1303 7619 1309
rect 2866 1272 2872 1284
rect 2240 1244 2872 1272
rect 2866 1232 2872 1244
rect 2924 1232 2930 1284
rect 3053 1275 3111 1281
rect 3053 1241 3065 1275
rect 3099 1272 3111 1275
rect 4246 1272 4252 1284
rect 3099 1244 4252 1272
rect 3099 1241 3111 1244
rect 3053 1235 3111 1241
rect 4246 1232 4252 1244
rect 4304 1232 4310 1284
rect 5258 1232 5264 1284
rect 5316 1232 5322 1284
rect 5442 1232 5448 1284
rect 5500 1232 5506 1284
rect 5629 1275 5687 1281
rect 5629 1241 5641 1275
rect 5675 1272 5687 1275
rect 5902 1272 5908 1284
rect 5675 1244 5908 1272
rect 5675 1241 5687 1244
rect 5629 1235 5687 1241
rect 5902 1232 5908 1244
rect 5960 1232 5966 1284
rect 1044 1204 1072 1232
rect 1673 1207 1731 1213
rect 1673 1204 1685 1207
rect 1044 1176 1685 1204
rect 1673 1173 1685 1176
rect 1719 1173 1731 1207
rect 1673 1167 1731 1173
rect 2041 1207 2099 1213
rect 2041 1173 2053 1207
rect 2087 1204 2099 1207
rect 2130 1204 2136 1216
rect 2087 1176 2136 1204
rect 2087 1173 2099 1176
rect 2041 1167 2099 1173
rect 2130 1164 2136 1176
rect 2188 1164 2194 1216
rect 2406 1164 2412 1216
rect 2464 1164 2470 1216
rect 2774 1164 2780 1216
rect 2832 1164 2838 1216
rect 3145 1207 3203 1213
rect 3145 1173 3157 1207
rect 3191 1204 3203 1207
rect 3418 1204 3424 1216
rect 3191 1176 3424 1204
rect 3191 1173 3203 1176
rect 3145 1167 3203 1173
rect 3418 1164 3424 1176
rect 3476 1164 3482 1216
rect 3513 1207 3571 1213
rect 3513 1173 3525 1207
rect 3559 1204 3571 1207
rect 3878 1204 3884 1216
rect 3559 1176 3884 1204
rect 3559 1173 3571 1176
rect 3513 1167 3571 1173
rect 3878 1164 3884 1176
rect 3936 1164 3942 1216
rect 3973 1207 4031 1213
rect 3973 1173 3985 1207
rect 4019 1204 4031 1207
rect 4062 1204 4068 1216
rect 4019 1176 4068 1204
rect 4019 1173 4031 1176
rect 3973 1167 4031 1173
rect 4062 1164 4068 1176
rect 4120 1164 4126 1216
rect 4798 1164 4804 1216
rect 4856 1204 4862 1216
rect 7300 1204 7328 1303
rect 7576 1272 7604 1303
rect 7926 1300 7932 1352
rect 7984 1300 7990 1352
rect 9030 1300 9036 1352
rect 9088 1300 9094 1352
rect 9600 1330 9628 1371
rect 12066 1368 12072 1420
rect 12124 1368 12130 1420
rect 12526 1368 12532 1420
rect 12584 1368 12590 1420
rect 15838 1368 15844 1420
rect 15896 1408 15902 1420
rect 17512 1408 17540 1439
rect 18230 1436 18236 1488
rect 18288 1436 18294 1488
rect 18708 1448 19932 1476
rect 18248 1408 18276 1436
rect 15896 1380 17540 1408
rect 17604 1380 18276 1408
rect 15896 1368 15902 1380
rect 9827 1343 9885 1349
rect 9600 1302 9674 1330
rect 9827 1309 9839 1343
rect 9873 1340 9885 1343
rect 9950 1340 9956 1352
rect 9873 1312 9956 1340
rect 9873 1309 9885 1312
rect 9827 1303 9885 1309
rect 8389 1275 8447 1281
rect 7576 1244 8248 1272
rect 4856 1176 7328 1204
rect 4856 1164 4862 1176
rect 7466 1164 7472 1216
rect 7524 1164 7530 1216
rect 7742 1164 7748 1216
rect 7800 1164 7806 1216
rect 8110 1164 8116 1216
rect 8168 1164 8174 1216
rect 8220 1204 8248 1244
rect 8389 1241 8401 1275
rect 8435 1272 8447 1275
rect 9214 1272 9220 1284
rect 8435 1244 9220 1272
rect 8435 1241 8447 1244
rect 8389 1235 8447 1241
rect 9214 1232 9220 1244
rect 9272 1232 9278 1284
rect 9646 1272 9674 1302
rect 9950 1300 9956 1312
rect 10008 1300 10014 1352
rect 10226 1300 10232 1352
rect 10284 1300 10290 1352
rect 11054 1300 11060 1352
rect 11112 1300 11118 1352
rect 11698 1300 11704 1352
rect 11756 1300 11762 1352
rect 11790 1300 11796 1352
rect 11848 1300 11854 1352
rect 12084 1340 12112 1368
rect 12084 1312 12204 1340
rect 10244 1272 10272 1300
rect 9646 1244 10272 1272
rect 12176 1272 12204 1312
rect 12250 1300 12256 1352
rect 12308 1300 12314 1352
rect 12710 1300 12716 1352
rect 12768 1300 12774 1352
rect 13081 1343 13139 1349
rect 13081 1309 13093 1343
rect 13127 1340 13139 1343
rect 13354 1340 13360 1352
rect 13127 1312 13360 1340
rect 13127 1309 13139 1312
rect 13081 1303 13139 1309
rect 13354 1300 13360 1312
rect 13412 1300 13418 1352
rect 13446 1300 13452 1352
rect 13504 1300 13510 1352
rect 14090 1300 14096 1352
rect 14148 1300 14154 1352
rect 14550 1300 14556 1352
rect 14608 1300 14614 1352
rect 15194 1300 15200 1352
rect 15252 1340 15258 1352
rect 15289 1343 15347 1349
rect 15289 1340 15301 1343
rect 15252 1312 15301 1340
rect 15252 1300 15258 1312
rect 15289 1309 15301 1312
rect 15335 1309 15347 1343
rect 15289 1303 15347 1309
rect 16114 1300 16120 1352
rect 16172 1300 16178 1352
rect 16482 1300 16488 1352
rect 16540 1300 16546 1352
rect 16758 1300 16764 1352
rect 16816 1300 16822 1352
rect 17402 1300 17408 1352
rect 17460 1340 17466 1352
rect 17604 1340 17632 1380
rect 17460 1312 17632 1340
rect 17773 1343 17831 1349
rect 17460 1300 17466 1312
rect 17773 1309 17785 1343
rect 17819 1309 17831 1343
rect 17773 1303 17831 1309
rect 15841 1275 15899 1281
rect 15841 1272 15853 1275
rect 12176 1244 15853 1272
rect 15841 1241 15853 1244
rect 15887 1241 15899 1275
rect 16132 1272 16160 1300
rect 17313 1275 17371 1281
rect 17313 1272 17325 1275
rect 16132 1244 17325 1272
rect 15841 1235 15899 1241
rect 17313 1241 17325 1244
rect 17359 1241 17371 1275
rect 17788 1272 17816 1303
rect 18230 1300 18236 1352
rect 18288 1300 18294 1352
rect 18414 1300 18420 1352
rect 18472 1340 18478 1352
rect 18708 1340 18736 1448
rect 19904 1417 19932 1448
rect 20162 1436 20168 1488
rect 20220 1476 20226 1488
rect 23474 1476 23480 1488
rect 20220 1448 23480 1476
rect 20220 1436 20226 1448
rect 23474 1436 23480 1448
rect 23532 1436 23538 1488
rect 19889 1411 19947 1417
rect 19168 1380 19840 1408
rect 19168 1340 19196 1380
rect 18472 1312 18736 1340
rect 18800 1312 19196 1340
rect 19245 1343 19303 1349
rect 18472 1300 18478 1312
rect 18800 1272 18828 1312
rect 19245 1309 19257 1343
rect 19291 1309 19303 1343
rect 19245 1303 19303 1309
rect 19337 1343 19395 1349
rect 19337 1309 19349 1343
rect 19383 1340 19395 1343
rect 19426 1340 19432 1352
rect 19383 1312 19432 1340
rect 19383 1309 19395 1312
rect 19337 1303 19395 1309
rect 17788 1244 18828 1272
rect 18877 1275 18935 1281
rect 17313 1235 17371 1241
rect 18877 1241 18889 1275
rect 18923 1241 18935 1275
rect 19260 1272 19288 1303
rect 19426 1300 19432 1312
rect 19484 1300 19490 1352
rect 19705 1343 19763 1349
rect 19705 1309 19717 1343
rect 19751 1309 19763 1343
rect 19812 1340 19840 1380
rect 19889 1377 19901 1411
rect 19935 1377 19947 1411
rect 19889 1371 19947 1377
rect 23860 1380 24164 1408
rect 20714 1340 20720 1352
rect 19812 1312 20720 1340
rect 19705 1303 19763 1309
rect 19610 1272 19616 1284
rect 19260 1244 19616 1272
rect 18877 1235 18935 1241
rect 9306 1204 9312 1216
rect 8220 1176 9312 1204
rect 9306 1164 9312 1176
rect 9364 1164 9370 1216
rect 11514 1164 11520 1216
rect 11572 1164 11578 1216
rect 11977 1207 12035 1213
rect 11977 1173 11989 1207
rect 12023 1204 12035 1207
rect 12250 1204 12256 1216
rect 12023 1176 12256 1204
rect 12023 1173 12035 1176
rect 11977 1167 12035 1173
rect 12250 1164 12256 1176
rect 12308 1164 12314 1216
rect 12894 1164 12900 1216
rect 12952 1164 12958 1216
rect 13262 1164 13268 1216
rect 13320 1164 13326 1216
rect 13354 1164 13360 1216
rect 13412 1204 13418 1216
rect 13633 1207 13691 1213
rect 13633 1204 13645 1207
rect 13412 1176 13645 1204
rect 13412 1164 13418 1176
rect 13633 1173 13645 1176
rect 13679 1173 13691 1207
rect 13633 1167 13691 1173
rect 13906 1164 13912 1216
rect 13964 1204 13970 1216
rect 14277 1207 14335 1213
rect 14277 1204 14289 1207
rect 13964 1176 14289 1204
rect 13964 1164 13970 1176
rect 14277 1173 14289 1176
rect 14323 1173 14335 1207
rect 14277 1167 14335 1173
rect 15102 1164 15108 1216
rect 15160 1204 15166 1216
rect 16853 1207 16911 1213
rect 16853 1204 16865 1207
rect 15160 1176 16865 1204
rect 15160 1164 15166 1176
rect 16853 1173 16865 1176
rect 16899 1173 16911 1207
rect 16853 1167 16911 1173
rect 17954 1164 17960 1216
rect 18012 1164 18018 1216
rect 18892 1204 18920 1235
rect 19610 1232 19616 1244
rect 19668 1232 19674 1284
rect 19334 1204 19340 1216
rect 18892 1176 19340 1204
rect 19334 1164 19340 1176
rect 19392 1164 19398 1216
rect 19720 1204 19748 1303
rect 20714 1300 20720 1312
rect 20772 1300 20778 1352
rect 20809 1343 20867 1349
rect 20809 1309 20821 1343
rect 20855 1340 20867 1343
rect 21910 1340 21916 1352
rect 20855 1312 21916 1340
rect 20855 1309 20867 1312
rect 20809 1303 20867 1309
rect 21910 1300 21916 1312
rect 21968 1300 21974 1352
rect 22186 1300 22192 1352
rect 22244 1340 22250 1352
rect 23860 1340 23888 1380
rect 22244 1312 23888 1340
rect 24136 1340 24164 1380
rect 24213 1343 24271 1349
rect 24213 1340 24225 1343
rect 24136 1312 24225 1340
rect 22244 1300 22250 1312
rect 24213 1309 24225 1312
rect 24259 1309 24271 1343
rect 24213 1303 24271 1309
rect 20990 1232 20996 1284
rect 21048 1272 21054 1284
rect 21453 1275 21511 1281
rect 21453 1272 21465 1275
rect 21048 1244 21465 1272
rect 21048 1232 21054 1244
rect 21453 1241 21465 1244
rect 21499 1241 21511 1275
rect 21453 1235 21511 1241
rect 21542 1232 21548 1284
rect 21600 1272 21606 1284
rect 21821 1275 21879 1281
rect 21821 1272 21833 1275
rect 21600 1244 21833 1272
rect 21600 1232 21606 1244
rect 21821 1241 21833 1244
rect 21867 1241 21879 1275
rect 21821 1235 21879 1241
rect 23753 1275 23811 1281
rect 23753 1241 23765 1275
rect 23799 1272 23811 1275
rect 24302 1272 24308 1284
rect 23799 1244 24308 1272
rect 23799 1241 23811 1244
rect 23753 1235 23811 1241
rect 24302 1232 24308 1244
rect 24360 1232 24366 1284
rect 22186 1204 22192 1216
rect 19720 1176 22192 1204
rect 22186 1164 22192 1176
rect 22244 1164 22250 1216
rect 22278 1164 22284 1216
rect 22336 1204 22342 1216
rect 24029 1207 24087 1213
rect 24029 1204 24041 1207
rect 22336 1176 24041 1204
rect 22336 1164 22342 1176
rect 24029 1173 24041 1176
rect 24075 1173 24087 1207
rect 24029 1167 24087 1173
rect 1104 1114 24723 1136
rect 1104 1062 6814 1114
rect 6866 1062 6878 1114
rect 6930 1062 6942 1114
rect 6994 1062 7006 1114
rect 7058 1062 7070 1114
rect 7122 1062 12679 1114
rect 12731 1062 12743 1114
rect 12795 1062 12807 1114
rect 12859 1062 12871 1114
rect 12923 1062 12935 1114
rect 12987 1062 18544 1114
rect 18596 1062 18608 1114
rect 18660 1062 18672 1114
rect 18724 1062 18736 1114
rect 18788 1062 18800 1114
rect 18852 1062 24409 1114
rect 24461 1062 24473 1114
rect 24525 1062 24537 1114
rect 24589 1062 24601 1114
rect 24653 1062 24665 1114
rect 24717 1062 24723 1114
rect 1104 1040 24723 1062
rect 6270 1000 6276 1012
rect 2746 972 6276 1000
rect 474 620 480 672
rect 532 660 538 672
rect 2746 660 2774 972
rect 6270 960 6276 972
rect 6328 960 6334 1012
rect 7760 972 17080 1000
rect 3418 892 3424 944
rect 3476 892 3482 944
rect 5626 892 5632 944
rect 5684 932 5690 944
rect 6086 932 6092 944
rect 5684 904 6092 932
rect 5684 892 5690 904
rect 6086 892 6092 904
rect 6144 892 6150 944
rect 3436 864 3464 892
rect 7760 864 7788 972
rect 3436 836 7788 864
rect 8036 904 12434 932
rect 3326 756 3332 808
rect 3384 796 3390 808
rect 5718 796 5724 808
rect 3384 768 5724 796
rect 3384 756 3390 768
rect 5718 756 5724 768
rect 5776 756 5782 808
rect 8036 796 8064 904
rect 8110 824 8116 876
rect 8168 864 8174 876
rect 11422 864 11428 876
rect 8168 836 11428 864
rect 8168 824 8174 836
rect 11422 824 11428 836
rect 11480 824 11486 876
rect 6564 768 8064 796
rect 5442 688 5448 740
rect 5500 728 5506 740
rect 6564 728 6592 768
rect 8938 756 8944 808
rect 8996 796 9002 808
rect 9858 796 9864 808
rect 8996 768 9864 796
rect 8996 756 9002 768
rect 9858 756 9864 768
rect 9916 756 9922 808
rect 9950 756 9956 808
rect 10008 796 10014 808
rect 10778 796 10784 808
rect 10008 768 10784 796
rect 10008 756 10014 768
rect 10778 756 10784 768
rect 10836 756 10842 808
rect 12406 796 12434 904
rect 16574 796 16580 808
rect 12406 768 16580 796
rect 16574 756 16580 768
rect 16632 756 16638 808
rect 17052 796 17080 972
rect 19610 960 19616 1012
rect 19668 1000 19674 1012
rect 22094 1000 22100 1012
rect 19668 972 22100 1000
rect 19668 960 19674 972
rect 22094 960 22100 972
rect 22152 960 22158 1012
rect 18230 892 18236 944
rect 18288 932 18294 944
rect 18288 904 22508 932
rect 18288 892 18294 904
rect 17126 824 17132 876
rect 17184 864 17190 876
rect 17184 836 19288 864
rect 17184 824 17190 836
rect 17052 768 17264 796
rect 5500 700 6592 728
rect 5500 688 5506 700
rect 6638 688 6644 740
rect 6696 728 6702 740
rect 10318 728 10324 740
rect 6696 700 10324 728
rect 6696 688 6702 700
rect 10318 688 10324 700
rect 10376 688 10382 740
rect 17126 728 17132 740
rect 12406 700 17132 728
rect 12406 660 12434 700
rect 17126 688 17132 700
rect 17184 688 17190 740
rect 532 632 2774 660
rect 7576 632 12434 660
rect 17236 660 17264 768
rect 17954 756 17960 808
rect 18012 756 18018 808
rect 19260 796 19288 836
rect 19334 824 19340 876
rect 19392 864 19398 876
rect 20530 864 20536 876
rect 19392 836 20536 864
rect 19392 824 19398 836
rect 20530 824 20536 836
rect 20588 824 20594 876
rect 22278 864 22284 876
rect 22066 836 22284 864
rect 22066 796 22094 836
rect 22278 824 22284 836
rect 22336 824 22342 876
rect 22480 808 22508 904
rect 19260 768 22094 796
rect 22462 756 22468 808
rect 22520 756 22526 808
rect 17972 728 18000 756
rect 22922 728 22928 740
rect 17972 700 22928 728
rect 22922 688 22928 700
rect 22980 688 22986 740
rect 23842 660 23848 672
rect 17236 632 23848 660
rect 532 620 538 632
rect 2406 552 2412 604
rect 2464 592 2470 604
rect 7576 592 7604 632
rect 23842 620 23848 632
rect 23900 620 23906 672
rect 2464 564 7604 592
rect 2464 552 2470 564
rect 11238 552 11244 604
rect 11296 592 11302 604
rect 11974 592 11980 604
rect 11296 564 11980 592
rect 11296 552 11302 564
rect 11974 552 11980 564
rect 12032 552 12038 604
rect 14366 592 14372 604
rect 12406 564 14372 592
rect 3878 484 3884 536
rect 3936 524 3942 536
rect 12406 524 12434 564
rect 14366 552 14372 564
rect 14424 552 14430 604
rect 14642 552 14648 604
rect 14700 592 14706 604
rect 20990 592 20996 604
rect 14700 564 20996 592
rect 14700 552 14706 564
rect 20990 552 20996 564
rect 21048 552 21054 604
rect 3936 496 12434 524
rect 3936 484 3942 496
rect 16482 484 16488 536
rect 16540 524 16546 536
rect 25590 524 25596 536
rect 16540 496 25596 524
rect 16540 484 16546 496
rect 25590 484 25596 496
rect 25648 484 25654 536
rect 106 416 112 468
rect 164 456 170 468
rect 5534 456 5540 468
rect 164 428 5540 456
rect 164 416 170 428
rect 5534 416 5540 428
rect 5592 416 5598 468
<< via1 >>
rect 664 44276 716 44328
rect 7748 44276 7800 44328
rect 6184 44208 6236 44260
rect 6552 44208 6604 44260
rect 3056 44140 3108 44192
rect 4528 44140 4580 44192
rect 5448 44140 5500 44192
rect 3516 44072 3568 44124
rect 10692 44072 10744 44124
rect 5816 44004 5868 44056
rect 6276 43936 6328 43988
rect 1400 43800 1452 43852
rect 2688 43800 2740 43852
rect 3240 43800 3292 43852
rect 6000 43800 6052 43852
rect 112 43732 164 43784
rect 1584 43664 1636 43716
rect 6184 43664 6236 43716
rect 9864 43664 9916 43716
rect 2320 43596 2372 43648
rect 5540 43596 5592 43648
rect 5724 43596 5776 43648
rect 11060 43596 11112 43648
rect 18052 44072 18104 44124
rect 19156 44072 19208 44124
rect 17960 44004 18012 44056
rect 19064 44004 19116 44056
rect 17776 43936 17828 43988
rect 18420 43936 18472 43988
rect 16856 43596 16908 43648
rect 6814 43494 6866 43546
rect 6878 43494 6930 43546
rect 6942 43494 6994 43546
rect 7006 43494 7058 43546
rect 7070 43494 7122 43546
rect 12679 43494 12731 43546
rect 12743 43494 12795 43546
rect 12807 43494 12859 43546
rect 12871 43494 12923 43546
rect 12935 43494 12987 43546
rect 18544 43494 18596 43546
rect 18608 43494 18660 43546
rect 18672 43494 18724 43546
rect 18736 43494 18788 43546
rect 18800 43494 18852 43546
rect 24409 43494 24461 43546
rect 24473 43494 24525 43546
rect 24537 43494 24589 43546
rect 24601 43494 24653 43546
rect 24665 43494 24717 43546
rect 1584 43435 1636 43444
rect 1584 43401 1593 43435
rect 1593 43401 1627 43435
rect 1627 43401 1636 43435
rect 1584 43392 1636 43401
rect 3148 43392 3200 43444
rect 2688 43367 2740 43376
rect 2688 43333 2697 43367
rect 2697 43333 2731 43367
rect 2731 43333 2740 43367
rect 2688 43324 2740 43333
rect 5632 43392 5684 43444
rect 5908 43392 5960 43444
rect 6736 43392 6788 43444
rect 7196 43435 7248 43444
rect 7196 43401 7205 43435
rect 7205 43401 7239 43435
rect 7239 43401 7248 43435
rect 7196 43392 7248 43401
rect 1400 43299 1452 43308
rect 1400 43265 1409 43299
rect 1409 43265 1443 43299
rect 1443 43265 1452 43299
rect 1400 43256 1452 43265
rect 2964 43256 3016 43308
rect 3240 43299 3292 43308
rect 3240 43265 3249 43299
rect 3249 43265 3283 43299
rect 3283 43265 3292 43299
rect 3240 43256 3292 43265
rect 4712 43256 4764 43308
rect 5724 43256 5776 43308
rect 7748 43324 7800 43376
rect 3332 43188 3384 43240
rect 5540 43231 5592 43240
rect 5540 43197 5549 43231
rect 5549 43197 5583 43231
rect 5583 43197 5592 43231
rect 5540 43188 5592 43197
rect 2504 43120 2556 43172
rect 6644 43256 6696 43308
rect 8944 43392 8996 43444
rect 9496 43392 9548 43444
rect 9772 43392 9824 43444
rect 9864 43392 9916 43444
rect 12164 43392 12216 43444
rect 16120 43392 16172 43444
rect 7564 43188 7616 43240
rect 9128 43188 9180 43240
rect 8668 43120 8720 43172
rect 9588 43256 9640 43308
rect 9772 43256 9824 43308
rect 10232 43256 10284 43308
rect 10968 43299 11020 43308
rect 10968 43265 10977 43299
rect 10977 43265 11011 43299
rect 11011 43265 11020 43299
rect 10968 43256 11020 43265
rect 11152 43256 11204 43308
rect 12072 43299 12124 43308
rect 12072 43265 12081 43299
rect 12081 43265 12115 43299
rect 12115 43265 12124 43299
rect 12072 43256 12124 43265
rect 12256 43324 12308 43376
rect 13176 43367 13228 43376
rect 13176 43333 13185 43367
rect 13185 43333 13219 43367
rect 13219 43333 13228 43367
rect 13176 43324 13228 43333
rect 13544 43367 13596 43376
rect 13544 43333 13553 43367
rect 13553 43333 13587 43367
rect 13587 43333 13596 43367
rect 13544 43324 13596 43333
rect 15292 43324 15344 43376
rect 16028 43324 16080 43376
rect 16856 43324 16908 43376
rect 17316 43392 17368 43444
rect 20260 43392 20312 43444
rect 20536 43392 20588 43444
rect 21364 43392 21416 43444
rect 23756 43435 23808 43444
rect 23756 43401 23765 43435
rect 23765 43401 23799 43435
rect 23799 43401 23808 43435
rect 23756 43392 23808 43401
rect 25504 43392 25556 43444
rect 17224 43324 17276 43376
rect 12348 43256 12400 43308
rect 13084 43256 13136 43308
rect 14096 43299 14148 43308
rect 14096 43265 14105 43299
rect 14105 43265 14139 43299
rect 14139 43265 14148 43299
rect 14096 43256 14148 43265
rect 14464 43299 14516 43308
rect 14464 43265 14473 43299
rect 14473 43265 14507 43299
rect 14507 43265 14516 43299
rect 14464 43256 14516 43265
rect 14832 43299 14884 43308
rect 14832 43265 14841 43299
rect 14841 43265 14875 43299
rect 14875 43265 14884 43299
rect 14832 43256 14884 43265
rect 15568 43256 15620 43308
rect 16396 43256 16448 43308
rect 18420 43324 18472 43376
rect 18880 43324 18932 43376
rect 10508 43188 10560 43240
rect 10416 43120 10468 43172
rect 13176 43188 13228 43240
rect 15016 43188 15068 43240
rect 16672 43188 16724 43240
rect 18052 43188 18104 43240
rect 19064 43299 19116 43308
rect 19064 43265 19073 43299
rect 19073 43265 19107 43299
rect 19107 43265 19116 43299
rect 19064 43256 19116 43265
rect 19156 43256 19208 43308
rect 18696 43188 18748 43240
rect 20168 43299 20220 43308
rect 20168 43265 20177 43299
rect 20177 43265 20211 43299
rect 20211 43265 20220 43299
rect 20168 43256 20220 43265
rect 20076 43188 20128 43240
rect 21272 43299 21324 43308
rect 21272 43265 21281 43299
rect 21281 43265 21315 43299
rect 21315 43265 21324 43299
rect 21272 43256 21324 43265
rect 20812 43188 20864 43240
rect 22376 43256 22428 43308
rect 22836 43299 22888 43308
rect 22836 43265 22845 43299
rect 22845 43265 22879 43299
rect 22879 43265 22888 43299
rect 22836 43256 22888 43265
rect 23664 43299 23716 43308
rect 23664 43265 23673 43299
rect 23673 43265 23707 43299
rect 23707 43265 23716 43299
rect 23664 43256 23716 43265
rect 11888 43120 11940 43172
rect 13360 43163 13412 43172
rect 13360 43129 13369 43163
rect 13369 43129 13403 43163
rect 13403 43129 13412 43163
rect 13360 43120 13412 43129
rect 14188 43120 14240 43172
rect 9680 43052 9732 43104
rect 9772 43052 9824 43104
rect 10876 43052 10928 43104
rect 11796 43052 11848 43104
rect 11980 43052 12032 43104
rect 12532 43095 12584 43104
rect 12532 43061 12541 43095
rect 12541 43061 12575 43095
rect 12575 43061 12584 43095
rect 12532 43052 12584 43061
rect 13636 43095 13688 43104
rect 13636 43061 13645 43095
rect 13645 43061 13679 43095
rect 13679 43061 13688 43095
rect 13636 43052 13688 43061
rect 14648 43095 14700 43104
rect 14648 43061 14657 43095
rect 14657 43061 14691 43095
rect 14691 43061 14700 43095
rect 14648 43052 14700 43061
rect 15476 43052 15528 43104
rect 16304 43095 16356 43104
rect 16304 43061 16313 43095
rect 16313 43061 16347 43095
rect 16347 43061 16356 43095
rect 16304 43052 16356 43061
rect 17868 43120 17920 43172
rect 19616 43120 19668 43172
rect 20536 43120 20588 43172
rect 24216 43188 24268 43240
rect 17592 43095 17644 43104
rect 17592 43061 17601 43095
rect 17601 43061 17635 43095
rect 17635 43061 17644 43095
rect 17592 43052 17644 43061
rect 17776 43095 17828 43104
rect 17776 43061 17785 43095
rect 17785 43061 17819 43095
rect 17819 43061 17828 43095
rect 17776 43052 17828 43061
rect 18052 43095 18104 43104
rect 18052 43061 18061 43095
rect 18061 43061 18095 43095
rect 18095 43061 18104 43095
rect 18052 43052 18104 43061
rect 18604 43095 18656 43104
rect 18604 43061 18613 43095
rect 18613 43061 18647 43095
rect 18647 43061 18656 43095
rect 18604 43052 18656 43061
rect 19248 43095 19300 43104
rect 19248 43061 19257 43095
rect 19257 43061 19291 43095
rect 19291 43061 19300 43095
rect 19248 43052 19300 43061
rect 19432 43052 19484 43104
rect 19800 43095 19852 43104
rect 19800 43061 19809 43095
rect 19809 43061 19843 43095
rect 19843 43061 19852 43095
rect 19800 43052 19852 43061
rect 21916 43052 21968 43104
rect 3882 42950 3934 43002
rect 3946 42950 3998 43002
rect 4010 42950 4062 43002
rect 4074 42950 4126 43002
rect 4138 42950 4190 43002
rect 9747 42950 9799 43002
rect 9811 42950 9863 43002
rect 9875 42950 9927 43002
rect 9939 42950 9991 43002
rect 10003 42950 10055 43002
rect 15612 42950 15664 43002
rect 15676 42950 15728 43002
rect 15740 42950 15792 43002
rect 15804 42950 15856 43002
rect 15868 42950 15920 43002
rect 21477 42950 21529 43002
rect 21541 42950 21593 43002
rect 21605 42950 21657 43002
rect 21669 42950 21721 43002
rect 21733 42950 21785 43002
rect 3056 42848 3108 42900
rect 3240 42780 3292 42832
rect 3516 42780 3568 42832
rect 3424 42712 3476 42764
rect 940 42644 992 42696
rect 1952 42576 2004 42628
rect 2688 42619 2740 42628
rect 2688 42585 2697 42619
rect 2697 42585 2731 42619
rect 2731 42585 2740 42619
rect 2688 42576 2740 42585
rect 3240 42619 3292 42628
rect 3240 42585 3249 42619
rect 3249 42585 3283 42619
rect 3283 42585 3292 42619
rect 3240 42576 3292 42585
rect 7932 42891 7984 42900
rect 7932 42857 7941 42891
rect 7941 42857 7975 42891
rect 7975 42857 7984 42891
rect 7932 42848 7984 42857
rect 8484 42891 8536 42900
rect 8484 42857 8493 42891
rect 8493 42857 8527 42891
rect 8527 42857 8536 42891
rect 8484 42848 8536 42857
rect 8024 42780 8076 42832
rect 9496 42891 9548 42900
rect 9496 42857 9505 42891
rect 9505 42857 9539 42891
rect 9539 42857 9548 42891
rect 9496 42848 9548 42857
rect 9588 42848 9640 42900
rect 14924 42848 14976 42900
rect 10232 42780 10284 42832
rect 9496 42712 9548 42764
rect 13084 42712 13136 42764
rect 3976 42687 4028 42696
rect 3976 42653 3985 42687
rect 3985 42653 4019 42687
rect 4019 42653 4028 42687
rect 3976 42644 4028 42653
rect 4252 42644 4304 42696
rect 4436 42644 4488 42696
rect 4712 42644 4764 42696
rect 4896 42644 4948 42696
rect 5356 42644 5408 42696
rect 5724 42687 5776 42696
rect 5724 42653 5731 42687
rect 5731 42653 5765 42687
rect 5765 42653 5776 42687
rect 5724 42644 5776 42653
rect 8944 42687 8996 42696
rect 8944 42653 8953 42687
rect 8953 42653 8987 42687
rect 8987 42653 8996 42687
rect 8944 42644 8996 42653
rect 10140 42644 10192 42696
rect 10232 42687 10284 42696
rect 10232 42653 10241 42687
rect 10241 42653 10275 42687
rect 10275 42653 10284 42687
rect 10232 42644 10284 42653
rect 10600 42687 10652 42696
rect 10600 42653 10609 42687
rect 10609 42653 10643 42687
rect 10643 42653 10652 42687
rect 10600 42644 10652 42653
rect 11428 42644 11480 42696
rect 11796 42687 11848 42696
rect 11796 42653 11805 42687
rect 11805 42653 11839 42687
rect 11839 42653 11848 42687
rect 11796 42644 11848 42653
rect 12624 42687 12676 42696
rect 12624 42653 12633 42687
rect 12633 42653 12667 42687
rect 12667 42653 12676 42687
rect 12624 42644 12676 42653
rect 13728 42687 13780 42696
rect 13728 42653 13737 42687
rect 13737 42653 13771 42687
rect 13771 42653 13780 42687
rect 13728 42644 13780 42653
rect 14280 42687 14332 42696
rect 14280 42653 14289 42687
rect 14289 42653 14323 42687
rect 14323 42653 14332 42687
rect 14280 42644 14332 42653
rect 15108 42687 15160 42696
rect 15108 42653 15117 42687
rect 15117 42653 15151 42687
rect 15151 42653 15160 42687
rect 15108 42644 15160 42653
rect 17776 42780 17828 42832
rect 18604 42848 18656 42900
rect 19156 42848 19208 42900
rect 17316 42644 17368 42696
rect 17868 42644 17920 42696
rect 18052 42644 18104 42696
rect 19248 42780 19300 42832
rect 19800 42780 19852 42832
rect 18328 42687 18380 42696
rect 18328 42653 18337 42687
rect 18337 42653 18371 42687
rect 18371 42653 18380 42687
rect 18328 42644 18380 42653
rect 20168 42848 20220 42900
rect 20628 42848 20680 42900
rect 22100 42848 22152 42900
rect 22652 42848 22704 42900
rect 20352 42780 20404 42832
rect 22836 42780 22888 42832
rect 20260 42712 20312 42764
rect 20444 42687 20496 42696
rect 20444 42653 20453 42687
rect 20453 42653 20487 42687
rect 20487 42653 20496 42687
rect 20444 42644 20496 42653
rect 20536 42644 20588 42696
rect 1216 42508 1268 42560
rect 3424 42508 3476 42560
rect 4804 42508 4856 42560
rect 5080 42551 5132 42560
rect 5080 42517 5089 42551
rect 5089 42517 5123 42551
rect 5123 42517 5132 42551
rect 5080 42508 5132 42517
rect 5264 42508 5316 42560
rect 7012 42576 7064 42628
rect 7564 42576 7616 42628
rect 8300 42576 8352 42628
rect 9220 42576 9272 42628
rect 9404 42619 9456 42628
rect 9404 42585 9413 42619
rect 9413 42585 9447 42619
rect 9447 42585 9456 42619
rect 9404 42576 9456 42585
rect 6460 42551 6512 42560
rect 6460 42517 6469 42551
rect 6469 42517 6503 42551
rect 6503 42517 6512 42551
rect 6460 42508 6512 42517
rect 10784 42576 10836 42628
rect 12072 42576 12124 42628
rect 10140 42508 10192 42560
rect 11520 42551 11572 42560
rect 11520 42517 11529 42551
rect 11529 42517 11563 42551
rect 11563 42517 11572 42551
rect 11520 42508 11572 42517
rect 11612 42508 11664 42560
rect 12440 42508 12492 42560
rect 16488 42619 16540 42628
rect 16488 42585 16497 42619
rect 16497 42585 16531 42619
rect 16531 42585 16540 42619
rect 16488 42576 16540 42585
rect 14096 42508 14148 42560
rect 16764 42551 16816 42560
rect 16764 42517 16773 42551
rect 16773 42517 16807 42551
rect 16807 42517 16816 42551
rect 16764 42508 16816 42517
rect 17132 42551 17184 42560
rect 17132 42517 17141 42551
rect 17141 42517 17175 42551
rect 17175 42517 17184 42551
rect 17132 42508 17184 42517
rect 17500 42551 17552 42560
rect 17500 42517 17509 42551
rect 17509 42517 17543 42551
rect 17543 42517 17552 42551
rect 17500 42508 17552 42517
rect 17960 42619 18012 42628
rect 17960 42585 17969 42619
rect 17969 42585 18003 42619
rect 18003 42585 18012 42619
rect 17960 42576 18012 42585
rect 19432 42576 19484 42628
rect 19524 42619 19576 42628
rect 19524 42585 19533 42619
rect 19533 42585 19567 42619
rect 19567 42585 19576 42619
rect 19524 42576 19576 42585
rect 20628 42576 20680 42628
rect 21916 42712 21968 42764
rect 22008 42712 22060 42764
rect 23020 42712 23072 42764
rect 18328 42508 18380 42560
rect 18696 42508 18748 42560
rect 19800 42551 19852 42560
rect 19800 42517 19809 42551
rect 19809 42517 19843 42551
rect 19843 42517 19852 42551
rect 19800 42508 19852 42517
rect 20168 42508 20220 42560
rect 20720 42508 20772 42560
rect 20812 42551 20864 42560
rect 20812 42517 20821 42551
rect 20821 42517 20855 42551
rect 20855 42517 20864 42551
rect 20812 42508 20864 42517
rect 21272 42508 21324 42560
rect 23480 42644 23532 42696
rect 23756 42644 23808 42696
rect 22284 42619 22336 42628
rect 22284 42585 22293 42619
rect 22293 42585 22327 42619
rect 22327 42585 22336 42619
rect 22284 42576 22336 42585
rect 22652 42576 22704 42628
rect 22192 42508 22244 42560
rect 24124 42551 24176 42560
rect 24124 42517 24133 42551
rect 24133 42517 24167 42551
rect 24167 42517 24176 42551
rect 24124 42508 24176 42517
rect 6814 42406 6866 42458
rect 6878 42406 6930 42458
rect 6942 42406 6994 42458
rect 7006 42406 7058 42458
rect 7070 42406 7122 42458
rect 12679 42406 12731 42458
rect 12743 42406 12795 42458
rect 12807 42406 12859 42458
rect 12871 42406 12923 42458
rect 12935 42406 12987 42458
rect 18544 42406 18596 42458
rect 18608 42406 18660 42458
rect 18672 42406 18724 42458
rect 18736 42406 18788 42458
rect 18800 42406 18852 42458
rect 24409 42406 24461 42458
rect 24473 42406 24525 42458
rect 24537 42406 24589 42458
rect 24601 42406 24653 42458
rect 24665 42406 24717 42458
rect 2596 42304 2648 42356
rect 3424 42304 3476 42356
rect 7288 42304 7340 42356
rect 7748 42304 7800 42356
rect 2228 42236 2280 42288
rect 1676 42168 1728 42220
rect 2044 42211 2096 42220
rect 2044 42177 2053 42211
rect 2053 42177 2087 42211
rect 2087 42177 2096 42211
rect 2044 42168 2096 42177
rect 3148 42236 3200 42288
rect 4160 42236 4212 42288
rect 4252 42236 4304 42288
rect 4804 42236 4856 42288
rect 4896 42236 4948 42288
rect 5172 42236 5224 42288
rect 5356 42236 5408 42288
rect 9128 42347 9180 42356
rect 9128 42313 9137 42347
rect 9137 42313 9171 42347
rect 9171 42313 9180 42347
rect 9128 42304 9180 42313
rect 9956 42347 10008 42356
rect 9956 42313 9965 42347
rect 9965 42313 9999 42347
rect 9999 42313 10008 42347
rect 9956 42304 10008 42313
rect 16488 42304 16540 42356
rect 16764 42304 16816 42356
rect 3056 42211 3108 42220
rect 3056 42177 3065 42211
rect 3065 42177 3099 42211
rect 3099 42177 3108 42211
rect 3056 42168 3108 42177
rect 4344 42168 4396 42220
rect 5448 42168 5500 42220
rect 1584 42143 1636 42152
rect 1584 42109 1593 42143
rect 1593 42109 1627 42143
rect 1627 42109 1636 42143
rect 1584 42100 1636 42109
rect 2504 42100 2556 42152
rect 3884 42100 3936 42152
rect 6368 42168 6420 42220
rect 7472 42168 7524 42220
rect 8300 42211 8352 42220
rect 8300 42177 8309 42211
rect 8309 42177 8343 42211
rect 8343 42177 8352 42211
rect 8300 42168 8352 42177
rect 6828 42143 6880 42152
rect 6828 42109 6837 42143
rect 6837 42109 6871 42143
rect 6871 42109 6880 42143
rect 6828 42100 6880 42109
rect 7564 42100 7616 42152
rect 4436 41964 4488 42016
rect 4620 41964 4672 42016
rect 6644 42032 6696 42084
rect 5172 42007 5224 42016
rect 5172 41973 5181 42007
rect 5181 41973 5215 42007
rect 5215 41973 5224 42007
rect 5172 41964 5224 41973
rect 5448 41964 5500 42016
rect 6920 41964 6972 42016
rect 7656 41964 7708 42016
rect 7840 42007 7892 42016
rect 7840 41973 7849 42007
rect 7849 41973 7883 42007
rect 7883 41973 7892 42007
rect 7840 41964 7892 41973
rect 7932 41964 7984 42016
rect 9036 42211 9088 42220
rect 9036 42177 9045 42211
rect 9045 42177 9079 42211
rect 9079 42177 9088 42211
rect 9036 42168 9088 42177
rect 9312 42211 9364 42220
rect 9312 42177 9321 42211
rect 9321 42177 9355 42211
rect 9355 42177 9364 42211
rect 9312 42168 9364 42177
rect 10140 42211 10192 42220
rect 10140 42177 10149 42211
rect 10149 42177 10183 42211
rect 10183 42177 10192 42211
rect 10140 42168 10192 42177
rect 10416 42211 10468 42220
rect 10416 42177 10425 42211
rect 10425 42177 10459 42211
rect 10459 42177 10468 42211
rect 10416 42168 10468 42177
rect 16396 42236 16448 42288
rect 20812 42304 20864 42356
rect 21088 42304 21140 42356
rect 22744 42304 22796 42356
rect 22928 42304 22980 42356
rect 24860 42304 24912 42356
rect 20168 42236 20220 42288
rect 24032 42236 24084 42288
rect 18696 42211 18748 42220
rect 18696 42177 18705 42211
rect 18705 42177 18739 42211
rect 18739 42177 18748 42211
rect 18696 42168 18748 42177
rect 19064 42168 19116 42220
rect 20260 42168 20312 42220
rect 20168 42100 20220 42152
rect 18512 42007 18564 42016
rect 18512 41973 18521 42007
rect 18521 41973 18555 42007
rect 18555 41973 18564 42007
rect 18512 41964 18564 41973
rect 19340 42032 19392 42084
rect 20996 42211 21048 42220
rect 20996 42177 21005 42211
rect 21005 42177 21039 42211
rect 21039 42177 21048 42211
rect 20996 42168 21048 42177
rect 21088 42168 21140 42220
rect 21364 42211 21416 42220
rect 21364 42177 21373 42211
rect 21373 42177 21407 42211
rect 21407 42177 21416 42211
rect 21364 42168 21416 42177
rect 20628 42100 20680 42152
rect 22560 42211 22612 42220
rect 22560 42177 22569 42211
rect 22569 42177 22603 42211
rect 22603 42177 22612 42211
rect 22560 42168 22612 42177
rect 23112 42211 23164 42220
rect 23112 42177 23121 42211
rect 23121 42177 23155 42211
rect 23155 42177 23164 42211
rect 23112 42168 23164 42177
rect 23572 42168 23624 42220
rect 22928 42100 22980 42152
rect 20260 41964 20312 42016
rect 20904 41964 20956 42016
rect 21456 41964 21508 42016
rect 3882 41862 3934 41914
rect 3946 41862 3998 41914
rect 4010 41862 4062 41914
rect 4074 41862 4126 41914
rect 4138 41862 4190 41914
rect 9747 41862 9799 41914
rect 9811 41862 9863 41914
rect 9875 41862 9927 41914
rect 9939 41862 9991 41914
rect 10003 41862 10055 41914
rect 15612 41862 15664 41914
rect 15676 41862 15728 41914
rect 15740 41862 15792 41914
rect 15804 41862 15856 41914
rect 15868 41862 15920 41914
rect 21477 41862 21529 41914
rect 21541 41862 21593 41914
rect 21605 41862 21657 41914
rect 21669 41862 21721 41914
rect 21733 41862 21785 41914
rect 3056 41760 3108 41812
rect 4896 41760 4948 41812
rect 6460 41760 6512 41812
rect 6552 41760 6604 41812
rect 3240 41692 3292 41744
rect 3424 41692 3476 41744
rect 4620 41692 4672 41744
rect 3148 41624 3200 41676
rect 4712 41624 4764 41676
rect 4804 41624 4856 41676
rect 5080 41624 5132 41676
rect 1400 41599 1452 41608
rect 1400 41565 1409 41599
rect 1409 41565 1443 41599
rect 1443 41565 1452 41599
rect 1400 41556 1452 41565
rect 2044 41531 2096 41540
rect 2044 41497 2053 41531
rect 2053 41497 2087 41531
rect 2087 41497 2096 41531
rect 2044 41488 2096 41497
rect 2504 41556 2556 41608
rect 6736 41692 6788 41744
rect 8944 41803 8996 41812
rect 8944 41769 8953 41803
rect 8953 41769 8987 41803
rect 8987 41769 8996 41803
rect 8944 41760 8996 41769
rect 9220 41803 9272 41812
rect 9220 41769 9229 41803
rect 9229 41769 9263 41803
rect 9263 41769 9272 41803
rect 9220 41760 9272 41769
rect 15200 41760 15252 41812
rect 19340 41760 19392 41812
rect 20444 41760 20496 41812
rect 6368 41624 6420 41676
rect 6828 41624 6880 41676
rect 10232 41692 10284 41744
rect 13912 41624 13964 41676
rect 2780 41488 2832 41540
rect 2964 41488 3016 41540
rect 3516 41488 3568 41540
rect 4712 41488 4764 41540
rect 5264 41488 5316 41540
rect 5540 41488 5592 41540
rect 5908 41488 5960 41540
rect 4988 41420 5040 41472
rect 5448 41420 5500 41472
rect 5632 41420 5684 41472
rect 6368 41463 6420 41472
rect 6368 41429 6377 41463
rect 6377 41429 6411 41463
rect 6411 41429 6420 41463
rect 6368 41420 6420 41429
rect 6644 41531 6696 41540
rect 6644 41497 6653 41531
rect 6653 41497 6687 41531
rect 6687 41497 6696 41531
rect 6644 41488 6696 41497
rect 7104 41599 7156 41608
rect 7104 41565 7113 41599
rect 7113 41565 7147 41599
rect 7147 41565 7156 41599
rect 7104 41556 7156 41565
rect 7656 41556 7708 41608
rect 9128 41599 9180 41608
rect 9128 41565 9137 41599
rect 9137 41565 9171 41599
rect 9171 41565 9180 41599
rect 9128 41556 9180 41565
rect 9220 41556 9272 41608
rect 13820 41556 13872 41608
rect 19432 41556 19484 41608
rect 10968 41488 11020 41540
rect 19340 41531 19392 41540
rect 19340 41497 19349 41531
rect 19349 41497 19383 41531
rect 19383 41497 19392 41531
rect 19340 41488 19392 41497
rect 8484 41463 8536 41472
rect 8484 41429 8493 41463
rect 8493 41429 8527 41463
rect 8527 41429 8536 41463
rect 8484 41420 8536 41429
rect 19432 41463 19484 41472
rect 19432 41429 19441 41463
rect 19441 41429 19475 41463
rect 19475 41429 19484 41463
rect 19432 41420 19484 41429
rect 19616 41463 19668 41472
rect 19616 41429 19625 41463
rect 19625 41429 19659 41463
rect 19659 41429 19668 41463
rect 19616 41420 19668 41429
rect 20076 41692 20128 41744
rect 20352 41735 20404 41744
rect 20352 41701 20361 41735
rect 20361 41701 20395 41735
rect 20395 41701 20404 41735
rect 20352 41692 20404 41701
rect 21272 41760 21324 41812
rect 22560 41760 22612 41812
rect 23296 41760 23348 41812
rect 23940 41803 23992 41812
rect 23940 41769 23949 41803
rect 23949 41769 23983 41803
rect 23983 41769 23992 41803
rect 23940 41760 23992 41769
rect 24308 41760 24360 41812
rect 22376 41692 22428 41744
rect 20904 41624 20956 41676
rect 20536 41599 20588 41608
rect 20536 41565 20545 41599
rect 20545 41565 20579 41599
rect 20579 41565 20588 41599
rect 20536 41556 20588 41565
rect 25136 41624 25188 41676
rect 21272 41556 21324 41608
rect 21640 41599 21692 41608
rect 21640 41565 21649 41599
rect 21649 41565 21683 41599
rect 21683 41565 21692 41599
rect 21640 41556 21692 41565
rect 21824 41556 21876 41608
rect 24952 41556 25004 41608
rect 20628 41420 20680 41472
rect 22100 41488 22152 41540
rect 22192 41531 22244 41540
rect 22192 41497 22201 41531
rect 22201 41497 22235 41531
rect 22235 41497 22244 41531
rect 22192 41488 22244 41497
rect 21548 41420 21600 41472
rect 22376 41420 22428 41472
rect 23296 41531 23348 41540
rect 23296 41497 23305 41531
rect 23305 41497 23339 41531
rect 23339 41497 23348 41531
rect 23296 41488 23348 41497
rect 23848 41531 23900 41540
rect 23848 41497 23857 41531
rect 23857 41497 23891 41531
rect 23891 41497 23900 41531
rect 23848 41488 23900 41497
rect 24032 41420 24084 41472
rect 6814 41318 6866 41370
rect 6878 41318 6930 41370
rect 6942 41318 6994 41370
rect 7006 41318 7058 41370
rect 7070 41318 7122 41370
rect 12679 41318 12731 41370
rect 12743 41318 12795 41370
rect 12807 41318 12859 41370
rect 12871 41318 12923 41370
rect 12935 41318 12987 41370
rect 18544 41318 18596 41370
rect 18608 41318 18660 41370
rect 18672 41318 18724 41370
rect 18736 41318 18788 41370
rect 18800 41318 18852 41370
rect 24409 41318 24461 41370
rect 24473 41318 24525 41370
rect 24537 41318 24589 41370
rect 24601 41318 24653 41370
rect 24665 41318 24717 41370
rect 3700 41216 3752 41268
rect 2412 41148 2464 41200
rect 4436 41216 4488 41268
rect 4712 41216 4764 41268
rect 4344 41148 4396 41200
rect 5172 41148 5224 41200
rect 5540 41148 5592 41200
rect 5632 41191 5684 41200
rect 5632 41157 5641 41191
rect 5641 41157 5675 41191
rect 5675 41157 5684 41191
rect 5632 41148 5684 41157
rect 6000 41259 6052 41268
rect 6000 41225 6009 41259
rect 6009 41225 6043 41259
rect 6043 41225 6052 41259
rect 6000 41216 6052 41225
rect 7656 41216 7708 41268
rect 1400 41123 1452 41132
rect 1400 41089 1409 41123
rect 1409 41089 1443 41123
rect 1443 41089 1452 41123
rect 1400 41080 1452 41089
rect 2504 41123 2556 41132
rect 2504 41089 2513 41123
rect 2513 41089 2547 41123
rect 2547 41089 2556 41123
rect 2504 41080 2556 41089
rect 4436 41080 4488 41132
rect 5080 41080 5132 41132
rect 5448 41080 5500 41132
rect 848 41012 900 41064
rect 2320 41012 2372 41064
rect 2964 41055 3016 41064
rect 2964 41021 2973 41055
rect 2973 41021 3007 41055
rect 3007 41021 3016 41055
rect 2964 41012 3016 41021
rect 5816 41080 5868 41132
rect 7564 41191 7616 41200
rect 7564 41157 7573 41191
rect 7573 41157 7607 41191
rect 7607 41157 7616 41191
rect 7564 41148 7616 41157
rect 8484 41148 8536 41200
rect 13912 41148 13964 41200
rect 21088 41216 21140 41268
rect 5724 41012 5776 41064
rect 8116 41080 8168 41132
rect 8668 41080 8720 41132
rect 19248 41123 19300 41132
rect 19248 41089 19257 41123
rect 19257 41089 19291 41123
rect 19291 41089 19300 41123
rect 19248 41080 19300 41089
rect 20996 41148 21048 41200
rect 22192 41216 22244 41268
rect 22652 41216 22704 41268
rect 23112 41216 23164 41268
rect 23388 41259 23440 41268
rect 23388 41225 23397 41259
rect 23397 41225 23431 41259
rect 23431 41225 23440 41259
rect 23388 41216 23440 41225
rect 23480 41216 23532 41268
rect 23848 41216 23900 41268
rect 24768 41216 24820 41268
rect 7748 41012 7800 41064
rect 16212 41012 16264 41064
rect 6000 40944 6052 40996
rect 21272 41080 21324 41132
rect 21456 41080 21508 41132
rect 22008 41080 22060 41132
rect 22192 41123 22244 41132
rect 22192 41089 22201 41123
rect 22201 41089 22235 41123
rect 22235 41089 22244 41123
rect 22192 41080 22244 41089
rect 22468 41123 22520 41132
rect 22468 41089 22477 41123
rect 22477 41089 22511 41123
rect 22511 41089 22520 41123
rect 22468 41080 22520 41089
rect 21916 41012 21968 41064
rect 23112 41123 23164 41132
rect 23112 41089 23121 41123
rect 23121 41089 23155 41123
rect 23155 41089 23164 41123
rect 23112 41080 23164 41089
rect 23848 41080 23900 41132
rect 2136 40876 2188 40928
rect 2688 40876 2740 40928
rect 3240 40876 3292 40928
rect 4344 40876 4396 40928
rect 6552 40919 6604 40928
rect 6552 40885 6561 40919
rect 6561 40885 6595 40919
rect 6595 40885 6604 40919
rect 6552 40876 6604 40885
rect 17040 40876 17092 40928
rect 23664 40876 23716 40928
rect 23756 40876 23808 40928
rect 3882 40774 3934 40826
rect 3946 40774 3998 40826
rect 4010 40774 4062 40826
rect 4074 40774 4126 40826
rect 4138 40774 4190 40826
rect 9747 40774 9799 40826
rect 9811 40774 9863 40826
rect 9875 40774 9927 40826
rect 9939 40774 9991 40826
rect 10003 40774 10055 40826
rect 15612 40774 15664 40826
rect 15676 40774 15728 40826
rect 15740 40774 15792 40826
rect 15804 40774 15856 40826
rect 15868 40774 15920 40826
rect 21477 40774 21529 40826
rect 21541 40774 21593 40826
rect 21605 40774 21657 40826
rect 21669 40774 21721 40826
rect 21733 40774 21785 40826
rect 2688 40672 2740 40724
rect 3424 40715 3476 40724
rect 3424 40681 3433 40715
rect 3433 40681 3467 40715
rect 3467 40681 3476 40715
rect 3424 40672 3476 40681
rect 4068 40672 4120 40724
rect 4712 40672 4764 40724
rect 5724 40672 5776 40724
rect 5908 40672 5960 40724
rect 6092 40672 6144 40724
rect 7196 40715 7248 40724
rect 7196 40681 7205 40715
rect 7205 40681 7239 40715
rect 7239 40681 7248 40715
rect 7196 40672 7248 40681
rect 19248 40672 19300 40724
rect 19984 40672 20036 40724
rect 21824 40672 21876 40724
rect 21916 40715 21968 40724
rect 21916 40681 21925 40715
rect 21925 40681 21959 40715
rect 21959 40681 21968 40715
rect 21916 40672 21968 40681
rect 22468 40672 22520 40724
rect 23296 40672 23348 40724
rect 25228 40672 25280 40724
rect 2136 40579 2188 40588
rect 2136 40545 2145 40579
rect 2145 40545 2179 40579
rect 2179 40545 2188 40579
rect 2136 40536 2188 40545
rect 2412 40579 2464 40588
rect 2412 40545 2421 40579
rect 2421 40545 2455 40579
rect 2455 40545 2464 40579
rect 2412 40536 2464 40545
rect 3240 40536 3292 40588
rect 7472 40604 7524 40656
rect 7840 40604 7892 40656
rect 21088 40647 21140 40656
rect 21088 40613 21097 40647
rect 21097 40613 21131 40647
rect 21131 40613 21140 40647
rect 21088 40604 21140 40613
rect 22376 40604 22428 40656
rect 23020 40604 23072 40656
rect 24952 40604 25004 40656
rect 6276 40536 6328 40588
rect 9496 40536 9548 40588
rect 20812 40536 20864 40588
rect 1676 40511 1728 40520
rect 1676 40477 1685 40511
rect 1685 40477 1719 40511
rect 1719 40477 1728 40511
rect 1676 40468 1728 40477
rect 2688 40511 2740 40520
rect 2688 40477 2697 40511
rect 2697 40477 2731 40511
rect 2731 40477 2740 40511
rect 2688 40468 2740 40477
rect 3608 40511 3660 40520
rect 3608 40477 3617 40511
rect 3617 40477 3651 40511
rect 3651 40477 3660 40511
rect 3608 40468 3660 40477
rect 4252 40468 4304 40520
rect 3240 40400 3292 40452
rect 4436 40443 4488 40452
rect 4436 40409 4445 40443
rect 4445 40409 4479 40443
rect 4479 40409 4488 40443
rect 4436 40400 4488 40409
rect 6184 40511 6236 40520
rect 6184 40477 6193 40511
rect 6193 40477 6227 40511
rect 6227 40477 6236 40511
rect 6184 40468 6236 40477
rect 5540 40443 5592 40452
rect 5540 40409 5549 40443
rect 5549 40409 5583 40443
rect 5583 40409 5592 40443
rect 5540 40400 5592 40409
rect 5632 40400 5684 40452
rect 5908 40400 5960 40452
rect 2320 40332 2372 40384
rect 2964 40332 3016 40384
rect 5724 40332 5776 40384
rect 7196 40468 7248 40520
rect 10508 40468 10560 40520
rect 21916 40536 21968 40588
rect 23664 40536 23716 40588
rect 13544 40400 13596 40452
rect 20812 40400 20864 40452
rect 22100 40511 22152 40520
rect 22100 40477 22109 40511
rect 22109 40477 22143 40511
rect 22143 40477 22152 40511
rect 22100 40468 22152 40477
rect 22468 40468 22520 40520
rect 23296 40511 23348 40520
rect 23296 40477 23305 40511
rect 23305 40477 23339 40511
rect 23339 40477 23348 40511
rect 23296 40468 23348 40477
rect 19708 40332 19760 40384
rect 23204 40400 23256 40452
rect 23756 40400 23808 40452
rect 22652 40375 22704 40384
rect 22652 40341 22661 40375
rect 22661 40341 22695 40375
rect 22695 40341 22704 40375
rect 22652 40332 22704 40341
rect 6814 40230 6866 40282
rect 6878 40230 6930 40282
rect 6942 40230 6994 40282
rect 7006 40230 7058 40282
rect 7070 40230 7122 40282
rect 12679 40230 12731 40282
rect 12743 40230 12795 40282
rect 12807 40230 12859 40282
rect 12871 40230 12923 40282
rect 12935 40230 12987 40282
rect 18544 40230 18596 40282
rect 18608 40230 18660 40282
rect 18672 40230 18724 40282
rect 18736 40230 18788 40282
rect 18800 40230 18852 40282
rect 24409 40230 24461 40282
rect 24473 40230 24525 40282
rect 24537 40230 24589 40282
rect 24601 40230 24653 40282
rect 24665 40230 24717 40282
rect 2688 40128 2740 40180
rect 388 40060 440 40112
rect 6552 40128 6604 40180
rect 19340 40128 19392 40180
rect 22008 40171 22060 40180
rect 22008 40137 22017 40171
rect 22017 40137 22051 40171
rect 22051 40137 22060 40171
rect 22008 40128 22060 40137
rect 2964 40103 3016 40112
rect 2964 40069 2973 40103
rect 2973 40069 3007 40103
rect 3007 40069 3016 40103
rect 2964 40060 3016 40069
rect 3516 40060 3568 40112
rect 6460 40060 6512 40112
rect 2320 39992 2372 40044
rect 3424 39992 3476 40044
rect 4804 39992 4856 40044
rect 6736 39992 6788 40044
rect 19892 40060 19944 40112
rect 22652 40128 22704 40180
rect 22928 40171 22980 40180
rect 22928 40137 22937 40171
rect 22937 40137 22971 40171
rect 22971 40137 22980 40171
rect 22928 40128 22980 40137
rect 23572 40128 23624 40180
rect 23664 40128 23716 40180
rect 10508 39992 10560 40044
rect 10968 39992 11020 40044
rect 16580 39992 16632 40044
rect 22376 39992 22428 40044
rect 23020 39992 23072 40044
rect 25504 40060 25556 40112
rect 1584 39967 1636 39976
rect 1584 39933 1593 39967
rect 1593 39933 1627 39967
rect 1627 39933 1636 39967
rect 1584 39924 1636 39933
rect 3700 39924 3752 39976
rect 3792 39967 3844 39976
rect 3792 39933 3801 39967
rect 3801 39933 3835 39967
rect 3835 39933 3844 39967
rect 3792 39924 3844 39933
rect 3976 39967 4028 39976
rect 3976 39933 3985 39967
rect 3985 39933 4019 39967
rect 4019 39933 4028 39967
rect 3976 39924 4028 39933
rect 3516 39788 3568 39840
rect 4988 39831 5040 39840
rect 4988 39797 4997 39831
rect 4997 39797 5031 39831
rect 5031 39797 5040 39831
rect 4988 39788 5040 39797
rect 5632 39899 5684 39908
rect 5632 39865 5641 39899
rect 5641 39865 5675 39899
rect 5675 39865 5684 39899
rect 5632 39856 5684 39865
rect 6184 39856 6236 39908
rect 7656 39924 7708 39976
rect 13636 39856 13688 39908
rect 7380 39831 7432 39840
rect 7380 39797 7389 39831
rect 7389 39797 7423 39831
rect 7423 39797 7432 39831
rect 7380 39788 7432 39797
rect 8300 39788 8352 39840
rect 10784 39788 10836 39840
rect 21272 39788 21324 39840
rect 23572 39788 23624 39840
rect 24124 39831 24176 39840
rect 24124 39797 24133 39831
rect 24133 39797 24167 39831
rect 24167 39797 24176 39831
rect 24124 39788 24176 39797
rect 3882 39686 3934 39738
rect 3946 39686 3998 39738
rect 4010 39686 4062 39738
rect 4074 39686 4126 39738
rect 4138 39686 4190 39738
rect 9747 39686 9799 39738
rect 9811 39686 9863 39738
rect 9875 39686 9927 39738
rect 9939 39686 9991 39738
rect 10003 39686 10055 39738
rect 15612 39686 15664 39738
rect 15676 39686 15728 39738
rect 15740 39686 15792 39738
rect 15804 39686 15856 39738
rect 15868 39686 15920 39738
rect 21477 39686 21529 39738
rect 21541 39686 21593 39738
rect 21605 39686 21657 39738
rect 21669 39686 21721 39738
rect 21733 39686 21785 39738
rect 2228 39584 2280 39636
rect 2596 39584 2648 39636
rect 1492 39516 1544 39568
rect 1860 39355 1912 39364
rect 1860 39321 1869 39355
rect 1869 39321 1903 39355
rect 1903 39321 1912 39355
rect 1860 39312 1912 39321
rect 2504 39380 2556 39432
rect 2688 39380 2740 39432
rect 3792 39423 3844 39432
rect 3792 39389 3801 39423
rect 3801 39389 3835 39423
rect 3835 39389 3844 39423
rect 3792 39380 3844 39389
rect 3056 39312 3108 39364
rect 4988 39448 5040 39500
rect 4528 39423 4580 39432
rect 4528 39389 4537 39423
rect 4537 39389 4571 39423
rect 4571 39389 4580 39423
rect 4528 39380 4580 39389
rect 4712 39380 4764 39432
rect 3332 39287 3384 39296
rect 3332 39253 3341 39287
rect 3341 39253 3375 39287
rect 3375 39253 3384 39287
rect 3332 39244 3384 39253
rect 4896 39244 4948 39296
rect 5080 39355 5132 39364
rect 5080 39321 5089 39355
rect 5089 39321 5123 39355
rect 5123 39321 5132 39355
rect 5080 39312 5132 39321
rect 5172 39355 5224 39364
rect 5172 39321 5181 39355
rect 5181 39321 5215 39355
rect 5215 39321 5224 39355
rect 5172 39312 5224 39321
rect 5908 39380 5960 39432
rect 8208 39584 8260 39636
rect 9404 39584 9456 39636
rect 10232 39584 10284 39636
rect 21364 39584 21416 39636
rect 23204 39584 23256 39636
rect 23296 39584 23348 39636
rect 21916 39516 21968 39568
rect 20352 39448 20404 39500
rect 6184 39380 6236 39432
rect 8116 39380 8168 39432
rect 7288 39312 7340 39364
rect 5632 39244 5684 39296
rect 6000 39244 6052 39296
rect 6092 39287 6144 39296
rect 6092 39253 6101 39287
rect 6101 39253 6135 39287
rect 6135 39253 6144 39287
rect 6092 39244 6144 39253
rect 6460 39244 6512 39296
rect 7472 39244 7524 39296
rect 7932 39244 7984 39296
rect 9496 39423 9548 39432
rect 9496 39389 9505 39423
rect 9505 39389 9539 39423
rect 9539 39389 9548 39423
rect 9496 39380 9548 39389
rect 9588 39423 9640 39432
rect 9588 39389 9597 39423
rect 9597 39389 9631 39423
rect 9631 39389 9640 39423
rect 9588 39380 9640 39389
rect 9312 39244 9364 39296
rect 9404 39244 9456 39296
rect 9496 39244 9548 39296
rect 12440 39380 12492 39432
rect 19524 39423 19576 39432
rect 19524 39389 19533 39423
rect 19533 39389 19567 39423
rect 19567 39389 19576 39423
rect 19524 39380 19576 39389
rect 9772 39312 9824 39364
rect 22560 39423 22612 39432
rect 22560 39389 22569 39423
rect 22569 39389 22603 39423
rect 22603 39389 22612 39423
rect 22560 39380 22612 39389
rect 23204 39380 23256 39432
rect 23572 39423 23624 39432
rect 23572 39389 23581 39423
rect 23581 39389 23615 39423
rect 23615 39389 23624 39423
rect 23572 39380 23624 39389
rect 25228 39448 25280 39500
rect 10416 39244 10468 39296
rect 12072 39244 12124 39296
rect 23480 39244 23532 39296
rect 24860 39244 24912 39296
rect 6814 39142 6866 39194
rect 6878 39142 6930 39194
rect 6942 39142 6994 39194
rect 7006 39142 7058 39194
rect 7070 39142 7122 39194
rect 12679 39142 12731 39194
rect 12743 39142 12795 39194
rect 12807 39142 12859 39194
rect 12871 39142 12923 39194
rect 12935 39142 12987 39194
rect 18544 39142 18596 39194
rect 18608 39142 18660 39194
rect 18672 39142 18724 39194
rect 18736 39142 18788 39194
rect 18800 39142 18852 39194
rect 24409 39142 24461 39194
rect 24473 39142 24525 39194
rect 24537 39142 24589 39194
rect 24601 39142 24653 39194
rect 24665 39142 24717 39194
rect 3424 39040 3476 39092
rect 5172 39040 5224 39092
rect 2320 38972 2372 39024
rect 2044 38904 2096 38956
rect 2688 38904 2740 38956
rect 2780 38947 2832 38956
rect 2780 38913 2789 38947
rect 2789 38913 2823 38947
rect 2823 38913 2832 38947
rect 2780 38904 2832 38913
rect 3056 38904 3108 38956
rect 3976 38904 4028 38956
rect 4344 38947 4396 38956
rect 4344 38913 4353 38947
rect 4353 38913 4387 38947
rect 4387 38913 4396 38947
rect 4344 38904 4396 38913
rect 9588 39040 9640 39092
rect 9772 39083 9824 39092
rect 9772 39049 9781 39083
rect 9781 39049 9815 39083
rect 9815 39049 9824 39083
rect 9772 39040 9824 39049
rect 9496 38972 9548 39024
rect 10048 39015 10100 39024
rect 10048 38981 10057 39015
rect 10057 38981 10091 39015
rect 10091 38981 10100 39015
rect 10048 38972 10100 38981
rect 10416 39040 10468 39092
rect 20352 39083 20404 39092
rect 20352 39049 20361 39083
rect 20361 39049 20395 39083
rect 20395 39049 20404 39083
rect 20352 39040 20404 39049
rect 22560 39040 22612 39092
rect 23940 39040 23992 39092
rect 10692 38972 10744 39024
rect 10968 38972 11020 39024
rect 21088 38972 21140 39024
rect 7656 38947 7708 38956
rect 7656 38913 7665 38947
rect 7665 38913 7699 38947
rect 7699 38913 7708 38947
rect 7656 38904 7708 38913
rect 7748 38947 7800 38956
rect 7748 38913 7782 38947
rect 7782 38913 7800 38947
rect 7748 38904 7800 38913
rect 7932 38947 7984 38956
rect 7932 38913 7941 38947
rect 7941 38913 7975 38947
rect 7975 38913 7984 38947
rect 7932 38904 7984 38913
rect 8944 38947 8996 38956
rect 8944 38913 8953 38947
rect 8953 38913 8987 38947
rect 8987 38913 8996 38947
rect 8944 38904 8996 38913
rect 12072 38904 12124 38956
rect 20536 38947 20588 38956
rect 20536 38913 20545 38947
rect 20545 38913 20579 38947
rect 20579 38913 20588 38947
rect 20536 38904 20588 38913
rect 22008 38947 22060 38956
rect 22008 38913 22017 38947
rect 22017 38913 22051 38947
rect 22051 38913 22060 38947
rect 22008 38904 22060 38913
rect 23204 38972 23256 39024
rect 3608 38879 3660 38888
rect 3608 38845 3617 38879
rect 3617 38845 3651 38879
rect 3651 38845 3660 38879
rect 3608 38836 3660 38845
rect 3700 38836 3752 38888
rect 4528 38836 4580 38888
rect 4712 38836 4764 38888
rect 6368 38836 6420 38888
rect 6552 38836 6604 38888
rect 2136 38768 2188 38820
rect 2504 38768 2556 38820
rect 4804 38768 4856 38820
rect 7380 38879 7432 38888
rect 7380 38845 7389 38879
rect 7389 38845 7423 38879
rect 7423 38845 7432 38879
rect 7380 38836 7432 38845
rect 10232 38836 10284 38888
rect 20996 38836 21048 38888
rect 14648 38768 14700 38820
rect 1492 38700 1544 38752
rect 3424 38700 3476 38752
rect 3608 38700 3660 38752
rect 3700 38700 3752 38752
rect 8024 38700 8076 38752
rect 8576 38743 8628 38752
rect 8576 38709 8585 38743
rect 8585 38709 8619 38743
rect 8619 38709 8628 38743
rect 8576 38700 8628 38709
rect 10968 38700 11020 38752
rect 11704 38743 11756 38752
rect 11704 38709 11713 38743
rect 11713 38709 11747 38743
rect 11747 38709 11756 38743
rect 11704 38700 11756 38709
rect 23112 38768 23164 38820
rect 24308 38768 24360 38820
rect 24124 38743 24176 38752
rect 24124 38709 24133 38743
rect 24133 38709 24167 38743
rect 24167 38709 24176 38743
rect 24124 38700 24176 38709
rect 3882 38598 3934 38650
rect 3946 38598 3998 38650
rect 4010 38598 4062 38650
rect 4074 38598 4126 38650
rect 4138 38598 4190 38650
rect 9747 38598 9799 38650
rect 9811 38598 9863 38650
rect 9875 38598 9927 38650
rect 9939 38598 9991 38650
rect 10003 38598 10055 38650
rect 15612 38598 15664 38650
rect 15676 38598 15728 38650
rect 15740 38598 15792 38650
rect 15804 38598 15856 38650
rect 15868 38598 15920 38650
rect 21477 38598 21529 38650
rect 21541 38598 21593 38650
rect 21605 38598 21657 38650
rect 21669 38598 21721 38650
rect 21733 38598 21785 38650
rect 1032 38496 1084 38548
rect 5724 38496 5776 38548
rect 3700 38428 3752 38480
rect 4712 38428 4764 38480
rect 5448 38428 5500 38480
rect 7380 38496 7432 38548
rect 7472 38496 7524 38548
rect 3240 38360 3292 38412
rect 2780 38292 2832 38344
rect 2964 38335 3016 38344
rect 2964 38301 2973 38335
rect 2973 38301 3007 38335
rect 3007 38301 3016 38335
rect 2964 38292 3016 38301
rect 4068 38335 4120 38344
rect 4068 38301 4075 38335
rect 4075 38301 4109 38335
rect 4109 38301 4120 38335
rect 4068 38292 4120 38301
rect 4988 38292 5040 38344
rect 756 38224 808 38276
rect 2596 38224 2648 38276
rect 2872 38224 2924 38276
rect 4160 38224 4212 38276
rect 5264 38224 5316 38276
rect 5448 38267 5500 38276
rect 5448 38233 5457 38267
rect 5457 38233 5491 38267
rect 5491 38233 5500 38267
rect 5448 38224 5500 38233
rect 5816 38360 5868 38412
rect 6092 38360 6144 38412
rect 8944 38496 8996 38548
rect 10140 38496 10192 38548
rect 10232 38539 10284 38548
rect 10232 38505 10241 38539
rect 10241 38505 10275 38539
rect 10275 38505 10284 38539
rect 10232 38496 10284 38505
rect 19524 38496 19576 38548
rect 20536 38496 20588 38548
rect 23204 38496 23256 38548
rect 10416 38428 10468 38480
rect 10784 38428 10836 38480
rect 10968 38428 11020 38480
rect 10232 38360 10284 38412
rect 22008 38360 22060 38412
rect 6460 38335 6512 38344
rect 6460 38301 6469 38335
rect 6469 38301 6503 38335
rect 6503 38301 6512 38335
rect 6460 38292 6512 38301
rect 7472 38335 7524 38344
rect 7472 38301 7506 38335
rect 7506 38301 7524 38335
rect 7472 38292 7524 38301
rect 8576 38292 8628 38344
rect 9496 38335 9548 38344
rect 9496 38301 9503 38335
rect 9503 38301 9537 38335
rect 9537 38301 9548 38335
rect 9496 38292 9548 38301
rect 8208 38224 8260 38276
rect 3608 38156 3660 38208
rect 3976 38156 4028 38208
rect 7196 38156 7248 38208
rect 9220 38156 9272 38208
rect 15476 38224 15528 38276
rect 22836 38335 22888 38344
rect 22836 38301 22845 38335
rect 22845 38301 22879 38335
rect 22879 38301 22888 38335
rect 22836 38292 22888 38301
rect 23940 38335 23992 38344
rect 23940 38301 23949 38335
rect 23949 38301 23983 38335
rect 23983 38301 23992 38335
rect 23940 38292 23992 38301
rect 24860 38156 24912 38208
rect 6814 38054 6866 38106
rect 6878 38054 6930 38106
rect 6942 38054 6994 38106
rect 7006 38054 7058 38106
rect 7070 38054 7122 38106
rect 12679 38054 12731 38106
rect 12743 38054 12795 38106
rect 12807 38054 12859 38106
rect 12871 38054 12923 38106
rect 12935 38054 12987 38106
rect 18544 38054 18596 38106
rect 18608 38054 18660 38106
rect 18672 38054 18724 38106
rect 18736 38054 18788 38106
rect 18800 38054 18852 38106
rect 24409 38054 24461 38106
rect 24473 38054 24525 38106
rect 24537 38054 24589 38106
rect 24601 38054 24653 38106
rect 24665 38054 24717 38106
rect 20 37952 72 38004
rect 3976 37952 4028 38004
rect 4068 37952 4120 38004
rect 2320 37884 2372 37936
rect 2596 37816 2648 37868
rect 3148 37816 3200 37868
rect 3608 37884 3660 37936
rect 5172 37884 5224 37936
rect 1492 37791 1544 37800
rect 1492 37757 1501 37791
rect 1501 37757 1535 37791
rect 1535 37757 1544 37791
rect 1492 37748 1544 37757
rect 2596 37612 2648 37664
rect 3240 37612 3292 37664
rect 3424 37612 3476 37664
rect 4528 37816 4580 37868
rect 5632 37952 5684 38004
rect 9404 37995 9456 38004
rect 9404 37961 9413 37995
rect 9413 37961 9447 37995
rect 9447 37961 9456 37995
rect 9404 37952 9456 37961
rect 22836 37952 22888 38004
rect 23388 37995 23440 38004
rect 23388 37961 23397 37995
rect 23397 37961 23431 37995
rect 23431 37961 23440 37995
rect 23388 37952 23440 37961
rect 23940 37952 23992 38004
rect 11336 37816 11388 37868
rect 15476 37816 15528 37868
rect 5724 37748 5776 37800
rect 7656 37748 7708 37800
rect 5356 37655 5408 37664
rect 5356 37621 5365 37655
rect 5365 37621 5399 37655
rect 5399 37621 5408 37655
rect 5356 37612 5408 37621
rect 5448 37612 5500 37664
rect 7656 37612 7708 37664
rect 13544 37748 13596 37800
rect 13820 37748 13872 37800
rect 23572 37859 23624 37868
rect 23572 37825 23581 37859
rect 23581 37825 23615 37859
rect 23615 37825 23624 37859
rect 23572 37816 23624 37825
rect 23388 37748 23440 37800
rect 9128 37612 9180 37664
rect 11520 37612 11572 37664
rect 23020 37680 23072 37732
rect 12532 37655 12584 37664
rect 12532 37621 12541 37655
rect 12541 37621 12575 37655
rect 12575 37621 12584 37655
rect 12532 37612 12584 37621
rect 24124 37655 24176 37664
rect 24124 37621 24133 37655
rect 24133 37621 24167 37655
rect 24167 37621 24176 37655
rect 24124 37612 24176 37621
rect 3882 37510 3934 37562
rect 3946 37510 3998 37562
rect 4010 37510 4062 37562
rect 4074 37510 4126 37562
rect 4138 37510 4190 37562
rect 9747 37510 9799 37562
rect 9811 37510 9863 37562
rect 9875 37510 9927 37562
rect 9939 37510 9991 37562
rect 10003 37510 10055 37562
rect 15612 37510 15664 37562
rect 15676 37510 15728 37562
rect 15740 37510 15792 37562
rect 15804 37510 15856 37562
rect 15868 37510 15920 37562
rect 21477 37510 21529 37562
rect 21541 37510 21593 37562
rect 21605 37510 21657 37562
rect 21669 37510 21721 37562
rect 21733 37510 21785 37562
rect 1860 37408 1912 37460
rect 4528 37408 4580 37460
rect 4988 37408 5040 37460
rect 6184 37408 6236 37460
rect 10508 37408 10560 37460
rect 23388 37451 23440 37460
rect 23388 37417 23397 37451
rect 23397 37417 23431 37451
rect 23431 37417 23440 37451
rect 23388 37408 23440 37417
rect 23572 37408 23624 37460
rect 6552 37340 6604 37392
rect 7656 37340 7708 37392
rect 10232 37340 10284 37392
rect 12164 37340 12216 37392
rect 664 37204 716 37256
rect 2044 37315 2096 37324
rect 2044 37281 2053 37315
rect 2053 37281 2087 37315
rect 2087 37281 2096 37315
rect 2044 37272 2096 37281
rect 2320 37315 2372 37324
rect 2320 37281 2329 37315
rect 2329 37281 2363 37315
rect 2363 37281 2372 37315
rect 2320 37272 2372 37281
rect 2412 37315 2464 37324
rect 2412 37281 2446 37315
rect 2446 37281 2464 37315
rect 2412 37272 2464 37281
rect 2596 37315 2648 37324
rect 2596 37281 2605 37315
rect 2605 37281 2639 37315
rect 2639 37281 2648 37315
rect 2596 37272 2648 37281
rect 5448 37272 5500 37324
rect 10968 37272 11020 37324
rect 3240 37204 3292 37256
rect 5080 37204 5132 37256
rect 6920 37247 6972 37256
rect 6920 37213 6929 37247
rect 6929 37213 6963 37247
rect 6963 37213 6972 37247
rect 6920 37204 6972 37213
rect 3976 37136 4028 37188
rect 4896 37136 4948 37188
rect 5356 37179 5408 37188
rect 5356 37145 5365 37179
rect 5365 37145 5399 37179
rect 5399 37145 5408 37179
rect 5356 37136 5408 37145
rect 5632 37136 5684 37188
rect 5908 37136 5960 37188
rect 6000 37136 6052 37188
rect 6092 37179 6144 37188
rect 6092 37145 6101 37179
rect 6101 37145 6135 37179
rect 6135 37145 6144 37179
rect 6092 37136 6144 37145
rect 2504 37068 2556 37120
rect 2596 37068 2648 37120
rect 3884 37068 3936 37120
rect 5264 37068 5316 37120
rect 8852 37204 8904 37256
rect 9220 37204 9272 37256
rect 10232 37204 10284 37256
rect 7472 37136 7524 37188
rect 7748 37136 7800 37188
rect 8024 37136 8076 37188
rect 9404 37136 9456 37188
rect 12532 37204 12584 37256
rect 20996 37247 21048 37256
rect 20996 37213 21005 37247
rect 21005 37213 21039 37247
rect 21039 37213 21048 37247
rect 20996 37204 21048 37213
rect 21916 37247 21968 37256
rect 21916 37213 21925 37247
rect 21925 37213 21959 37247
rect 21959 37213 21968 37247
rect 21916 37204 21968 37213
rect 7932 37111 7984 37120
rect 7932 37077 7941 37111
rect 7941 37077 7975 37111
rect 7975 37077 7984 37111
rect 7932 37068 7984 37077
rect 8208 37068 8260 37120
rect 10784 37136 10836 37188
rect 11428 37179 11480 37188
rect 11428 37145 11437 37179
rect 11437 37145 11471 37179
rect 11471 37145 11480 37179
rect 11428 37136 11480 37145
rect 23572 37247 23624 37256
rect 23572 37213 23581 37247
rect 23581 37213 23615 37247
rect 23615 37213 23624 37247
rect 23572 37204 23624 37213
rect 25596 37204 25648 37256
rect 10508 37068 10560 37120
rect 23020 37068 23072 37120
rect 24860 37068 24912 37120
rect 6814 36966 6866 37018
rect 6878 36966 6930 37018
rect 6942 36966 6994 37018
rect 7006 36966 7058 37018
rect 7070 36966 7122 37018
rect 12679 36966 12731 37018
rect 12743 36966 12795 37018
rect 12807 36966 12859 37018
rect 12871 36966 12923 37018
rect 12935 36966 12987 37018
rect 18544 36966 18596 37018
rect 18608 36966 18660 37018
rect 18672 36966 18724 37018
rect 18736 36966 18788 37018
rect 18800 36966 18852 37018
rect 24409 36966 24461 37018
rect 24473 36966 24525 37018
rect 24537 36966 24589 37018
rect 24601 36966 24653 37018
rect 24665 36966 24717 37018
rect 2044 36864 2096 36916
rect 3056 36864 3108 36916
rect 4896 36864 4948 36916
rect 5264 36864 5316 36916
rect 5356 36864 5408 36916
rect 6276 36864 6328 36916
rect 10508 36864 10560 36916
rect 10968 36907 11020 36916
rect 10968 36873 10977 36907
rect 10977 36873 11011 36907
rect 11011 36873 11020 36907
rect 10968 36864 11020 36873
rect 20996 36864 21048 36916
rect 21916 36864 21968 36916
rect 4160 36839 4212 36848
rect 4160 36805 4169 36839
rect 4169 36805 4203 36839
rect 4203 36805 4212 36839
rect 4160 36796 4212 36805
rect 4436 36796 4488 36848
rect 5080 36796 5132 36848
rect 7104 36796 7156 36848
rect 7472 36839 7524 36848
rect 7472 36805 7481 36839
rect 7481 36805 7515 36839
rect 7515 36805 7524 36839
rect 7472 36796 7524 36805
rect 7564 36796 7616 36848
rect 8392 36796 8444 36848
rect 8668 36796 8720 36848
rect 2780 36771 2832 36780
rect 2780 36737 2789 36771
rect 2789 36737 2823 36771
rect 2823 36737 2832 36771
rect 2780 36728 2832 36737
rect 3056 36728 3108 36780
rect 3608 36728 3660 36780
rect 5172 36771 5224 36780
rect 5172 36737 5179 36771
rect 5179 36737 5213 36771
rect 5213 36737 5224 36771
rect 5172 36728 5224 36737
rect 7380 36728 7432 36780
rect 8208 36771 8260 36780
rect 8208 36737 8217 36771
rect 8217 36737 8251 36771
rect 8251 36737 8260 36771
rect 8208 36728 8260 36737
rect 9128 36728 9180 36780
rect 11520 36796 11572 36848
rect 13820 36796 13872 36848
rect 10140 36728 10192 36780
rect 14188 36728 14240 36780
rect 20352 36771 20404 36780
rect 20352 36737 20361 36771
rect 20361 36737 20395 36771
rect 20395 36737 20404 36771
rect 20352 36728 20404 36737
rect 1400 36703 1452 36712
rect 1400 36669 1409 36703
rect 1409 36669 1443 36703
rect 1443 36669 1452 36703
rect 1400 36660 1452 36669
rect 664 36524 716 36576
rect 2596 36592 2648 36644
rect 3700 36660 3752 36712
rect 3976 36660 4028 36712
rect 4436 36660 4488 36712
rect 4712 36660 4764 36712
rect 7932 36660 7984 36712
rect 18144 36660 18196 36712
rect 4896 36524 4948 36576
rect 10692 36592 10744 36644
rect 10968 36592 11020 36644
rect 7288 36524 7340 36576
rect 8944 36524 8996 36576
rect 9036 36524 9088 36576
rect 10232 36524 10284 36576
rect 13268 36524 13320 36576
rect 13544 36524 13596 36576
rect 19340 36524 19392 36576
rect 23572 36864 23624 36916
rect 23664 36771 23716 36780
rect 23664 36737 23673 36771
rect 23673 36737 23707 36771
rect 23707 36737 23716 36771
rect 23664 36728 23716 36737
rect 23940 36771 23992 36780
rect 23940 36737 23949 36771
rect 23949 36737 23983 36771
rect 23983 36737 23992 36771
rect 23940 36728 23992 36737
rect 24032 36660 24084 36712
rect 24952 36592 25004 36644
rect 25228 36592 25280 36644
rect 24124 36567 24176 36576
rect 24124 36533 24133 36567
rect 24133 36533 24167 36567
rect 24167 36533 24176 36567
rect 24124 36524 24176 36533
rect 3882 36422 3934 36474
rect 3946 36422 3998 36474
rect 4010 36422 4062 36474
rect 4074 36422 4126 36474
rect 4138 36422 4190 36474
rect 9747 36422 9799 36474
rect 9811 36422 9863 36474
rect 9875 36422 9927 36474
rect 9939 36422 9991 36474
rect 10003 36422 10055 36474
rect 15612 36422 15664 36474
rect 15676 36422 15728 36474
rect 15740 36422 15792 36474
rect 15804 36422 15856 36474
rect 15868 36422 15920 36474
rect 21477 36422 21529 36474
rect 21541 36422 21593 36474
rect 21605 36422 21657 36474
rect 21669 36422 21721 36474
rect 21733 36422 21785 36474
rect 2136 36184 2188 36236
rect 2596 36320 2648 36372
rect 3148 36320 3200 36372
rect 7196 36320 7248 36372
rect 7380 36184 7432 36236
rect 9128 36320 9180 36372
rect 9404 36320 9456 36372
rect 10232 36184 10284 36236
rect 23940 36320 23992 36372
rect 23848 36252 23900 36304
rect 1400 36159 1452 36168
rect 1400 36125 1409 36159
rect 1409 36125 1443 36159
rect 1443 36125 1452 36159
rect 1400 36116 1452 36125
rect 2320 36048 2372 36100
rect 5448 36159 5500 36168
rect 5448 36125 5457 36159
rect 5457 36125 5491 36159
rect 5491 36125 5500 36159
rect 5448 36116 5500 36125
rect 6644 36116 6696 36168
rect 7748 36159 7800 36168
rect 7748 36125 7757 36159
rect 7757 36125 7800 36159
rect 7748 36116 7800 36125
rect 8300 36116 8352 36168
rect 3148 35980 3200 36032
rect 4068 35980 4120 36032
rect 4436 35980 4488 36032
rect 4528 35980 4580 36032
rect 5724 36091 5776 36100
rect 5724 36057 5733 36091
rect 5733 36057 5767 36091
rect 5767 36057 5776 36091
rect 11428 36184 11480 36236
rect 14556 36159 14608 36168
rect 14556 36125 14565 36159
rect 14565 36125 14599 36159
rect 14599 36125 14608 36159
rect 14556 36116 14608 36125
rect 15016 36116 15068 36168
rect 5724 36048 5776 36057
rect 4896 35980 4948 36032
rect 5080 36023 5132 36032
rect 5080 35989 5089 36023
rect 5089 35989 5123 36023
rect 5123 35989 5132 36023
rect 5080 35980 5132 35989
rect 5448 35980 5500 36032
rect 8484 36023 8536 36032
rect 8484 35989 8493 36023
rect 8493 35989 8527 36023
rect 8527 35989 8536 36023
rect 8484 35980 8536 35989
rect 9772 35980 9824 36032
rect 10784 36048 10836 36100
rect 13176 36048 13228 36100
rect 19984 36184 20036 36236
rect 23296 36159 23348 36168
rect 23296 36125 23305 36159
rect 23305 36125 23339 36159
rect 23339 36125 23348 36159
rect 23296 36116 23348 36125
rect 23572 36159 23624 36168
rect 23572 36125 23581 36159
rect 23581 36125 23615 36159
rect 23615 36125 23624 36159
rect 23572 36116 23624 36125
rect 11796 35980 11848 36032
rect 12440 35980 12492 36032
rect 13820 35980 13872 36032
rect 14740 36023 14792 36032
rect 14740 35989 14749 36023
rect 14749 35989 14783 36023
rect 14783 35989 14792 36023
rect 14740 35980 14792 35989
rect 24952 36048 25004 36100
rect 6814 35878 6866 35930
rect 6878 35878 6930 35930
rect 6942 35878 6994 35930
rect 7006 35878 7058 35930
rect 7070 35878 7122 35930
rect 12679 35878 12731 35930
rect 12743 35878 12795 35930
rect 12807 35878 12859 35930
rect 12871 35878 12923 35930
rect 12935 35878 12987 35930
rect 18544 35878 18596 35930
rect 18608 35878 18660 35930
rect 18672 35878 18724 35930
rect 18736 35878 18788 35930
rect 18800 35878 18852 35930
rect 24409 35878 24461 35930
rect 24473 35878 24525 35930
rect 24537 35878 24589 35930
rect 24601 35878 24653 35930
rect 24665 35878 24717 35930
rect 2044 35776 2096 35828
rect 2964 35776 3016 35828
rect 3148 35776 3200 35828
rect 1768 35708 1820 35760
rect 2412 35708 2464 35760
rect 3976 35776 4028 35828
rect 6184 35776 6236 35828
rect 6736 35776 6788 35828
rect 8392 35819 8444 35828
rect 8392 35785 8401 35819
rect 8401 35785 8435 35819
rect 8435 35785 8444 35819
rect 8392 35776 8444 35785
rect 3424 35751 3476 35760
rect 3424 35717 3433 35751
rect 3433 35717 3467 35751
rect 3467 35717 3476 35751
rect 3424 35708 3476 35717
rect 4988 35708 5040 35760
rect 8944 35751 8996 35760
rect 8944 35717 8953 35751
rect 8953 35717 8987 35751
rect 8987 35717 8996 35751
rect 8944 35708 8996 35717
rect 9772 35708 9824 35760
rect 10048 35751 10100 35760
rect 10048 35717 10057 35751
rect 10057 35717 10091 35751
rect 10091 35717 10100 35751
rect 10048 35708 10100 35717
rect 2964 35640 3016 35692
rect 5080 35640 5132 35692
rect 5264 35640 5316 35692
rect 7288 35640 7340 35692
rect 7656 35683 7708 35692
rect 7656 35649 7665 35683
rect 7665 35649 7708 35683
rect 7656 35640 7708 35649
rect 9220 35683 9272 35692
rect 3332 35572 3384 35624
rect 4804 35572 4856 35624
rect 7380 35615 7432 35624
rect 7380 35581 7389 35615
rect 7389 35581 7423 35615
rect 7423 35581 7432 35615
rect 7380 35572 7432 35581
rect 1492 35436 1544 35488
rect 2412 35479 2464 35488
rect 2412 35445 2421 35479
rect 2421 35445 2455 35479
rect 2455 35445 2464 35479
rect 2412 35436 2464 35445
rect 4344 35479 4396 35488
rect 4344 35445 4353 35479
rect 4353 35445 4387 35479
rect 4387 35445 4396 35479
rect 4344 35436 4396 35445
rect 5908 35479 5960 35488
rect 5908 35445 5917 35479
rect 5917 35445 5951 35479
rect 5951 35445 5960 35479
rect 5908 35436 5960 35445
rect 9220 35649 9229 35683
rect 9229 35649 9263 35683
rect 9263 35649 9272 35683
rect 9220 35640 9272 35649
rect 10140 35640 10192 35692
rect 10232 35640 10284 35692
rect 10692 35640 10744 35692
rect 8484 35572 8536 35624
rect 13636 35776 13688 35828
rect 14556 35776 14608 35828
rect 14924 35776 14976 35828
rect 22560 35776 22612 35828
rect 23296 35776 23348 35828
rect 23664 35819 23716 35828
rect 23664 35785 23673 35819
rect 23673 35785 23707 35819
rect 23707 35785 23716 35819
rect 23664 35776 23716 35785
rect 13820 35708 13872 35760
rect 24216 35776 24268 35828
rect 14924 35640 14976 35692
rect 19340 35640 19392 35692
rect 10232 35547 10284 35556
rect 10232 35513 10241 35547
rect 10241 35513 10275 35547
rect 10275 35513 10284 35547
rect 10232 35504 10284 35513
rect 11796 35572 11848 35624
rect 12532 35615 12584 35624
rect 12532 35581 12566 35615
rect 12566 35581 12584 35615
rect 12532 35572 12584 35581
rect 12716 35615 12768 35624
rect 12716 35581 12725 35615
rect 12725 35581 12759 35615
rect 12759 35581 12768 35615
rect 12716 35572 12768 35581
rect 14740 35572 14792 35624
rect 17224 35572 17276 35624
rect 22560 35683 22612 35692
rect 22560 35649 22569 35683
rect 22569 35649 22603 35683
rect 22603 35649 22612 35683
rect 22560 35640 22612 35649
rect 22836 35683 22888 35692
rect 22836 35649 22845 35683
rect 22845 35649 22879 35683
rect 22879 35649 22888 35683
rect 22836 35640 22888 35649
rect 23204 35640 23256 35692
rect 17316 35436 17368 35488
rect 23296 35479 23348 35488
rect 23296 35445 23305 35479
rect 23305 35445 23339 35479
rect 23339 35445 23348 35479
rect 23296 35436 23348 35445
rect 23388 35479 23440 35488
rect 23388 35445 23397 35479
rect 23397 35445 23431 35479
rect 23431 35445 23440 35479
rect 23388 35436 23440 35445
rect 24124 35479 24176 35488
rect 24124 35445 24133 35479
rect 24133 35445 24167 35479
rect 24167 35445 24176 35479
rect 24124 35436 24176 35445
rect 3882 35334 3934 35386
rect 3946 35334 3998 35386
rect 4010 35334 4062 35386
rect 4074 35334 4126 35386
rect 4138 35334 4190 35386
rect 9747 35334 9799 35386
rect 9811 35334 9863 35386
rect 9875 35334 9927 35386
rect 9939 35334 9991 35386
rect 10003 35334 10055 35386
rect 15612 35334 15664 35386
rect 15676 35334 15728 35386
rect 15740 35334 15792 35386
rect 15804 35334 15856 35386
rect 15868 35334 15920 35386
rect 21477 35334 21529 35386
rect 21541 35334 21593 35386
rect 21605 35334 21657 35386
rect 21669 35334 21721 35386
rect 21733 35334 21785 35386
rect 2412 35232 2464 35284
rect 2964 35232 3016 35284
rect 3332 35232 3384 35284
rect 3608 35232 3660 35284
rect 2412 35096 2464 35148
rect 1768 35028 1820 35080
rect 2872 35071 2924 35080
rect 2872 35037 2881 35071
rect 2881 35037 2915 35071
rect 2915 35037 2924 35071
rect 2872 35028 2924 35037
rect 3516 35071 3568 35080
rect 3516 35037 3525 35071
rect 3525 35037 3559 35071
rect 3559 35037 3568 35071
rect 3516 35028 3568 35037
rect 3608 35028 3660 35080
rect 3792 35071 3844 35080
rect 3792 35037 3801 35071
rect 3801 35037 3835 35071
rect 3835 35037 3844 35071
rect 3792 35028 3844 35037
rect 3884 35028 3936 35080
rect 5724 35096 5776 35148
rect 5908 35028 5960 35080
rect 6000 35071 6052 35080
rect 6000 35037 6009 35071
rect 6009 35037 6043 35071
rect 6043 35037 6052 35071
rect 6000 35028 6052 35037
rect 4620 35003 4672 35012
rect 4620 34969 4629 35003
rect 4629 34969 4663 35003
rect 4663 34969 4672 35003
rect 4620 34960 4672 34969
rect 5448 34960 5500 35012
rect 6644 35028 6696 35080
rect 7840 35164 7892 35216
rect 8944 35164 8996 35216
rect 10692 35096 10744 35148
rect 11520 35232 11572 35284
rect 12716 35232 12768 35284
rect 14924 35232 14976 35284
rect 15016 35275 15068 35284
rect 15016 35241 15025 35275
rect 15025 35241 15059 35275
rect 15059 35241 15068 35275
rect 15016 35232 15068 35241
rect 17224 35232 17276 35284
rect 19248 35232 19300 35284
rect 7748 35028 7800 35080
rect 3424 34892 3476 34944
rect 4528 34892 4580 34944
rect 4896 34892 4948 34944
rect 4988 34892 5040 34944
rect 5172 34892 5224 34944
rect 5264 34935 5316 34944
rect 5264 34901 5273 34935
rect 5273 34901 5307 34935
rect 5307 34901 5316 34935
rect 5264 34892 5316 34901
rect 5632 34892 5684 34944
rect 6276 34892 6328 34944
rect 7472 34960 7524 35012
rect 11336 35028 11388 35080
rect 11796 35028 11848 35080
rect 14924 35071 14976 35080
rect 14924 35037 14933 35071
rect 14933 35037 14967 35071
rect 14967 35037 14976 35071
rect 14924 35028 14976 35037
rect 15200 35071 15252 35080
rect 15200 35037 15209 35071
rect 15209 35037 15243 35071
rect 15243 35037 15252 35071
rect 15200 35028 15252 35037
rect 17316 35028 17368 35080
rect 19156 35028 19208 35080
rect 20260 35028 20312 35080
rect 23204 35232 23256 35284
rect 23388 35232 23440 35284
rect 23572 35232 23624 35284
rect 6736 34892 6788 34944
rect 15108 34892 15160 34944
rect 16488 34892 16540 34944
rect 20076 34935 20128 34944
rect 20076 34901 20085 34935
rect 20085 34901 20119 34935
rect 20119 34901 20128 34935
rect 20076 34892 20128 34901
rect 20352 34935 20404 34944
rect 20352 34901 20361 34935
rect 20361 34901 20395 34935
rect 20395 34901 20404 34935
rect 20352 34892 20404 34901
rect 21732 34892 21784 34944
rect 22928 34892 22980 34944
rect 24860 34892 24912 34944
rect 6814 34790 6866 34842
rect 6878 34790 6930 34842
rect 6942 34790 6994 34842
rect 7006 34790 7058 34842
rect 7070 34790 7122 34842
rect 12679 34790 12731 34842
rect 12743 34790 12795 34842
rect 12807 34790 12859 34842
rect 12871 34790 12923 34842
rect 12935 34790 12987 34842
rect 18544 34790 18596 34842
rect 18608 34790 18660 34842
rect 18672 34790 18724 34842
rect 18736 34790 18788 34842
rect 18800 34790 18852 34842
rect 24409 34790 24461 34842
rect 24473 34790 24525 34842
rect 24537 34790 24589 34842
rect 24601 34790 24653 34842
rect 24665 34790 24717 34842
rect 2780 34731 2832 34740
rect 2780 34697 2789 34731
rect 2789 34697 2823 34731
rect 2823 34697 2832 34731
rect 2780 34688 2832 34697
rect 4988 34688 5040 34740
rect 5724 34731 5776 34740
rect 5724 34697 5733 34731
rect 5733 34697 5767 34731
rect 5767 34697 5776 34731
rect 5724 34688 5776 34697
rect 7472 34688 7524 34740
rect 9588 34688 9640 34740
rect 10324 34688 10376 34740
rect 10784 34688 10836 34740
rect 12256 34688 12308 34740
rect 4620 34620 4672 34672
rect 4804 34620 4856 34672
rect 9220 34620 9272 34672
rect 12532 34688 12584 34740
rect 20076 34688 20128 34740
rect 20260 34731 20312 34740
rect 20260 34697 20269 34731
rect 20269 34697 20303 34731
rect 20303 34697 20312 34731
rect 20260 34688 20312 34697
rect 20352 34688 20404 34740
rect 19156 34663 19208 34672
rect 19156 34629 19190 34663
rect 19190 34629 19208 34663
rect 19156 34620 19208 34629
rect 1492 34484 1544 34536
rect 2964 34484 3016 34536
rect 4896 34552 4948 34604
rect 5908 34552 5960 34604
rect 6184 34552 6236 34604
rect 10324 34552 10376 34604
rect 12256 34552 12308 34604
rect 13820 34552 13872 34604
rect 16672 34552 16724 34604
rect 18880 34595 18932 34604
rect 18880 34561 18889 34595
rect 18889 34561 18923 34595
rect 18923 34561 18932 34595
rect 18880 34552 18932 34561
rect 6092 34484 6144 34536
rect 6644 34527 6696 34536
rect 6644 34493 6653 34527
rect 6653 34493 6687 34527
rect 6687 34493 6696 34527
rect 6644 34484 6696 34493
rect 10784 34484 10836 34536
rect 20628 34552 20680 34604
rect 21824 34731 21876 34740
rect 21824 34697 21833 34731
rect 21833 34697 21867 34731
rect 21867 34697 21876 34731
rect 21824 34688 21876 34697
rect 22008 34595 22060 34604
rect 22008 34561 22017 34595
rect 22017 34561 22051 34595
rect 22051 34561 22060 34595
rect 22008 34552 22060 34561
rect 3608 34348 3660 34400
rect 4252 34348 4304 34400
rect 4620 34348 4672 34400
rect 5448 34348 5500 34400
rect 20536 34459 20588 34468
rect 20536 34425 20545 34459
rect 20545 34425 20579 34459
rect 20579 34425 20588 34459
rect 20536 34416 20588 34425
rect 21732 34416 21784 34468
rect 24124 34527 24176 34536
rect 24124 34493 24133 34527
rect 24133 34493 24167 34527
rect 24167 34493 24176 34527
rect 24124 34484 24176 34493
rect 7656 34391 7708 34400
rect 7656 34357 7665 34391
rect 7665 34357 7699 34391
rect 7699 34357 7708 34391
rect 7656 34348 7708 34357
rect 8668 34348 8720 34400
rect 11336 34348 11388 34400
rect 15108 34348 15160 34400
rect 17224 34348 17276 34400
rect 21364 34348 21416 34400
rect 22836 34348 22888 34400
rect 3882 34246 3934 34298
rect 3946 34246 3998 34298
rect 4010 34246 4062 34298
rect 4074 34246 4126 34298
rect 4138 34246 4190 34298
rect 9747 34246 9799 34298
rect 9811 34246 9863 34298
rect 9875 34246 9927 34298
rect 9939 34246 9991 34298
rect 10003 34246 10055 34298
rect 15612 34246 15664 34298
rect 15676 34246 15728 34298
rect 15740 34246 15792 34298
rect 15804 34246 15856 34298
rect 15868 34246 15920 34298
rect 21477 34246 21529 34298
rect 21541 34246 21593 34298
rect 21605 34246 21657 34298
rect 21669 34246 21721 34298
rect 21733 34246 21785 34298
rect 3608 34144 3660 34196
rect 4068 34144 4120 34196
rect 5264 34144 5316 34196
rect 8668 34187 8720 34196
rect 8668 34153 8677 34187
rect 8677 34153 8711 34187
rect 8711 34153 8720 34187
rect 8668 34144 8720 34153
rect 7840 34076 7892 34128
rect 9404 34144 9456 34196
rect 10324 34187 10376 34196
rect 10324 34153 10333 34187
rect 10333 34153 10367 34187
rect 10367 34153 10376 34187
rect 10324 34144 10376 34153
rect 10784 34187 10836 34196
rect 10784 34153 10793 34187
rect 10793 34153 10827 34187
rect 10827 34153 10836 34187
rect 10784 34144 10836 34153
rect 13268 34144 13320 34196
rect 1308 34008 1360 34060
rect 1400 33983 1452 33992
rect 1400 33949 1409 33983
rect 1409 33949 1443 33983
rect 1443 33949 1452 33983
rect 1400 33940 1452 33949
rect 1952 33983 2004 33992
rect 1952 33949 1961 33983
rect 1961 33949 1995 33983
rect 1995 33949 2004 33983
rect 1952 33940 2004 33949
rect 3700 34008 3752 34060
rect 4252 34008 4304 34060
rect 6736 34008 6788 34060
rect 1676 33915 1728 33924
rect 1676 33881 1685 33915
rect 1685 33881 1719 33915
rect 1719 33881 1728 33915
rect 1676 33872 1728 33881
rect 2228 33915 2280 33924
rect 2228 33881 2237 33915
rect 2237 33881 2271 33915
rect 2271 33881 2280 33915
rect 2228 33872 2280 33881
rect 1124 33804 1176 33856
rect 6276 33940 6328 33992
rect 6460 33940 6512 33992
rect 6644 33940 6696 33992
rect 7656 33940 7708 33992
rect 12164 34076 12216 34128
rect 12348 34076 12400 34128
rect 10324 34008 10376 34060
rect 10416 34008 10468 34060
rect 9128 33940 9180 33992
rect 9312 33983 9364 33992
rect 9312 33949 9321 33983
rect 9321 33949 9355 33983
rect 9355 33949 9364 33983
rect 9312 33940 9364 33949
rect 9496 33940 9548 33992
rect 10784 33940 10836 33992
rect 15936 34008 15988 34060
rect 19708 34144 19760 34196
rect 20628 34144 20680 34196
rect 22008 34144 22060 34196
rect 3608 33872 3660 33924
rect 4344 33915 4396 33924
rect 4344 33881 4353 33915
rect 4353 33881 4387 33915
rect 4387 33881 4396 33915
rect 4344 33872 4396 33881
rect 3240 33804 3292 33856
rect 4160 33804 4212 33856
rect 4712 33872 4764 33924
rect 4620 33804 4672 33856
rect 5080 33804 5132 33856
rect 6184 33804 6236 33856
rect 7288 33915 7340 33924
rect 7288 33881 7297 33915
rect 7297 33881 7331 33915
rect 7331 33881 7340 33915
rect 7288 33872 7340 33881
rect 10324 33872 10376 33924
rect 7932 33804 7984 33856
rect 15016 33940 15068 33992
rect 15108 33983 15160 33992
rect 15108 33949 15115 33983
rect 15115 33949 15149 33983
rect 15149 33949 15160 33983
rect 15108 33940 15160 33949
rect 19616 33940 19668 33992
rect 20076 33940 20128 33992
rect 13084 33872 13136 33924
rect 17960 33872 18012 33924
rect 18052 33872 18104 33924
rect 23848 33983 23900 33992
rect 23848 33949 23857 33983
rect 23857 33949 23891 33983
rect 23891 33949 23900 33983
rect 23848 33940 23900 33949
rect 12256 33847 12308 33856
rect 12256 33813 12265 33847
rect 12265 33813 12299 33847
rect 12299 33813 12308 33847
rect 12256 33804 12308 33813
rect 15384 33804 15436 33856
rect 17224 33804 17276 33856
rect 22744 33804 22796 33856
rect 24860 33804 24912 33856
rect 6814 33702 6866 33754
rect 6878 33702 6930 33754
rect 6942 33702 6994 33754
rect 7006 33702 7058 33754
rect 7070 33702 7122 33754
rect 12679 33702 12731 33754
rect 12743 33702 12795 33754
rect 12807 33702 12859 33754
rect 12871 33702 12923 33754
rect 12935 33702 12987 33754
rect 18544 33702 18596 33754
rect 18608 33702 18660 33754
rect 18672 33702 18724 33754
rect 18736 33702 18788 33754
rect 18800 33702 18852 33754
rect 24409 33702 24461 33754
rect 24473 33702 24525 33754
rect 24537 33702 24589 33754
rect 24601 33702 24653 33754
rect 24665 33702 24717 33754
rect 4344 33600 4396 33652
rect 4896 33600 4948 33652
rect 5632 33600 5684 33652
rect 6368 33600 6420 33652
rect 6644 33600 6696 33652
rect 7012 33600 7064 33652
rect 7472 33600 7524 33652
rect 7656 33600 7708 33652
rect 9312 33600 9364 33652
rect 10784 33600 10836 33652
rect 11704 33643 11756 33652
rect 11704 33609 11713 33643
rect 11713 33609 11747 33643
rect 11747 33609 11756 33643
rect 11704 33600 11756 33609
rect 12256 33600 12308 33652
rect 1308 33532 1360 33584
rect 1584 33464 1636 33516
rect 2136 33464 2188 33516
rect 2596 33464 2648 33516
rect 6000 33532 6052 33584
rect 6184 33532 6236 33584
rect 8208 33532 8260 33584
rect 3976 33507 4028 33516
rect 3976 33473 3985 33507
rect 3985 33473 4019 33507
rect 4019 33473 4028 33507
rect 3976 33464 4028 33473
rect 4068 33464 4120 33516
rect 4436 33464 4488 33516
rect 7932 33507 7984 33516
rect 7932 33473 7941 33507
rect 7941 33473 7984 33507
rect 7932 33464 7984 33473
rect 9404 33464 9456 33516
rect 11336 33532 11388 33584
rect 11980 33575 12032 33584
rect 11980 33541 11989 33575
rect 11989 33541 12023 33575
rect 12023 33541 12032 33575
rect 11980 33532 12032 33541
rect 13084 33600 13136 33652
rect 848 33396 900 33448
rect 1124 33396 1176 33448
rect 1492 33260 1544 33312
rect 2136 33260 2188 33312
rect 3792 33396 3844 33448
rect 7472 33396 7524 33448
rect 7656 33439 7708 33448
rect 7656 33405 7665 33439
rect 7665 33405 7699 33439
rect 7699 33405 7708 33439
rect 7656 33396 7708 33405
rect 8852 33396 8904 33448
rect 12808 33575 12860 33584
rect 12808 33541 12817 33575
rect 12817 33541 12851 33575
rect 12851 33541 12860 33575
rect 12808 33532 12860 33541
rect 10048 33439 10100 33448
rect 10048 33405 10057 33439
rect 10057 33405 10091 33439
rect 10091 33405 10100 33439
rect 10048 33396 10100 33405
rect 3332 33328 3384 33380
rect 4252 33328 4304 33380
rect 5540 33328 5592 33380
rect 7288 33328 7340 33380
rect 9496 33328 9548 33380
rect 8760 33260 8812 33312
rect 8852 33260 8904 33312
rect 12440 33507 12492 33516
rect 12440 33473 12449 33507
rect 12449 33473 12483 33507
rect 12483 33473 12492 33507
rect 12440 33464 12492 33473
rect 12532 33464 12584 33516
rect 13636 33600 13688 33652
rect 13268 33532 13320 33584
rect 16396 33600 16448 33652
rect 15568 33507 15620 33516
rect 15568 33473 15577 33507
rect 15577 33473 15611 33507
rect 15611 33473 15620 33507
rect 15568 33464 15620 33473
rect 16764 33532 16816 33584
rect 16856 33464 16908 33516
rect 17960 33464 18012 33516
rect 18880 33464 18932 33516
rect 23848 33600 23900 33652
rect 14648 33439 14700 33448
rect 14648 33405 14657 33439
rect 14657 33405 14691 33439
rect 14691 33405 14700 33439
rect 14648 33396 14700 33405
rect 14832 33439 14884 33448
rect 14832 33405 14841 33439
rect 14841 33405 14875 33439
rect 14875 33405 14884 33439
rect 14832 33396 14884 33405
rect 15292 33439 15344 33448
rect 15292 33405 15301 33439
rect 15301 33405 15335 33439
rect 15335 33405 15344 33439
rect 15292 33396 15344 33405
rect 13084 33260 13136 33312
rect 13268 33260 13320 33312
rect 14372 33260 14424 33312
rect 15108 33260 15160 33312
rect 16488 33396 16540 33448
rect 22744 33464 22796 33516
rect 21272 33260 21324 33312
rect 22192 33303 22244 33312
rect 22192 33269 22201 33303
rect 22201 33269 22235 33303
rect 22235 33269 22244 33303
rect 22192 33260 22244 33269
rect 23020 33260 23072 33312
rect 24124 33303 24176 33312
rect 24124 33269 24133 33303
rect 24133 33269 24167 33303
rect 24167 33269 24176 33303
rect 24124 33260 24176 33269
rect 3882 33158 3934 33210
rect 3946 33158 3998 33210
rect 4010 33158 4062 33210
rect 4074 33158 4126 33210
rect 4138 33158 4190 33210
rect 9747 33158 9799 33210
rect 9811 33158 9863 33210
rect 9875 33158 9927 33210
rect 9939 33158 9991 33210
rect 10003 33158 10055 33210
rect 15612 33158 15664 33210
rect 15676 33158 15728 33210
rect 15740 33158 15792 33210
rect 15804 33158 15856 33210
rect 15868 33158 15920 33210
rect 21477 33158 21529 33210
rect 21541 33158 21593 33210
rect 21605 33158 21657 33210
rect 21669 33158 21721 33210
rect 21733 33158 21785 33210
rect 6184 33056 6236 33108
rect 6736 33056 6788 33108
rect 3424 32988 3476 33040
rect 7012 32988 7064 33040
rect 8300 32988 8352 33040
rect 9220 32988 9272 33040
rect 10692 32988 10744 33040
rect 11888 32988 11940 33040
rect 1492 32852 1544 32904
rect 3332 32920 3384 32972
rect 7104 32963 7156 32972
rect 7104 32929 7113 32963
rect 7113 32929 7147 32963
rect 7147 32929 7156 32963
rect 7104 32920 7156 32929
rect 12532 32963 12584 32972
rect 12532 32929 12541 32963
rect 12541 32929 12575 32963
rect 12575 32929 12584 32963
rect 12532 32920 12584 32929
rect 13820 33056 13872 33108
rect 13636 32988 13688 33040
rect 15200 33056 15252 33108
rect 16488 33056 16540 33108
rect 17224 33056 17276 33108
rect 19064 33056 19116 33108
rect 19708 33056 19760 33108
rect 22192 33056 22244 33108
rect 25596 33056 25648 33108
rect 2044 32784 2096 32836
rect 7748 32852 7800 32904
rect 11704 32852 11756 32904
rect 12348 32852 12400 32904
rect 3148 32784 3200 32836
rect 5172 32784 5224 32836
rect 6184 32784 6236 32836
rect 6276 32784 6328 32836
rect 2596 32759 2648 32768
rect 2596 32725 2605 32759
rect 2605 32725 2639 32759
rect 2639 32725 2648 32759
rect 2596 32716 2648 32725
rect 3056 32716 3108 32768
rect 5356 32716 5408 32768
rect 6000 32716 6052 32768
rect 8116 32759 8168 32768
rect 8116 32725 8125 32759
rect 8125 32725 8159 32759
rect 8159 32725 8168 32759
rect 8116 32716 8168 32725
rect 9312 32716 9364 32768
rect 9680 32716 9732 32768
rect 11704 32716 11756 32768
rect 13084 32784 13136 32836
rect 13636 32784 13688 32836
rect 14004 32716 14056 32768
rect 14280 32895 14332 32904
rect 14280 32861 14289 32895
rect 14289 32861 14323 32895
rect 14323 32861 14332 32895
rect 14280 32852 14332 32861
rect 15108 32963 15160 32972
rect 15108 32929 15142 32963
rect 15142 32929 15160 32963
rect 15108 32920 15160 32929
rect 15844 32920 15896 32972
rect 20720 32920 20772 32972
rect 20996 32920 21048 32972
rect 14464 32852 14516 32904
rect 15292 32895 15344 32904
rect 15292 32861 15301 32895
rect 15301 32861 15335 32895
rect 15335 32861 15344 32895
rect 15292 32852 15344 32861
rect 15936 32852 15988 32904
rect 19248 32852 19300 32904
rect 21364 32895 21416 32904
rect 21364 32861 21371 32895
rect 21371 32861 21405 32895
rect 21405 32861 21416 32895
rect 21364 32852 21416 32861
rect 23020 32895 23072 32904
rect 23020 32861 23029 32895
rect 23029 32861 23063 32895
rect 23063 32861 23072 32895
rect 23020 32852 23072 32861
rect 16120 32716 16172 32768
rect 16672 32716 16724 32768
rect 17224 32716 17276 32768
rect 24860 32716 24912 32768
rect 6814 32614 6866 32666
rect 6878 32614 6930 32666
rect 6942 32614 6994 32666
rect 7006 32614 7058 32666
rect 7070 32614 7122 32666
rect 12679 32614 12731 32666
rect 12743 32614 12795 32666
rect 12807 32614 12859 32666
rect 12871 32614 12923 32666
rect 12935 32614 12987 32666
rect 18544 32614 18596 32666
rect 18608 32614 18660 32666
rect 18672 32614 18724 32666
rect 18736 32614 18788 32666
rect 18800 32614 18852 32666
rect 24409 32614 24461 32666
rect 24473 32614 24525 32666
rect 24537 32614 24589 32666
rect 24601 32614 24653 32666
rect 24665 32614 24717 32666
rect 2320 32512 2372 32564
rect 5172 32512 5224 32564
rect 5264 32512 5316 32564
rect 3608 32487 3660 32496
rect 3608 32453 3617 32487
rect 3617 32453 3651 32487
rect 3651 32453 3660 32487
rect 3608 32444 3660 32453
rect 6000 32444 6052 32496
rect 1584 32419 1636 32428
rect 1584 32385 1593 32419
rect 1593 32385 1627 32419
rect 1627 32385 1636 32419
rect 1584 32376 1636 32385
rect 2320 32419 2372 32428
rect 2320 32385 2329 32419
rect 2329 32385 2363 32419
rect 2363 32385 2372 32419
rect 2320 32376 2372 32385
rect 2596 32419 2648 32428
rect 2596 32385 2605 32419
rect 2605 32385 2639 32419
rect 2639 32385 2648 32419
rect 2596 32376 2648 32385
rect 1400 32351 1452 32360
rect 1400 32317 1409 32351
rect 1409 32317 1443 32351
rect 1443 32317 1452 32351
rect 1400 32308 1452 32317
rect 2136 32308 2188 32360
rect 2780 32308 2832 32360
rect 3424 32376 3476 32428
rect 4344 32376 4396 32428
rect 6184 32376 6236 32428
rect 9404 32555 9456 32564
rect 9404 32521 9413 32555
rect 9413 32521 9447 32555
rect 9447 32521 9456 32555
rect 9404 32512 9456 32521
rect 14924 32512 14976 32564
rect 17408 32512 17460 32564
rect 19340 32512 19392 32564
rect 6920 32376 6972 32428
rect 8760 32419 8812 32428
rect 8760 32385 8769 32419
rect 8769 32385 8803 32419
rect 8803 32385 8812 32419
rect 8760 32376 8812 32385
rect 13268 32376 13320 32428
rect 14372 32419 14424 32428
rect 14372 32385 14381 32419
rect 14381 32385 14415 32419
rect 14415 32385 14424 32419
rect 14372 32376 14424 32385
rect 3608 32308 3660 32360
rect 3792 32308 3844 32360
rect 4804 32308 4856 32360
rect 4896 32351 4948 32360
rect 4896 32317 4905 32351
rect 4905 32317 4939 32351
rect 4939 32317 4948 32351
rect 4896 32308 4948 32317
rect 7656 32308 7708 32360
rect 8116 32308 8168 32360
rect 1308 32172 1360 32224
rect 6276 32240 6328 32292
rect 8024 32240 8076 32292
rect 5908 32215 5960 32224
rect 5908 32181 5917 32215
rect 5917 32181 5951 32215
rect 5951 32181 5960 32215
rect 5908 32172 5960 32181
rect 6368 32172 6420 32224
rect 8944 32308 8996 32360
rect 9404 32308 9456 32360
rect 8484 32172 8536 32224
rect 8760 32172 8812 32224
rect 11336 32172 11388 32224
rect 13820 32351 13872 32360
rect 13820 32317 13829 32351
rect 13829 32317 13863 32351
rect 13863 32317 13872 32351
rect 13820 32308 13872 32317
rect 13636 32240 13688 32292
rect 14188 32351 14240 32360
rect 14188 32317 14222 32351
rect 14222 32317 14240 32351
rect 14188 32308 14240 32317
rect 20720 32444 20772 32496
rect 17040 32376 17092 32428
rect 18880 32419 18932 32428
rect 18880 32385 18889 32419
rect 18889 32385 18923 32419
rect 18923 32385 18932 32419
rect 18880 32376 18932 32385
rect 19156 32419 19208 32428
rect 19156 32385 19179 32419
rect 19179 32385 19208 32419
rect 19156 32376 19208 32385
rect 22652 32376 22704 32428
rect 23664 32419 23716 32428
rect 23664 32385 23673 32419
rect 23673 32385 23707 32419
rect 23707 32385 23716 32419
rect 23664 32376 23716 32385
rect 14280 32172 14332 32224
rect 14740 32172 14792 32224
rect 16856 32172 16908 32224
rect 23756 32240 23808 32292
rect 20260 32215 20312 32224
rect 20260 32181 20269 32215
rect 20269 32181 20303 32215
rect 20303 32181 20312 32215
rect 20260 32172 20312 32181
rect 24124 32215 24176 32224
rect 24124 32181 24133 32215
rect 24133 32181 24167 32215
rect 24167 32181 24176 32215
rect 24124 32172 24176 32181
rect 3882 32070 3934 32122
rect 3946 32070 3998 32122
rect 4010 32070 4062 32122
rect 4074 32070 4126 32122
rect 4138 32070 4190 32122
rect 9747 32070 9799 32122
rect 9811 32070 9863 32122
rect 9875 32070 9927 32122
rect 9939 32070 9991 32122
rect 10003 32070 10055 32122
rect 15612 32070 15664 32122
rect 15676 32070 15728 32122
rect 15740 32070 15792 32122
rect 15804 32070 15856 32122
rect 15868 32070 15920 32122
rect 21477 32070 21529 32122
rect 21541 32070 21593 32122
rect 21605 32070 21657 32122
rect 21669 32070 21721 32122
rect 21733 32070 21785 32122
rect 3700 31968 3752 32020
rect 3792 31968 3844 32020
rect 5172 31968 5224 32020
rect 5448 31968 5500 32020
rect 6736 32011 6788 32020
rect 6736 31977 6745 32011
rect 6745 31977 6779 32011
rect 6779 31977 6788 32011
rect 6736 31968 6788 31977
rect 1400 31807 1452 31816
rect 1400 31773 1409 31807
rect 1409 31773 1443 31807
rect 1443 31773 1452 31807
rect 1400 31764 1452 31773
rect 1676 31807 1728 31816
rect 1676 31773 1685 31807
rect 1685 31773 1719 31807
rect 1719 31773 1728 31807
rect 1676 31764 1728 31773
rect 2044 31807 2096 31816
rect 2044 31773 2053 31807
rect 2053 31773 2087 31807
rect 2087 31773 2096 31807
rect 2044 31764 2096 31773
rect 2596 31807 2648 31816
rect 1492 31696 1544 31748
rect 2596 31773 2603 31807
rect 2603 31773 2637 31807
rect 2637 31773 2648 31807
rect 2596 31764 2648 31773
rect 3148 31764 3200 31816
rect 3608 31832 3660 31884
rect 5356 31900 5408 31952
rect 8116 31968 8168 32020
rect 8484 31968 8536 32020
rect 9128 31968 9180 32020
rect 12624 31968 12676 32020
rect 13636 31968 13688 32020
rect 16028 31968 16080 32020
rect 5908 31832 5960 31884
rect 3332 31764 3384 31816
rect 4988 31764 5040 31816
rect 5724 31807 5776 31816
rect 5724 31773 5733 31807
rect 5733 31773 5767 31807
rect 5767 31773 5776 31807
rect 5724 31764 5776 31773
rect 7196 31832 7248 31884
rect 8668 31832 8720 31884
rect 1676 31628 1728 31680
rect 2320 31628 2372 31680
rect 5356 31696 5408 31748
rect 3332 31671 3384 31680
rect 3332 31637 3341 31671
rect 3341 31637 3375 31671
rect 3375 31637 3384 31671
rect 3332 31628 3384 31637
rect 3700 31628 3752 31680
rect 5264 31628 5316 31680
rect 5908 31696 5960 31748
rect 6460 31696 6512 31748
rect 5816 31628 5868 31680
rect 6644 31628 6696 31680
rect 6920 31628 6972 31680
rect 7104 31807 7156 31816
rect 7104 31773 7113 31807
rect 7113 31773 7147 31807
rect 7147 31773 7156 31807
rect 7104 31764 7156 31773
rect 7840 31807 7892 31816
rect 7840 31773 7849 31807
rect 7849 31773 7883 31807
rect 7883 31773 7892 31807
rect 7840 31764 7892 31773
rect 8024 31764 8076 31816
rect 14188 31900 14240 31952
rect 14924 31900 14976 31952
rect 8944 31832 8996 31884
rect 12348 31875 12400 31884
rect 12348 31841 12357 31875
rect 12357 31841 12391 31875
rect 12391 31841 12400 31875
rect 12348 31832 12400 31841
rect 14004 31832 14056 31884
rect 14740 31832 14792 31884
rect 17408 31968 17460 32020
rect 17960 31968 18012 32020
rect 18880 31968 18932 32020
rect 9864 31807 9916 31816
rect 9864 31773 9873 31807
rect 9873 31773 9907 31807
rect 9907 31773 9916 31807
rect 9864 31764 9916 31773
rect 11336 31764 11388 31816
rect 13176 31764 13228 31816
rect 13636 31764 13688 31816
rect 14372 31764 14424 31816
rect 9496 31739 9548 31748
rect 9496 31705 9505 31739
rect 9505 31705 9539 31739
rect 9539 31705 9548 31739
rect 9496 31696 9548 31705
rect 10784 31696 10836 31748
rect 7288 31628 7340 31680
rect 7380 31628 7432 31680
rect 7932 31628 7984 31680
rect 8024 31628 8076 31680
rect 10140 31628 10192 31680
rect 10232 31671 10284 31680
rect 10232 31637 10241 31671
rect 10241 31637 10275 31671
rect 10275 31637 10284 31671
rect 10232 31628 10284 31637
rect 13176 31628 13228 31680
rect 14464 31628 14516 31680
rect 15200 31807 15252 31816
rect 15200 31773 15207 31807
rect 15207 31773 15241 31807
rect 15241 31773 15252 31807
rect 15200 31764 15252 31773
rect 16672 31764 16724 31816
rect 17408 31764 17460 31816
rect 19800 31968 19852 32020
rect 20260 31968 20312 32020
rect 19156 31832 19208 31884
rect 20352 31943 20404 31952
rect 20352 31909 20361 31943
rect 20361 31909 20395 31943
rect 20395 31909 20404 31943
rect 20352 31900 20404 31909
rect 18788 31764 18840 31816
rect 18972 31807 19024 31816
rect 18972 31773 18981 31807
rect 18981 31773 19015 31807
rect 19015 31773 19024 31807
rect 18972 31764 19024 31773
rect 20168 31807 20220 31816
rect 20168 31773 20177 31807
rect 20177 31773 20211 31807
rect 20211 31773 20220 31807
rect 20168 31764 20220 31773
rect 23664 31968 23716 32020
rect 23388 31807 23440 31816
rect 23388 31773 23397 31807
rect 23397 31773 23431 31807
rect 23431 31773 23440 31807
rect 23388 31764 23440 31773
rect 25044 31764 25096 31816
rect 15936 31671 15988 31680
rect 15936 31637 15945 31671
rect 15945 31637 15979 31671
rect 15979 31637 15988 31671
rect 15936 31628 15988 31637
rect 17316 31671 17368 31680
rect 17316 31637 17325 31671
rect 17325 31637 17359 31671
rect 17359 31637 17368 31671
rect 17316 31628 17368 31637
rect 17500 31628 17552 31680
rect 20720 31628 20772 31680
rect 21824 31628 21876 31680
rect 6814 31526 6866 31578
rect 6878 31526 6930 31578
rect 6942 31526 6994 31578
rect 7006 31526 7058 31578
rect 7070 31526 7122 31578
rect 12679 31526 12731 31578
rect 12743 31526 12795 31578
rect 12807 31526 12859 31578
rect 12871 31526 12923 31578
rect 12935 31526 12987 31578
rect 18544 31526 18596 31578
rect 18608 31526 18660 31578
rect 18672 31526 18724 31578
rect 18736 31526 18788 31578
rect 18800 31526 18852 31578
rect 24409 31526 24461 31578
rect 24473 31526 24525 31578
rect 24537 31526 24589 31578
rect 24601 31526 24653 31578
rect 24665 31526 24717 31578
rect 4436 31424 4488 31476
rect 4528 31467 4580 31476
rect 4528 31433 4537 31467
rect 4537 31433 4571 31467
rect 4571 31433 4580 31467
rect 4528 31424 4580 31433
rect 7748 31424 7800 31476
rect 8760 31424 8812 31476
rect 9496 31424 9548 31476
rect 9772 31424 9824 31476
rect 9956 31424 10008 31476
rect 11704 31424 11756 31476
rect 12072 31424 12124 31476
rect 13268 31424 13320 31476
rect 13728 31424 13780 31476
rect 14464 31424 14516 31476
rect 1400 31399 1452 31408
rect 1400 31365 1409 31399
rect 1409 31365 1443 31399
rect 1443 31365 1452 31399
rect 1400 31356 1452 31365
rect 1308 31288 1360 31340
rect 3240 31356 3292 31408
rect 3608 31288 3660 31340
rect 3976 31288 4028 31340
rect 4620 31288 4672 31340
rect 1768 31220 1820 31272
rect 2228 31220 2280 31272
rect 2872 31220 2924 31272
rect 3332 31220 3384 31272
rect 4804 31356 4856 31408
rect 5448 31356 5500 31408
rect 6000 31356 6052 31408
rect 5172 31331 5224 31340
rect 5172 31297 5179 31331
rect 5179 31297 5213 31331
rect 5213 31297 5224 31331
rect 5172 31288 5224 31297
rect 5264 31288 5316 31340
rect 4804 31152 4856 31204
rect 7104 31152 7156 31204
rect 5908 31127 5960 31136
rect 5908 31093 5917 31127
rect 5917 31093 5951 31127
rect 5951 31093 5960 31127
rect 5908 31084 5960 31093
rect 7472 31331 7524 31340
rect 7472 31297 7481 31331
rect 7481 31297 7515 31331
rect 7515 31297 7524 31331
rect 7472 31288 7524 31297
rect 8208 31288 8260 31340
rect 8576 31288 8628 31340
rect 9128 31356 9180 31408
rect 9036 31288 9088 31340
rect 9680 31331 9732 31340
rect 9680 31297 9689 31331
rect 9689 31297 9732 31331
rect 9680 31288 9732 31297
rect 10324 31288 10376 31340
rect 10968 31288 11020 31340
rect 11704 31331 11756 31340
rect 11704 31297 11713 31331
rect 11713 31297 11747 31331
rect 11747 31297 11756 31331
rect 11704 31288 11756 31297
rect 12348 31288 12400 31340
rect 13636 31356 13688 31408
rect 18972 31424 19024 31476
rect 20168 31424 20220 31476
rect 14556 31356 14608 31408
rect 18144 31356 18196 31408
rect 18880 31356 18932 31408
rect 12072 31220 12124 31272
rect 12808 31263 12860 31272
rect 12808 31229 12817 31263
rect 12817 31229 12851 31263
rect 12851 31229 12860 31263
rect 12808 31220 12860 31229
rect 14096 31220 14148 31272
rect 9036 31127 9088 31136
rect 9036 31093 9045 31127
rect 9045 31093 9079 31127
rect 9079 31093 9088 31127
rect 9036 31084 9088 31093
rect 11060 31152 11112 31204
rect 11888 31195 11940 31204
rect 11888 31161 11897 31195
rect 11897 31161 11931 31195
rect 11931 31161 11940 31195
rect 11888 31152 11940 31161
rect 12256 31084 12308 31136
rect 13636 31084 13688 31136
rect 13820 31127 13872 31136
rect 13820 31093 13829 31127
rect 13829 31093 13863 31127
rect 13863 31093 13872 31127
rect 13820 31084 13872 31093
rect 14464 31084 14516 31136
rect 17500 31331 17552 31340
rect 17500 31297 17534 31331
rect 17534 31297 17552 31331
rect 17500 31288 17552 31297
rect 17960 31288 18012 31340
rect 18420 31220 18472 31272
rect 19064 31288 19116 31340
rect 19248 31288 19300 31340
rect 23572 31331 23624 31340
rect 23572 31297 23581 31331
rect 23581 31297 23615 31331
rect 23615 31297 23624 31331
rect 23572 31288 23624 31297
rect 23848 31331 23900 31340
rect 23848 31297 23857 31331
rect 23857 31297 23891 31331
rect 23891 31297 23900 31331
rect 23848 31288 23900 31297
rect 20444 31084 20496 31136
rect 23204 31084 23256 31136
rect 23664 31127 23716 31136
rect 23664 31093 23673 31127
rect 23673 31093 23707 31127
rect 23707 31093 23716 31127
rect 23664 31084 23716 31093
rect 24124 31127 24176 31136
rect 24124 31093 24133 31127
rect 24133 31093 24167 31127
rect 24167 31093 24176 31127
rect 24124 31084 24176 31093
rect 3882 30982 3934 31034
rect 3946 30982 3998 31034
rect 4010 30982 4062 31034
rect 4074 30982 4126 31034
rect 4138 30982 4190 31034
rect 9747 30982 9799 31034
rect 9811 30982 9863 31034
rect 9875 30982 9927 31034
rect 9939 30982 9991 31034
rect 10003 30982 10055 31034
rect 15612 30982 15664 31034
rect 15676 30982 15728 31034
rect 15740 30982 15792 31034
rect 15804 30982 15856 31034
rect 15868 30982 15920 31034
rect 21477 30982 21529 31034
rect 21541 30982 21593 31034
rect 21605 30982 21657 31034
rect 21669 30982 21721 31034
rect 21733 30982 21785 31034
rect 1676 30880 1728 30932
rect 2872 30880 2924 30932
rect 3976 30880 4028 30932
rect 4436 30880 4488 30932
rect 5908 30880 5960 30932
rect 6000 30880 6052 30932
rect 7196 30880 7248 30932
rect 1400 30787 1452 30796
rect 1400 30753 1409 30787
rect 1409 30753 1443 30787
rect 1443 30753 1452 30787
rect 1400 30744 1452 30753
rect 2412 30676 2464 30728
rect 2780 30719 2832 30728
rect 2780 30685 2789 30719
rect 2789 30685 2823 30719
rect 2823 30685 2832 30719
rect 2780 30676 2832 30685
rect 2044 30540 2096 30592
rect 4160 30583 4212 30592
rect 4160 30549 4169 30583
rect 4169 30549 4203 30583
rect 4203 30549 4212 30583
rect 4160 30540 4212 30549
rect 4896 30744 4948 30796
rect 7472 30812 7524 30864
rect 10784 30880 10836 30932
rect 17500 30880 17552 30932
rect 19340 30923 19392 30932
rect 19340 30889 19349 30923
rect 19349 30889 19383 30923
rect 19383 30889 19392 30923
rect 19340 30880 19392 30889
rect 10232 30812 10284 30864
rect 7104 30744 7156 30796
rect 10508 30744 10560 30796
rect 14832 30812 14884 30864
rect 15108 30812 15160 30864
rect 15200 30812 15252 30864
rect 15568 30812 15620 30864
rect 15936 30812 15988 30864
rect 6184 30676 6236 30728
rect 7380 30676 7432 30728
rect 8116 30676 8168 30728
rect 10048 30676 10100 30728
rect 13084 30744 13136 30796
rect 17316 30744 17368 30796
rect 10968 30719 11020 30728
rect 10968 30685 10977 30719
rect 10977 30685 11020 30719
rect 10968 30676 11020 30685
rect 12072 30676 12124 30728
rect 13176 30676 13228 30728
rect 13636 30676 13688 30728
rect 14924 30676 14976 30728
rect 15200 30719 15252 30728
rect 15200 30685 15209 30719
rect 15209 30685 15243 30719
rect 15243 30685 15252 30719
rect 15200 30676 15252 30685
rect 5264 30608 5316 30660
rect 4436 30540 4488 30592
rect 4620 30583 4672 30592
rect 4620 30549 4629 30583
rect 4629 30549 4663 30583
rect 4663 30549 4672 30583
rect 4620 30540 4672 30549
rect 4804 30540 4856 30592
rect 5724 30651 5776 30660
rect 5724 30617 5733 30651
rect 5733 30617 5767 30651
rect 5767 30617 5776 30651
rect 5724 30608 5776 30617
rect 12256 30608 12308 30660
rect 5908 30583 5960 30592
rect 5908 30549 5917 30583
rect 5917 30549 5951 30583
rect 5951 30549 5960 30583
rect 5908 30540 5960 30549
rect 6368 30540 6420 30592
rect 7564 30540 7616 30592
rect 7932 30540 7984 30592
rect 9588 30540 9640 30592
rect 11152 30540 11204 30592
rect 11336 30540 11388 30592
rect 11520 30540 11572 30592
rect 11704 30583 11756 30592
rect 11704 30549 11713 30583
rect 11713 30549 11747 30583
rect 11747 30549 11756 30583
rect 11704 30540 11756 30549
rect 12072 30540 12124 30592
rect 12992 30608 13044 30660
rect 12532 30540 12584 30592
rect 13452 30583 13504 30592
rect 13452 30549 13461 30583
rect 13461 30549 13495 30583
rect 13495 30549 13504 30583
rect 13452 30540 13504 30549
rect 13636 30583 13688 30592
rect 13636 30549 13645 30583
rect 13645 30549 13679 30583
rect 13679 30549 13688 30583
rect 13636 30540 13688 30549
rect 14280 30540 14332 30592
rect 14832 30540 14884 30592
rect 16120 30719 16172 30728
rect 16120 30685 16129 30719
rect 16129 30685 16163 30719
rect 16163 30685 16172 30719
rect 16120 30676 16172 30685
rect 17500 30608 17552 30660
rect 18144 30676 18196 30728
rect 20444 30812 20496 30864
rect 19800 30719 19852 30728
rect 19800 30685 19809 30719
rect 19809 30685 19843 30719
rect 19843 30685 19852 30719
rect 19800 30676 19852 30685
rect 20996 30744 21048 30796
rect 21824 30608 21876 30660
rect 21088 30583 21140 30592
rect 21088 30549 21097 30583
rect 21097 30549 21131 30583
rect 21131 30549 21140 30583
rect 21088 30540 21140 30549
rect 22192 30540 22244 30592
rect 22836 30583 22888 30592
rect 22836 30549 22845 30583
rect 22845 30549 22879 30583
rect 22879 30549 22888 30583
rect 22836 30540 22888 30549
rect 23572 30880 23624 30932
rect 23664 30880 23716 30932
rect 23204 30719 23256 30728
rect 23204 30685 23213 30719
rect 23213 30685 23247 30719
rect 23247 30685 23256 30719
rect 23204 30676 23256 30685
rect 24032 30608 24084 30660
rect 24860 30608 24912 30660
rect 25504 30540 25556 30592
rect 6814 30438 6866 30490
rect 6878 30438 6930 30490
rect 6942 30438 6994 30490
rect 7006 30438 7058 30490
rect 7070 30438 7122 30490
rect 12679 30438 12731 30490
rect 12743 30438 12795 30490
rect 12807 30438 12859 30490
rect 12871 30438 12923 30490
rect 12935 30438 12987 30490
rect 18544 30438 18596 30490
rect 18608 30438 18660 30490
rect 18672 30438 18724 30490
rect 18736 30438 18788 30490
rect 18800 30438 18852 30490
rect 24409 30438 24461 30490
rect 24473 30438 24525 30490
rect 24537 30438 24589 30490
rect 24601 30438 24653 30490
rect 24665 30438 24717 30490
rect 2596 30243 2648 30252
rect 2596 30209 2605 30243
rect 2605 30209 2639 30243
rect 2639 30209 2648 30243
rect 2596 30200 2648 30209
rect 1860 30175 1912 30184
rect 1860 30141 1869 30175
rect 1869 30141 1903 30175
rect 1903 30141 1912 30175
rect 1860 30132 1912 30141
rect 2044 30132 2096 30184
rect 2228 30064 2280 30116
rect 2872 30175 2924 30184
rect 2872 30141 2881 30175
rect 2881 30141 2915 30175
rect 2915 30141 2924 30175
rect 2872 30132 2924 30141
rect 3056 30132 3108 30184
rect 3516 30311 3568 30320
rect 3516 30277 3525 30311
rect 3525 30277 3559 30311
rect 3559 30277 3568 30311
rect 3516 30268 3568 30277
rect 4896 30336 4948 30388
rect 5540 30336 5592 30388
rect 5908 30336 5960 30388
rect 6644 30336 6696 30388
rect 13452 30336 13504 30388
rect 15016 30336 15068 30388
rect 15108 30336 15160 30388
rect 16856 30336 16908 30388
rect 23848 30336 23900 30388
rect 10784 30268 10836 30320
rect 10968 30268 11020 30320
rect 4252 30219 4259 30252
rect 4259 30219 4293 30252
rect 4293 30219 4304 30252
rect 4252 30200 4304 30219
rect 4804 30200 4856 30252
rect 5080 30200 5132 30252
rect 5356 30243 5408 30252
rect 5356 30209 5365 30243
rect 5365 30209 5399 30243
rect 5399 30209 5408 30243
rect 5356 30200 5408 30209
rect 5908 30243 5960 30252
rect 5908 30209 5917 30243
rect 5917 30209 5951 30243
rect 5951 30209 5960 30243
rect 5908 30200 5960 30209
rect 7656 30243 7708 30252
rect 7656 30209 7663 30243
rect 7663 30209 7697 30243
rect 7697 30209 7708 30243
rect 7656 30200 7708 30209
rect 10048 30243 10100 30252
rect 10048 30209 10057 30243
rect 10057 30209 10091 30243
rect 10091 30209 10100 30243
rect 10048 30200 10100 30209
rect 10232 30200 10284 30252
rect 3976 30175 4028 30184
rect 3976 30141 3985 30175
rect 3985 30141 4019 30175
rect 4019 30141 4028 30175
rect 3976 30132 4028 30141
rect 6828 30132 6880 30184
rect 7380 30175 7432 30184
rect 7380 30141 7389 30175
rect 7389 30141 7423 30175
rect 7423 30141 7432 30175
rect 7380 30132 7432 30141
rect 1308 29996 1360 30048
rect 11520 30200 11572 30252
rect 11888 30243 11940 30252
rect 11888 30209 11897 30243
rect 11897 30209 11931 30243
rect 11931 30209 11940 30243
rect 11888 30200 11940 30209
rect 12440 30268 12492 30320
rect 13176 30268 13228 30320
rect 13268 30268 13320 30320
rect 14280 30268 14332 30320
rect 14464 30311 14516 30320
rect 14464 30277 14473 30311
rect 14473 30277 14507 30311
rect 14507 30277 14516 30311
rect 14464 30268 14516 30277
rect 14924 30200 14976 30252
rect 15384 30200 15436 30252
rect 13820 30132 13872 30184
rect 15936 30132 15988 30184
rect 22284 30268 22336 30320
rect 22376 30268 22428 30320
rect 21088 30200 21140 30252
rect 22192 30243 22244 30252
rect 22192 30209 22201 30243
rect 22201 30209 22235 30243
rect 22235 30209 22244 30243
rect 22192 30200 22244 30209
rect 17408 30132 17460 30184
rect 22836 30200 22888 30252
rect 3516 29996 3568 30048
rect 4068 29996 4120 30048
rect 6368 29996 6420 30048
rect 8392 30039 8444 30048
rect 8392 30005 8401 30039
rect 8401 30005 8435 30039
rect 8435 30005 8444 30039
rect 8392 29996 8444 30005
rect 10968 30064 11020 30116
rect 11244 30064 11296 30116
rect 13084 30064 13136 30116
rect 23572 30200 23624 30252
rect 10784 29996 10836 30048
rect 11060 30039 11112 30048
rect 11060 30005 11069 30039
rect 11069 30005 11103 30039
rect 11103 30005 11112 30039
rect 11060 29996 11112 30005
rect 11428 29996 11480 30048
rect 12348 29996 12400 30048
rect 13452 30039 13504 30048
rect 13452 30005 13461 30039
rect 13461 30005 13495 30039
rect 13495 30005 13504 30039
rect 13452 29996 13504 30005
rect 16488 29996 16540 30048
rect 16672 29996 16724 30048
rect 20904 29996 20956 30048
rect 22928 29996 22980 30048
rect 23664 30039 23716 30048
rect 23664 30005 23673 30039
rect 23673 30005 23707 30039
rect 23707 30005 23716 30039
rect 23664 29996 23716 30005
rect 24124 30039 24176 30048
rect 24124 30005 24133 30039
rect 24133 30005 24167 30039
rect 24167 30005 24176 30039
rect 24124 29996 24176 30005
rect 3882 29894 3934 29946
rect 3946 29894 3998 29946
rect 4010 29894 4062 29946
rect 4074 29894 4126 29946
rect 4138 29894 4190 29946
rect 9747 29894 9799 29946
rect 9811 29894 9863 29946
rect 9875 29894 9927 29946
rect 9939 29894 9991 29946
rect 10003 29894 10055 29946
rect 15612 29894 15664 29946
rect 15676 29894 15728 29946
rect 15740 29894 15792 29946
rect 15804 29894 15856 29946
rect 15868 29894 15920 29946
rect 21477 29894 21529 29946
rect 21541 29894 21593 29946
rect 21605 29894 21657 29946
rect 21669 29894 21721 29946
rect 21733 29894 21785 29946
rect 2872 29835 2924 29844
rect 2872 29801 2881 29835
rect 2881 29801 2915 29835
rect 2915 29801 2924 29835
rect 2872 29792 2924 29801
rect 6368 29792 6420 29844
rect 9956 29792 10008 29844
rect 10232 29792 10284 29844
rect 12532 29792 12584 29844
rect 21456 29792 21508 29844
rect 22928 29792 22980 29844
rect 23572 29792 23624 29844
rect 23664 29792 23716 29844
rect 2688 29724 2740 29776
rect 4436 29724 4488 29776
rect 1400 29656 1452 29708
rect 11796 29724 11848 29776
rect 14924 29724 14976 29776
rect 15752 29724 15804 29776
rect 16764 29767 16816 29776
rect 16764 29733 16773 29767
rect 16773 29733 16807 29767
rect 16807 29733 16816 29767
rect 16764 29724 16816 29733
rect 20720 29724 20772 29776
rect 11060 29656 11112 29708
rect 11612 29656 11664 29708
rect 12532 29656 12584 29708
rect 16672 29656 16724 29708
rect 756 29588 808 29640
rect 2136 29631 2188 29640
rect 2136 29597 2143 29631
rect 2143 29597 2177 29631
rect 2177 29597 2188 29631
rect 2136 29588 2188 29597
rect 1308 29520 1360 29572
rect 2412 29452 2464 29504
rect 2504 29452 2556 29504
rect 3424 29495 3476 29504
rect 3424 29461 3433 29495
rect 3433 29461 3467 29495
rect 3467 29461 3476 29495
rect 3424 29452 3476 29461
rect 3516 29452 3568 29504
rect 7380 29588 7432 29640
rect 8760 29588 8812 29640
rect 9220 29631 9272 29640
rect 9220 29597 9227 29631
rect 9227 29597 9261 29631
rect 9261 29597 9272 29631
rect 9220 29588 9272 29597
rect 10600 29588 10652 29640
rect 10692 29588 10744 29640
rect 11704 29588 11756 29640
rect 15660 29588 15712 29640
rect 5172 29567 5197 29572
rect 5197 29567 5224 29572
rect 5172 29520 5224 29567
rect 5632 29520 5684 29572
rect 6092 29520 6144 29572
rect 6276 29520 6328 29572
rect 6552 29520 6604 29572
rect 6828 29563 6880 29572
rect 6828 29529 6837 29563
rect 6837 29529 6871 29563
rect 6871 29529 6880 29563
rect 6828 29520 6880 29529
rect 6368 29452 6420 29504
rect 7288 29520 7340 29572
rect 10232 29520 10284 29572
rect 8944 29452 8996 29504
rect 11060 29520 11112 29572
rect 11244 29563 11296 29572
rect 11244 29529 11253 29563
rect 11253 29529 11287 29563
rect 11287 29529 11296 29563
rect 11244 29520 11296 29529
rect 13268 29520 13320 29572
rect 15568 29520 15620 29572
rect 11520 29452 11572 29504
rect 11796 29495 11848 29504
rect 11796 29461 11805 29495
rect 11805 29461 11839 29495
rect 11839 29461 11848 29495
rect 11796 29452 11848 29461
rect 12072 29452 12124 29504
rect 15476 29452 15528 29504
rect 17408 29631 17460 29640
rect 17408 29597 17415 29631
rect 17415 29597 17449 29631
rect 17449 29597 17460 29631
rect 17408 29588 17460 29597
rect 16764 29520 16816 29572
rect 17316 29520 17368 29572
rect 18880 29588 18932 29640
rect 22376 29656 22428 29708
rect 17684 29520 17736 29572
rect 19248 29520 19300 29572
rect 20352 29588 20404 29640
rect 20076 29520 20128 29572
rect 21364 29520 21416 29572
rect 23112 29588 23164 29640
rect 23480 29588 23532 29640
rect 23756 29520 23808 29572
rect 17868 29452 17920 29504
rect 21088 29452 21140 29504
rect 23664 29495 23716 29504
rect 23664 29461 23673 29495
rect 23673 29461 23707 29495
rect 23707 29461 23716 29495
rect 23664 29452 23716 29461
rect 24860 29452 24912 29504
rect 6814 29350 6866 29402
rect 6878 29350 6930 29402
rect 6942 29350 6994 29402
rect 7006 29350 7058 29402
rect 7070 29350 7122 29402
rect 12679 29350 12731 29402
rect 12743 29350 12795 29402
rect 12807 29350 12859 29402
rect 12871 29350 12923 29402
rect 12935 29350 12987 29402
rect 18544 29350 18596 29402
rect 18608 29350 18660 29402
rect 18672 29350 18724 29402
rect 18736 29350 18788 29402
rect 18800 29350 18852 29402
rect 24409 29350 24461 29402
rect 24473 29350 24525 29402
rect 24537 29350 24589 29402
rect 24601 29350 24653 29402
rect 24665 29350 24717 29402
rect 1584 29248 1636 29300
rect 3424 29248 3476 29300
rect 7288 29248 7340 29300
rect 1308 29180 1360 29232
rect 2688 29180 2740 29232
rect 2412 29155 2464 29164
rect 2412 29121 2421 29155
rect 2421 29121 2455 29155
rect 2455 29121 2464 29155
rect 2412 29112 2464 29121
rect 1400 29087 1452 29096
rect 1400 29053 1409 29087
rect 1409 29053 1443 29087
rect 1443 29053 1452 29087
rect 1400 29044 1452 29053
rect 1676 29087 1728 29096
rect 1676 29053 1685 29087
rect 1685 29053 1719 29087
rect 1719 29053 1728 29087
rect 4804 29180 4856 29232
rect 5264 29180 5316 29232
rect 3148 29112 3200 29164
rect 6092 29112 6144 29164
rect 6184 29112 6236 29164
rect 7196 29180 7248 29232
rect 10232 29248 10284 29300
rect 16672 29248 16724 29300
rect 8116 29112 8168 29164
rect 8668 29155 8720 29164
rect 8668 29121 8677 29155
rect 8677 29121 8711 29155
rect 8711 29121 8720 29155
rect 8668 29112 8720 29121
rect 8944 29155 8996 29164
rect 8944 29121 8953 29155
rect 8953 29121 8987 29155
rect 8987 29121 8996 29155
rect 8944 29112 8996 29121
rect 15384 29180 15436 29232
rect 17684 29248 17736 29300
rect 17960 29248 18012 29300
rect 1676 29044 1728 29053
rect 4252 29044 4304 29096
rect 4436 29044 4488 29096
rect 6276 29044 6328 29096
rect 7472 29044 7524 29096
rect 8024 29044 8076 29096
rect 8392 29087 8444 29096
rect 8392 29053 8401 29087
rect 8401 29053 8435 29087
rect 8435 29053 8444 29087
rect 8392 29044 8444 29053
rect 2228 28976 2280 29028
rect 2688 28976 2740 29028
rect 7196 28976 7248 29028
rect 10140 29044 10192 29096
rect 10508 29044 10560 29096
rect 10784 29112 10836 29164
rect 13084 29087 13136 29096
rect 13084 29053 13093 29087
rect 13093 29053 13127 29087
rect 13127 29053 13136 29087
rect 13084 29044 13136 29053
rect 13820 29087 13872 29096
rect 13820 29053 13829 29087
rect 13829 29053 13863 29087
rect 13863 29053 13872 29087
rect 13820 29044 13872 29053
rect 13912 29087 13964 29096
rect 13912 29053 13946 29087
rect 13946 29053 13964 29087
rect 13912 29044 13964 29053
rect 14096 29087 14148 29096
rect 14096 29053 14105 29087
rect 14105 29053 14139 29087
rect 14139 29053 14148 29087
rect 14096 29044 14148 29053
rect 14280 29044 14332 29096
rect 3700 28908 3752 28960
rect 4160 28908 4212 28960
rect 4436 28951 4488 28960
rect 4436 28917 4445 28951
rect 4445 28917 4479 28951
rect 4479 28917 4488 28951
rect 4436 28908 4488 28917
rect 5264 28908 5316 28960
rect 7840 28908 7892 28960
rect 8668 28908 8720 28960
rect 9496 28908 9548 28960
rect 10048 28908 10100 28960
rect 10508 28951 10560 28960
rect 10508 28917 10517 28951
rect 10517 28917 10551 28951
rect 10551 28917 10560 28951
rect 10508 28908 10560 28917
rect 10784 28951 10836 28960
rect 10784 28917 10793 28951
rect 10793 28917 10827 28951
rect 10827 28917 10836 28951
rect 10784 28908 10836 28917
rect 11060 28908 11112 28960
rect 11428 28908 11480 28960
rect 13544 29019 13596 29028
rect 13544 28985 13553 29019
rect 13553 28985 13587 29019
rect 13587 28985 13596 29019
rect 13544 28976 13596 28985
rect 15936 28976 15988 29028
rect 16672 29087 16724 29096
rect 16672 29053 16681 29087
rect 16681 29053 16715 29087
rect 16715 29053 16724 29087
rect 16672 29044 16724 29053
rect 16856 29155 16908 29164
rect 16856 29121 16865 29155
rect 16865 29121 16899 29155
rect 16899 29121 16908 29155
rect 16856 29112 16908 29121
rect 17684 29155 17736 29164
rect 17684 29121 17718 29155
rect 17718 29121 17736 29155
rect 17684 29112 17736 29121
rect 17868 29155 17920 29164
rect 17868 29121 17877 29155
rect 17877 29121 17911 29155
rect 17911 29121 17920 29155
rect 17868 29112 17920 29121
rect 20352 29291 20404 29300
rect 20352 29257 20361 29291
rect 20361 29257 20395 29291
rect 20395 29257 20404 29291
rect 20352 29248 20404 29257
rect 19248 29223 19300 29232
rect 19248 29189 19282 29223
rect 19282 29189 19300 29223
rect 19248 29180 19300 29189
rect 20352 29112 20404 29164
rect 17316 29087 17368 29096
rect 17316 29053 17325 29087
rect 17325 29053 17359 29087
rect 17359 29053 17368 29087
rect 17316 29044 17368 29053
rect 21088 29248 21140 29300
rect 22284 29248 22336 29300
rect 22928 29248 22980 29300
rect 23112 29248 23164 29300
rect 23480 29291 23532 29300
rect 23480 29257 23489 29291
rect 23489 29257 23523 29291
rect 23523 29257 23532 29291
rect 23480 29248 23532 29257
rect 23664 29248 23716 29300
rect 20720 29180 20772 29232
rect 21088 29155 21140 29164
rect 21088 29121 21097 29155
rect 21097 29121 21131 29155
rect 21131 29121 21140 29155
rect 21088 29112 21140 29121
rect 21456 29180 21508 29232
rect 21364 29112 21416 29164
rect 14556 28908 14608 28960
rect 16212 28908 16264 28960
rect 18972 28976 19024 29028
rect 17040 28908 17092 28960
rect 21916 28976 21968 29028
rect 23204 29019 23256 29028
rect 23204 28985 23213 29019
rect 23213 28985 23247 29019
rect 23247 28985 23256 29019
rect 23204 28976 23256 28985
rect 24124 29019 24176 29028
rect 24124 28985 24133 29019
rect 24133 28985 24167 29019
rect 24167 28985 24176 29019
rect 24124 28976 24176 28985
rect 3882 28806 3934 28858
rect 3946 28806 3998 28858
rect 4010 28806 4062 28858
rect 4074 28806 4126 28858
rect 4138 28806 4190 28858
rect 9747 28806 9799 28858
rect 9811 28806 9863 28858
rect 9875 28806 9927 28858
rect 9939 28806 9991 28858
rect 10003 28806 10055 28858
rect 15612 28806 15664 28858
rect 15676 28806 15728 28858
rect 15740 28806 15792 28858
rect 15804 28806 15856 28858
rect 15868 28806 15920 28858
rect 21477 28806 21529 28858
rect 21541 28806 21593 28858
rect 21605 28806 21657 28858
rect 21669 28806 21721 28858
rect 21733 28806 21785 28858
rect 3148 28704 3200 28756
rect 8760 28704 8812 28756
rect 1216 28500 1268 28552
rect 756 28432 808 28484
rect 2320 28432 2372 28484
rect 3700 28500 3752 28552
rect 4436 28500 4488 28552
rect 4528 28500 4580 28552
rect 3240 28432 3292 28484
rect 3792 28432 3844 28484
rect 4712 28475 4764 28484
rect 4712 28441 4721 28475
rect 4721 28441 4755 28475
rect 4755 28441 4764 28475
rect 4712 28432 4764 28441
rect 5448 28543 5500 28552
rect 5448 28509 5457 28543
rect 5457 28509 5491 28543
rect 5491 28509 5500 28543
rect 5448 28500 5500 28509
rect 9496 28568 9548 28620
rect 10692 28704 10744 28756
rect 11520 28704 11572 28756
rect 12072 28679 12124 28688
rect 12072 28645 12081 28679
rect 12081 28645 12115 28679
rect 12115 28645 12124 28679
rect 12072 28636 12124 28645
rect 8944 28500 8996 28552
rect 10600 28500 10652 28552
rect 11244 28500 11296 28552
rect 11428 28500 11480 28552
rect 13544 28704 13596 28756
rect 13820 28704 13872 28756
rect 6092 28432 6144 28484
rect 3332 28364 3384 28416
rect 4620 28364 4672 28416
rect 4896 28364 4948 28416
rect 5264 28407 5316 28416
rect 5264 28373 5273 28407
rect 5273 28373 5307 28407
rect 5307 28373 5316 28407
rect 5264 28364 5316 28373
rect 6184 28364 6236 28416
rect 7656 28364 7708 28416
rect 11612 28364 11664 28416
rect 13176 28432 13228 28484
rect 13636 28500 13688 28552
rect 13912 28500 13964 28552
rect 14188 28500 14240 28552
rect 14556 28500 14608 28552
rect 13820 28432 13872 28484
rect 14372 28432 14424 28484
rect 20628 28747 20680 28756
rect 20628 28713 20637 28747
rect 20637 28713 20671 28747
rect 20671 28713 20680 28747
rect 20628 28704 20680 28713
rect 17960 28500 18012 28552
rect 20720 28636 20772 28688
rect 20996 28568 21048 28620
rect 17592 28475 17644 28484
rect 17592 28441 17626 28475
rect 17626 28441 17644 28475
rect 19984 28500 20036 28552
rect 17592 28432 17644 28441
rect 15384 28364 15436 28416
rect 16488 28364 16540 28416
rect 18972 28364 19024 28416
rect 20076 28432 20128 28484
rect 22100 28543 22152 28552
rect 22100 28509 22109 28543
rect 22109 28509 22143 28543
rect 22143 28509 22152 28543
rect 22100 28500 22152 28509
rect 22192 28407 22244 28416
rect 22192 28373 22201 28407
rect 22201 28373 22235 28407
rect 22235 28373 22244 28407
rect 22192 28364 22244 28373
rect 24860 28364 24912 28416
rect 6814 28262 6866 28314
rect 6878 28262 6930 28314
rect 6942 28262 6994 28314
rect 7006 28262 7058 28314
rect 7070 28262 7122 28314
rect 12679 28262 12731 28314
rect 12743 28262 12795 28314
rect 12807 28262 12859 28314
rect 12871 28262 12923 28314
rect 12935 28262 12987 28314
rect 18544 28262 18596 28314
rect 18608 28262 18660 28314
rect 18672 28262 18724 28314
rect 18736 28262 18788 28314
rect 18800 28262 18852 28314
rect 24409 28262 24461 28314
rect 24473 28262 24525 28314
rect 24537 28262 24589 28314
rect 24601 28262 24653 28314
rect 24665 28262 24717 28314
rect 2320 28160 2372 28212
rect 3240 28203 3292 28212
rect 3240 28169 3249 28203
rect 3249 28169 3283 28203
rect 3283 28169 3292 28203
rect 3240 28160 3292 28169
rect 4528 28092 4580 28144
rect 4804 28135 4856 28144
rect 4804 28101 4813 28135
rect 4813 28101 4847 28135
rect 4847 28101 4856 28135
rect 4804 28092 4856 28101
rect 5816 28092 5868 28144
rect 6092 28203 6144 28212
rect 6092 28169 6101 28203
rect 6101 28169 6135 28203
rect 6135 28169 6144 28203
rect 6092 28160 6144 28169
rect 10140 28160 10192 28212
rect 11060 28160 11112 28212
rect 2320 28067 2372 28076
rect 2320 28033 2329 28067
rect 2329 28033 2363 28067
rect 2363 28033 2372 28067
rect 2320 28024 2372 28033
rect 2412 28067 2464 28076
rect 2412 28033 2446 28067
rect 2446 28033 2464 28067
rect 2412 28024 2464 28033
rect 2136 27956 2188 28008
rect 2596 27999 2648 28008
rect 2596 27965 2605 27999
rect 2605 27965 2639 27999
rect 2639 27965 2648 27999
rect 2596 27956 2648 27965
rect 1492 27888 1544 27940
rect 1768 27888 1820 27940
rect 2044 27931 2096 27940
rect 2044 27897 2053 27931
rect 2053 27897 2087 27931
rect 2087 27897 2096 27931
rect 2044 27888 2096 27897
rect 3700 28067 3752 28076
rect 3700 28033 3709 28067
rect 3709 28033 3743 28067
rect 3743 28033 3752 28067
rect 3700 28024 3752 28033
rect 5264 28024 5316 28076
rect 5632 28024 5684 28076
rect 10508 28092 10560 28144
rect 11612 28092 11664 28144
rect 11704 28135 11756 28144
rect 11704 28101 11713 28135
rect 11713 28101 11747 28135
rect 11747 28101 11756 28135
rect 11704 28092 11756 28101
rect 12900 28092 12952 28144
rect 14096 28160 14148 28212
rect 6368 28024 6420 28076
rect 6552 28024 6604 28076
rect 8208 28024 8260 28076
rect 8760 28067 8812 28076
rect 8760 28033 8769 28067
rect 8769 28033 8803 28067
rect 8803 28033 8812 28067
rect 8760 28024 8812 28033
rect 9036 28067 9088 28076
rect 9036 28033 9045 28067
rect 9045 28033 9079 28067
rect 9079 28033 9088 28067
rect 9036 28024 9088 28033
rect 10784 28024 10836 28076
rect 6184 27956 6236 28008
rect 6644 27956 6696 28008
rect 7656 27956 7708 28008
rect 1308 27820 1360 27872
rect 7748 27888 7800 27940
rect 8392 27956 8444 28008
rect 8576 27956 8628 28008
rect 9220 27956 9272 28008
rect 9404 27956 9456 28008
rect 10692 27999 10744 28008
rect 10692 27965 10701 27999
rect 10701 27965 10735 27999
rect 10735 27965 10744 27999
rect 10692 27956 10744 27965
rect 11796 28024 11848 28076
rect 12072 28067 12124 28076
rect 12072 28033 12081 28067
rect 12081 28033 12115 28067
rect 12115 28033 12124 28067
rect 12072 28024 12124 28033
rect 12440 28067 12492 28076
rect 12440 28033 12449 28067
rect 12449 28033 12483 28067
rect 12483 28033 12492 28067
rect 12440 28024 12492 28033
rect 13176 28067 13228 28076
rect 13176 28033 13185 28067
rect 13185 28033 13219 28067
rect 13219 28033 13228 28067
rect 13176 28024 13228 28033
rect 15200 28160 15252 28212
rect 16396 28160 16448 28212
rect 16764 28160 16816 28212
rect 18972 28160 19024 28212
rect 22100 28160 22152 28212
rect 22192 28160 22244 28212
rect 11612 27956 11664 28008
rect 12992 27931 13044 27940
rect 12992 27897 13001 27931
rect 13001 27897 13035 27931
rect 13035 27897 13044 27931
rect 12992 27888 13044 27897
rect 3332 27820 3384 27872
rect 6092 27820 6144 27872
rect 8760 27820 8812 27872
rect 10140 27820 10192 27872
rect 10784 27820 10836 27872
rect 15752 28024 15804 28076
rect 17592 28024 17644 28076
rect 20720 28092 20772 28144
rect 21088 28092 21140 28144
rect 20996 28024 21048 28076
rect 22652 28024 22704 28076
rect 13912 27956 13964 28008
rect 14832 27999 14884 28008
rect 14832 27965 14841 27999
rect 14841 27965 14875 27999
rect 14875 27965 14884 27999
rect 14832 27956 14884 27965
rect 15384 27956 15436 28008
rect 15568 27999 15620 28008
rect 15568 27965 15577 27999
rect 15577 27965 15611 27999
rect 15611 27965 15620 27999
rect 15568 27956 15620 27965
rect 16488 27956 16540 28008
rect 18604 27956 18656 28008
rect 18236 27888 18288 27940
rect 19708 27888 19760 27940
rect 14832 27820 14884 27872
rect 15568 27820 15620 27872
rect 16028 27820 16080 27872
rect 16396 27820 16448 27872
rect 16764 27820 16816 27872
rect 17592 27820 17644 27872
rect 22008 27820 22060 27872
rect 22744 27820 22796 27872
rect 23940 28067 23992 28076
rect 23940 28033 23949 28067
rect 23949 28033 23983 28067
rect 23983 28033 23992 28067
rect 23940 28024 23992 28033
rect 23112 27956 23164 28008
rect 23572 27863 23624 27872
rect 23572 27829 23581 27863
rect 23581 27829 23615 27863
rect 23615 27829 23624 27863
rect 23572 27820 23624 27829
rect 24124 27863 24176 27872
rect 24124 27829 24133 27863
rect 24133 27829 24167 27863
rect 24167 27829 24176 27863
rect 24124 27820 24176 27829
rect 3882 27718 3934 27770
rect 3946 27718 3998 27770
rect 4010 27718 4062 27770
rect 4074 27718 4126 27770
rect 4138 27718 4190 27770
rect 9747 27718 9799 27770
rect 9811 27718 9863 27770
rect 9875 27718 9927 27770
rect 9939 27718 9991 27770
rect 10003 27718 10055 27770
rect 15612 27718 15664 27770
rect 15676 27718 15728 27770
rect 15740 27718 15792 27770
rect 15804 27718 15856 27770
rect 15868 27718 15920 27770
rect 21477 27718 21529 27770
rect 21541 27718 21593 27770
rect 21605 27718 21657 27770
rect 21669 27718 21721 27770
rect 21733 27718 21785 27770
rect 848 27548 900 27600
rect 2596 27659 2648 27668
rect 2596 27625 2605 27659
rect 2605 27625 2639 27659
rect 2639 27625 2648 27659
rect 2596 27616 2648 27625
rect 1400 27412 1452 27464
rect 2872 27412 2924 27464
rect 2964 27455 3016 27464
rect 2964 27421 2973 27455
rect 2973 27421 3007 27455
rect 3007 27421 3016 27455
rect 2964 27412 3016 27421
rect 5448 27616 5500 27668
rect 5816 27616 5868 27668
rect 6552 27616 6604 27668
rect 15200 27616 15252 27668
rect 16488 27659 16540 27668
rect 16488 27625 16497 27659
rect 16497 27625 16531 27659
rect 16531 27625 16540 27659
rect 16488 27616 16540 27625
rect 18604 27659 18656 27668
rect 18604 27625 18613 27659
rect 18613 27625 18647 27659
rect 18647 27625 18656 27659
rect 18604 27616 18656 27625
rect 1768 27344 1820 27396
rect 4068 27412 4120 27464
rect 4988 27412 5040 27464
rect 7288 27455 7340 27464
rect 7288 27421 7295 27455
rect 7295 27421 7329 27455
rect 7329 27421 7340 27455
rect 7288 27412 7340 27421
rect 8576 27548 8628 27600
rect 11612 27548 11664 27600
rect 23112 27616 23164 27668
rect 23940 27616 23992 27668
rect 8116 27480 8168 27532
rect 9404 27480 9456 27532
rect 10140 27480 10192 27532
rect 10416 27480 10468 27532
rect 10508 27480 10560 27532
rect 17500 27480 17552 27532
rect 1308 27276 1360 27328
rect 11796 27412 11848 27464
rect 10416 27344 10468 27396
rect 13452 27344 13504 27396
rect 14096 27455 14148 27464
rect 14096 27421 14105 27455
rect 14105 27421 14139 27455
rect 14139 27421 14148 27455
rect 14096 27412 14148 27421
rect 14188 27344 14240 27396
rect 3976 27319 4028 27328
rect 3976 27285 3985 27319
rect 3985 27285 4019 27319
rect 4019 27285 4028 27319
rect 3976 27276 4028 27285
rect 5080 27276 5132 27328
rect 6368 27276 6420 27328
rect 6644 27276 6696 27328
rect 7196 27276 7248 27328
rect 7288 27276 7340 27328
rect 7748 27276 7800 27328
rect 8024 27319 8076 27328
rect 8024 27285 8033 27319
rect 8033 27285 8067 27319
rect 8067 27285 8076 27319
rect 8024 27276 8076 27285
rect 8116 27276 8168 27328
rect 8668 27276 8720 27328
rect 9036 27276 9088 27328
rect 14096 27276 14148 27328
rect 15292 27344 15344 27396
rect 16028 27344 16080 27396
rect 17224 27344 17276 27396
rect 17960 27412 18012 27464
rect 21088 27455 21140 27464
rect 21088 27421 21122 27455
rect 21122 27421 21140 27455
rect 21088 27412 21140 27421
rect 22744 27412 22796 27464
rect 23204 27480 23256 27532
rect 23296 27412 23348 27464
rect 14556 27276 14608 27328
rect 15108 27319 15160 27328
rect 15108 27285 15117 27319
rect 15117 27285 15151 27319
rect 15151 27285 15160 27319
rect 15108 27276 15160 27285
rect 16212 27276 16264 27328
rect 19340 27276 19392 27328
rect 20996 27276 21048 27328
rect 24860 27276 24912 27328
rect 6814 27174 6866 27226
rect 6878 27174 6930 27226
rect 6942 27174 6994 27226
rect 7006 27174 7058 27226
rect 7070 27174 7122 27226
rect 12679 27174 12731 27226
rect 12743 27174 12795 27226
rect 12807 27174 12859 27226
rect 12871 27174 12923 27226
rect 12935 27174 12987 27226
rect 18544 27174 18596 27226
rect 18608 27174 18660 27226
rect 18672 27174 18724 27226
rect 18736 27174 18788 27226
rect 18800 27174 18852 27226
rect 24409 27174 24461 27226
rect 24473 27174 24525 27226
rect 24537 27174 24589 27226
rect 24601 27174 24653 27226
rect 24665 27174 24717 27226
rect 2044 27072 2096 27124
rect 1216 27004 1268 27056
rect 2964 27072 3016 27124
rect 6552 27072 6604 27124
rect 6644 27072 6696 27124
rect 5632 27004 5684 27056
rect 6828 27004 6880 27056
rect 7840 27072 7892 27124
rect 7288 27047 7340 27056
rect 7288 27013 7297 27047
rect 7297 27013 7331 27047
rect 7331 27013 7340 27047
rect 7288 27004 7340 27013
rect 8024 27004 8076 27056
rect 8392 27072 8444 27124
rect 8760 27072 8812 27124
rect 11336 27072 11388 27124
rect 14188 27072 14240 27124
rect 2688 26936 2740 26988
rect 2780 26979 2832 26988
rect 2780 26945 2789 26979
rect 2789 26945 2823 26979
rect 2823 26945 2832 26979
rect 2780 26936 2832 26945
rect 2872 26936 2924 26988
rect 1400 26911 1452 26920
rect 1400 26877 1409 26911
rect 1409 26877 1443 26911
rect 1443 26877 1452 26911
rect 1400 26868 1452 26877
rect 3608 26979 3660 26988
rect 3608 26945 3617 26979
rect 3617 26945 3651 26979
rect 3651 26945 3660 26979
rect 3608 26936 3660 26945
rect 3884 26979 3936 26988
rect 3884 26945 3891 26979
rect 3891 26945 3925 26979
rect 3925 26945 3936 26979
rect 3884 26936 3936 26945
rect 3976 26936 4028 26988
rect 7472 26936 7524 26988
rect 8668 27004 8720 27056
rect 9404 26936 9456 26988
rect 7196 26868 7248 26920
rect 8392 26868 8444 26920
rect 8668 26868 8720 26920
rect 13820 27004 13872 27056
rect 15936 27004 15988 27056
rect 16212 27004 16264 27056
rect 1308 26732 1360 26784
rect 3516 26732 3568 26784
rect 4068 26732 4120 26784
rect 5356 26800 5408 26852
rect 11428 26868 11480 26920
rect 20444 27004 20496 27056
rect 17500 26936 17552 26988
rect 18144 26936 18196 26988
rect 19156 26936 19208 26988
rect 4988 26732 5040 26784
rect 5172 26732 5224 26784
rect 6368 26732 6420 26784
rect 9496 26732 9548 26784
rect 11612 26800 11664 26852
rect 16488 26800 16540 26852
rect 16856 26800 16908 26852
rect 13176 26732 13228 26784
rect 15016 26732 15068 26784
rect 17408 26732 17460 26784
rect 19800 26732 19852 26784
rect 20536 26979 20588 26988
rect 20536 26945 20545 26979
rect 20545 26945 20579 26979
rect 20579 26945 20588 26979
rect 20536 26936 20588 26945
rect 20996 27004 21048 27056
rect 23204 27004 23256 27056
rect 25136 27072 25188 27124
rect 25136 26868 25188 26920
rect 20168 26732 20220 26784
rect 20720 26775 20772 26784
rect 20720 26741 20729 26775
rect 20729 26741 20763 26775
rect 20763 26741 20772 26775
rect 20720 26732 20772 26741
rect 24124 26775 24176 26784
rect 24124 26741 24133 26775
rect 24133 26741 24167 26775
rect 24167 26741 24176 26775
rect 24124 26732 24176 26741
rect 24216 26732 24268 26784
rect 25228 26732 25280 26784
rect 3882 26630 3934 26682
rect 3946 26630 3998 26682
rect 4010 26630 4062 26682
rect 4074 26630 4126 26682
rect 4138 26630 4190 26682
rect 9747 26630 9799 26682
rect 9811 26630 9863 26682
rect 9875 26630 9927 26682
rect 9939 26630 9991 26682
rect 10003 26630 10055 26682
rect 15612 26630 15664 26682
rect 15676 26630 15728 26682
rect 15740 26630 15792 26682
rect 15804 26630 15856 26682
rect 15868 26630 15920 26682
rect 21477 26630 21529 26682
rect 21541 26630 21593 26682
rect 21605 26630 21657 26682
rect 21669 26630 21721 26682
rect 21733 26630 21785 26682
rect 6828 26528 6880 26580
rect 7196 26528 7248 26580
rect 10416 26571 10468 26580
rect 10416 26537 10425 26571
rect 10425 26537 10459 26571
rect 10459 26537 10468 26571
rect 10416 26528 10468 26537
rect 1400 26460 1452 26512
rect 2044 26460 2096 26512
rect 4436 26503 4488 26512
rect 4436 26469 4445 26503
rect 4445 26469 4479 26503
rect 4479 26469 4488 26503
rect 4436 26460 4488 26469
rect 5448 26460 5500 26512
rect 3056 26392 3108 26444
rect 3792 26435 3844 26444
rect 3792 26401 3801 26435
rect 3801 26401 3835 26435
rect 3835 26401 3844 26435
rect 3792 26392 3844 26401
rect 4344 26392 4396 26444
rect 13084 26528 13136 26580
rect 13452 26528 13504 26580
rect 19892 26528 19944 26580
rect 1216 26324 1268 26376
rect 1400 26367 1452 26376
rect 1400 26333 1409 26367
rect 1409 26333 1443 26367
rect 1443 26333 1452 26367
rect 1400 26324 1452 26333
rect 1676 26367 1728 26376
rect 1676 26333 1685 26367
rect 1685 26333 1719 26367
rect 1719 26333 1728 26367
rect 1676 26324 1728 26333
rect 2504 26324 2556 26376
rect 1952 26188 2004 26240
rect 3148 26188 3200 26240
rect 4988 26367 5040 26376
rect 4988 26333 4997 26367
rect 4997 26333 5031 26367
rect 5031 26333 5040 26367
rect 4988 26324 5040 26333
rect 5724 26324 5776 26376
rect 5816 26324 5868 26376
rect 5632 26299 5684 26308
rect 5632 26265 5641 26299
rect 5641 26265 5675 26299
rect 5675 26265 5684 26299
rect 5632 26256 5684 26265
rect 4712 26188 4764 26240
rect 6000 26188 6052 26240
rect 6276 26188 6328 26240
rect 6644 26188 6696 26240
rect 7380 26392 7432 26444
rect 7840 26324 7892 26376
rect 8484 26256 8536 26308
rect 9220 26256 9272 26308
rect 9496 26299 9548 26308
rect 9496 26265 9505 26299
rect 9505 26265 9539 26299
rect 9539 26265 9548 26299
rect 9496 26256 9548 26265
rect 14556 26435 14608 26444
rect 7380 26188 7432 26240
rect 7748 26188 7800 26240
rect 8208 26188 8260 26240
rect 10968 26367 11020 26376
rect 10968 26333 10977 26367
rect 10977 26333 11011 26367
rect 11011 26333 11020 26367
rect 10968 26324 11020 26333
rect 10692 26256 10744 26308
rect 11428 26367 11480 26376
rect 11428 26333 11437 26367
rect 11437 26333 11471 26367
rect 11471 26333 11480 26367
rect 11428 26324 11480 26333
rect 11520 26256 11572 26308
rect 12256 26324 12308 26376
rect 14556 26401 14565 26435
rect 14565 26401 14599 26435
rect 14599 26401 14608 26435
rect 14556 26392 14608 26401
rect 16304 26392 16356 26444
rect 16672 26435 16724 26444
rect 16672 26401 16681 26435
rect 16681 26401 16715 26435
rect 16715 26401 16724 26435
rect 16672 26392 16724 26401
rect 14188 26324 14240 26376
rect 15200 26324 15252 26376
rect 15292 26324 15344 26376
rect 10876 26231 10928 26240
rect 10876 26197 10885 26231
rect 10885 26197 10919 26231
rect 10919 26197 10928 26231
rect 10876 26188 10928 26197
rect 13084 26188 13136 26240
rect 13820 26188 13872 26240
rect 14188 26188 14240 26240
rect 15476 26188 15528 26240
rect 16948 26367 17000 26376
rect 17408 26392 17460 26444
rect 17960 26392 18012 26444
rect 20168 26392 20220 26444
rect 16948 26333 16975 26367
rect 16975 26333 17000 26367
rect 16948 26324 17000 26333
rect 17224 26367 17276 26376
rect 17224 26333 17233 26367
rect 17233 26333 17267 26367
rect 17267 26333 17276 26367
rect 17224 26324 17276 26333
rect 18420 26324 18472 26376
rect 19800 26367 19852 26376
rect 19800 26333 19809 26367
rect 19809 26333 19843 26367
rect 19843 26333 19852 26367
rect 19800 26324 19852 26333
rect 22376 26460 22428 26512
rect 22008 26324 22060 26376
rect 17684 26188 17736 26240
rect 20444 26256 20496 26308
rect 24124 26256 24176 26308
rect 24860 26256 24912 26308
rect 6814 26086 6866 26138
rect 6878 26086 6930 26138
rect 6942 26086 6994 26138
rect 7006 26086 7058 26138
rect 7070 26086 7122 26138
rect 12679 26086 12731 26138
rect 12743 26086 12795 26138
rect 12807 26086 12859 26138
rect 12871 26086 12923 26138
rect 12935 26086 12987 26138
rect 18544 26086 18596 26138
rect 18608 26086 18660 26138
rect 18672 26086 18724 26138
rect 18736 26086 18788 26138
rect 18800 26086 18852 26138
rect 24409 26086 24461 26138
rect 24473 26086 24525 26138
rect 24537 26086 24589 26138
rect 24601 26086 24653 26138
rect 24665 26086 24717 26138
rect 1860 25984 1912 26036
rect 2504 25984 2556 26036
rect 848 25916 900 25968
rect 4436 25984 4488 26036
rect 6276 25984 6328 26036
rect 9036 25984 9088 26036
rect 9680 25984 9732 26036
rect 10324 25984 10376 26036
rect 10692 26027 10744 26036
rect 10692 25993 10701 26027
rect 10701 25993 10735 26027
rect 10735 25993 10744 26027
rect 10692 25984 10744 25993
rect 11428 25984 11480 26036
rect 11612 25984 11664 26036
rect 13820 25984 13872 26036
rect 15200 25984 15252 26036
rect 16488 25984 16540 26036
rect 16672 25984 16724 26036
rect 17224 25984 17276 26036
rect 2412 25848 2464 25900
rect 1216 25780 1268 25832
rect 4160 25848 4212 25900
rect 5172 25887 5197 25900
rect 5197 25887 5224 25900
rect 5172 25848 5224 25887
rect 7380 25848 7432 25900
rect 8944 25848 8996 25900
rect 9864 25848 9916 25900
rect 10324 25848 10376 25900
rect 10876 25848 10928 25900
rect 11520 25891 11572 25900
rect 11520 25857 11529 25891
rect 11529 25857 11563 25891
rect 11563 25857 11572 25891
rect 11520 25848 11572 25857
rect 11704 25848 11756 25900
rect 12348 25848 12400 25900
rect 13820 25848 13872 25900
rect 14464 25916 14516 25968
rect 14740 25916 14792 25968
rect 14832 25916 14884 25968
rect 14556 25848 14608 25900
rect 18420 25916 18472 25968
rect 17224 25858 17276 25910
rect 17960 25848 18012 25900
rect 20536 25984 20588 26036
rect 21824 25984 21876 26036
rect 2412 25687 2464 25696
rect 2412 25653 2421 25687
rect 2421 25653 2455 25687
rect 2455 25653 2464 25687
rect 2412 25644 2464 25653
rect 2780 25644 2832 25696
rect 4896 25823 4948 25832
rect 4896 25789 4905 25823
rect 4905 25789 4939 25823
rect 4939 25789 4948 25823
rect 4896 25780 4948 25789
rect 9312 25780 9364 25832
rect 9496 25780 9548 25832
rect 9588 25780 9640 25832
rect 16488 25780 16540 25832
rect 3516 25644 3568 25696
rect 3608 25644 3660 25696
rect 5908 25687 5960 25696
rect 5908 25653 5917 25687
rect 5917 25653 5951 25687
rect 5951 25653 5960 25687
rect 5908 25644 5960 25653
rect 6092 25712 6144 25764
rect 6828 25712 6880 25764
rect 13820 25712 13872 25764
rect 14648 25712 14700 25764
rect 12532 25687 12584 25696
rect 12532 25653 12541 25687
rect 12541 25653 12575 25687
rect 12575 25653 12584 25687
rect 12532 25644 12584 25653
rect 14832 25644 14884 25696
rect 17592 25712 17644 25764
rect 19340 25712 19392 25764
rect 20076 25712 20128 25764
rect 22376 25891 22428 25900
rect 22376 25857 22385 25891
rect 22385 25857 22419 25891
rect 22419 25857 22428 25891
rect 22376 25848 22428 25857
rect 24032 25916 24084 25968
rect 23572 25891 23624 25900
rect 23572 25857 23581 25891
rect 23581 25857 23615 25891
rect 23615 25857 23624 25891
rect 23572 25848 23624 25857
rect 23756 25848 23808 25900
rect 23664 25780 23716 25832
rect 23940 25712 23992 25764
rect 21824 25644 21876 25696
rect 21916 25687 21968 25696
rect 21916 25653 21925 25687
rect 21925 25653 21959 25687
rect 21959 25653 21968 25687
rect 21916 25644 21968 25653
rect 22652 25687 22704 25696
rect 22652 25653 22661 25687
rect 22661 25653 22695 25687
rect 22695 25653 22704 25687
rect 22652 25644 22704 25653
rect 23388 25687 23440 25696
rect 23388 25653 23397 25687
rect 23397 25653 23431 25687
rect 23431 25653 23440 25687
rect 23388 25644 23440 25653
rect 23756 25687 23808 25696
rect 23756 25653 23765 25687
rect 23765 25653 23799 25687
rect 23799 25653 23808 25687
rect 23756 25644 23808 25653
rect 24860 25644 24912 25696
rect 3882 25542 3934 25594
rect 3946 25542 3998 25594
rect 4010 25542 4062 25594
rect 4074 25542 4126 25594
rect 4138 25542 4190 25594
rect 9747 25542 9799 25594
rect 9811 25542 9863 25594
rect 9875 25542 9927 25594
rect 9939 25542 9991 25594
rect 10003 25542 10055 25594
rect 15612 25542 15664 25594
rect 15676 25542 15728 25594
rect 15740 25542 15792 25594
rect 15804 25542 15856 25594
rect 15868 25542 15920 25594
rect 21477 25542 21529 25594
rect 21541 25542 21593 25594
rect 21605 25542 21657 25594
rect 21669 25542 21721 25594
rect 21733 25542 21785 25594
rect 3332 25440 3384 25492
rect 6552 25372 6604 25424
rect 10968 25440 11020 25492
rect 12072 25372 12124 25424
rect 12532 25440 12584 25492
rect 14648 25440 14700 25492
rect 15108 25440 15160 25492
rect 2412 25304 2464 25356
rect 1308 25236 1360 25288
rect 4896 25236 4948 25288
rect 5448 25236 5500 25288
rect 6828 25304 6880 25356
rect 8944 25304 8996 25356
rect 9956 25304 10008 25356
rect 11336 25304 11388 25356
rect 11520 25347 11572 25356
rect 6368 25236 6420 25288
rect 7380 25236 7432 25288
rect 8300 25236 8352 25288
rect 10692 25236 10744 25288
rect 10968 25279 11020 25288
rect 10968 25245 10977 25279
rect 10977 25245 11011 25279
rect 11011 25245 11020 25279
rect 10968 25236 11020 25245
rect 11520 25313 11529 25347
rect 11529 25313 11563 25347
rect 11563 25313 11572 25347
rect 11520 25304 11572 25313
rect 12256 25304 12308 25356
rect 12532 25347 12584 25356
rect 12532 25313 12566 25347
rect 12566 25313 12584 25347
rect 12532 25304 12584 25313
rect 13084 25304 13136 25356
rect 15476 25304 15528 25356
rect 15844 25304 15896 25356
rect 16488 25440 16540 25492
rect 16764 25440 16816 25492
rect 21916 25440 21968 25492
rect 23388 25440 23440 25492
rect 16948 25372 17000 25424
rect 17408 25372 17460 25424
rect 1584 25211 1636 25220
rect 1584 25177 1593 25211
rect 1593 25177 1627 25211
rect 1627 25177 1636 25211
rect 1584 25168 1636 25177
rect 1860 25211 1912 25220
rect 1860 25177 1869 25211
rect 1869 25177 1903 25211
rect 1903 25177 1912 25211
rect 1860 25168 1912 25177
rect 1952 25211 2004 25220
rect 1952 25177 1961 25211
rect 1961 25177 1995 25211
rect 1995 25177 2004 25211
rect 1952 25168 2004 25177
rect 2320 25211 2372 25220
rect 2320 25177 2329 25211
rect 2329 25177 2363 25211
rect 2363 25177 2372 25211
rect 2320 25168 2372 25177
rect 2964 25168 3016 25220
rect 11704 25279 11756 25288
rect 11704 25245 11713 25279
rect 11713 25245 11747 25279
rect 11747 25245 11756 25279
rect 11704 25236 11756 25245
rect 13820 25236 13872 25288
rect 2872 25143 2924 25152
rect 2872 25109 2881 25143
rect 2881 25109 2915 25143
rect 2915 25109 2924 25143
rect 2872 25100 2924 25109
rect 4252 25100 4304 25152
rect 5172 25100 5224 25152
rect 7196 25100 7248 25152
rect 8576 25100 8628 25152
rect 15016 25279 15068 25288
rect 15016 25245 15025 25279
rect 15025 25245 15059 25279
rect 15059 25245 15068 25279
rect 15016 25236 15068 25245
rect 15108 25279 15160 25288
rect 15108 25245 15142 25279
rect 15142 25245 15160 25279
rect 15108 25236 15160 25245
rect 15936 25236 15988 25288
rect 20720 25236 20772 25288
rect 21824 25236 21876 25288
rect 22100 25279 22152 25288
rect 22100 25245 22109 25279
rect 22109 25245 22143 25279
rect 22143 25245 22152 25279
rect 22100 25236 22152 25245
rect 22652 25236 22704 25288
rect 23664 25279 23716 25288
rect 23664 25245 23673 25279
rect 23673 25245 23707 25279
rect 23707 25245 23716 25279
rect 23664 25236 23716 25245
rect 14004 25100 14056 25152
rect 14648 25100 14700 25152
rect 15384 25100 15436 25152
rect 17776 25100 17828 25152
rect 20260 25100 20312 25152
rect 20720 25100 20772 25152
rect 23480 25143 23532 25152
rect 23480 25109 23489 25143
rect 23489 25109 23523 25143
rect 23523 25109 23532 25143
rect 23480 25100 23532 25109
rect 23664 25100 23716 25152
rect 6814 24998 6866 25050
rect 6878 24998 6930 25050
rect 6942 24998 6994 25050
rect 7006 24998 7058 25050
rect 7070 24998 7122 25050
rect 12679 24998 12731 25050
rect 12743 24998 12795 25050
rect 12807 24998 12859 25050
rect 12871 24998 12923 25050
rect 12935 24998 12987 25050
rect 18544 24998 18596 25050
rect 18608 24998 18660 25050
rect 18672 24998 18724 25050
rect 18736 24998 18788 25050
rect 18800 24998 18852 25050
rect 24409 24998 24461 25050
rect 24473 24998 24525 25050
rect 24537 24998 24589 25050
rect 24601 24998 24653 25050
rect 24665 24998 24717 25050
rect 1952 24896 2004 24948
rect 3424 24896 3476 24948
rect 2780 24828 2832 24880
rect 5080 24828 5132 24880
rect 848 24760 900 24812
rect 1584 24760 1636 24812
rect 6184 24896 6236 24948
rect 7104 24896 7156 24948
rect 5356 24828 5408 24880
rect 6552 24871 6604 24880
rect 6552 24837 6561 24871
rect 6561 24837 6595 24871
rect 6595 24837 6604 24871
rect 6552 24828 6604 24837
rect 7196 24828 7248 24880
rect 7472 24896 7524 24948
rect 7656 24939 7708 24948
rect 7656 24905 7665 24939
rect 7665 24905 7699 24939
rect 7699 24905 7708 24939
rect 7656 24896 7708 24905
rect 8668 24896 8720 24948
rect 1216 24692 1268 24744
rect 1584 24667 1636 24676
rect 1584 24633 1593 24667
rect 1593 24633 1627 24667
rect 1627 24633 1636 24667
rect 1584 24624 1636 24633
rect 3792 24735 3844 24744
rect 3792 24701 3801 24735
rect 3801 24701 3835 24735
rect 3835 24701 3844 24735
rect 3792 24692 3844 24701
rect 6736 24760 6788 24812
rect 9128 24828 9180 24880
rect 9588 24828 9640 24880
rect 11428 24828 11480 24880
rect 11888 24828 11940 24880
rect 12256 24828 12308 24880
rect 13452 24828 13504 24880
rect 8668 24760 8720 24812
rect 2044 24556 2096 24608
rect 5908 24692 5960 24744
rect 8760 24692 8812 24744
rect 9956 24760 10008 24812
rect 11612 24692 11664 24744
rect 11980 24692 12032 24744
rect 14280 24896 14332 24948
rect 23480 24896 23532 24948
rect 23572 24896 23624 24948
rect 24032 24939 24084 24948
rect 24032 24905 24041 24939
rect 24041 24905 24075 24939
rect 24075 24905 24084 24939
rect 24032 24896 24084 24905
rect 13820 24828 13872 24880
rect 14648 24803 14700 24812
rect 14648 24769 14682 24803
rect 14682 24769 14700 24803
rect 14648 24760 14700 24769
rect 14832 24803 14884 24812
rect 14832 24769 14841 24803
rect 14841 24769 14875 24803
rect 14875 24769 14884 24803
rect 14832 24760 14884 24769
rect 17408 24803 17460 24812
rect 17408 24769 17442 24803
rect 17442 24769 17460 24803
rect 17408 24760 17460 24769
rect 17960 24760 18012 24812
rect 6276 24624 6328 24676
rect 7840 24667 7892 24676
rect 7840 24633 7849 24667
rect 7849 24633 7883 24667
rect 7883 24633 7892 24667
rect 7840 24624 7892 24633
rect 13912 24692 13964 24744
rect 14556 24735 14608 24744
rect 14556 24701 14565 24735
rect 14565 24701 14599 24735
rect 14599 24701 14608 24735
rect 14556 24692 14608 24701
rect 15016 24692 15068 24744
rect 4804 24599 4856 24608
rect 4804 24565 4813 24599
rect 4813 24565 4847 24599
rect 4847 24565 4856 24599
rect 4804 24556 4856 24565
rect 9036 24599 9088 24608
rect 9036 24565 9045 24599
rect 9045 24565 9079 24599
rect 9079 24565 9088 24599
rect 9036 24556 9088 24565
rect 9312 24556 9364 24608
rect 10508 24556 10560 24608
rect 14188 24556 14240 24608
rect 14924 24556 14976 24608
rect 18328 24692 18380 24744
rect 19156 24803 19208 24812
rect 19156 24769 19165 24803
rect 19165 24769 19199 24803
rect 19199 24769 19208 24803
rect 19156 24760 19208 24769
rect 19524 24760 19576 24812
rect 21180 24760 21232 24812
rect 22652 24735 22704 24744
rect 22652 24701 22661 24735
rect 22661 24701 22695 24735
rect 22695 24701 22704 24735
rect 22652 24692 22704 24701
rect 18788 24556 18840 24608
rect 24216 24624 24268 24676
rect 19248 24599 19300 24608
rect 19248 24565 19257 24599
rect 19257 24565 19291 24599
rect 19291 24565 19300 24599
rect 19248 24556 19300 24565
rect 20168 24599 20220 24608
rect 20168 24565 20177 24599
rect 20177 24565 20211 24599
rect 20211 24565 20220 24599
rect 20168 24556 20220 24565
rect 3882 24454 3934 24506
rect 3946 24454 3998 24506
rect 4010 24454 4062 24506
rect 4074 24454 4126 24506
rect 4138 24454 4190 24506
rect 9747 24454 9799 24506
rect 9811 24454 9863 24506
rect 9875 24454 9927 24506
rect 9939 24454 9991 24506
rect 10003 24454 10055 24506
rect 15612 24454 15664 24506
rect 15676 24454 15728 24506
rect 15740 24454 15792 24506
rect 15804 24454 15856 24506
rect 15868 24454 15920 24506
rect 21477 24454 21529 24506
rect 21541 24454 21593 24506
rect 21605 24454 21657 24506
rect 21669 24454 21721 24506
rect 21733 24454 21785 24506
rect 756 24216 808 24268
rect 3608 24352 3660 24404
rect 2780 24327 2832 24336
rect 2780 24293 2789 24327
rect 2789 24293 2823 24327
rect 2823 24293 2832 24327
rect 2780 24284 2832 24293
rect 2136 24216 2188 24268
rect 4620 24284 4672 24336
rect 4804 24284 4856 24336
rect 5172 24352 5224 24404
rect 6092 24395 6144 24404
rect 6092 24361 6101 24395
rect 6101 24361 6135 24395
rect 6135 24361 6144 24395
rect 6092 24352 6144 24361
rect 9036 24352 9088 24404
rect 10876 24352 10928 24404
rect 12348 24352 12400 24404
rect 7380 24216 7432 24268
rect 1216 24148 1268 24200
rect 1308 24080 1360 24132
rect 4068 24148 4120 24200
rect 5172 24191 5224 24200
rect 5172 24157 5181 24191
rect 5181 24157 5215 24191
rect 5215 24157 5224 24191
rect 5172 24148 5224 24157
rect 5448 24191 5500 24200
rect 5448 24157 5457 24191
rect 5457 24157 5491 24191
rect 5491 24157 5500 24191
rect 5448 24148 5500 24157
rect 9588 24284 9640 24336
rect 9312 24259 9364 24268
rect 9312 24225 9321 24259
rect 9321 24225 9355 24259
rect 9355 24225 9364 24259
rect 9312 24216 9364 24225
rect 9680 24216 9732 24268
rect 9772 24259 9824 24268
rect 9772 24225 9781 24259
rect 9781 24225 9815 24259
rect 9815 24225 9824 24259
rect 9772 24216 9824 24225
rect 10232 24216 10284 24268
rect 9128 24191 9180 24200
rect 9128 24157 9137 24191
rect 9137 24157 9171 24191
rect 9171 24157 9180 24191
rect 9128 24148 9180 24157
rect 10508 24216 10560 24268
rect 10876 24216 10928 24268
rect 11520 24216 11572 24268
rect 12348 24216 12400 24268
rect 12440 24259 12492 24268
rect 12440 24225 12449 24259
rect 12449 24225 12483 24259
rect 12483 24225 12492 24259
rect 12440 24216 12492 24225
rect 13176 24216 13228 24268
rect 11060 24148 11112 24200
rect 11704 24148 11756 24200
rect 12716 24191 12768 24200
rect 12716 24157 12725 24191
rect 12725 24157 12759 24191
rect 12759 24157 12768 24191
rect 12716 24148 12768 24157
rect 6276 24012 6328 24064
rect 6644 24012 6696 24064
rect 7104 24012 7156 24064
rect 7472 24123 7524 24132
rect 7472 24089 7481 24123
rect 7481 24089 7515 24123
rect 7515 24089 7524 24123
rect 7472 24080 7524 24089
rect 7656 24080 7708 24132
rect 18328 24352 18380 24404
rect 19156 24352 19208 24404
rect 20168 24352 20220 24404
rect 21180 24352 21232 24404
rect 23848 24352 23900 24404
rect 17500 24284 17552 24336
rect 14280 24216 14332 24268
rect 14464 24216 14516 24268
rect 17408 24148 17460 24200
rect 8392 24012 8444 24064
rect 8484 24055 8536 24064
rect 8484 24021 8493 24055
rect 8493 24021 8527 24055
rect 8527 24021 8536 24055
rect 8484 24012 8536 24021
rect 14280 24080 14332 24132
rect 17960 24148 18012 24200
rect 19524 24191 19576 24200
rect 19524 24157 19558 24191
rect 19558 24157 19576 24191
rect 19524 24148 19576 24157
rect 13820 24012 13872 24064
rect 14464 24012 14516 24064
rect 20444 24012 20496 24064
rect 22376 24080 22428 24132
rect 23664 24148 23716 24200
rect 24124 24148 24176 24200
rect 21824 24012 21876 24064
rect 23204 24012 23256 24064
rect 24860 24012 24912 24064
rect 6814 23910 6866 23962
rect 6878 23910 6930 23962
rect 6942 23910 6994 23962
rect 7006 23910 7058 23962
rect 7070 23910 7122 23962
rect 12679 23910 12731 23962
rect 12743 23910 12795 23962
rect 12807 23910 12859 23962
rect 12871 23910 12923 23962
rect 12935 23910 12987 23962
rect 18544 23910 18596 23962
rect 18608 23910 18660 23962
rect 18672 23910 18724 23962
rect 18736 23910 18788 23962
rect 18800 23910 18852 23962
rect 24409 23910 24461 23962
rect 24473 23910 24525 23962
rect 24537 23910 24589 23962
rect 24601 23910 24653 23962
rect 24665 23910 24717 23962
rect 2504 23740 2556 23792
rect 2596 23783 2648 23792
rect 2596 23749 2605 23783
rect 2605 23749 2639 23783
rect 2639 23749 2648 23783
rect 2596 23740 2648 23749
rect 3148 23808 3200 23860
rect 756 23672 808 23724
rect 1676 23715 1728 23724
rect 1676 23681 1685 23715
rect 1685 23681 1719 23715
rect 1719 23681 1728 23715
rect 1676 23672 1728 23681
rect 1952 23715 2004 23724
rect 1952 23681 1961 23715
rect 1961 23681 1995 23715
rect 1995 23681 2004 23715
rect 1952 23672 2004 23681
rect 2136 23672 2188 23724
rect 2780 23672 2832 23724
rect 3148 23672 3200 23724
rect 3700 23783 3752 23792
rect 3700 23749 3709 23783
rect 3709 23749 3743 23783
rect 3743 23749 3752 23783
rect 3700 23740 3752 23749
rect 4068 23740 4120 23792
rect 4804 23740 4856 23792
rect 7196 23808 7248 23860
rect 8392 23808 8444 23860
rect 9128 23808 9180 23860
rect 3792 23672 3844 23724
rect 4160 23672 4212 23724
rect 5080 23672 5132 23724
rect 7564 23672 7616 23724
rect 7656 23672 7708 23724
rect 8208 23740 8260 23792
rect 10968 23851 11020 23860
rect 10968 23817 10977 23851
rect 10977 23817 11011 23851
rect 11011 23817 11020 23851
rect 10968 23808 11020 23817
rect 11244 23808 11296 23860
rect 11704 23808 11756 23860
rect 12440 23808 12492 23860
rect 13084 23808 13136 23860
rect 20444 23851 20496 23860
rect 20444 23817 20453 23851
rect 20453 23817 20487 23851
rect 20487 23817 20496 23851
rect 20444 23808 20496 23817
rect 8392 23672 8444 23724
rect 3056 23604 3108 23656
rect 3884 23604 3936 23656
rect 6276 23604 6328 23656
rect 9312 23647 9364 23656
rect 9312 23613 9321 23647
rect 9321 23613 9355 23647
rect 9355 23613 9364 23647
rect 9312 23604 9364 23613
rect 11612 23715 11664 23724
rect 11612 23681 11621 23715
rect 11621 23681 11655 23715
rect 11655 23681 11664 23715
rect 11612 23672 11664 23681
rect 11888 23715 11940 23724
rect 11888 23681 11895 23715
rect 11895 23681 11929 23715
rect 11929 23681 11940 23715
rect 11888 23672 11940 23681
rect 9864 23604 9916 23656
rect 10048 23647 10100 23656
rect 10048 23613 10057 23647
rect 10057 23613 10091 23647
rect 10091 23613 10100 23647
rect 10048 23604 10100 23613
rect 10232 23604 10284 23656
rect 10876 23604 10928 23656
rect 4436 23468 4488 23520
rect 5448 23511 5500 23520
rect 5448 23477 5457 23511
rect 5457 23477 5491 23511
rect 5491 23477 5500 23511
rect 5448 23468 5500 23477
rect 7104 23536 7156 23588
rect 7288 23536 7340 23588
rect 7380 23579 7432 23588
rect 7380 23545 7389 23579
rect 7389 23545 7423 23579
rect 7423 23545 7432 23579
rect 7380 23536 7432 23545
rect 9772 23579 9824 23588
rect 9772 23545 9795 23579
rect 9795 23545 9824 23579
rect 9772 23536 9824 23545
rect 9588 23468 9640 23520
rect 9864 23468 9916 23520
rect 11060 23468 11112 23520
rect 14648 23468 14700 23520
rect 15200 23468 15252 23520
rect 16304 23672 16356 23724
rect 16764 23672 16816 23724
rect 17684 23715 17736 23724
rect 17684 23681 17718 23715
rect 17718 23681 17736 23715
rect 17684 23672 17736 23681
rect 17040 23604 17092 23656
rect 17408 23604 17460 23656
rect 17868 23647 17920 23656
rect 17868 23613 17877 23647
rect 17877 23613 17911 23647
rect 17911 23613 17920 23647
rect 17868 23604 17920 23613
rect 18420 23604 18472 23656
rect 18788 23672 18840 23724
rect 21088 23740 21140 23792
rect 22376 23740 22428 23792
rect 23940 23740 23992 23792
rect 21364 23715 21416 23724
rect 21364 23681 21373 23715
rect 21373 23681 21407 23715
rect 21407 23681 21416 23715
rect 21364 23672 21416 23681
rect 19248 23604 19300 23656
rect 19340 23604 19392 23656
rect 20260 23604 20312 23656
rect 22100 23672 22152 23724
rect 19156 23536 19208 23588
rect 16764 23468 16816 23520
rect 17592 23468 17644 23520
rect 18420 23468 18472 23520
rect 20536 23468 20588 23520
rect 21916 23468 21968 23520
rect 23296 23468 23348 23520
rect 24124 23511 24176 23520
rect 24124 23477 24133 23511
rect 24133 23477 24167 23511
rect 24167 23477 24176 23511
rect 24124 23468 24176 23477
rect 3882 23366 3934 23418
rect 3946 23366 3998 23418
rect 4010 23366 4062 23418
rect 4074 23366 4126 23418
rect 4138 23366 4190 23418
rect 9747 23366 9799 23418
rect 9811 23366 9863 23418
rect 9875 23366 9927 23418
rect 9939 23366 9991 23418
rect 10003 23366 10055 23418
rect 15612 23366 15664 23418
rect 15676 23366 15728 23418
rect 15740 23366 15792 23418
rect 15804 23366 15856 23418
rect 15868 23366 15920 23418
rect 21477 23366 21529 23418
rect 21541 23366 21593 23418
rect 21605 23366 21657 23418
rect 21669 23366 21721 23418
rect 21733 23366 21785 23418
rect 2596 23264 2648 23316
rect 3148 23264 3200 23316
rect 5632 23264 5684 23316
rect 5816 23264 5868 23316
rect 7104 23264 7156 23316
rect 7380 23264 7432 23316
rect 8392 23264 8444 23316
rect 10692 23264 10744 23316
rect 10968 23264 11020 23316
rect 11520 23264 11572 23316
rect 14464 23264 14516 23316
rect 17868 23264 17920 23316
rect 21364 23264 21416 23316
rect 22652 23264 22704 23316
rect 8668 23196 8720 23248
rect 8944 23196 8996 23248
rect 10232 23196 10284 23248
rect 12348 23196 12400 23248
rect 17776 23196 17828 23248
rect 2044 23128 2096 23180
rect 6460 23128 6512 23180
rect 9496 23128 9548 23180
rect 10692 23128 10744 23180
rect 15200 23128 15252 23180
rect 756 22992 808 23044
rect 848 22924 900 22976
rect 2504 23060 2556 23112
rect 2688 23060 2740 23112
rect 3792 23060 3844 23112
rect 12532 23060 12584 23112
rect 13820 23060 13872 23112
rect 14004 23060 14056 23112
rect 2780 22992 2832 23044
rect 7932 22992 7984 23044
rect 9404 22992 9456 23044
rect 10232 22992 10284 23044
rect 3608 22924 3660 22976
rect 6276 22924 6328 22976
rect 6552 22924 6604 22976
rect 7564 22924 7616 22976
rect 7748 22924 7800 22976
rect 11612 22992 11664 23044
rect 14832 23060 14884 23112
rect 10600 22924 10652 22976
rect 12256 22924 12308 22976
rect 12440 22924 12492 22976
rect 14004 22924 14056 22976
rect 15200 22924 15252 22976
rect 19340 23128 19392 23180
rect 16120 22992 16172 23044
rect 16304 22992 16356 23044
rect 20444 23060 20496 23112
rect 18144 22992 18196 23044
rect 21272 23103 21324 23112
rect 21272 23069 21279 23103
rect 21279 23069 21313 23103
rect 21313 23069 21324 23103
rect 21272 23060 21324 23069
rect 22836 23103 22888 23112
rect 22836 23069 22845 23103
rect 22845 23069 22888 23103
rect 22836 23060 22888 23069
rect 23112 22992 23164 23044
rect 16488 22924 16540 22976
rect 22008 22967 22060 22976
rect 22008 22933 22017 22967
rect 22017 22933 22051 22967
rect 22051 22933 22060 22967
rect 22008 22924 22060 22933
rect 23480 22924 23532 22976
rect 24032 23103 24084 23112
rect 24032 23069 24041 23103
rect 24041 23069 24075 23103
rect 24075 23069 24084 23103
rect 24032 23060 24084 23069
rect 6814 22822 6866 22874
rect 6878 22822 6930 22874
rect 6942 22822 6994 22874
rect 7006 22822 7058 22874
rect 7070 22822 7122 22874
rect 12679 22822 12731 22874
rect 12743 22822 12795 22874
rect 12807 22822 12859 22874
rect 12871 22822 12923 22874
rect 12935 22822 12987 22874
rect 18544 22822 18596 22874
rect 18608 22822 18660 22874
rect 18672 22822 18724 22874
rect 18736 22822 18788 22874
rect 18800 22822 18852 22874
rect 24409 22822 24461 22874
rect 24473 22822 24525 22874
rect 24537 22822 24589 22874
rect 24601 22822 24653 22874
rect 24665 22822 24717 22874
rect 3240 22720 3292 22772
rect 3516 22720 3568 22772
rect 5816 22720 5868 22772
rect 1308 22652 1360 22704
rect 1768 22584 1820 22636
rect 1400 22559 1452 22568
rect 1400 22525 1409 22559
rect 1409 22525 1443 22559
rect 1443 22525 1452 22559
rect 1400 22516 1452 22525
rect 3608 22627 3660 22636
rect 3608 22593 3617 22627
rect 3617 22593 3660 22627
rect 3608 22584 3660 22593
rect 4712 22584 4764 22636
rect 6368 22652 6420 22704
rect 7196 22720 7248 22772
rect 8484 22720 8536 22772
rect 10508 22652 10560 22704
rect 10784 22652 10836 22704
rect 11520 22652 11572 22704
rect 12716 22657 12768 22704
rect 5724 22584 5776 22636
rect 6000 22584 6052 22636
rect 6184 22584 6236 22636
rect 6736 22627 6788 22636
rect 6736 22593 6745 22627
rect 6745 22593 6779 22627
rect 6779 22593 6788 22627
rect 6736 22584 6788 22593
rect 7564 22627 7616 22636
rect 7564 22593 7598 22627
rect 7598 22593 7616 22627
rect 7564 22584 7616 22593
rect 4896 22559 4948 22568
rect 4896 22525 4905 22559
rect 4905 22525 4939 22559
rect 4939 22525 4948 22559
rect 4896 22516 4948 22525
rect 5908 22516 5960 22568
rect 6644 22516 6696 22568
rect 2688 22380 2740 22432
rect 2872 22380 2924 22432
rect 3240 22380 3292 22432
rect 4344 22423 4396 22432
rect 4344 22389 4353 22423
rect 4353 22389 4387 22423
rect 4387 22389 4396 22423
rect 4344 22380 4396 22389
rect 5632 22448 5684 22500
rect 7932 22516 7984 22568
rect 7196 22491 7248 22500
rect 7196 22457 7205 22491
rect 7205 22457 7239 22491
rect 7239 22457 7248 22491
rect 7196 22448 7248 22457
rect 8208 22448 8260 22500
rect 11796 22584 11848 22636
rect 12348 22584 12400 22636
rect 12440 22627 12492 22636
rect 12440 22593 12449 22627
rect 12449 22593 12483 22627
rect 12483 22593 12492 22627
rect 12440 22584 12492 22593
rect 12716 22652 12741 22657
rect 12741 22652 12768 22657
rect 14740 22720 14792 22772
rect 14832 22720 14884 22772
rect 15108 22720 15160 22772
rect 16856 22720 16908 22772
rect 17408 22720 17460 22772
rect 20444 22720 20496 22772
rect 22008 22720 22060 22772
rect 23112 22763 23164 22772
rect 23112 22729 23121 22763
rect 23121 22729 23155 22763
rect 23155 22729 23164 22763
rect 23112 22720 23164 22729
rect 23296 22720 23348 22772
rect 24032 22720 24084 22772
rect 13452 22584 13504 22636
rect 9588 22516 9640 22568
rect 13820 22559 13872 22568
rect 13820 22525 13829 22559
rect 13829 22525 13863 22559
rect 13863 22525 13872 22559
rect 13820 22516 13872 22525
rect 13912 22516 13964 22568
rect 14832 22627 14884 22636
rect 14832 22593 14866 22627
rect 14866 22593 14884 22627
rect 14832 22584 14884 22593
rect 17960 22584 18012 22636
rect 19248 22652 19300 22704
rect 18420 22627 18472 22636
rect 18420 22593 18454 22627
rect 18454 22593 18472 22627
rect 18420 22584 18472 22593
rect 15200 22516 15252 22568
rect 10600 22448 10652 22500
rect 11520 22448 11572 22500
rect 12164 22448 12216 22500
rect 14464 22491 14516 22500
rect 14464 22457 14473 22491
rect 14473 22457 14507 22491
rect 14507 22457 14516 22491
rect 14464 22448 14516 22457
rect 20260 22627 20312 22636
rect 20260 22593 20276 22627
rect 20276 22593 20310 22627
rect 20310 22593 20312 22627
rect 20260 22584 20312 22593
rect 21916 22627 21968 22636
rect 21916 22593 21925 22627
rect 21925 22593 21959 22627
rect 21959 22593 21968 22627
rect 21916 22584 21968 22593
rect 23204 22627 23256 22636
rect 23204 22593 23213 22627
rect 23213 22593 23247 22627
rect 23247 22593 23256 22627
rect 23204 22584 23256 22593
rect 23480 22516 23532 22568
rect 22928 22448 22980 22500
rect 23388 22448 23440 22500
rect 8576 22380 8628 22432
rect 8668 22423 8720 22432
rect 8668 22389 8677 22423
rect 8677 22389 8711 22423
rect 8711 22389 8720 22423
rect 8668 22380 8720 22389
rect 9036 22380 9088 22432
rect 10784 22423 10836 22432
rect 10784 22389 10793 22423
rect 10793 22389 10827 22423
rect 10827 22389 10836 22423
rect 10784 22380 10836 22389
rect 10968 22380 11020 22432
rect 14832 22380 14884 22432
rect 17316 22380 17368 22432
rect 20904 22380 20956 22432
rect 23756 22423 23808 22432
rect 23756 22389 23765 22423
rect 23765 22389 23799 22423
rect 23799 22389 23808 22423
rect 23756 22380 23808 22389
rect 24860 22380 24912 22432
rect 3882 22278 3934 22330
rect 3946 22278 3998 22330
rect 4010 22278 4062 22330
rect 4074 22278 4126 22330
rect 4138 22278 4190 22330
rect 9747 22278 9799 22330
rect 9811 22278 9863 22330
rect 9875 22278 9927 22330
rect 9939 22278 9991 22330
rect 10003 22278 10055 22330
rect 15612 22278 15664 22330
rect 15676 22278 15728 22330
rect 15740 22278 15792 22330
rect 15804 22278 15856 22330
rect 15868 22278 15920 22330
rect 21477 22278 21529 22330
rect 21541 22278 21593 22330
rect 21605 22278 21657 22330
rect 21669 22278 21721 22330
rect 21733 22278 21785 22330
rect 24860 22244 24912 22296
rect 25136 22244 25188 22296
rect 3424 22176 3476 22228
rect 3608 22176 3660 22228
rect 4896 22176 4948 22228
rect 5356 22176 5408 22228
rect 7748 22176 7800 22228
rect 1860 22040 1912 22092
rect 2136 22083 2188 22092
rect 2136 22049 2145 22083
rect 2145 22049 2179 22083
rect 2179 22049 2188 22083
rect 2136 22040 2188 22049
rect 6276 22108 6328 22160
rect 7288 22108 7340 22160
rect 11520 22219 11572 22228
rect 11520 22185 11529 22219
rect 11529 22185 11563 22219
rect 11563 22185 11572 22219
rect 11520 22176 11572 22185
rect 14832 22176 14884 22228
rect 21456 22176 21508 22228
rect 2596 22040 2648 22092
rect 2688 22083 2740 22092
rect 2688 22049 2697 22083
rect 2697 22049 2731 22083
rect 2731 22049 2740 22083
rect 2688 22040 2740 22049
rect 296 21904 348 21956
rect 940 21904 992 21956
rect 1492 21836 1544 21888
rect 3608 21972 3660 22024
rect 4436 21904 4488 21956
rect 1952 21836 2004 21888
rect 3332 21879 3384 21888
rect 3332 21845 3341 21879
rect 3341 21845 3375 21879
rect 3375 21845 3384 21879
rect 3332 21836 3384 21845
rect 4160 21836 4212 21888
rect 4988 21972 5040 22024
rect 4896 21904 4948 21956
rect 6184 21972 6236 22024
rect 4988 21879 5040 21888
rect 4988 21845 4997 21879
rect 4997 21845 5031 21879
rect 5031 21845 5040 21879
rect 4988 21836 5040 21845
rect 6000 21836 6052 21888
rect 7196 22040 7248 22092
rect 8760 22108 8812 22160
rect 13268 22151 13320 22160
rect 13268 22117 13277 22151
rect 13277 22117 13311 22151
rect 13311 22117 13320 22151
rect 13268 22108 13320 22117
rect 14464 22108 14516 22160
rect 19156 22108 19208 22160
rect 6552 21972 6604 22024
rect 6644 21972 6696 22024
rect 7748 22015 7800 22024
rect 7748 21981 7757 22015
rect 7757 21981 7791 22015
rect 7791 21981 7800 22015
rect 7748 21972 7800 21981
rect 9312 22040 9364 22092
rect 8024 22015 8076 22024
rect 8024 21981 8033 22015
rect 8033 21981 8067 22015
rect 8067 21981 8076 22015
rect 8024 21972 8076 21981
rect 9404 22015 9456 22024
rect 9404 21981 9413 22015
rect 9413 21981 9447 22015
rect 9447 21981 9456 22015
rect 9404 21972 9456 21981
rect 10784 22040 10836 22092
rect 12440 22040 12492 22092
rect 13084 22040 13136 22092
rect 13452 22040 13504 22092
rect 14188 22040 14240 22092
rect 10324 21904 10376 21956
rect 10600 21947 10652 21956
rect 10600 21913 10609 21947
rect 10609 21913 10643 21947
rect 10643 21913 10652 21947
rect 10600 21904 10652 21913
rect 10968 22015 11020 22024
rect 10968 21981 10977 22015
rect 10977 21981 11011 22015
rect 11011 21981 11020 22015
rect 10968 21972 11020 21981
rect 12256 22015 12308 22024
rect 12256 21981 12265 22015
rect 12265 21981 12299 22015
rect 12299 21981 12308 22015
rect 14832 22040 14884 22092
rect 15108 22083 15160 22092
rect 15108 22049 15142 22083
rect 15142 22049 15160 22083
rect 15108 22040 15160 22049
rect 15292 22083 15344 22092
rect 15292 22049 15301 22083
rect 15301 22049 15335 22083
rect 15335 22049 15344 22083
rect 15292 22040 15344 22049
rect 12256 21972 12308 21981
rect 15016 22015 15068 22024
rect 15016 21981 15025 22015
rect 15025 21981 15059 22015
rect 15059 21981 15068 22015
rect 15016 21972 15068 21981
rect 17040 21972 17092 22024
rect 17316 21972 17368 22024
rect 17868 21972 17920 22024
rect 12348 21947 12400 21956
rect 12348 21913 12357 21947
rect 12357 21913 12391 21947
rect 12391 21913 12400 21947
rect 12348 21904 12400 21913
rect 12532 21904 12584 21956
rect 9588 21879 9640 21888
rect 9588 21845 9597 21879
rect 9597 21845 9631 21879
rect 9631 21845 9640 21879
rect 9588 21836 9640 21845
rect 10416 21836 10468 21888
rect 10692 21836 10744 21888
rect 11428 21836 11480 21888
rect 11796 21836 11848 21888
rect 12072 21836 12124 21888
rect 14188 21904 14240 21956
rect 18512 21972 18564 22024
rect 13176 21836 13228 21888
rect 15016 21836 15068 21888
rect 18328 21879 18380 21888
rect 18328 21845 18337 21879
rect 18337 21845 18371 21879
rect 18371 21845 18380 21879
rect 18328 21836 18380 21845
rect 18972 21879 19024 21888
rect 18972 21845 18981 21879
rect 18981 21845 19015 21879
rect 19015 21845 19024 21879
rect 18972 21836 19024 21845
rect 19156 21836 19208 21888
rect 19340 21836 19392 21888
rect 19616 21836 19668 21888
rect 20812 22015 20864 22024
rect 20812 21981 20821 22015
rect 20821 21981 20855 22015
rect 20855 21981 20864 22015
rect 20812 21972 20864 21981
rect 21180 22015 21232 22024
rect 21180 21981 21189 22015
rect 21189 21981 21223 22015
rect 21223 21981 21232 22015
rect 21180 21972 21232 21981
rect 25504 22040 25556 22092
rect 24860 21972 24912 22024
rect 25136 21972 25188 22024
rect 25596 21972 25648 22024
rect 20720 21879 20772 21888
rect 20720 21845 20729 21879
rect 20729 21845 20763 21879
rect 20763 21845 20772 21879
rect 20720 21836 20772 21845
rect 21364 21879 21416 21888
rect 21364 21845 21373 21879
rect 21373 21845 21407 21879
rect 21407 21845 21416 21879
rect 21364 21836 21416 21845
rect 24860 21836 24912 21888
rect 25596 21836 25648 21888
rect 6814 21734 6866 21786
rect 6878 21734 6930 21786
rect 6942 21734 6994 21786
rect 7006 21734 7058 21786
rect 7070 21734 7122 21786
rect 12679 21734 12731 21786
rect 12743 21734 12795 21786
rect 12807 21734 12859 21786
rect 12871 21734 12923 21786
rect 12935 21734 12987 21786
rect 18544 21734 18596 21786
rect 18608 21734 18660 21786
rect 18672 21734 18724 21786
rect 18736 21734 18788 21786
rect 18800 21734 18852 21786
rect 24409 21734 24461 21786
rect 24473 21734 24525 21786
rect 24537 21734 24589 21786
rect 24601 21734 24653 21786
rect 24665 21734 24717 21786
rect 2136 21632 2188 21684
rect 3792 21632 3844 21684
rect 1124 21564 1176 21616
rect 2044 21496 2096 21548
rect 2412 21496 2464 21548
rect 5540 21564 5592 21616
rect 7932 21632 7984 21684
rect 10416 21632 10468 21684
rect 10600 21632 10652 21684
rect 12072 21632 12124 21684
rect 1400 21471 1452 21480
rect 1400 21437 1409 21471
rect 1409 21437 1443 21471
rect 1443 21437 1452 21471
rect 1400 21428 1452 21437
rect 4988 21539 5040 21548
rect 4988 21505 4997 21539
rect 4997 21505 5031 21539
rect 5031 21505 5040 21539
rect 4988 21496 5040 21505
rect 1308 21292 1360 21344
rect 3240 21428 3292 21480
rect 3976 21471 4028 21480
rect 3976 21437 3985 21471
rect 3985 21437 4019 21471
rect 4019 21437 4028 21471
rect 3976 21428 4028 21437
rect 2136 21360 2188 21412
rect 4436 21403 4488 21412
rect 4436 21369 4445 21403
rect 4445 21369 4479 21403
rect 4479 21369 4488 21403
rect 4436 21360 4488 21369
rect 2964 21335 3016 21344
rect 2964 21301 2973 21335
rect 2973 21301 3007 21335
rect 3007 21301 3016 21335
rect 2964 21292 3016 21301
rect 3700 21292 3752 21344
rect 4160 21292 4212 21344
rect 11704 21564 11756 21616
rect 12348 21632 12400 21684
rect 13912 21632 13964 21684
rect 15384 21632 15436 21684
rect 5448 21360 5500 21412
rect 6184 21496 6236 21548
rect 6552 21496 6604 21548
rect 8024 21496 8076 21548
rect 10968 21496 11020 21548
rect 11520 21496 11572 21548
rect 12072 21539 12124 21548
rect 12072 21505 12081 21539
rect 12081 21505 12115 21539
rect 12115 21505 12124 21539
rect 12072 21496 12124 21505
rect 6000 21428 6052 21480
rect 6276 21360 6328 21412
rect 6736 21360 6788 21412
rect 5172 21292 5224 21344
rect 6552 21292 6604 21344
rect 9680 21428 9732 21480
rect 9404 21292 9456 21344
rect 12164 21292 12216 21344
rect 14464 21496 14516 21548
rect 14648 21496 14700 21548
rect 16856 21632 16908 21684
rect 17684 21632 17736 21684
rect 17960 21632 18012 21684
rect 18420 21632 18472 21684
rect 18972 21632 19024 21684
rect 19156 21632 19208 21684
rect 20720 21632 20772 21684
rect 16028 21564 16080 21616
rect 16488 21428 16540 21480
rect 17316 21496 17368 21548
rect 18052 21471 18104 21480
rect 18052 21437 18061 21471
rect 18061 21437 18095 21471
rect 18095 21437 18104 21471
rect 18052 21428 18104 21437
rect 12900 21360 12952 21412
rect 15200 21292 15252 21344
rect 16212 21335 16264 21344
rect 16212 21301 16221 21335
rect 16221 21301 16255 21335
rect 16255 21301 16264 21335
rect 16212 21292 16264 21301
rect 17960 21360 18012 21412
rect 17684 21335 17736 21344
rect 17684 21301 17693 21335
rect 17693 21301 17727 21335
rect 17727 21301 17736 21335
rect 17684 21292 17736 21301
rect 19340 21496 19392 21548
rect 19616 21539 19668 21548
rect 19616 21505 19625 21539
rect 19625 21505 19659 21539
rect 19659 21505 19668 21539
rect 19616 21496 19668 21505
rect 21456 21496 21508 21548
rect 22008 21496 22060 21548
rect 23848 21539 23900 21548
rect 23848 21505 23857 21539
rect 23857 21505 23891 21539
rect 23891 21505 23900 21539
rect 23848 21496 23900 21505
rect 21916 21428 21968 21480
rect 18880 21360 18932 21412
rect 23204 21360 23256 21412
rect 23388 21360 23440 21412
rect 18420 21292 18472 21344
rect 18512 21292 18564 21344
rect 19524 21292 19576 21344
rect 22744 21292 22796 21344
rect 24032 21292 24084 21344
rect 24124 21335 24176 21344
rect 24124 21301 24133 21335
rect 24133 21301 24167 21335
rect 24167 21301 24176 21335
rect 24124 21292 24176 21301
rect 3882 21190 3934 21242
rect 3946 21190 3998 21242
rect 4010 21190 4062 21242
rect 4074 21190 4126 21242
rect 4138 21190 4190 21242
rect 9747 21190 9799 21242
rect 9811 21190 9863 21242
rect 9875 21190 9927 21242
rect 9939 21190 9991 21242
rect 10003 21190 10055 21242
rect 15612 21190 15664 21242
rect 15676 21190 15728 21242
rect 15740 21190 15792 21242
rect 15804 21190 15856 21242
rect 15868 21190 15920 21242
rect 21477 21190 21529 21242
rect 21541 21190 21593 21242
rect 21605 21190 21657 21242
rect 21669 21190 21721 21242
rect 21733 21190 21785 21242
rect 4252 21088 4304 21140
rect 3700 21020 3752 21072
rect 5448 21088 5500 21140
rect 5540 21088 5592 21140
rect 5816 21088 5868 21140
rect 940 20952 992 21004
rect 756 20884 808 20936
rect 2688 20952 2740 21004
rect 4344 20952 4396 21004
rect 2136 20884 2188 20936
rect 2320 20884 2372 20936
rect 2964 20927 3016 20936
rect 2964 20893 2973 20927
rect 2973 20893 3007 20927
rect 3007 20893 3016 20927
rect 2964 20884 3016 20893
rect 940 20816 992 20868
rect 2596 20859 2648 20868
rect 2596 20825 2605 20859
rect 2605 20825 2639 20859
rect 2639 20825 2648 20859
rect 2596 20816 2648 20825
rect 3332 20859 3384 20868
rect 3332 20825 3341 20859
rect 3341 20825 3375 20859
rect 3375 20825 3384 20859
rect 3332 20816 3384 20825
rect 5724 21063 5776 21072
rect 5724 21029 5733 21063
rect 5733 21029 5767 21063
rect 5767 21029 5776 21063
rect 5724 21020 5776 21029
rect 5448 20952 5500 21004
rect 9588 21088 9640 21140
rect 10140 21088 10192 21140
rect 10784 21088 10836 21140
rect 11520 21088 11572 21140
rect 12440 21131 12492 21140
rect 12440 21097 12449 21131
rect 12449 21097 12483 21131
rect 12483 21097 12492 21131
rect 12440 21088 12492 21097
rect 16212 21088 16264 21140
rect 17684 21088 17736 21140
rect 17868 21088 17920 21140
rect 18328 21088 18380 21140
rect 19156 21088 19208 21140
rect 23848 21088 23900 21140
rect 6184 20884 6236 20936
rect 6920 20884 6972 20936
rect 7840 20884 7892 20936
rect 8208 20884 8260 20936
rect 8668 20884 8720 20936
rect 9404 20927 9456 20936
rect 9404 20893 9413 20927
rect 9413 20893 9447 20927
rect 9447 20893 9456 20927
rect 9404 20884 9456 20893
rect 12164 21020 12216 21072
rect 12900 21020 12952 21072
rect 14188 20952 14240 21004
rect 17040 20995 17092 21004
rect 17040 20961 17049 20995
rect 17049 20961 17083 20995
rect 17083 20961 17092 20995
rect 17040 20952 17092 20961
rect 11244 20884 11296 20936
rect 12532 20884 12584 20936
rect 17224 20884 17276 20936
rect 19340 20884 19392 20936
rect 22192 20927 22244 20936
rect 22192 20893 22201 20927
rect 22201 20893 22235 20927
rect 22235 20893 22244 20927
rect 22192 20884 22244 20893
rect 25136 20884 25188 20936
rect 1584 20791 1636 20800
rect 1584 20757 1593 20791
rect 1593 20757 1627 20791
rect 1627 20757 1636 20791
rect 1584 20748 1636 20757
rect 1860 20748 1912 20800
rect 2136 20748 2188 20800
rect 3424 20748 3476 20800
rect 10968 20816 11020 20868
rect 6092 20748 6144 20800
rect 6552 20748 6604 20800
rect 12440 20816 12492 20868
rect 13176 20816 13228 20868
rect 16028 20816 16080 20868
rect 16212 20816 16264 20868
rect 17316 20748 17368 20800
rect 19892 20816 19944 20868
rect 20352 20859 20404 20868
rect 20352 20825 20364 20859
rect 20364 20825 20404 20859
rect 20352 20816 20404 20825
rect 20720 20816 20772 20868
rect 21916 20816 21968 20868
rect 22008 20816 22060 20868
rect 24860 20816 24912 20868
rect 17960 20791 18012 20800
rect 17960 20757 17969 20791
rect 17969 20757 18003 20791
rect 18003 20757 18012 20791
rect 17960 20748 18012 20757
rect 18880 20748 18932 20800
rect 19616 20748 19668 20800
rect 21456 20791 21508 20800
rect 21456 20757 21465 20791
rect 21465 20757 21499 20791
rect 21499 20757 21508 20791
rect 21456 20748 21508 20757
rect 6814 20646 6866 20698
rect 6878 20646 6930 20698
rect 6942 20646 6994 20698
rect 7006 20646 7058 20698
rect 7070 20646 7122 20698
rect 12679 20646 12731 20698
rect 12743 20646 12795 20698
rect 12807 20646 12859 20698
rect 12871 20646 12923 20698
rect 12935 20646 12987 20698
rect 18544 20646 18596 20698
rect 18608 20646 18660 20698
rect 18672 20646 18724 20698
rect 18736 20646 18788 20698
rect 18800 20646 18852 20698
rect 24409 20646 24461 20698
rect 24473 20646 24525 20698
rect 24537 20646 24589 20698
rect 24601 20646 24653 20698
rect 24665 20646 24717 20698
rect 664 20544 716 20596
rect 1584 20587 1636 20596
rect 1584 20553 1593 20587
rect 1593 20553 1627 20587
rect 1627 20553 1636 20587
rect 1584 20544 1636 20553
rect 2044 20544 2096 20596
rect 2228 20544 2280 20596
rect 2596 20544 2648 20596
rect 940 20476 992 20528
rect 1492 20451 1544 20460
rect 1492 20417 1501 20451
rect 1501 20417 1535 20451
rect 1535 20417 1544 20451
rect 1492 20408 1544 20417
rect 1124 20340 1176 20392
rect 2504 20408 2556 20460
rect 3516 20476 3568 20528
rect 3700 20408 3752 20460
rect 5816 20544 5868 20596
rect 6368 20544 6420 20596
rect 6736 20544 6788 20596
rect 4804 20476 4856 20528
rect 8300 20544 8352 20596
rect 14372 20544 14424 20596
rect 20352 20544 20404 20596
rect 4344 20451 4396 20460
rect 4344 20417 4353 20451
rect 4353 20417 4387 20451
rect 4387 20417 4396 20451
rect 4344 20408 4396 20417
rect 5540 20408 5592 20460
rect 6644 20408 6696 20460
rect 1308 20204 1360 20256
rect 7196 20340 7248 20392
rect 8668 20476 8720 20528
rect 10232 20476 10284 20528
rect 11152 20476 11204 20528
rect 12256 20476 12308 20528
rect 13912 20476 13964 20528
rect 21456 20544 21508 20596
rect 7748 20408 7800 20460
rect 12348 20451 12400 20460
rect 12348 20417 12357 20451
rect 12357 20417 12391 20451
rect 12391 20417 12400 20451
rect 12348 20408 12400 20417
rect 13176 20408 13228 20460
rect 13360 20451 13412 20460
rect 13360 20417 13369 20451
rect 13369 20417 13403 20451
rect 13403 20417 13412 20451
rect 13360 20408 13412 20417
rect 13820 20408 13872 20460
rect 14464 20451 14516 20460
rect 14464 20417 14473 20451
rect 14473 20417 14507 20451
rect 14507 20417 14516 20451
rect 14464 20408 14516 20417
rect 15108 20408 15160 20460
rect 18880 20408 18932 20460
rect 20352 20451 20404 20460
rect 20352 20417 20361 20451
rect 20361 20417 20395 20451
rect 20395 20417 20404 20451
rect 20352 20408 20404 20417
rect 22100 20451 22152 20460
rect 22100 20417 22109 20451
rect 22109 20417 22143 20451
rect 22143 20417 22152 20451
rect 22100 20408 22152 20417
rect 8300 20340 8352 20392
rect 11520 20340 11572 20392
rect 13452 20340 13504 20392
rect 14280 20340 14332 20392
rect 14464 20272 14516 20324
rect 15200 20340 15252 20392
rect 20260 20272 20312 20324
rect 20720 20272 20772 20324
rect 22376 20272 22428 20324
rect 22560 20272 22612 20324
rect 8300 20204 8352 20256
rect 8576 20247 8628 20256
rect 8576 20213 8585 20247
rect 8585 20213 8619 20247
rect 8619 20213 8628 20247
rect 8576 20204 8628 20213
rect 11152 20204 11204 20256
rect 12532 20247 12584 20256
rect 12532 20213 12541 20247
rect 12541 20213 12575 20247
rect 12575 20213 12584 20247
rect 12532 20204 12584 20213
rect 14280 20247 14332 20256
rect 14280 20213 14289 20247
rect 14289 20213 14323 20247
rect 14323 20213 14332 20247
rect 14280 20204 14332 20213
rect 15384 20204 15436 20256
rect 16028 20247 16080 20256
rect 16028 20213 16037 20247
rect 16037 20213 16071 20247
rect 16071 20213 16080 20247
rect 16028 20204 16080 20213
rect 19800 20247 19852 20256
rect 19800 20213 19809 20247
rect 19809 20213 19843 20247
rect 19843 20213 19852 20247
rect 19800 20204 19852 20213
rect 20168 20247 20220 20256
rect 20168 20213 20177 20247
rect 20177 20213 20211 20247
rect 20211 20213 20220 20247
rect 20168 20204 20220 20213
rect 21364 20204 21416 20256
rect 22284 20204 22336 20256
rect 23848 20247 23900 20256
rect 23848 20213 23857 20247
rect 23857 20213 23891 20247
rect 23891 20213 23900 20247
rect 23848 20204 23900 20213
rect 3882 20102 3934 20154
rect 3946 20102 3998 20154
rect 4010 20102 4062 20154
rect 4074 20102 4126 20154
rect 4138 20102 4190 20154
rect 9747 20102 9799 20154
rect 9811 20102 9863 20154
rect 9875 20102 9927 20154
rect 9939 20102 9991 20154
rect 10003 20102 10055 20154
rect 15612 20102 15664 20154
rect 15676 20102 15728 20154
rect 15740 20102 15792 20154
rect 15804 20102 15856 20154
rect 15868 20102 15920 20154
rect 21477 20102 21529 20154
rect 21541 20102 21593 20154
rect 21605 20102 21657 20154
rect 21669 20102 21721 20154
rect 21733 20102 21785 20154
rect 1216 20000 1268 20052
rect 1676 19975 1728 19984
rect 1676 19941 1685 19975
rect 1685 19941 1719 19975
rect 1719 19941 1728 19975
rect 1676 19932 1728 19941
rect 2412 20000 2464 20052
rect 2688 20000 2740 20052
rect 3056 20000 3108 20052
rect 4068 20000 4120 20052
rect 3240 19932 3292 19984
rect 756 19796 808 19848
rect 2688 19864 2740 19916
rect 2136 19796 2188 19848
rect 1308 19728 1360 19780
rect 4896 19864 4948 19916
rect 5356 19864 5408 19916
rect 2228 19660 2280 19712
rect 5356 19728 5408 19780
rect 8576 20000 8628 20052
rect 8760 20000 8812 20052
rect 8944 20000 8996 20052
rect 12256 20000 12308 20052
rect 7932 19864 7984 19916
rect 5908 19728 5960 19780
rect 6460 19728 6512 19780
rect 6828 19703 6880 19712
rect 6828 19669 6837 19703
rect 6837 19669 6871 19703
rect 6871 19669 6880 19703
rect 6828 19660 6880 19669
rect 7380 19771 7432 19780
rect 7380 19737 7389 19771
rect 7389 19737 7423 19771
rect 7423 19737 7432 19771
rect 7380 19728 7432 19737
rect 7656 19839 7708 19848
rect 7656 19805 7665 19839
rect 7665 19805 7699 19839
rect 7699 19805 7708 19839
rect 7656 19796 7708 19805
rect 13360 20000 13412 20052
rect 13820 20000 13872 20052
rect 12072 19864 12124 19916
rect 18880 20043 18932 20052
rect 18880 20009 18889 20043
rect 18889 20009 18923 20043
rect 18923 20009 18932 20043
rect 18880 20000 18932 20009
rect 15384 19932 15436 19984
rect 19984 20000 20036 20052
rect 20260 20000 20312 20052
rect 20352 20000 20404 20052
rect 22100 20000 22152 20052
rect 22284 20000 22336 20052
rect 23756 20043 23808 20052
rect 23756 20009 23765 20043
rect 23765 20009 23799 20043
rect 23799 20009 23808 20043
rect 23756 20000 23808 20009
rect 24032 20043 24084 20052
rect 24032 20009 24041 20043
rect 24041 20009 24075 20043
rect 24075 20009 24084 20043
rect 24032 20000 24084 20009
rect 16028 19864 16080 19916
rect 9312 19839 9364 19848
rect 9312 19805 9321 19839
rect 9321 19805 9355 19839
rect 9355 19805 9364 19839
rect 9312 19796 9364 19805
rect 9588 19839 9640 19848
rect 9588 19805 9613 19839
rect 9613 19805 9640 19839
rect 9588 19796 9640 19805
rect 11152 19839 11204 19848
rect 11152 19805 11161 19839
rect 11161 19805 11195 19839
rect 11195 19805 11204 19839
rect 11152 19796 11204 19805
rect 11612 19839 11664 19848
rect 11612 19805 11621 19839
rect 11621 19805 11655 19839
rect 11655 19805 11664 19839
rect 11612 19796 11664 19805
rect 7840 19728 7892 19780
rect 8116 19771 8168 19780
rect 8116 19737 8125 19771
rect 8125 19737 8159 19771
rect 8159 19737 8168 19771
rect 8116 19728 8168 19737
rect 8300 19728 8352 19780
rect 10140 19728 10192 19780
rect 9588 19660 9640 19712
rect 10508 19660 10560 19712
rect 11244 19771 11296 19780
rect 11244 19737 11253 19771
rect 11253 19737 11287 19771
rect 11287 19737 11296 19771
rect 11244 19728 11296 19737
rect 12256 19728 12308 19780
rect 15660 19839 15712 19848
rect 15660 19805 15694 19839
rect 15694 19805 15712 19839
rect 15660 19796 15712 19805
rect 15844 19839 15896 19848
rect 15844 19805 15853 19839
rect 15853 19805 15887 19839
rect 15887 19805 15896 19839
rect 15844 19796 15896 19805
rect 19248 19907 19300 19916
rect 19248 19873 19257 19907
rect 19257 19873 19291 19907
rect 19291 19873 19300 19907
rect 19248 19864 19300 19873
rect 18880 19796 18932 19848
rect 19064 19839 19116 19848
rect 19064 19805 19073 19839
rect 19073 19805 19107 19839
rect 19107 19805 19116 19839
rect 19064 19796 19116 19805
rect 20628 19864 20680 19916
rect 21364 19796 21416 19848
rect 23848 19864 23900 19916
rect 23388 19796 23440 19848
rect 23572 19728 23624 19780
rect 22100 19660 22152 19712
rect 22652 19660 22704 19712
rect 24216 19703 24268 19712
rect 24216 19669 24225 19703
rect 24225 19669 24259 19703
rect 24259 19669 24268 19703
rect 24216 19660 24268 19669
rect 6814 19558 6866 19610
rect 6878 19558 6930 19610
rect 6942 19558 6994 19610
rect 7006 19558 7058 19610
rect 7070 19558 7122 19610
rect 12679 19558 12731 19610
rect 12743 19558 12795 19610
rect 12807 19558 12859 19610
rect 12871 19558 12923 19610
rect 12935 19558 12987 19610
rect 18544 19558 18596 19610
rect 18608 19558 18660 19610
rect 18672 19558 18724 19610
rect 18736 19558 18788 19610
rect 18800 19558 18852 19610
rect 24409 19558 24461 19610
rect 24473 19558 24525 19610
rect 24537 19558 24589 19610
rect 24601 19558 24653 19610
rect 24665 19558 24717 19610
rect 664 19456 716 19508
rect 1860 19388 1912 19440
rect 2136 19388 2188 19440
rect 2228 19388 2280 19440
rect 2780 19363 2832 19372
rect 2780 19329 2789 19363
rect 2789 19329 2823 19363
rect 2823 19329 2832 19363
rect 2780 19320 2832 19329
rect 3240 19388 3292 19440
rect 7656 19456 7708 19508
rect 7840 19456 7892 19508
rect 7932 19499 7984 19508
rect 7932 19465 7941 19499
rect 7941 19465 7975 19499
rect 7975 19465 7984 19499
rect 7932 19456 7984 19465
rect 4528 19388 4580 19440
rect 3056 19252 3108 19304
rect 1492 19116 1544 19168
rect 2412 19159 2464 19168
rect 2412 19125 2421 19159
rect 2421 19125 2455 19159
rect 2455 19125 2464 19159
rect 2412 19116 2464 19125
rect 4252 19159 4304 19168
rect 4252 19125 4261 19159
rect 4261 19125 4295 19159
rect 4295 19125 4304 19159
rect 4252 19116 4304 19125
rect 4896 19363 4948 19372
rect 4896 19329 4905 19363
rect 4905 19329 4939 19363
rect 4939 19329 4948 19363
rect 4896 19320 4948 19329
rect 5080 19320 5132 19372
rect 5632 19320 5684 19372
rect 6644 19320 6696 19372
rect 6920 19363 6972 19372
rect 6920 19329 6929 19363
rect 6929 19329 6963 19363
rect 6963 19329 6972 19363
rect 6920 19320 6972 19329
rect 7472 19388 7524 19440
rect 9312 19388 9364 19440
rect 9496 19388 9548 19440
rect 9588 19388 9640 19440
rect 12072 19320 12124 19372
rect 13176 19388 13228 19440
rect 13452 19499 13504 19508
rect 13452 19465 13461 19499
rect 13461 19465 13495 19499
rect 13495 19465 13504 19499
rect 13452 19456 13504 19465
rect 15844 19456 15896 19508
rect 16672 19456 16724 19508
rect 16856 19456 16908 19508
rect 18144 19456 18196 19508
rect 13452 19320 13504 19372
rect 9404 19252 9456 19304
rect 15660 19320 15712 19372
rect 16396 19320 16448 19372
rect 16212 19252 16264 19304
rect 18880 19456 18932 19508
rect 20628 19456 20680 19508
rect 22652 19456 22704 19508
rect 5632 19184 5684 19236
rect 6368 19184 6420 19236
rect 6552 19184 6604 19236
rect 6736 19184 6788 19236
rect 7932 19184 7984 19236
rect 5908 19159 5960 19168
rect 5908 19125 5917 19159
rect 5917 19125 5951 19159
rect 5951 19125 5960 19159
rect 5908 19116 5960 19125
rect 6092 19116 6144 19168
rect 9680 19159 9732 19168
rect 9680 19125 9689 19159
rect 9689 19125 9723 19159
rect 9723 19125 9732 19159
rect 9680 19116 9732 19125
rect 10968 19116 11020 19168
rect 12440 19116 12492 19168
rect 14280 19184 14332 19236
rect 16488 19184 16540 19236
rect 17040 19252 17092 19304
rect 19524 19320 19576 19372
rect 17684 19295 17736 19304
rect 17684 19261 17718 19295
rect 17718 19261 17736 19295
rect 17684 19252 17736 19261
rect 17868 19295 17920 19304
rect 17868 19261 17877 19295
rect 17877 19261 17911 19295
rect 17911 19261 17920 19295
rect 17868 19252 17920 19261
rect 18604 19295 18656 19304
rect 18604 19261 18613 19295
rect 18613 19261 18647 19295
rect 18647 19261 18656 19295
rect 18604 19252 18656 19261
rect 19892 19320 19944 19372
rect 20352 19320 20404 19372
rect 21272 19320 21324 19372
rect 22192 19388 22244 19440
rect 22100 19363 22152 19372
rect 22100 19329 22134 19363
rect 22134 19329 22152 19363
rect 22100 19320 22152 19329
rect 22376 19320 22428 19372
rect 23572 19456 23624 19508
rect 17316 19227 17368 19236
rect 17316 19193 17325 19227
rect 17325 19193 17359 19227
rect 17359 19193 17368 19227
rect 17316 19184 17368 19193
rect 14372 19116 14424 19168
rect 18512 19159 18564 19168
rect 18512 19125 18521 19159
rect 18521 19125 18555 19159
rect 18555 19125 18564 19159
rect 18512 19116 18564 19125
rect 19524 19116 19576 19168
rect 22836 19252 22888 19304
rect 23112 19252 23164 19304
rect 20076 19116 20128 19168
rect 20996 19159 21048 19168
rect 20996 19125 21005 19159
rect 21005 19125 21039 19159
rect 21039 19125 21048 19159
rect 20996 19116 21048 19125
rect 22836 19116 22888 19168
rect 23940 19159 23992 19168
rect 23940 19125 23949 19159
rect 23949 19125 23983 19159
rect 23983 19125 23992 19159
rect 23940 19116 23992 19125
rect 3882 19014 3934 19066
rect 3946 19014 3998 19066
rect 4010 19014 4062 19066
rect 4074 19014 4126 19066
rect 4138 19014 4190 19066
rect 9747 19014 9799 19066
rect 9811 19014 9863 19066
rect 9875 19014 9927 19066
rect 9939 19014 9991 19066
rect 10003 19014 10055 19066
rect 15612 19014 15664 19066
rect 15676 19014 15728 19066
rect 15740 19014 15792 19066
rect 15804 19014 15856 19066
rect 15868 19014 15920 19066
rect 21477 19014 21529 19066
rect 21541 19014 21593 19066
rect 21605 19014 21657 19066
rect 21669 19014 21721 19066
rect 21733 19014 21785 19066
rect 4804 18912 4856 18964
rect 6368 18912 6420 18964
rect 7288 18912 7340 18964
rect 8760 18912 8812 18964
rect 11244 18912 11296 18964
rect 12440 18912 12492 18964
rect 2412 18844 2464 18896
rect 5908 18844 5960 18896
rect 480 18776 532 18828
rect 3056 18776 3108 18828
rect 3608 18776 3660 18828
rect 5264 18776 5316 18828
rect 6092 18776 6144 18828
rect 1400 18751 1452 18760
rect 1400 18717 1409 18751
rect 1409 18717 1443 18751
rect 1443 18717 1452 18751
rect 1400 18708 1452 18717
rect 1584 18708 1636 18760
rect 2596 18751 2648 18760
rect 2596 18717 2605 18751
rect 2605 18717 2639 18751
rect 2639 18717 2648 18751
rect 2596 18708 2648 18717
rect 2872 18751 2924 18760
rect 2872 18717 2881 18751
rect 2881 18717 2915 18751
rect 2915 18717 2924 18751
rect 2872 18708 2924 18717
rect 4528 18708 4580 18760
rect 5448 18708 5500 18760
rect 6368 18819 6420 18828
rect 6368 18785 6402 18819
rect 6402 18785 6420 18819
rect 6368 18776 6420 18785
rect 6552 18819 6604 18828
rect 6552 18785 6561 18819
rect 6561 18785 6595 18819
rect 6595 18785 6604 18819
rect 6552 18776 6604 18785
rect 7564 18708 7616 18760
rect 8576 18708 8628 18760
rect 3608 18640 3660 18692
rect 9680 18776 9732 18828
rect 9404 18751 9456 18760
rect 9404 18717 9413 18751
rect 9413 18717 9447 18751
rect 9447 18717 9456 18751
rect 9404 18708 9456 18717
rect 9496 18751 9548 18760
rect 9496 18717 9505 18751
rect 9505 18717 9539 18751
rect 9539 18717 9548 18751
rect 9496 18708 9548 18717
rect 9956 18708 10008 18760
rect 10508 18708 10560 18760
rect 11244 18708 11296 18760
rect 12256 18708 12308 18760
rect 10232 18683 10284 18692
rect 10232 18649 10241 18683
rect 10241 18649 10275 18683
rect 10275 18649 10284 18683
rect 10232 18640 10284 18649
rect 3424 18572 3476 18624
rect 3516 18615 3568 18624
rect 3516 18581 3525 18615
rect 3525 18581 3559 18615
rect 3559 18581 3568 18615
rect 3516 18572 3568 18581
rect 4804 18615 4856 18624
rect 4804 18581 4813 18615
rect 4813 18581 4847 18615
rect 4847 18581 4856 18615
rect 4804 18572 4856 18581
rect 5356 18572 5408 18624
rect 5540 18572 5592 18624
rect 7288 18572 7340 18624
rect 8300 18572 8352 18624
rect 13360 18640 13412 18692
rect 16948 18844 17000 18896
rect 17684 18844 17736 18896
rect 18052 18776 18104 18828
rect 18144 18708 18196 18760
rect 18512 18776 18564 18828
rect 19800 18912 19852 18964
rect 22744 18912 22796 18964
rect 23388 18912 23440 18964
rect 18420 18708 18472 18760
rect 11980 18572 12032 18624
rect 13820 18572 13872 18624
rect 13912 18572 13964 18624
rect 15200 18572 15252 18624
rect 17684 18640 17736 18692
rect 19524 18751 19576 18760
rect 19524 18717 19533 18751
rect 19533 18717 19567 18751
rect 19567 18717 19576 18751
rect 19524 18708 19576 18717
rect 20168 18844 20220 18896
rect 22284 18708 22336 18760
rect 22376 18751 22428 18760
rect 22376 18717 22385 18751
rect 22385 18717 22419 18751
rect 22419 18717 22428 18751
rect 22376 18708 22428 18717
rect 22744 18751 22796 18760
rect 22744 18717 22753 18751
rect 22753 18717 22796 18751
rect 22744 18708 22796 18717
rect 20996 18640 21048 18692
rect 22560 18640 22612 18692
rect 18328 18572 18380 18624
rect 19248 18572 19300 18624
rect 20444 18615 20496 18624
rect 20444 18581 20453 18615
rect 20453 18581 20487 18615
rect 20487 18581 20496 18615
rect 20444 18572 20496 18581
rect 22192 18615 22244 18624
rect 22192 18581 22201 18615
rect 22201 18581 22235 18615
rect 22235 18581 22244 18615
rect 22192 18572 22244 18581
rect 22652 18572 22704 18624
rect 23940 18751 23992 18760
rect 23940 18717 23949 18751
rect 23949 18717 23983 18751
rect 23983 18717 23992 18751
rect 23940 18708 23992 18717
rect 23848 18572 23900 18624
rect 940 18436 992 18488
rect 6814 18470 6866 18522
rect 6878 18470 6930 18522
rect 6942 18470 6994 18522
rect 7006 18470 7058 18522
rect 7070 18470 7122 18522
rect 12679 18470 12731 18522
rect 12743 18470 12795 18522
rect 12807 18470 12859 18522
rect 12871 18470 12923 18522
rect 12935 18470 12987 18522
rect 18544 18470 18596 18522
rect 18608 18470 18660 18522
rect 18672 18470 18724 18522
rect 18736 18470 18788 18522
rect 18800 18470 18852 18522
rect 24409 18470 24461 18522
rect 24473 18470 24525 18522
rect 24537 18470 24589 18522
rect 24601 18470 24653 18522
rect 24665 18470 24717 18522
rect 2872 18368 2924 18420
rect 3424 18368 3476 18420
rect 756 18232 808 18284
rect 1584 18232 1636 18284
rect 1860 18232 1912 18284
rect 5448 18368 5500 18420
rect 6092 18368 6144 18420
rect 6552 18368 6604 18420
rect 7564 18368 7616 18420
rect 9036 18368 9088 18420
rect 9680 18368 9732 18420
rect 10968 18368 11020 18420
rect 16120 18368 16172 18420
rect 5356 18300 5408 18352
rect 1492 18164 1544 18216
rect 1400 18028 1452 18080
rect 3332 18096 3384 18148
rect 4804 18275 4856 18284
rect 4804 18241 4813 18275
rect 4813 18241 4847 18275
rect 4847 18241 4856 18275
rect 4804 18232 4856 18241
rect 5724 18232 5776 18284
rect 6368 18232 6420 18284
rect 6460 18232 6512 18284
rect 7196 18232 7248 18284
rect 4252 18207 4304 18216
rect 4252 18173 4261 18207
rect 4261 18173 4295 18207
rect 4295 18173 4304 18207
rect 4252 18164 4304 18173
rect 4344 18164 4396 18216
rect 3240 18071 3292 18080
rect 3240 18037 3249 18071
rect 3249 18037 3283 18071
rect 3283 18037 3292 18071
rect 3240 18028 3292 18037
rect 3608 18028 3660 18080
rect 4252 18028 4304 18080
rect 5264 18096 5316 18148
rect 7748 18096 7800 18148
rect 5448 18071 5500 18080
rect 5448 18037 5457 18071
rect 5457 18037 5491 18071
rect 5491 18037 5500 18071
rect 5448 18028 5500 18037
rect 5632 18028 5684 18080
rect 5908 18028 5960 18080
rect 7932 18232 7984 18284
rect 9588 18232 9640 18284
rect 11704 18300 11756 18352
rect 10600 18232 10652 18284
rect 11520 18232 11572 18284
rect 13452 18300 13504 18352
rect 11980 18275 12032 18284
rect 11980 18241 11989 18275
rect 11989 18241 12023 18275
rect 12023 18241 12032 18275
rect 11980 18232 12032 18241
rect 16580 18300 16632 18352
rect 17408 18368 17460 18420
rect 17684 18368 17736 18420
rect 18420 18368 18472 18420
rect 22192 18368 22244 18420
rect 22560 18368 22612 18420
rect 23940 18368 23992 18420
rect 25136 18368 25188 18420
rect 14372 18275 14424 18284
rect 14372 18241 14406 18275
rect 14406 18241 14424 18275
rect 14372 18232 14424 18241
rect 14556 18275 14608 18284
rect 14556 18241 14565 18275
rect 14565 18241 14599 18275
rect 14599 18241 14608 18275
rect 14556 18232 14608 18241
rect 16120 18232 16172 18284
rect 16304 18232 16356 18284
rect 20812 18300 20864 18352
rect 17868 18275 17920 18284
rect 17868 18241 17877 18275
rect 17877 18241 17911 18275
rect 17911 18241 17920 18275
rect 17868 18232 17920 18241
rect 22652 18275 22704 18284
rect 22652 18241 22661 18275
rect 22661 18241 22695 18275
rect 22695 18241 22704 18275
rect 22652 18232 22704 18241
rect 22836 18275 22888 18284
rect 22836 18241 22845 18275
rect 22845 18241 22879 18275
rect 22879 18241 22888 18275
rect 22836 18232 22888 18241
rect 9312 18164 9364 18216
rect 11704 18164 11756 18216
rect 11888 18164 11940 18216
rect 11888 18071 11940 18080
rect 11888 18037 11897 18071
rect 11897 18037 11931 18071
rect 11931 18037 11940 18071
rect 11888 18028 11940 18037
rect 13452 18164 13504 18216
rect 17316 18207 17368 18216
rect 17316 18173 17325 18207
rect 17325 18173 17359 18207
rect 17359 18173 17368 18207
rect 17316 18164 17368 18173
rect 17408 18164 17460 18216
rect 17684 18207 17736 18216
rect 17684 18173 17718 18207
rect 17718 18173 17736 18207
rect 17684 18164 17736 18173
rect 20720 18164 20772 18216
rect 17224 18096 17276 18148
rect 21824 18096 21876 18148
rect 23388 18232 23440 18284
rect 15200 18071 15252 18080
rect 15200 18037 15209 18071
rect 15209 18037 15243 18071
rect 15243 18037 15252 18071
rect 15200 18028 15252 18037
rect 18052 18028 18104 18080
rect 20168 18028 20220 18080
rect 22100 18028 22152 18080
rect 23572 18071 23624 18080
rect 23572 18037 23581 18071
rect 23581 18037 23615 18071
rect 23615 18037 23624 18071
rect 23572 18028 23624 18037
rect 24860 18028 24912 18080
rect 756 17960 808 18012
rect 940 17960 992 18012
rect 3882 17926 3934 17978
rect 3946 17926 3998 17978
rect 4010 17926 4062 17978
rect 4074 17926 4126 17978
rect 4138 17926 4190 17978
rect 9747 17926 9799 17978
rect 9811 17926 9863 17978
rect 9875 17926 9927 17978
rect 9939 17926 9991 17978
rect 10003 17926 10055 17978
rect 15612 17926 15664 17978
rect 15676 17926 15728 17978
rect 15740 17926 15792 17978
rect 15804 17926 15856 17978
rect 15868 17926 15920 17978
rect 21477 17926 21529 17978
rect 21541 17926 21593 17978
rect 21605 17926 21657 17978
rect 21669 17926 21721 17978
rect 21733 17926 21785 17978
rect 2136 17824 2188 17876
rect 5448 17824 5500 17876
rect 6276 17824 6328 17876
rect 7196 17824 7248 17876
rect 8208 17756 8260 17808
rect 9680 17756 9732 17808
rect 9864 17756 9916 17808
rect 1400 17663 1452 17672
rect 1400 17629 1409 17663
rect 1409 17629 1443 17663
rect 1443 17629 1452 17663
rect 1400 17620 1452 17629
rect 2780 17663 2832 17672
rect 2780 17629 2789 17663
rect 2789 17629 2823 17663
rect 2823 17629 2832 17663
rect 2780 17620 2832 17629
rect 3700 17620 3752 17672
rect 4252 17620 4304 17672
rect 4712 17620 4764 17672
rect 5540 17620 5592 17672
rect 1308 17552 1360 17604
rect 1860 17484 1912 17536
rect 3424 17484 3476 17536
rect 4344 17484 4396 17536
rect 6092 17484 6144 17536
rect 9128 17688 9180 17740
rect 11888 17824 11940 17876
rect 14556 17824 14608 17876
rect 7196 17663 7248 17672
rect 7196 17629 7205 17663
rect 7205 17629 7239 17663
rect 7239 17629 7248 17663
rect 7196 17620 7248 17629
rect 7380 17620 7432 17672
rect 8024 17620 8076 17672
rect 8944 17620 8996 17672
rect 9312 17620 9364 17672
rect 10140 17663 10192 17672
rect 10140 17629 10149 17663
rect 10149 17629 10192 17663
rect 10140 17620 10192 17629
rect 10600 17620 10652 17672
rect 11152 17620 11204 17672
rect 12256 17663 12308 17672
rect 12256 17629 12290 17663
rect 12290 17629 12308 17663
rect 12256 17620 12308 17629
rect 12440 17663 12492 17672
rect 12440 17629 12449 17663
rect 12449 17629 12483 17663
rect 12483 17629 12492 17663
rect 12440 17620 12492 17629
rect 13820 17620 13872 17672
rect 14740 17620 14792 17672
rect 7656 17484 7708 17536
rect 8116 17484 8168 17536
rect 16488 17688 16540 17740
rect 15568 17620 15620 17672
rect 16948 17663 17000 17672
rect 11152 17484 11204 17536
rect 11888 17484 11940 17536
rect 16948 17629 16955 17663
rect 16955 17629 16989 17663
rect 16989 17629 17000 17663
rect 16948 17620 17000 17629
rect 17868 17824 17920 17876
rect 22376 17824 22428 17876
rect 24860 17756 24912 17808
rect 21456 17688 21508 17740
rect 17960 17620 18012 17672
rect 19156 17620 19208 17672
rect 22008 17663 22060 17672
rect 22008 17629 22017 17663
rect 22017 17629 22051 17663
rect 22051 17629 22060 17663
rect 22008 17620 22060 17629
rect 23848 17620 23900 17672
rect 24216 17620 24268 17672
rect 20720 17595 20772 17604
rect 20720 17561 20732 17595
rect 20732 17561 20772 17595
rect 20720 17552 20772 17561
rect 20812 17552 20864 17604
rect 19340 17527 19392 17536
rect 19340 17493 19349 17527
rect 19349 17493 19383 17527
rect 19383 17493 19392 17527
rect 19340 17484 19392 17493
rect 20076 17484 20128 17536
rect 21456 17484 21508 17536
rect 21824 17527 21876 17536
rect 21824 17493 21833 17527
rect 21833 17493 21867 17527
rect 21867 17493 21876 17527
rect 21824 17484 21876 17493
rect 22744 17484 22796 17536
rect 23388 17527 23440 17536
rect 23388 17493 23397 17527
rect 23397 17493 23431 17527
rect 23431 17493 23440 17527
rect 23388 17484 23440 17493
rect 6814 17382 6866 17434
rect 6878 17382 6930 17434
rect 6942 17382 6994 17434
rect 7006 17382 7058 17434
rect 7070 17382 7122 17434
rect 12679 17382 12731 17434
rect 12743 17382 12795 17434
rect 12807 17382 12859 17434
rect 12871 17382 12923 17434
rect 12935 17382 12987 17434
rect 18544 17382 18596 17434
rect 18608 17382 18660 17434
rect 18672 17382 18724 17434
rect 18736 17382 18788 17434
rect 18800 17382 18852 17434
rect 24409 17382 24461 17434
rect 24473 17382 24525 17434
rect 24537 17382 24589 17434
rect 24601 17382 24653 17434
rect 24665 17382 24717 17434
rect 2596 17280 2648 17332
rect 4344 17280 4396 17332
rect 4620 17280 4672 17332
rect 1492 17187 1544 17196
rect 1492 17153 1501 17187
rect 1501 17153 1535 17187
rect 1535 17153 1544 17187
rect 1492 17144 1544 17153
rect 3056 17212 3108 17264
rect 5172 17280 5224 17332
rect 7288 17280 7340 17332
rect 2228 17187 2280 17196
rect 2228 17153 2235 17187
rect 2235 17153 2269 17187
rect 2269 17153 2280 17187
rect 2228 17144 2280 17153
rect 3240 17144 3292 17196
rect 4068 17144 4120 17196
rect 6644 17217 6696 17264
rect 5908 17144 5960 17196
rect 6368 17187 6420 17196
rect 6368 17153 6377 17187
rect 6377 17153 6411 17187
rect 6411 17153 6420 17187
rect 6368 17144 6420 17153
rect 6644 17212 6669 17217
rect 6669 17212 6696 17217
rect 7104 17212 7156 17264
rect 8300 17280 8352 17332
rect 8852 17280 8904 17332
rect 10416 17280 10468 17332
rect 8024 17144 8076 17196
rect 8576 17144 8628 17196
rect 8852 17144 8904 17196
rect 4712 17076 4764 17128
rect 8116 17076 8168 17128
rect 848 16940 900 16992
rect 3608 16940 3660 16992
rect 4436 16940 4488 16992
rect 5356 16940 5408 16992
rect 6184 17008 6236 17060
rect 7196 17008 7248 17060
rect 9128 17212 9180 17264
rect 12256 17280 12308 17332
rect 12440 17280 12492 17332
rect 11152 17212 11204 17264
rect 15292 17280 15344 17332
rect 16304 17280 16356 17332
rect 16580 17280 16632 17332
rect 17316 17280 17368 17332
rect 21824 17280 21876 17332
rect 19156 17255 19208 17264
rect 19156 17221 19190 17255
rect 19190 17221 19208 17255
rect 19156 17212 19208 17221
rect 9312 17144 9364 17196
rect 9864 17144 9916 17196
rect 13452 17144 13504 17196
rect 15016 17144 15068 17196
rect 15568 17187 15620 17196
rect 15568 17153 15577 17187
rect 15577 17153 15611 17187
rect 15611 17153 15620 17187
rect 15568 17144 15620 17153
rect 16488 17144 16540 17196
rect 16580 17144 16632 17196
rect 19616 17144 19668 17196
rect 20720 17144 20772 17196
rect 10600 17076 10652 17128
rect 5908 16983 5960 16992
rect 5908 16949 5917 16983
rect 5917 16949 5951 16983
rect 5951 16949 5960 16983
rect 5908 16940 5960 16949
rect 6092 16940 6144 16992
rect 7104 16940 7156 16992
rect 7380 16983 7432 16992
rect 7380 16949 7389 16983
rect 7389 16949 7423 16983
rect 7423 16949 7432 16983
rect 7380 16940 7432 16949
rect 7932 16940 7984 16992
rect 9220 16983 9272 16992
rect 9220 16949 9229 16983
rect 9229 16949 9263 16983
rect 9263 16949 9272 16983
rect 9220 16940 9272 16949
rect 9496 16940 9548 16992
rect 9588 16940 9640 16992
rect 10232 16940 10284 16992
rect 14372 17076 14424 17128
rect 14740 17076 14792 17128
rect 16028 17076 16080 17128
rect 17960 17076 18012 17128
rect 18880 17119 18932 17128
rect 18880 17085 18889 17119
rect 18889 17085 18923 17119
rect 18923 17085 18932 17119
rect 18880 17076 18932 17085
rect 20352 17119 20404 17128
rect 20352 17085 20361 17119
rect 20361 17085 20395 17119
rect 20395 17085 20404 17119
rect 20352 17076 20404 17085
rect 23388 17280 23440 17332
rect 22744 17187 22796 17196
rect 22744 17153 22753 17187
rect 22753 17153 22787 17187
rect 22787 17153 22796 17187
rect 22744 17144 22796 17153
rect 23756 17187 23808 17196
rect 23756 17153 23765 17187
rect 23765 17153 23799 17187
rect 23799 17153 23808 17187
rect 23756 17144 23808 17153
rect 23848 17144 23900 17196
rect 15292 17051 15344 17060
rect 15292 17017 15301 17051
rect 15301 17017 15335 17051
rect 15335 17017 15344 17051
rect 15292 17008 15344 17017
rect 12256 16940 12308 16992
rect 16488 16983 16540 16992
rect 16488 16949 16497 16983
rect 16497 16949 16531 16983
rect 16531 16949 16540 16983
rect 16488 16940 16540 16949
rect 20720 16940 20772 16992
rect 21088 16940 21140 16992
rect 22284 16940 22336 16992
rect 23480 16940 23532 16992
rect 23572 16983 23624 16992
rect 23572 16949 23581 16983
rect 23581 16949 23615 16983
rect 23615 16949 23624 16983
rect 23572 16940 23624 16949
rect 24124 16940 24176 16992
rect 3882 16838 3934 16890
rect 3946 16838 3998 16890
rect 4010 16838 4062 16890
rect 4074 16838 4126 16890
rect 4138 16838 4190 16890
rect 9747 16838 9799 16890
rect 9811 16838 9863 16890
rect 9875 16838 9927 16890
rect 9939 16838 9991 16890
rect 10003 16838 10055 16890
rect 15612 16838 15664 16890
rect 15676 16838 15728 16890
rect 15740 16838 15792 16890
rect 15804 16838 15856 16890
rect 15868 16838 15920 16890
rect 21477 16838 21529 16890
rect 21541 16838 21593 16890
rect 21605 16838 21657 16890
rect 21669 16838 21721 16890
rect 21733 16838 21785 16890
rect 1768 16668 1820 16720
rect 1860 16668 1912 16720
rect 2320 16600 2372 16652
rect 2596 16643 2648 16652
rect 2596 16609 2630 16643
rect 2630 16609 2648 16643
rect 2596 16600 2648 16609
rect 2964 16600 3016 16652
rect 4620 16668 4672 16720
rect 3424 16643 3476 16652
rect 3424 16609 3433 16643
rect 3433 16609 3467 16643
rect 3467 16609 3476 16643
rect 3424 16600 3476 16609
rect 5540 16736 5592 16788
rect 5908 16736 5960 16788
rect 5172 16643 5224 16652
rect 5172 16609 5181 16643
rect 5181 16609 5215 16643
rect 5215 16609 5224 16643
rect 5172 16600 5224 16609
rect 5356 16600 5408 16652
rect 7380 16736 7432 16788
rect 7932 16736 7984 16788
rect 9588 16736 9640 16788
rect 6092 16600 6144 16652
rect 6184 16643 6236 16652
rect 6184 16609 6193 16643
rect 6193 16609 6227 16643
rect 6227 16609 6236 16643
rect 6184 16600 6236 16609
rect 1952 16532 2004 16584
rect 2780 16575 2832 16584
rect 2780 16541 2789 16575
rect 2789 16541 2823 16575
rect 2823 16541 2832 16575
rect 2780 16532 2832 16541
rect 3792 16575 3844 16584
rect 3792 16541 3801 16575
rect 3801 16541 3835 16575
rect 3835 16541 3844 16575
rect 3792 16532 3844 16541
rect 3884 16532 3936 16584
rect 4344 16532 4396 16584
rect 6276 16532 6328 16584
rect 6736 16600 6788 16652
rect 8024 16600 8076 16652
rect 9680 16600 9732 16652
rect 10876 16668 10928 16720
rect 11612 16600 11664 16652
rect 12256 16736 12308 16788
rect 15292 16736 15344 16788
rect 21456 16736 21508 16788
rect 22284 16736 22336 16788
rect 7104 16575 7156 16584
rect 7104 16541 7113 16575
rect 7113 16541 7147 16575
rect 7147 16541 7156 16575
rect 7104 16532 7156 16541
rect 7378 16575 7430 16584
rect 7378 16541 7387 16575
rect 7387 16541 7421 16575
rect 7421 16541 7430 16575
rect 7378 16532 7430 16541
rect 10048 16532 10100 16584
rect 17960 16600 18012 16652
rect 19340 16600 19392 16652
rect 848 16396 900 16448
rect 1216 16396 1268 16448
rect 1676 16396 1728 16448
rect 4252 16396 4304 16448
rect 5908 16396 5960 16448
rect 6184 16396 6236 16448
rect 6552 16396 6604 16448
rect 9128 16464 9180 16516
rect 9404 16464 9456 16516
rect 8024 16439 8076 16448
rect 8024 16405 8033 16439
rect 8033 16405 8067 16439
rect 8067 16405 8076 16439
rect 8024 16396 8076 16405
rect 9496 16396 9548 16448
rect 11428 16396 11480 16448
rect 11980 16464 12032 16516
rect 13360 16532 13412 16584
rect 14096 16532 14148 16584
rect 14556 16464 14608 16516
rect 16488 16532 16540 16584
rect 18420 16532 18472 16584
rect 18880 16575 18932 16584
rect 18880 16541 18889 16575
rect 18889 16541 18923 16575
rect 18923 16541 18932 16575
rect 18880 16532 18932 16541
rect 19524 16575 19576 16584
rect 19524 16541 19533 16575
rect 19533 16541 19567 16575
rect 19567 16541 19576 16575
rect 19524 16532 19576 16541
rect 20996 16668 21048 16720
rect 20720 16532 20772 16584
rect 20996 16575 21048 16584
rect 20996 16541 21005 16575
rect 21005 16541 21039 16575
rect 21039 16541 21048 16575
rect 20996 16532 21048 16541
rect 12440 16396 12492 16448
rect 13084 16396 13136 16448
rect 14372 16396 14424 16448
rect 15108 16396 15160 16448
rect 20628 16507 20680 16516
rect 20628 16473 20637 16507
rect 20637 16473 20671 16507
rect 20671 16473 20680 16507
rect 20628 16464 20680 16473
rect 22100 16575 22152 16584
rect 22100 16541 22109 16575
rect 22109 16541 22143 16575
rect 22143 16541 22152 16575
rect 22100 16532 22152 16541
rect 23480 16736 23532 16788
rect 23756 16736 23808 16788
rect 24124 16779 24176 16788
rect 24124 16745 24133 16779
rect 24133 16745 24167 16779
rect 24167 16745 24176 16779
rect 24124 16736 24176 16745
rect 22468 16464 22520 16516
rect 22100 16396 22152 16448
rect 22192 16396 22244 16448
rect 22836 16396 22888 16448
rect 6814 16294 6866 16346
rect 6878 16294 6930 16346
rect 6942 16294 6994 16346
rect 7006 16294 7058 16346
rect 7070 16294 7122 16346
rect 12679 16294 12731 16346
rect 12743 16294 12795 16346
rect 12807 16294 12859 16346
rect 12871 16294 12923 16346
rect 12935 16294 12987 16346
rect 18544 16294 18596 16346
rect 18608 16294 18660 16346
rect 18672 16294 18724 16346
rect 18736 16294 18788 16346
rect 18800 16294 18852 16346
rect 24409 16294 24461 16346
rect 24473 16294 24525 16346
rect 24537 16294 24589 16346
rect 24601 16294 24653 16346
rect 24665 16294 24717 16346
rect 2044 16192 2096 16244
rect 2228 16192 2280 16244
rect 2780 16192 2832 16244
rect 2964 16124 3016 16176
rect 2320 16056 2372 16108
rect 4344 16192 4396 16244
rect 5908 16192 5960 16244
rect 7380 16192 7432 16244
rect 8852 16192 8904 16244
rect 4160 16099 4212 16108
rect 4160 16065 4169 16099
rect 4169 16065 4203 16099
rect 4203 16065 4212 16099
rect 4160 16056 4212 16065
rect 4436 16099 4488 16108
rect 4436 16065 4445 16099
rect 4445 16065 4479 16099
rect 4479 16065 4488 16099
rect 4436 16056 4488 16065
rect 5264 16056 5316 16108
rect 6092 16056 6144 16108
rect 6368 16056 6420 16108
rect 6828 16056 6880 16108
rect 7932 16056 7984 16108
rect 8300 16099 8352 16108
rect 8300 16065 8307 16099
rect 8307 16065 8341 16099
rect 8341 16065 8352 16099
rect 8300 16056 8352 16065
rect 9496 16099 9548 16108
rect 9496 16065 9505 16099
rect 9505 16065 9539 16099
rect 9539 16065 9548 16099
rect 9496 16056 9548 16065
rect 12992 16192 13044 16244
rect 13176 16192 13228 16244
rect 13452 16192 13504 16244
rect 13636 16192 13688 16244
rect 14096 16192 14148 16244
rect 13360 16099 13412 16108
rect 13360 16065 13369 16099
rect 13369 16065 13403 16099
rect 13403 16065 13412 16099
rect 13360 16056 13412 16065
rect 13636 16099 13688 16108
rect 13636 16065 13645 16099
rect 13645 16065 13679 16099
rect 13679 16065 13688 16099
rect 13636 16056 13688 16065
rect 1400 15988 1452 16040
rect 3608 15988 3660 16040
rect 6276 15988 6328 16040
rect 7656 15988 7708 16040
rect 1768 15852 1820 15904
rect 2780 15852 2832 15904
rect 3792 15852 3844 15904
rect 4252 15852 4304 15904
rect 9588 15988 9640 16040
rect 10048 15988 10100 16040
rect 10140 16031 10192 16040
rect 10140 15997 10149 16031
rect 10149 15997 10183 16031
rect 10183 15997 10192 16031
rect 10140 15988 10192 15997
rect 10554 16031 10606 16040
rect 10554 15997 10563 16031
rect 10563 15997 10597 16031
rect 10597 15997 10606 16031
rect 10554 15988 10606 15997
rect 10876 15988 10928 16040
rect 12440 16031 12492 16040
rect 12440 15997 12449 16031
rect 12449 15997 12483 16031
rect 12483 15997 12492 16031
rect 12440 15988 12492 15997
rect 13084 16031 13136 16040
rect 13084 15997 13093 16031
rect 13093 15997 13127 16031
rect 13127 15997 13136 16031
rect 13084 15988 13136 15997
rect 12348 15920 12400 15972
rect 15200 16124 15252 16176
rect 15292 16056 15344 16108
rect 15108 16031 15160 16040
rect 15108 15997 15117 16031
rect 15117 15997 15151 16031
rect 15151 15997 15160 16031
rect 15108 15988 15160 15997
rect 16028 16192 16080 16244
rect 16488 16192 16540 16244
rect 18420 16192 18472 16244
rect 19524 16192 19576 16244
rect 22100 16192 22152 16244
rect 18880 16124 18932 16176
rect 21456 16124 21508 16176
rect 22468 16192 22520 16244
rect 24860 16192 24912 16244
rect 18512 16056 18564 16108
rect 20352 15988 20404 16040
rect 9128 15852 9180 15904
rect 16580 15852 16632 15904
rect 17684 15852 17736 15904
rect 22192 15852 22244 15904
rect 23756 15895 23808 15904
rect 23756 15861 23765 15895
rect 23765 15861 23799 15895
rect 23799 15861 23808 15895
rect 23756 15852 23808 15861
rect 3882 15750 3934 15802
rect 3946 15750 3998 15802
rect 4010 15750 4062 15802
rect 4074 15750 4126 15802
rect 4138 15750 4190 15802
rect 9747 15750 9799 15802
rect 9811 15750 9863 15802
rect 9875 15750 9927 15802
rect 9939 15750 9991 15802
rect 10003 15750 10055 15802
rect 15612 15750 15664 15802
rect 15676 15750 15728 15802
rect 15740 15750 15792 15802
rect 15804 15750 15856 15802
rect 15868 15750 15920 15802
rect 21477 15750 21529 15802
rect 21541 15750 21593 15802
rect 21605 15750 21657 15802
rect 21669 15750 21721 15802
rect 21733 15750 21785 15802
rect 1124 15648 1176 15700
rect 1216 15580 1268 15632
rect 3332 15648 3384 15700
rect 5540 15691 5592 15700
rect 5540 15657 5549 15691
rect 5549 15657 5583 15691
rect 5583 15657 5592 15691
rect 5540 15648 5592 15657
rect 11336 15648 11388 15700
rect 12256 15648 12308 15700
rect 9588 15580 9640 15632
rect 11612 15580 11664 15632
rect 12164 15580 12216 15632
rect 13636 15691 13688 15700
rect 13636 15657 13645 15691
rect 13645 15657 13679 15691
rect 13679 15657 13688 15691
rect 13636 15648 13688 15657
rect 14372 15512 14424 15564
rect 1308 15376 1360 15428
rect 2964 15376 3016 15428
rect 4712 15444 4764 15496
rect 4804 15487 4856 15496
rect 4804 15453 4811 15487
rect 4811 15453 4845 15487
rect 4845 15453 4856 15487
rect 4804 15444 4856 15453
rect 7196 15444 7248 15496
rect 7288 15444 7340 15496
rect 8024 15444 8076 15496
rect 9404 15444 9456 15496
rect 10140 15444 10192 15496
rect 10508 15444 10560 15496
rect 11244 15376 11296 15428
rect 14096 15444 14148 15496
rect 15936 15648 15988 15700
rect 16212 15580 16264 15632
rect 14832 15487 14884 15496
rect 14832 15453 14839 15487
rect 14839 15453 14873 15487
rect 14873 15453 14884 15487
rect 14832 15444 14884 15453
rect 14740 15376 14792 15428
rect 16580 15444 16632 15496
rect 18512 15444 18564 15496
rect 15108 15376 15160 15428
rect 17224 15376 17276 15428
rect 19984 15444 20036 15496
rect 23848 15487 23900 15496
rect 23848 15453 23857 15487
rect 23857 15453 23891 15487
rect 23891 15453 23900 15487
rect 23848 15444 23900 15453
rect 22652 15376 22704 15428
rect 24860 15376 24912 15428
rect 5540 15308 5592 15360
rect 11428 15308 11480 15360
rect 13452 15308 13504 15360
rect 13912 15308 13964 15360
rect 14280 15308 14332 15360
rect 14832 15308 14884 15360
rect 15016 15308 15068 15360
rect 15476 15308 15528 15360
rect 18052 15308 18104 15360
rect 20352 15308 20404 15360
rect 20812 15308 20864 15360
rect 21364 15308 21416 15360
rect 6814 15206 6866 15258
rect 6878 15206 6930 15258
rect 6942 15206 6994 15258
rect 7006 15206 7058 15258
rect 7070 15206 7122 15258
rect 12679 15206 12731 15258
rect 12743 15206 12795 15258
rect 12807 15206 12859 15258
rect 12871 15206 12923 15258
rect 12935 15206 12987 15258
rect 18544 15206 18596 15258
rect 18608 15206 18660 15258
rect 18672 15206 18724 15258
rect 18736 15206 18788 15258
rect 18800 15206 18852 15258
rect 24409 15206 24461 15258
rect 24473 15206 24525 15258
rect 24537 15206 24589 15258
rect 24601 15206 24653 15258
rect 24665 15206 24717 15258
rect 1308 15104 1360 15156
rect 3700 15147 3752 15156
rect 3700 15113 3709 15147
rect 3709 15113 3743 15147
rect 3743 15113 3752 15147
rect 3700 15104 3752 15113
rect 4436 15104 4488 15156
rect 7196 15104 7248 15156
rect 8024 15104 8076 15156
rect 664 15036 716 15088
rect 4344 15036 4396 15088
rect 1400 14943 1452 14952
rect 1400 14909 1409 14943
rect 1409 14909 1443 14943
rect 1443 14909 1452 14943
rect 1400 14900 1452 14909
rect 2228 14764 2280 14816
rect 3700 14968 3752 15020
rect 4528 15036 4580 15088
rect 7472 14968 7524 15020
rect 8484 15011 8536 15020
rect 8484 14977 8493 15011
rect 8493 14977 8527 15011
rect 8527 14977 8536 15011
rect 8484 14968 8536 14977
rect 9404 15011 9456 15020
rect 9404 14977 9413 15011
rect 9413 14977 9447 15011
rect 9447 14977 9456 15011
rect 9404 14968 9456 14977
rect 4528 14900 4580 14952
rect 3792 14832 3844 14884
rect 4160 14832 4212 14884
rect 7104 14943 7156 14952
rect 7104 14909 7113 14943
rect 7113 14909 7147 14943
rect 7147 14909 7156 14943
rect 7104 14900 7156 14909
rect 8300 14900 8352 14952
rect 9036 14900 9088 14952
rect 10232 14900 10284 14952
rect 11980 14900 12032 14952
rect 13176 14900 13228 14952
rect 16580 15036 16632 15088
rect 18144 15104 18196 15156
rect 18972 15104 19024 15156
rect 5540 14764 5592 14816
rect 10140 14832 10192 14884
rect 10600 14764 10652 14816
rect 14464 14943 14516 14952
rect 14464 14909 14473 14943
rect 14473 14909 14507 14943
rect 14507 14909 14516 14943
rect 14464 14900 14516 14909
rect 15476 15011 15528 15020
rect 15476 14977 15485 15011
rect 15485 14977 15519 15011
rect 15519 14977 15528 15011
rect 15476 14968 15528 14977
rect 16304 14968 16356 15020
rect 18696 15011 18748 15020
rect 18696 14977 18705 15011
rect 18705 14977 18739 15011
rect 18739 14977 18748 15011
rect 18696 14968 18748 14977
rect 18880 15011 18932 15020
rect 18880 14977 18889 15011
rect 18889 14977 18923 15011
rect 18923 14977 18932 15011
rect 18880 14968 18932 14977
rect 19984 14968 20036 15020
rect 20628 15011 20680 15020
rect 20628 14977 20637 15011
rect 20637 14977 20671 15011
rect 20671 14977 20680 15011
rect 20628 14968 20680 14977
rect 14832 14900 14884 14952
rect 15200 14943 15252 14952
rect 15200 14909 15209 14943
rect 15209 14909 15243 14943
rect 15243 14909 15252 14943
rect 15200 14900 15252 14909
rect 14280 14832 14332 14884
rect 14924 14875 14976 14884
rect 14924 14841 14933 14875
rect 14933 14841 14967 14875
rect 14967 14841 14976 14875
rect 14924 14832 14976 14841
rect 22008 14968 22060 15020
rect 23020 14968 23072 15020
rect 21088 14832 21140 14884
rect 17960 14764 18012 14816
rect 18328 14807 18380 14816
rect 18328 14773 18337 14807
rect 18337 14773 18371 14807
rect 18371 14773 18380 14807
rect 18328 14764 18380 14773
rect 18788 14807 18840 14816
rect 18788 14773 18797 14807
rect 18797 14773 18831 14807
rect 18831 14773 18840 14807
rect 18788 14764 18840 14773
rect 19156 14764 19208 14816
rect 20812 14764 20864 14816
rect 20996 14807 21048 14816
rect 20996 14773 21005 14807
rect 21005 14773 21039 14807
rect 21039 14773 21048 14807
rect 20996 14764 21048 14773
rect 21364 14764 21416 14816
rect 23296 14764 23348 14816
rect 24124 14807 24176 14816
rect 24124 14773 24133 14807
rect 24133 14773 24167 14807
rect 24167 14773 24176 14807
rect 24124 14764 24176 14773
rect 3882 14662 3934 14714
rect 3946 14662 3998 14714
rect 4010 14662 4062 14714
rect 4074 14662 4126 14714
rect 4138 14662 4190 14714
rect 9747 14662 9799 14714
rect 9811 14662 9863 14714
rect 9875 14662 9927 14714
rect 9939 14662 9991 14714
rect 10003 14662 10055 14714
rect 15612 14662 15664 14714
rect 15676 14662 15728 14714
rect 15740 14662 15792 14714
rect 15804 14662 15856 14714
rect 15868 14662 15920 14714
rect 21477 14662 21529 14714
rect 21541 14662 21593 14714
rect 21605 14662 21657 14714
rect 21669 14662 21721 14714
rect 21733 14662 21785 14714
rect 1584 14603 1636 14612
rect 1584 14569 1593 14603
rect 1593 14569 1627 14603
rect 1627 14569 1636 14603
rect 1584 14560 1636 14569
rect 1124 14492 1176 14544
rect 3976 14603 4028 14612
rect 3976 14569 3985 14603
rect 3985 14569 4019 14603
rect 4019 14569 4028 14603
rect 3976 14560 4028 14569
rect 7104 14560 7156 14612
rect 4160 14492 4212 14544
rect 296 14424 348 14476
rect 940 14424 992 14476
rect 4988 14467 5040 14476
rect 4988 14433 4997 14467
rect 4997 14433 5031 14467
rect 5031 14433 5040 14467
rect 4988 14424 5040 14433
rect 5264 14467 5316 14476
rect 5264 14433 5273 14467
rect 5273 14433 5307 14467
rect 5307 14433 5316 14467
rect 5264 14424 5316 14433
rect 5540 14467 5592 14476
rect 5540 14433 5549 14467
rect 5549 14433 5583 14467
rect 5583 14433 5592 14467
rect 5540 14424 5592 14433
rect 6368 14424 6420 14476
rect 10140 14560 10192 14612
rect 11336 14560 11388 14612
rect 11888 14492 11940 14544
rect 11980 14492 12032 14544
rect 13084 14560 13136 14612
rect 14924 14560 14976 14612
rect 15200 14560 15252 14612
rect 15936 14560 15988 14612
rect 16580 14560 16632 14612
rect 17408 14560 17460 14612
rect 18696 14603 18748 14612
rect 18696 14569 18705 14603
rect 18705 14569 18739 14603
rect 18739 14569 18748 14603
rect 18696 14560 18748 14569
rect 18788 14560 18840 14612
rect 20628 14603 20680 14612
rect 20628 14569 20637 14603
rect 20637 14569 20671 14603
rect 20671 14569 20680 14603
rect 20628 14560 20680 14569
rect 20996 14560 21048 14612
rect 21088 14603 21140 14612
rect 21088 14569 21097 14603
rect 21097 14569 21131 14603
rect 21131 14569 21140 14603
rect 21088 14560 21140 14569
rect 21364 14603 21416 14612
rect 21364 14569 21373 14603
rect 21373 14569 21407 14603
rect 21407 14569 21416 14603
rect 21364 14560 21416 14569
rect 10876 14424 10928 14476
rect 2688 14356 2740 14408
rect 4436 14356 4488 14408
rect 5448 14356 5500 14408
rect 7564 14356 7616 14408
rect 8024 14356 8076 14408
rect 8760 14356 8812 14408
rect 1492 14331 1544 14340
rect 1492 14297 1501 14331
rect 1501 14297 1535 14331
rect 1535 14297 1544 14331
rect 1492 14288 1544 14297
rect 4528 14288 4580 14340
rect 7196 14288 7248 14340
rect 2320 14220 2372 14272
rect 4896 14220 4948 14272
rect 5080 14220 5132 14272
rect 8300 14220 8352 14272
rect 14096 14399 14148 14408
rect 14096 14365 14105 14399
rect 14105 14365 14139 14399
rect 14139 14365 14148 14399
rect 14096 14356 14148 14365
rect 15200 14356 15252 14408
rect 17500 14356 17552 14408
rect 17684 14399 17736 14408
rect 17684 14365 17693 14399
rect 17693 14365 17727 14399
rect 17727 14365 17736 14399
rect 17684 14356 17736 14365
rect 14188 14288 14240 14340
rect 18144 14288 18196 14340
rect 12440 14220 12492 14272
rect 13084 14263 13136 14272
rect 13084 14229 13093 14263
rect 13093 14229 13127 14263
rect 13127 14229 13136 14263
rect 13084 14220 13136 14229
rect 13452 14220 13504 14272
rect 14740 14220 14792 14272
rect 15016 14220 15068 14272
rect 16212 14220 16264 14272
rect 17684 14220 17736 14272
rect 19984 14356 20036 14408
rect 20352 14356 20404 14408
rect 23756 14560 23808 14612
rect 22836 14535 22888 14544
rect 22836 14501 22845 14535
rect 22845 14501 22879 14535
rect 22879 14501 22888 14535
rect 22836 14492 22888 14501
rect 23296 14492 23348 14544
rect 23020 14399 23072 14408
rect 23020 14365 23029 14399
rect 23029 14365 23063 14399
rect 23063 14365 23072 14399
rect 23020 14356 23072 14365
rect 20812 14288 20864 14340
rect 23756 14399 23808 14408
rect 23756 14365 23765 14399
rect 23765 14365 23799 14399
rect 23799 14365 23808 14399
rect 23756 14356 23808 14365
rect 23848 14399 23900 14408
rect 23848 14365 23857 14399
rect 23857 14365 23891 14399
rect 23891 14365 23900 14399
rect 23848 14356 23900 14365
rect 19800 14220 19852 14272
rect 21180 14220 21232 14272
rect 23020 14220 23072 14272
rect 24860 14220 24912 14272
rect 6814 14118 6866 14170
rect 6878 14118 6930 14170
rect 6942 14118 6994 14170
rect 7006 14118 7058 14170
rect 7070 14118 7122 14170
rect 12679 14118 12731 14170
rect 12743 14118 12795 14170
rect 12807 14118 12859 14170
rect 12871 14118 12923 14170
rect 12935 14118 12987 14170
rect 18544 14118 18596 14170
rect 18608 14118 18660 14170
rect 18672 14118 18724 14170
rect 18736 14118 18788 14170
rect 18800 14118 18852 14170
rect 24409 14118 24461 14170
rect 24473 14118 24525 14170
rect 24537 14118 24589 14170
rect 24601 14118 24653 14170
rect 24665 14118 24717 14170
rect 1492 14016 1544 14068
rect 7656 14016 7708 14068
rect 7748 14016 7800 14068
rect 1676 13948 1728 14000
rect 2412 13923 2464 13932
rect 2412 13889 2421 13923
rect 2421 13889 2455 13923
rect 2455 13889 2464 13923
rect 2412 13880 2464 13889
rect 2596 13880 2648 13932
rect 6368 13948 6420 14000
rect 12072 14016 12124 14068
rect 12164 14016 12216 14068
rect 13360 14016 13412 14068
rect 1492 13855 1544 13864
rect 1492 13821 1501 13855
rect 1501 13821 1535 13855
rect 1535 13821 1544 13855
rect 1492 13812 1544 13821
rect 2228 13812 2280 13864
rect 2688 13855 2740 13864
rect 2688 13821 2697 13855
rect 2697 13821 2731 13855
rect 2731 13821 2740 13855
rect 2688 13812 2740 13821
rect 2872 13812 2924 13864
rect 5172 13923 5224 13932
rect 5172 13889 5179 13923
rect 5179 13889 5213 13923
rect 5213 13889 5224 13923
rect 5172 13880 5224 13889
rect 5540 13880 5592 13932
rect 6552 13880 6604 13932
rect 7472 13880 7524 13932
rect 8300 13923 8352 13932
rect 8300 13889 8309 13923
rect 8309 13889 8343 13923
rect 8343 13889 8352 13923
rect 8300 13880 8352 13889
rect 9312 13880 9364 13932
rect 1860 13744 1912 13796
rect 1952 13676 2004 13728
rect 2872 13676 2924 13728
rect 3240 13676 3292 13728
rect 6460 13812 6512 13864
rect 6736 13812 6788 13864
rect 7196 13812 7248 13864
rect 8024 13855 8076 13864
rect 8024 13821 8033 13855
rect 8033 13821 8067 13855
rect 8067 13821 8076 13855
rect 8024 13812 8076 13821
rect 8208 13812 8260 13864
rect 3792 13676 3844 13728
rect 4436 13719 4488 13728
rect 4436 13685 4445 13719
rect 4445 13685 4479 13719
rect 4479 13685 4488 13719
rect 4436 13676 4488 13685
rect 4620 13676 4672 13728
rect 7472 13744 7524 13796
rect 7748 13787 7800 13796
rect 7748 13753 7757 13787
rect 7757 13753 7791 13787
rect 7791 13753 7800 13787
rect 7748 13744 7800 13753
rect 5908 13719 5960 13728
rect 5908 13685 5917 13719
rect 5917 13685 5951 13719
rect 5951 13685 5960 13719
rect 5908 13676 5960 13685
rect 9036 13676 9088 13728
rect 11336 13744 11388 13796
rect 11612 13812 11664 13864
rect 12440 13923 12492 13932
rect 12440 13889 12449 13923
rect 12449 13889 12483 13923
rect 12483 13889 12492 13923
rect 12440 13880 12492 13889
rect 12716 13923 12768 13932
rect 12716 13889 12725 13923
rect 12725 13889 12759 13923
rect 12759 13889 12768 13923
rect 12716 13880 12768 13889
rect 14740 13991 14792 14000
rect 14740 13957 14749 13991
rect 14749 13957 14783 13991
rect 14783 13957 14792 13991
rect 14740 13948 14792 13957
rect 15292 13948 15344 14000
rect 15568 13948 15620 14000
rect 13912 13923 13964 13932
rect 13912 13889 13921 13923
rect 13921 13889 13955 13923
rect 13955 13889 13964 13923
rect 13912 13880 13964 13889
rect 14004 13923 14056 13932
rect 14004 13889 14013 13923
rect 14013 13889 14047 13923
rect 14047 13889 14056 13923
rect 14004 13880 14056 13889
rect 14188 13880 14240 13932
rect 14556 13880 14608 13932
rect 11796 13744 11848 13796
rect 10876 13676 10928 13728
rect 11612 13676 11664 13728
rect 13084 13812 13136 13864
rect 15016 13812 15068 13864
rect 16212 13812 16264 13864
rect 18052 14016 18104 14068
rect 18144 14059 18196 14068
rect 18144 14025 18153 14059
rect 18153 14025 18187 14059
rect 18187 14025 18196 14059
rect 18144 14016 18196 14025
rect 18328 14016 18380 14068
rect 18880 14016 18932 14068
rect 19892 14016 19944 14068
rect 20168 14016 20220 14068
rect 22284 14016 22336 14068
rect 23848 14016 23900 14068
rect 18972 13948 19024 14000
rect 21180 13948 21232 14000
rect 19800 13880 19852 13932
rect 22192 13948 22244 14000
rect 13084 13676 13136 13728
rect 13544 13676 13596 13728
rect 14832 13676 14884 13728
rect 16212 13719 16264 13728
rect 16212 13685 16221 13719
rect 16221 13685 16255 13719
rect 16255 13685 16264 13719
rect 16212 13676 16264 13685
rect 16488 13676 16540 13728
rect 21088 13812 21140 13864
rect 22100 13923 22152 13932
rect 22100 13889 22109 13923
rect 22109 13889 22143 13923
rect 22143 13889 22152 13923
rect 22100 13880 22152 13889
rect 22284 13923 22336 13932
rect 22284 13889 22293 13923
rect 22293 13889 22327 13923
rect 22327 13889 22336 13923
rect 22284 13880 22336 13889
rect 22560 13923 22612 13932
rect 22560 13889 22569 13923
rect 22569 13889 22603 13923
rect 22603 13889 22612 13923
rect 22560 13880 22612 13889
rect 23020 13948 23072 14000
rect 23756 13948 23808 14000
rect 22836 13812 22888 13864
rect 18328 13744 18380 13796
rect 19156 13744 19208 13796
rect 20352 13744 20404 13796
rect 17684 13719 17736 13728
rect 17684 13685 17693 13719
rect 17693 13685 17727 13719
rect 17727 13685 17736 13719
rect 17684 13676 17736 13685
rect 21364 13719 21416 13728
rect 21364 13685 21373 13719
rect 21373 13685 21407 13719
rect 21407 13685 21416 13719
rect 21364 13676 21416 13685
rect 22192 13719 22244 13728
rect 22192 13685 22201 13719
rect 22201 13685 22235 13719
rect 22235 13685 22244 13719
rect 22192 13676 22244 13685
rect 22652 13676 22704 13728
rect 3882 13574 3934 13626
rect 3946 13574 3998 13626
rect 4010 13574 4062 13626
rect 4074 13574 4126 13626
rect 4138 13574 4190 13626
rect 9747 13574 9799 13626
rect 9811 13574 9863 13626
rect 9875 13574 9927 13626
rect 9939 13574 9991 13626
rect 10003 13574 10055 13626
rect 15612 13574 15664 13626
rect 15676 13574 15728 13626
rect 15740 13574 15792 13626
rect 15804 13574 15856 13626
rect 15868 13574 15920 13626
rect 21477 13574 21529 13626
rect 21541 13574 21593 13626
rect 21605 13574 21657 13626
rect 21669 13574 21721 13626
rect 21733 13574 21785 13626
rect 2688 13472 2740 13524
rect 4988 13472 5040 13524
rect 7656 13515 7708 13524
rect 7656 13481 7665 13515
rect 7665 13481 7699 13515
rect 7699 13481 7708 13515
rect 7656 13472 7708 13481
rect 5908 13404 5960 13456
rect 3700 13336 3752 13388
rect 3792 13336 3844 13388
rect 4896 13336 4948 13388
rect 5172 13336 5224 13388
rect 6092 13336 6144 13388
rect 1400 13268 1452 13320
rect 4344 13281 4396 13320
rect 1952 13200 2004 13252
rect 2044 13200 2096 13252
rect 2596 13200 2648 13252
rect 2688 13200 2740 13252
rect 3700 13200 3752 13252
rect 4344 13268 4369 13281
rect 4369 13268 4396 13281
rect 5724 13268 5776 13320
rect 5172 13200 5224 13252
rect 6736 13311 6788 13320
rect 6736 13277 6745 13311
rect 6745 13277 6779 13311
rect 6779 13277 6788 13311
rect 6736 13268 6788 13277
rect 7380 13336 7432 13388
rect 7656 13336 7708 13388
rect 11888 13472 11940 13524
rect 12716 13472 12768 13524
rect 14004 13472 14056 13524
rect 14372 13472 14424 13524
rect 16028 13472 16080 13524
rect 16488 13472 16540 13524
rect 17040 13472 17092 13524
rect 22560 13472 22612 13524
rect 24124 13515 24176 13524
rect 24124 13481 24133 13515
rect 24133 13481 24167 13515
rect 24167 13481 24176 13515
rect 24124 13472 24176 13481
rect 16212 13404 16264 13456
rect 8668 13336 8720 13388
rect 10876 13336 10928 13388
rect 10232 13268 10284 13320
rect 10508 13311 10560 13320
rect 10508 13277 10517 13311
rect 10517 13277 10551 13311
rect 10551 13277 10560 13311
rect 10508 13268 10560 13277
rect 11980 13336 12032 13388
rect 14464 13336 14516 13388
rect 8576 13200 8628 13252
rect 11704 13268 11756 13320
rect 14280 13268 14332 13320
rect 15292 13268 15344 13320
rect 2228 13132 2280 13184
rect 6184 13132 6236 13184
rect 9956 13175 10008 13184
rect 9956 13141 9965 13175
rect 9965 13141 9999 13175
rect 9999 13141 10008 13175
rect 9956 13132 10008 13141
rect 12072 13200 12124 13252
rect 14004 13200 14056 13252
rect 11612 13132 11664 13184
rect 11980 13132 12032 13184
rect 13360 13132 13412 13184
rect 14188 13132 14240 13184
rect 16396 13379 16448 13388
rect 16396 13345 16405 13379
rect 16405 13345 16439 13379
rect 16439 13345 16448 13379
rect 16396 13336 16448 13345
rect 16488 13379 16540 13388
rect 16488 13345 16522 13379
rect 16522 13345 16540 13379
rect 16488 13336 16540 13345
rect 17684 13336 17736 13388
rect 22008 13336 22060 13388
rect 22560 13301 22612 13320
rect 22560 13268 22569 13301
rect 22569 13268 22612 13301
rect 21088 13243 21140 13252
rect 21088 13209 21122 13243
rect 21122 13209 21140 13243
rect 21088 13200 21140 13209
rect 21180 13200 21232 13252
rect 22376 13200 22428 13252
rect 22836 13200 22888 13252
rect 16396 13132 16448 13184
rect 17316 13175 17368 13184
rect 17316 13141 17325 13175
rect 17325 13141 17359 13175
rect 17359 13141 17368 13175
rect 17316 13132 17368 13141
rect 22284 13132 22336 13184
rect 6814 13030 6866 13082
rect 6878 13030 6930 13082
rect 6942 13030 6994 13082
rect 7006 13030 7058 13082
rect 7070 13030 7122 13082
rect 12679 13030 12731 13082
rect 12743 13030 12795 13082
rect 12807 13030 12859 13082
rect 12871 13030 12923 13082
rect 12935 13030 12987 13082
rect 18544 13030 18596 13082
rect 18608 13030 18660 13082
rect 18672 13030 18724 13082
rect 18736 13030 18788 13082
rect 18800 13030 18852 13082
rect 24409 13030 24461 13082
rect 24473 13030 24525 13082
rect 24537 13030 24589 13082
rect 24601 13030 24653 13082
rect 24665 13030 24717 13082
rect 1216 12928 1268 12980
rect 3608 12928 3660 12980
rect 6184 12928 6236 12980
rect 6736 12928 6788 12980
rect 7748 12928 7800 12980
rect 2136 12860 2188 12912
rect 2228 12903 2280 12912
rect 2228 12869 2237 12903
rect 2237 12869 2271 12903
rect 2271 12869 2280 12903
rect 2228 12860 2280 12869
rect 17316 12928 17368 12980
rect 18972 12928 19024 12980
rect 9496 12903 9548 12912
rect 9496 12869 9505 12903
rect 9505 12869 9539 12903
rect 9539 12869 9548 12903
rect 9496 12860 9548 12869
rect 10508 12860 10560 12912
rect 10600 12903 10652 12912
rect 10600 12869 10609 12903
rect 10609 12869 10643 12903
rect 10643 12869 10652 12903
rect 10600 12860 10652 12869
rect 11336 12860 11388 12912
rect 11612 12860 11664 12912
rect 2412 12792 2464 12844
rect 2688 12835 2740 12844
rect 2688 12801 2697 12835
rect 2697 12801 2731 12835
rect 2731 12801 2740 12835
rect 2688 12792 2740 12801
rect 2872 12835 2924 12844
rect 2872 12801 2881 12835
rect 2881 12801 2915 12835
rect 2915 12801 2924 12835
rect 2872 12792 2924 12801
rect 3700 12835 3752 12844
rect 3700 12801 3734 12835
rect 3734 12801 3752 12835
rect 3700 12792 3752 12801
rect 6368 12792 6420 12844
rect 6736 12792 6788 12844
rect 7656 12792 7708 12844
rect 10140 12792 10192 12844
rect 4436 12724 4488 12776
rect 4528 12724 4580 12776
rect 6276 12724 6328 12776
rect 9956 12724 10008 12776
rect 10784 12724 10836 12776
rect 11152 12724 11204 12776
rect 11888 12792 11940 12844
rect 15936 12792 15988 12844
rect 16120 12792 16172 12844
rect 17408 12792 17460 12844
rect 19616 12835 19668 12844
rect 19616 12801 19625 12835
rect 19625 12801 19659 12835
rect 19659 12801 19668 12835
rect 19616 12792 19668 12801
rect 20720 12860 20772 12912
rect 20352 12835 20404 12844
rect 20352 12801 20361 12835
rect 20361 12801 20395 12835
rect 20395 12801 20404 12835
rect 20352 12792 20404 12801
rect 21364 12928 21416 12980
rect 23296 12928 23348 12980
rect 24860 12928 24912 12980
rect 21456 12860 21508 12912
rect 22192 12792 22244 12844
rect 22284 12792 22336 12844
rect 22652 12792 22704 12844
rect 3332 12699 3384 12708
rect 3332 12665 3341 12699
rect 3341 12665 3375 12699
rect 3375 12665 3384 12699
rect 3332 12656 3384 12665
rect 4344 12656 4396 12708
rect 1400 12588 1452 12640
rect 2872 12588 2924 12640
rect 4528 12631 4580 12640
rect 4528 12597 4537 12631
rect 4537 12597 4571 12631
rect 4571 12597 4580 12631
rect 4528 12588 4580 12597
rect 11520 12767 11572 12776
rect 11520 12733 11529 12767
rect 11529 12733 11563 12767
rect 11563 12733 11572 12767
rect 11520 12724 11572 12733
rect 12440 12724 12492 12776
rect 12992 12724 13044 12776
rect 14280 12724 14332 12776
rect 20260 12724 20312 12776
rect 12532 12631 12584 12640
rect 12532 12597 12541 12631
rect 12541 12597 12575 12631
rect 12575 12597 12584 12631
rect 12532 12588 12584 12597
rect 13544 12588 13596 12640
rect 13820 12588 13872 12640
rect 14096 12588 14148 12640
rect 14832 12588 14884 12640
rect 17040 12588 17092 12640
rect 18052 12631 18104 12640
rect 18052 12597 18061 12631
rect 18061 12597 18095 12631
rect 18095 12597 18104 12631
rect 18052 12588 18104 12597
rect 19156 12588 19208 12640
rect 19800 12588 19852 12640
rect 20444 12588 20496 12640
rect 21364 12631 21416 12640
rect 21364 12597 21373 12631
rect 21373 12597 21407 12631
rect 21407 12597 21416 12631
rect 21364 12588 21416 12597
rect 22744 12588 22796 12640
rect 23940 12631 23992 12640
rect 23940 12597 23949 12631
rect 23949 12597 23983 12631
rect 23983 12597 23992 12631
rect 23940 12588 23992 12597
rect 3882 12486 3934 12538
rect 3946 12486 3998 12538
rect 4010 12486 4062 12538
rect 4074 12486 4126 12538
rect 4138 12486 4190 12538
rect 9747 12486 9799 12538
rect 9811 12486 9863 12538
rect 9875 12486 9927 12538
rect 9939 12486 9991 12538
rect 10003 12486 10055 12538
rect 15612 12486 15664 12538
rect 15676 12486 15728 12538
rect 15740 12486 15792 12538
rect 15804 12486 15856 12538
rect 15868 12486 15920 12538
rect 21477 12486 21529 12538
rect 21541 12486 21593 12538
rect 21605 12486 21657 12538
rect 21669 12486 21721 12538
rect 21733 12486 21785 12538
rect 1584 12427 1636 12436
rect 1584 12393 1593 12427
rect 1593 12393 1627 12427
rect 1627 12393 1636 12427
rect 1584 12384 1636 12393
rect 3332 12427 3384 12436
rect 3332 12393 3341 12427
rect 3341 12393 3375 12427
rect 3375 12393 3384 12427
rect 3332 12384 3384 12393
rect 3700 12384 3752 12436
rect 5172 12384 5224 12436
rect 3792 12248 3844 12300
rect 1492 12223 1544 12232
rect 1492 12189 1501 12223
rect 1501 12189 1535 12223
rect 1535 12189 1544 12223
rect 1492 12180 1544 12189
rect 2596 12223 2648 12232
rect 2596 12189 2603 12223
rect 2603 12189 2637 12223
rect 2637 12189 2648 12223
rect 2596 12180 2648 12189
rect 4712 12180 4764 12232
rect 5264 12180 5316 12232
rect 3424 12044 3476 12096
rect 5540 12044 5592 12096
rect 6368 12044 6420 12096
rect 6460 12087 6512 12096
rect 6460 12053 6469 12087
rect 6469 12053 6503 12087
rect 6503 12053 6512 12087
rect 6460 12044 6512 12053
rect 6644 12044 6696 12096
rect 10048 12384 10100 12436
rect 11888 12384 11940 12436
rect 12164 12384 12216 12436
rect 12440 12384 12492 12436
rect 14004 12384 14056 12436
rect 14188 12384 14240 12436
rect 19616 12384 19668 12436
rect 19708 12384 19760 12436
rect 8668 12248 8720 12300
rect 12348 12316 12400 12368
rect 12532 12316 12584 12368
rect 15568 12316 15620 12368
rect 15936 12316 15988 12368
rect 12164 12248 12216 12300
rect 12992 12291 13044 12300
rect 12992 12257 13001 12291
rect 13001 12257 13035 12291
rect 13035 12257 13044 12291
rect 12992 12248 13044 12257
rect 14924 12248 14976 12300
rect 15752 12248 15804 12300
rect 11244 12180 11296 12232
rect 13084 12223 13136 12232
rect 13084 12189 13118 12223
rect 13118 12189 13136 12223
rect 13084 12180 13136 12189
rect 13268 12223 13320 12232
rect 13268 12189 13277 12223
rect 13277 12189 13311 12223
rect 13311 12189 13320 12223
rect 13268 12180 13320 12189
rect 14740 12223 14792 12232
rect 14740 12189 14749 12223
rect 14749 12189 14783 12223
rect 14783 12189 14792 12223
rect 14740 12180 14792 12189
rect 8760 12112 8812 12164
rect 11980 12112 12032 12164
rect 14004 12044 14056 12096
rect 14372 12087 14424 12096
rect 14372 12053 14381 12087
rect 14381 12053 14415 12087
rect 14415 12053 14424 12087
rect 14372 12044 14424 12053
rect 14556 12112 14608 12164
rect 16304 12180 16356 12232
rect 18052 12180 18104 12232
rect 18144 12223 18196 12232
rect 18144 12189 18153 12223
rect 18153 12189 18187 12223
rect 18187 12189 18196 12223
rect 18144 12180 18196 12189
rect 15016 12044 15068 12096
rect 15568 12044 15620 12096
rect 15660 12087 15712 12096
rect 15660 12053 15669 12087
rect 15669 12053 15703 12087
rect 15703 12053 15712 12087
rect 15660 12044 15712 12053
rect 18144 12044 18196 12096
rect 19156 12248 19208 12300
rect 18880 12223 18932 12232
rect 18880 12189 18889 12223
rect 18889 12189 18923 12223
rect 18923 12189 18932 12223
rect 18880 12180 18932 12189
rect 19432 12180 19484 12232
rect 20260 12427 20312 12436
rect 20260 12393 20269 12427
rect 20269 12393 20303 12427
rect 20303 12393 20312 12427
rect 20260 12384 20312 12393
rect 20720 12427 20772 12436
rect 20720 12393 20729 12427
rect 20729 12393 20763 12427
rect 20763 12393 20772 12427
rect 20720 12384 20772 12393
rect 21916 12248 21968 12300
rect 22192 12291 22244 12300
rect 22192 12257 22201 12291
rect 22201 12257 22235 12291
rect 22235 12257 22244 12291
rect 22192 12248 22244 12257
rect 20812 12223 20864 12232
rect 20812 12189 20821 12223
rect 20821 12189 20855 12223
rect 20855 12189 20864 12223
rect 20812 12180 20864 12189
rect 21456 12223 21508 12232
rect 21456 12189 21465 12223
rect 21465 12189 21499 12223
rect 21499 12189 21508 12223
rect 21456 12180 21508 12189
rect 21824 12223 21876 12232
rect 21824 12189 21833 12223
rect 21833 12189 21867 12223
rect 21867 12189 21876 12223
rect 21824 12180 21876 12189
rect 22100 12223 22152 12232
rect 22100 12189 22109 12223
rect 22109 12189 22143 12223
rect 22143 12189 22152 12223
rect 22100 12180 22152 12189
rect 24860 12316 24912 12368
rect 23480 12180 23532 12232
rect 24032 12155 24084 12164
rect 24032 12121 24041 12155
rect 24041 12121 24075 12155
rect 24075 12121 24084 12155
rect 24032 12112 24084 12121
rect 19156 12044 19208 12096
rect 19432 12044 19484 12096
rect 6814 11942 6866 11994
rect 6878 11942 6930 11994
rect 6942 11942 6994 11994
rect 7006 11942 7058 11994
rect 7070 11942 7122 11994
rect 12679 11942 12731 11994
rect 12743 11942 12795 11994
rect 12807 11942 12859 11994
rect 12871 11942 12923 11994
rect 12935 11942 12987 11994
rect 18544 11942 18596 11994
rect 18608 11942 18660 11994
rect 18672 11942 18724 11994
rect 18736 11942 18788 11994
rect 18800 11942 18852 11994
rect 24409 11942 24461 11994
rect 24473 11942 24525 11994
rect 24537 11942 24589 11994
rect 24601 11942 24653 11994
rect 24665 11942 24717 11994
rect 1860 11840 1912 11892
rect 3516 11840 3568 11892
rect 5632 11840 5684 11892
rect 2412 11747 2464 11756
rect 2412 11713 2421 11747
rect 2421 11713 2455 11747
rect 2455 11713 2464 11747
rect 2412 11704 2464 11713
rect 2504 11747 2556 11756
rect 2504 11713 2538 11747
rect 2538 11713 2556 11747
rect 2504 11704 2556 11713
rect 1492 11679 1544 11688
rect 1492 11645 1501 11679
rect 1501 11645 1535 11679
rect 1535 11645 1544 11679
rect 1492 11636 1544 11645
rect 1860 11636 1912 11688
rect 2688 11679 2740 11688
rect 2688 11645 2697 11679
rect 2697 11645 2731 11679
rect 2731 11645 2740 11679
rect 2688 11636 2740 11645
rect 3700 11636 3752 11688
rect 4804 11747 4856 11756
rect 4804 11713 4813 11747
rect 4813 11713 4847 11747
rect 4847 11713 4856 11747
rect 4804 11704 4856 11713
rect 6736 11840 6788 11892
rect 7104 11840 7156 11892
rect 7380 11883 7432 11892
rect 7380 11849 7389 11883
rect 7389 11849 7423 11883
rect 7423 11849 7432 11883
rect 7380 11840 7432 11849
rect 7472 11840 7524 11892
rect 6644 11777 6696 11824
rect 6644 11772 6669 11777
rect 6669 11772 6696 11777
rect 6828 11772 6880 11824
rect 8208 11704 8260 11756
rect 9036 11747 9088 11756
rect 9036 11713 9045 11747
rect 9045 11713 9079 11747
rect 9079 11713 9088 11747
rect 9036 11704 9088 11713
rect 12440 11840 12492 11892
rect 12716 11840 12768 11892
rect 13084 11772 13136 11824
rect 13268 11840 13320 11892
rect 14188 11840 14240 11892
rect 14924 11883 14976 11892
rect 14924 11849 14933 11883
rect 14933 11849 14967 11883
rect 14967 11849 14976 11883
rect 14924 11840 14976 11849
rect 15016 11840 15068 11892
rect 15752 11840 15804 11892
rect 13912 11772 13964 11824
rect 12624 11704 12676 11756
rect 13544 11704 13596 11756
rect 13820 11704 13872 11756
rect 16856 11704 16908 11756
rect 20812 11840 20864 11892
rect 22100 11840 22152 11892
rect 22284 11840 22336 11892
rect 22652 11840 22704 11892
rect 2136 11611 2188 11620
rect 2136 11577 2145 11611
rect 2145 11577 2179 11611
rect 2179 11577 2188 11611
rect 2136 11568 2188 11577
rect 2780 11500 2832 11552
rect 3332 11543 3384 11552
rect 3332 11509 3341 11543
rect 3341 11509 3375 11543
rect 3375 11509 3384 11543
rect 3332 11500 3384 11509
rect 4528 11679 4580 11688
rect 4528 11645 4537 11679
rect 4537 11645 4571 11679
rect 4571 11645 4580 11679
rect 4528 11636 4580 11645
rect 5724 11636 5776 11688
rect 8484 11611 8536 11620
rect 8484 11577 8493 11611
rect 8493 11577 8527 11611
rect 8527 11577 8536 11611
rect 8484 11568 8536 11577
rect 4620 11500 4672 11552
rect 5172 11500 5224 11552
rect 5448 11543 5500 11552
rect 5448 11509 5457 11543
rect 5457 11509 5491 11543
rect 5491 11509 5500 11543
rect 5448 11500 5500 11509
rect 7932 11500 7984 11552
rect 8300 11500 8352 11552
rect 9588 11636 9640 11688
rect 11520 11636 11572 11688
rect 13268 11636 13320 11688
rect 17960 11704 18012 11756
rect 18144 11704 18196 11756
rect 18788 11704 18840 11756
rect 24308 11772 24360 11824
rect 19708 11704 19760 11756
rect 9496 11500 9548 11552
rect 11980 11500 12032 11552
rect 12900 11500 12952 11552
rect 14280 11500 14332 11552
rect 14924 11500 14976 11552
rect 17316 11500 17368 11552
rect 18788 11611 18840 11620
rect 18788 11577 18797 11611
rect 18797 11577 18831 11611
rect 18831 11577 18840 11611
rect 18788 11568 18840 11577
rect 21456 11704 21508 11756
rect 22376 11747 22428 11756
rect 22376 11713 22385 11747
rect 22385 11713 22419 11747
rect 22419 11713 22428 11747
rect 22376 11704 22428 11713
rect 21088 11500 21140 11552
rect 22652 11636 22704 11688
rect 23848 11543 23900 11552
rect 23848 11509 23857 11543
rect 23857 11509 23891 11543
rect 23891 11509 23900 11543
rect 23848 11500 23900 11509
rect 3882 11398 3934 11450
rect 3946 11398 3998 11450
rect 4010 11398 4062 11450
rect 4074 11398 4126 11450
rect 4138 11398 4190 11450
rect 9747 11398 9799 11450
rect 9811 11398 9863 11450
rect 9875 11398 9927 11450
rect 9939 11398 9991 11450
rect 10003 11398 10055 11450
rect 15612 11398 15664 11450
rect 15676 11398 15728 11450
rect 15740 11398 15792 11450
rect 15804 11398 15856 11450
rect 15868 11398 15920 11450
rect 21477 11398 21529 11450
rect 21541 11398 21593 11450
rect 21605 11398 21657 11450
rect 21669 11398 21721 11450
rect 21733 11398 21785 11450
rect 1308 11296 1360 11348
rect 2688 11339 2740 11348
rect 2688 11305 2697 11339
rect 2697 11305 2731 11339
rect 2731 11305 2740 11339
rect 2688 11296 2740 11305
rect 3608 11296 3660 11348
rect 5540 11296 5592 11348
rect 2504 11160 2556 11212
rect 3608 11160 3660 11212
rect 2320 11092 2372 11144
rect 3148 11092 3200 11144
rect 4252 11024 4304 11076
rect 5448 11160 5500 11212
rect 5724 11203 5776 11212
rect 5724 11169 5733 11203
rect 5733 11169 5767 11203
rect 5767 11169 5776 11203
rect 5724 11160 5776 11169
rect 6092 11203 6144 11212
rect 6092 11169 6126 11203
rect 6126 11169 6144 11203
rect 6092 11160 6144 11169
rect 6460 11160 6512 11212
rect 6644 11160 6696 11212
rect 8300 11296 8352 11348
rect 8484 11339 8536 11348
rect 8484 11305 8493 11339
rect 8493 11305 8527 11339
rect 8527 11305 8536 11339
rect 8484 11296 8536 11305
rect 9036 11296 9088 11348
rect 10692 11296 10744 11348
rect 12440 11296 12492 11348
rect 14924 11296 14976 11348
rect 16304 11296 16356 11348
rect 16856 11296 16908 11348
rect 12072 11228 12124 11280
rect 14556 11228 14608 11280
rect 14648 11228 14700 11280
rect 18052 11339 18104 11348
rect 18052 11305 18061 11339
rect 18061 11305 18095 11339
rect 18095 11305 18104 11339
rect 18052 11296 18104 11305
rect 18880 11296 18932 11348
rect 22376 11296 22428 11348
rect 7104 11160 7156 11212
rect 5172 11092 5224 11144
rect 7840 11092 7892 11144
rect 10232 11160 10284 11212
rect 8576 11092 8628 11144
rect 8760 11092 8812 11144
rect 10140 11092 10192 11144
rect 10968 11160 11020 11212
rect 11060 11203 11112 11212
rect 11060 11169 11069 11203
rect 11069 11169 11103 11203
rect 11103 11169 11112 11203
rect 11060 11160 11112 11169
rect 11336 11135 11388 11144
rect 11336 11101 11345 11135
rect 11345 11101 11379 11135
rect 11379 11101 11388 11135
rect 11336 11092 11388 11101
rect 11612 11135 11664 11144
rect 11612 11101 11621 11135
rect 11621 11101 11655 11135
rect 11655 11101 11664 11135
rect 11612 11092 11664 11101
rect 14280 11160 14332 11212
rect 15936 11160 15988 11212
rect 16304 11203 16356 11212
rect 16304 11169 16313 11203
rect 16313 11169 16347 11203
rect 16347 11169 16356 11203
rect 16304 11160 16356 11169
rect 17408 11160 17460 11212
rect 19800 11203 19852 11212
rect 12348 11092 12400 11144
rect 12900 11092 12952 11144
rect 15016 11092 15068 11144
rect 1952 10956 2004 11008
rect 3148 10956 3200 11008
rect 3884 10956 3936 11008
rect 3976 10999 4028 11008
rect 3976 10965 3985 10999
rect 3985 10965 4019 10999
rect 4019 10965 4028 10999
rect 3976 10956 4028 10965
rect 4344 10956 4396 11008
rect 6092 10956 6144 11008
rect 16580 11135 16632 11144
rect 16580 11101 16589 11135
rect 16589 11101 16623 11135
rect 16623 11101 16632 11135
rect 16580 11092 16632 11101
rect 16856 11135 16908 11144
rect 16856 11101 16865 11135
rect 16865 11101 16899 11135
rect 16899 11101 16908 11135
rect 16856 11092 16908 11101
rect 17408 11024 17460 11076
rect 18236 11024 18288 11076
rect 18880 11024 18932 11076
rect 13268 10956 13320 11008
rect 15844 10956 15896 11008
rect 16948 10956 17000 11008
rect 18052 10956 18104 11008
rect 19800 11169 19809 11203
rect 19809 11169 19843 11203
rect 19843 11169 19852 11203
rect 19800 11160 19852 11169
rect 22560 11160 22612 11212
rect 22744 11203 22796 11212
rect 22744 11169 22753 11203
rect 22753 11169 22787 11203
rect 22787 11169 22796 11203
rect 22744 11160 22796 11169
rect 19708 11135 19760 11144
rect 19708 11101 19717 11135
rect 19717 11101 19751 11135
rect 19751 11101 19760 11135
rect 19708 11092 19760 11101
rect 20076 11135 20128 11144
rect 20076 11101 20085 11135
rect 20085 11101 20128 11135
rect 20076 11092 20128 11101
rect 21272 11092 21324 11144
rect 22928 11092 22980 11144
rect 22560 11024 22612 11076
rect 23204 11024 23256 11076
rect 20352 10956 20404 11008
rect 20812 10999 20864 11008
rect 20812 10965 20821 10999
rect 20821 10965 20855 10999
rect 20855 10965 20864 10999
rect 20812 10956 20864 10965
rect 20996 10956 21048 11008
rect 22376 10956 22428 11008
rect 6814 10854 6866 10906
rect 6878 10854 6930 10906
rect 6942 10854 6994 10906
rect 7006 10854 7058 10906
rect 7070 10854 7122 10906
rect 12679 10854 12731 10906
rect 12743 10854 12795 10906
rect 12807 10854 12859 10906
rect 12871 10854 12923 10906
rect 12935 10854 12987 10906
rect 18544 10854 18596 10906
rect 18608 10854 18660 10906
rect 18672 10854 18724 10906
rect 18736 10854 18788 10906
rect 18800 10854 18852 10906
rect 24409 10854 24461 10906
rect 24473 10854 24525 10906
rect 24537 10854 24589 10906
rect 24601 10854 24653 10906
rect 24665 10854 24717 10906
rect 664 10752 716 10804
rect 2780 10752 2832 10804
rect 2228 10659 2280 10668
rect 2228 10625 2235 10659
rect 2235 10625 2269 10659
rect 2269 10625 2280 10659
rect 2228 10616 2280 10625
rect 2412 10684 2464 10736
rect 4160 10752 4212 10804
rect 4804 10752 4856 10804
rect 5724 10795 5776 10804
rect 5724 10761 5733 10795
rect 5733 10761 5767 10795
rect 5767 10761 5776 10795
rect 5724 10752 5776 10761
rect 11060 10795 11112 10804
rect 11060 10761 11069 10795
rect 11069 10761 11103 10795
rect 11103 10761 11112 10795
rect 11060 10752 11112 10761
rect 11612 10752 11664 10804
rect 3148 10616 3200 10668
rect 3884 10684 3936 10736
rect 5264 10684 5316 10736
rect 4896 10616 4948 10668
rect 7104 10616 7156 10668
rect 7932 10616 7984 10668
rect 7380 10548 7432 10600
rect 10324 10659 10376 10668
rect 10324 10625 10331 10659
rect 10331 10625 10365 10659
rect 10365 10625 10376 10659
rect 10324 10616 10376 10625
rect 10968 10616 11020 10668
rect 11520 10684 11572 10736
rect 11244 10616 11296 10668
rect 12164 10616 12216 10668
rect 13912 10684 13964 10736
rect 13820 10616 13872 10668
rect 15200 10684 15252 10736
rect 16304 10752 16356 10804
rect 16856 10752 16908 10804
rect 21824 10752 21876 10804
rect 23848 10752 23900 10804
rect 18328 10684 18380 10736
rect 22468 10684 22520 10736
rect 22744 10684 22796 10736
rect 23112 10684 23164 10736
rect 16948 10659 17000 10668
rect 16948 10625 16955 10659
rect 16955 10625 16989 10659
rect 16989 10625 17000 10659
rect 16948 10616 17000 10625
rect 7012 10480 7064 10532
rect 7472 10480 7524 10532
rect 8760 10412 8812 10464
rect 13268 10480 13320 10532
rect 13452 10480 13504 10532
rect 14924 10480 14976 10532
rect 19432 10480 19484 10532
rect 21824 10480 21876 10532
rect 22560 10616 22612 10668
rect 22836 10616 22888 10668
rect 14464 10455 14516 10464
rect 14464 10421 14473 10455
rect 14473 10421 14507 10455
rect 14507 10421 14516 10455
rect 14464 10412 14516 10421
rect 14740 10412 14792 10464
rect 16948 10412 17000 10464
rect 22652 10412 22704 10464
rect 24032 10455 24084 10464
rect 24032 10421 24041 10455
rect 24041 10421 24075 10455
rect 24075 10421 24084 10455
rect 24032 10412 24084 10421
rect 3882 10310 3934 10362
rect 3946 10310 3998 10362
rect 4010 10310 4062 10362
rect 4074 10310 4126 10362
rect 4138 10310 4190 10362
rect 9747 10310 9799 10362
rect 9811 10310 9863 10362
rect 9875 10310 9927 10362
rect 9939 10310 9991 10362
rect 10003 10310 10055 10362
rect 15612 10310 15664 10362
rect 15676 10310 15728 10362
rect 15740 10310 15792 10362
rect 15804 10310 15856 10362
rect 15868 10310 15920 10362
rect 21477 10310 21529 10362
rect 21541 10310 21593 10362
rect 21605 10310 21657 10362
rect 21669 10310 21721 10362
rect 21733 10310 21785 10362
rect 2136 10208 2188 10260
rect 2872 10208 2924 10260
rect 2964 10251 3016 10260
rect 2964 10217 2973 10251
rect 2973 10217 3007 10251
rect 3007 10217 3016 10251
rect 2964 10208 3016 10217
rect 3608 10208 3660 10260
rect 3700 10140 3752 10192
rect 8484 10208 8536 10260
rect 8760 10251 8812 10260
rect 8760 10217 8769 10251
rect 8769 10217 8803 10251
rect 8803 10217 8812 10251
rect 8760 10208 8812 10217
rect 9220 10208 9272 10260
rect 11980 10208 12032 10260
rect 14464 10208 14516 10260
rect 4344 10072 4396 10124
rect 7012 10072 7064 10124
rect 7104 10115 7156 10124
rect 7104 10081 7113 10115
rect 7113 10081 7147 10115
rect 7147 10081 7156 10115
rect 7104 10072 7156 10081
rect 14556 10140 14608 10192
rect 8300 10072 8352 10124
rect 12440 10072 12492 10124
rect 14280 10115 14332 10124
rect 14280 10081 14289 10115
rect 14289 10081 14323 10115
rect 14323 10081 14332 10115
rect 14280 10072 14332 10081
rect 14740 10208 14792 10260
rect 15752 10140 15804 10192
rect 20812 10115 20864 10124
rect 20812 10081 20821 10115
rect 20821 10081 20855 10115
rect 20855 10081 20864 10115
rect 20812 10072 20864 10081
rect 22376 10072 22428 10124
rect 3240 10004 3292 10056
rect 1952 9936 2004 9988
rect 3792 9936 3844 9988
rect 5632 10004 5684 10056
rect 6460 10004 6512 10056
rect 7288 10004 7340 10056
rect 8024 10004 8076 10056
rect 8760 10004 8812 10056
rect 4160 9868 4212 9920
rect 10508 9936 10560 9988
rect 11888 9936 11940 9988
rect 12072 9936 12124 9988
rect 9496 9868 9548 9920
rect 12624 10004 12676 10056
rect 13360 10004 13412 10056
rect 14464 10004 14516 10056
rect 15016 10047 15068 10056
rect 15016 10013 15025 10047
rect 15025 10013 15059 10047
rect 15059 10013 15068 10047
rect 15016 10004 15068 10013
rect 15200 10004 15252 10056
rect 15292 10047 15344 10056
rect 15292 10013 15301 10047
rect 15301 10013 15335 10047
rect 15335 10013 15344 10047
rect 15292 10004 15344 10013
rect 18144 10004 18196 10056
rect 18236 10047 18288 10056
rect 18236 10013 18245 10047
rect 18245 10013 18279 10047
rect 18279 10013 18288 10047
rect 18236 10004 18288 10013
rect 18328 10004 18380 10056
rect 12532 9979 12584 9988
rect 12532 9945 12541 9979
rect 12541 9945 12575 9979
rect 12575 9945 12584 9979
rect 12532 9936 12584 9945
rect 13084 9936 13136 9988
rect 14188 9936 14240 9988
rect 13268 9911 13320 9920
rect 13268 9877 13281 9911
rect 13281 9877 13315 9911
rect 13315 9877 13320 9911
rect 13268 9868 13320 9877
rect 15016 9868 15068 9920
rect 16488 9936 16540 9988
rect 19984 10047 20036 10056
rect 19984 10013 19993 10047
rect 19993 10013 20027 10047
rect 20027 10013 20036 10047
rect 19984 10004 20036 10013
rect 20904 10047 20956 10056
rect 20904 10013 20913 10047
rect 20913 10013 20947 10047
rect 20947 10013 20956 10047
rect 20904 10004 20956 10013
rect 22652 10004 22704 10056
rect 21548 9936 21600 9988
rect 24860 10208 24912 10260
rect 24032 10004 24084 10056
rect 25136 10004 25188 10056
rect 24860 9936 24912 9988
rect 15936 9911 15988 9920
rect 15936 9877 15945 9911
rect 15945 9877 15979 9911
rect 15979 9877 15988 9911
rect 15936 9868 15988 9877
rect 17224 9868 17276 9920
rect 18972 9868 19024 9920
rect 19800 9868 19852 9920
rect 20720 9868 20772 9920
rect 6814 9766 6866 9818
rect 6878 9766 6930 9818
rect 6942 9766 6994 9818
rect 7006 9766 7058 9818
rect 7070 9766 7122 9818
rect 12679 9766 12731 9818
rect 12743 9766 12795 9818
rect 12807 9766 12859 9818
rect 12871 9766 12923 9818
rect 12935 9766 12987 9818
rect 18544 9766 18596 9818
rect 18608 9766 18660 9818
rect 18672 9766 18724 9818
rect 18736 9766 18788 9818
rect 18800 9766 18852 9818
rect 24409 9766 24461 9818
rect 24473 9766 24525 9818
rect 24537 9766 24589 9818
rect 24601 9766 24653 9818
rect 24665 9766 24717 9818
rect 1768 9707 1820 9716
rect 1768 9673 1777 9707
rect 1777 9673 1811 9707
rect 1811 9673 1820 9707
rect 1768 9664 1820 9673
rect 2872 9664 2924 9716
rect 3240 9664 3292 9716
rect 3516 9664 3568 9716
rect 4068 9664 4120 9716
rect 5540 9664 5592 9716
rect 7380 9664 7432 9716
rect 8024 9664 8076 9716
rect 8208 9664 8260 9716
rect 8300 9707 8352 9716
rect 8300 9673 8309 9707
rect 8309 9673 8343 9707
rect 8343 9673 8352 9707
rect 8300 9664 8352 9673
rect 756 9596 808 9648
rect 2136 9528 2188 9580
rect 5264 9596 5316 9648
rect 6552 9596 6604 9648
rect 3608 9571 3660 9580
rect 3608 9537 3617 9571
rect 3617 9537 3651 9571
rect 3651 9537 3660 9571
rect 3608 9528 3660 9537
rect 4528 9528 4580 9580
rect 2320 9460 2372 9512
rect 2780 9460 2832 9512
rect 3516 9460 3568 9512
rect 2872 9392 2924 9444
rect 3056 9435 3108 9444
rect 3056 9401 3065 9435
rect 3065 9401 3099 9435
rect 3099 9401 3108 9435
rect 3056 9392 3108 9401
rect 4344 9324 4396 9376
rect 4896 9503 4948 9512
rect 4896 9469 4905 9503
rect 4905 9469 4939 9503
rect 4939 9469 4948 9503
rect 4896 9460 4948 9469
rect 5632 9460 5684 9512
rect 6736 9460 6788 9512
rect 4804 9392 4856 9444
rect 6184 9392 6236 9444
rect 5908 9367 5960 9376
rect 5908 9333 5917 9367
rect 5917 9333 5951 9367
rect 5951 9333 5960 9367
rect 5908 9324 5960 9333
rect 12532 9664 12584 9716
rect 14004 9664 14056 9716
rect 15016 9664 15068 9716
rect 15292 9664 15344 9716
rect 17868 9664 17920 9716
rect 20628 9664 20680 9716
rect 20812 9664 20864 9716
rect 20904 9664 20956 9716
rect 21548 9707 21600 9716
rect 21548 9673 21557 9707
rect 21557 9673 21591 9707
rect 21591 9673 21600 9707
rect 21548 9664 21600 9673
rect 21824 9664 21876 9716
rect 23940 9664 23992 9716
rect 9220 9596 9272 9648
rect 9404 9596 9456 9648
rect 10324 9596 10376 9648
rect 10600 9639 10652 9648
rect 10600 9605 10609 9639
rect 10609 9605 10643 9639
rect 10643 9605 10652 9639
rect 10600 9596 10652 9605
rect 7564 9571 7616 9580
rect 7564 9537 7571 9571
rect 7571 9537 7605 9571
rect 7605 9537 7616 9571
rect 7564 9528 7616 9537
rect 10140 9528 10192 9580
rect 10232 9571 10284 9580
rect 10232 9537 10241 9571
rect 10241 9537 10275 9571
rect 10275 9537 10284 9571
rect 10232 9528 10284 9537
rect 14556 9596 14608 9648
rect 16028 9596 16080 9648
rect 16488 9596 16540 9648
rect 18052 9596 18104 9648
rect 13912 9528 13964 9580
rect 14372 9571 14424 9580
rect 14372 9537 14379 9571
rect 14379 9537 14413 9571
rect 14413 9537 14424 9571
rect 14372 9528 14424 9537
rect 15016 9528 15068 9580
rect 9496 9460 9548 9512
rect 11428 9460 11480 9512
rect 15108 9460 15160 9512
rect 15384 9460 15436 9512
rect 15844 9460 15896 9512
rect 16028 9460 16080 9512
rect 17316 9571 17368 9580
rect 17316 9537 17323 9571
rect 17323 9537 17357 9571
rect 17357 9537 17368 9571
rect 17316 9528 17368 9537
rect 17684 9528 17736 9580
rect 17960 9528 18012 9580
rect 19156 9596 19208 9648
rect 19432 9528 19484 9580
rect 19616 9528 19668 9580
rect 20720 9528 20772 9580
rect 21180 9571 21232 9580
rect 21180 9537 21189 9571
rect 21189 9537 21223 9571
rect 21223 9537 21232 9571
rect 21180 9528 21232 9537
rect 16856 9460 16908 9512
rect 18604 9503 18656 9512
rect 7656 9324 7708 9376
rect 10692 9324 10744 9376
rect 14924 9324 14976 9376
rect 16488 9324 16540 9376
rect 17408 9324 17460 9376
rect 18604 9469 18613 9503
rect 18613 9469 18647 9503
rect 18647 9469 18656 9503
rect 18604 9460 18656 9469
rect 19800 9460 19852 9512
rect 20260 9460 20312 9512
rect 18144 9324 18196 9376
rect 18512 9324 18564 9376
rect 22008 9571 22060 9580
rect 22008 9537 22017 9571
rect 22017 9537 22051 9571
rect 22051 9537 22060 9571
rect 22008 9528 22060 9537
rect 22744 9460 22796 9512
rect 23848 9367 23900 9376
rect 23848 9333 23857 9367
rect 23857 9333 23891 9367
rect 23891 9333 23900 9367
rect 23848 9324 23900 9333
rect 3882 9222 3934 9274
rect 3946 9222 3998 9274
rect 4010 9222 4062 9274
rect 4074 9222 4126 9274
rect 4138 9222 4190 9274
rect 9747 9222 9799 9274
rect 9811 9222 9863 9274
rect 9875 9222 9927 9274
rect 9939 9222 9991 9274
rect 10003 9222 10055 9274
rect 15612 9222 15664 9274
rect 15676 9222 15728 9274
rect 15740 9222 15792 9274
rect 15804 9222 15856 9274
rect 15868 9222 15920 9274
rect 21477 9222 21529 9274
rect 21541 9222 21593 9274
rect 21605 9222 21657 9274
rect 21669 9222 21721 9274
rect 21733 9222 21785 9274
rect 3056 9120 3108 9172
rect 3792 9120 3844 9172
rect 4896 9052 4948 9104
rect 5724 9052 5776 9104
rect 5632 8984 5684 9036
rect 5908 9120 5960 9172
rect 6092 9120 6144 9172
rect 8484 9163 8536 9172
rect 8484 9129 8493 9163
rect 8493 9129 8527 9163
rect 8527 9129 8536 9163
rect 8484 9120 8536 9129
rect 10048 9120 10100 9172
rect 10324 9120 10376 9172
rect 10508 9052 10560 9104
rect 12440 9163 12492 9172
rect 12440 9129 12449 9163
rect 12449 9129 12483 9163
rect 12483 9129 12492 9163
rect 12440 9120 12492 9129
rect 15108 9052 15160 9104
rect 8484 8984 8536 9036
rect 11428 9027 11480 9036
rect 11428 8993 11437 9027
rect 11437 8993 11471 9027
rect 11471 8993 11480 9027
rect 11428 8984 11480 8993
rect 16212 9052 16264 9104
rect 17592 9120 17644 9172
rect 20260 9120 20312 9172
rect 20536 9120 20588 9172
rect 18604 9052 18656 9104
rect 19156 9052 19208 9104
rect 22008 9120 22060 9172
rect 23848 9120 23900 9172
rect 24124 9163 24176 9172
rect 24124 9129 24133 9163
rect 24133 9129 24167 9163
rect 24167 9129 24176 9163
rect 24124 9120 24176 9129
rect 22744 9052 22796 9104
rect 16304 9027 16356 9036
rect 16304 8993 16313 9027
rect 16313 8993 16347 9027
rect 16347 8993 16356 9027
rect 16304 8984 16356 8993
rect 16396 8984 16448 9036
rect 16764 8984 16816 9036
rect 1860 8959 1912 8968
rect 1860 8925 1869 8959
rect 1869 8925 1903 8959
rect 1903 8925 1912 8959
rect 1860 8916 1912 8925
rect 2228 8916 2280 8968
rect 3332 8916 3384 8968
rect 4068 8916 4120 8968
rect 4436 8959 4488 8968
rect 3056 8848 3108 8900
rect 3516 8848 3568 8900
rect 4436 8925 4443 8959
rect 4443 8925 4477 8959
rect 4477 8925 4488 8959
rect 4436 8916 4488 8925
rect 22100 8984 22152 9036
rect 5908 8916 5960 8968
rect 6460 8959 6512 8968
rect 6460 8925 6469 8959
rect 6469 8925 6503 8959
rect 6503 8925 6512 8959
rect 6460 8916 6512 8925
rect 6552 8959 6604 8968
rect 6552 8925 6586 8959
rect 6586 8925 6604 8959
rect 6552 8916 6604 8925
rect 6736 8959 6788 8968
rect 6736 8925 6745 8959
rect 6745 8925 6779 8959
rect 6779 8925 6788 8959
rect 6736 8916 6788 8925
rect 7656 8916 7708 8968
rect 8760 8916 8812 8968
rect 2044 8780 2096 8832
rect 2780 8780 2832 8832
rect 4252 8780 4304 8832
rect 4528 8780 4580 8832
rect 5080 8780 5132 8832
rect 7380 8848 7432 8900
rect 12348 8916 12400 8968
rect 14832 8916 14884 8968
rect 14924 8916 14976 8968
rect 16856 8959 16908 8968
rect 16856 8925 16865 8959
rect 16865 8925 16899 8959
rect 16899 8925 16908 8959
rect 16856 8916 16908 8925
rect 17500 8916 17552 8968
rect 17684 8916 17736 8968
rect 21272 8916 21324 8968
rect 22192 8916 22244 8968
rect 22284 8959 22336 8968
rect 22284 8925 22293 8959
rect 22293 8925 22327 8959
rect 22327 8925 22336 8959
rect 22284 8916 22336 8925
rect 23020 8959 23072 8968
rect 23020 8925 23029 8959
rect 23029 8925 23063 8959
rect 23063 8925 23072 8959
rect 23020 8916 23072 8925
rect 15200 8848 15252 8900
rect 19340 8848 19392 8900
rect 10324 8780 10376 8832
rect 11152 8780 11204 8832
rect 14464 8780 14516 8832
rect 16396 8780 16448 8832
rect 19156 8780 19208 8832
rect 19708 8848 19760 8900
rect 20996 8891 21048 8900
rect 19892 8780 19944 8832
rect 20628 8823 20680 8832
rect 20628 8789 20637 8823
rect 20637 8789 20671 8823
rect 20671 8789 20680 8823
rect 20628 8780 20680 8789
rect 20996 8857 21030 8891
rect 21030 8857 21048 8891
rect 20996 8848 21048 8857
rect 23572 8959 23624 8968
rect 23572 8925 23581 8959
rect 23581 8925 23615 8959
rect 23615 8925 23624 8959
rect 23572 8916 23624 8925
rect 23388 8823 23440 8832
rect 23388 8789 23397 8823
rect 23397 8789 23431 8823
rect 23431 8789 23440 8823
rect 23388 8780 23440 8789
rect 6814 8678 6866 8730
rect 6878 8678 6930 8730
rect 6942 8678 6994 8730
rect 7006 8678 7058 8730
rect 7070 8678 7122 8730
rect 12679 8678 12731 8730
rect 12743 8678 12795 8730
rect 12807 8678 12859 8730
rect 12871 8678 12923 8730
rect 12935 8678 12987 8730
rect 18544 8678 18596 8730
rect 18608 8678 18660 8730
rect 18672 8678 18724 8730
rect 18736 8678 18788 8730
rect 18800 8678 18852 8730
rect 24409 8678 24461 8730
rect 24473 8678 24525 8730
rect 24537 8678 24589 8730
rect 24601 8678 24653 8730
rect 24665 8678 24717 8730
rect 2320 8576 2372 8628
rect 6736 8576 6788 8628
rect 7656 8576 7708 8628
rect 11244 8576 11296 8628
rect 11336 8576 11388 8628
rect 13268 8576 13320 8628
rect 16764 8576 16816 8628
rect 16856 8576 16908 8628
rect 18236 8576 18288 8628
rect 18328 8576 18380 8628
rect 19616 8619 19668 8628
rect 19616 8585 19625 8619
rect 19625 8585 19659 8619
rect 19659 8585 19668 8619
rect 19616 8576 19668 8585
rect 19708 8576 19760 8628
rect 19984 8576 20036 8628
rect 20628 8576 20680 8628
rect 21180 8576 21232 8628
rect 23756 8619 23808 8628
rect 23756 8585 23765 8619
rect 23765 8585 23799 8619
rect 23799 8585 23808 8619
rect 23756 8576 23808 8585
rect 3240 8508 3292 8560
rect 1676 8483 1728 8492
rect 1676 8449 1685 8483
rect 1685 8449 1719 8483
rect 1719 8449 1728 8483
rect 1676 8440 1728 8449
rect 1308 8372 1360 8424
rect 1492 8415 1544 8424
rect 1492 8381 1501 8415
rect 1501 8381 1535 8415
rect 1535 8381 1544 8415
rect 1492 8372 1544 8381
rect 2044 8372 2096 8424
rect 2688 8483 2740 8492
rect 2688 8449 2697 8483
rect 2697 8449 2731 8483
rect 2731 8449 2740 8483
rect 2688 8440 2740 8449
rect 3700 8440 3752 8492
rect 5080 8483 5132 8492
rect 5080 8449 5089 8483
rect 5089 8449 5123 8483
rect 5123 8449 5132 8483
rect 5080 8440 5132 8449
rect 6000 8440 6052 8492
rect 10048 8508 10100 8560
rect 7564 8440 7616 8492
rect 8392 8440 8444 8492
rect 8852 8440 8904 8492
rect 10600 8440 10652 8492
rect 10968 8440 11020 8492
rect 15476 8483 15528 8492
rect 15476 8449 15483 8483
rect 15483 8449 15517 8483
rect 15517 8449 15528 8483
rect 15476 8440 15528 8449
rect 17316 8440 17368 8492
rect 3056 8372 3108 8424
rect 3792 8372 3844 8424
rect 4620 8372 4672 8424
rect 4896 8372 4948 8424
rect 6184 8372 6236 8424
rect 7380 8372 7432 8424
rect 14740 8372 14792 8424
rect 2136 8347 2188 8356
rect 2136 8313 2145 8347
rect 2145 8313 2179 8347
rect 2179 8313 2188 8347
rect 2136 8304 2188 8313
rect 2044 8236 2096 8288
rect 3884 8304 3936 8356
rect 4528 8347 4580 8356
rect 4528 8313 4537 8347
rect 4537 8313 4571 8347
rect 4571 8313 4580 8347
rect 4528 8304 4580 8313
rect 5724 8304 5776 8356
rect 4068 8236 4120 8288
rect 4988 8236 5040 8288
rect 5908 8236 5960 8288
rect 7656 8236 7708 8288
rect 7840 8236 7892 8288
rect 11060 8304 11112 8356
rect 8944 8236 8996 8288
rect 16304 8236 16356 8288
rect 18144 8440 18196 8492
rect 19156 8440 19208 8492
rect 19340 8372 19392 8424
rect 17868 8236 17920 8288
rect 19892 8440 19944 8492
rect 23204 8508 23256 8560
rect 20996 8483 21048 8492
rect 20996 8449 21005 8483
rect 21005 8449 21039 8483
rect 21039 8449 21048 8483
rect 20996 8440 21048 8449
rect 20720 8372 20772 8424
rect 22008 8481 22060 8492
rect 22008 8447 22017 8481
rect 22017 8447 22051 8481
rect 22051 8447 22060 8481
rect 22008 8440 22060 8447
rect 22376 8440 22428 8492
rect 22100 8415 22152 8424
rect 22100 8381 22109 8415
rect 22109 8381 22143 8415
rect 22143 8381 22152 8415
rect 22100 8372 22152 8381
rect 22192 8372 22244 8424
rect 21824 8304 21876 8356
rect 24216 8483 24268 8492
rect 24216 8449 24225 8483
rect 24225 8449 24259 8483
rect 24259 8449 24268 8483
rect 24216 8440 24268 8449
rect 3882 8134 3934 8186
rect 3946 8134 3998 8186
rect 4010 8134 4062 8186
rect 4074 8134 4126 8186
rect 4138 8134 4190 8186
rect 9747 8134 9799 8186
rect 9811 8134 9863 8186
rect 9875 8134 9927 8186
rect 9939 8134 9991 8186
rect 10003 8134 10055 8186
rect 15612 8134 15664 8186
rect 15676 8134 15728 8186
rect 15740 8134 15792 8186
rect 15804 8134 15856 8186
rect 15868 8134 15920 8186
rect 21477 8134 21529 8186
rect 21541 8134 21593 8186
rect 21605 8134 21657 8186
rect 21669 8134 21721 8186
rect 21733 8134 21785 8186
rect 1860 8032 1912 8084
rect 1952 8075 2004 8084
rect 1952 8041 1961 8075
rect 1961 8041 1995 8075
rect 1995 8041 2004 8075
rect 1952 8032 2004 8041
rect 3608 8032 3660 8084
rect 3608 7896 3660 7948
rect 4252 8032 4304 8084
rect 4528 8032 4580 8084
rect 5540 8032 5592 8084
rect 2504 7828 2556 7880
rect 4068 7871 4120 7880
rect 4068 7837 4075 7871
rect 4075 7837 4109 7871
rect 4109 7837 4120 7871
rect 4068 7828 4120 7837
rect 5172 7828 5224 7880
rect 6092 7828 6144 7880
rect 7380 8032 7432 8084
rect 8668 8032 8720 8084
rect 11336 8032 11388 8084
rect 12164 8032 12216 8084
rect 14004 8032 14056 8084
rect 22192 8032 22244 8084
rect 23020 8032 23072 8084
rect 23756 8032 23808 8084
rect 22284 7964 22336 8016
rect 9864 7896 9916 7948
rect 7656 7828 7708 7880
rect 8760 7828 8812 7880
rect 4344 7760 4396 7812
rect 4436 7760 4488 7812
rect 10600 7828 10652 7880
rect 10968 7939 11020 7948
rect 10968 7905 10977 7939
rect 10977 7905 11011 7939
rect 11011 7905 11020 7939
rect 10968 7896 11020 7905
rect 13544 7896 13596 7948
rect 22560 7964 22612 8016
rect 10324 7760 10376 7812
rect 11796 7760 11848 7812
rect 4068 7692 4120 7744
rect 6736 7692 6788 7744
rect 8300 7735 8352 7744
rect 8300 7701 8309 7735
rect 8309 7701 8343 7735
rect 8343 7701 8352 7735
rect 8300 7692 8352 7701
rect 8668 7692 8720 7744
rect 9312 7692 9364 7744
rect 9404 7692 9456 7744
rect 9680 7692 9732 7744
rect 10048 7692 10100 7744
rect 11888 7692 11940 7744
rect 12072 7692 12124 7744
rect 12532 7735 12584 7744
rect 12532 7701 12541 7735
rect 12541 7701 12575 7735
rect 12575 7701 12584 7735
rect 12532 7692 12584 7701
rect 13084 7760 13136 7812
rect 13360 7760 13412 7812
rect 13912 7828 13964 7880
rect 14740 7828 14792 7880
rect 15108 7871 15160 7880
rect 15108 7837 15115 7871
rect 15115 7837 15149 7871
rect 15149 7837 15160 7871
rect 15108 7828 15160 7837
rect 15200 7828 15252 7880
rect 16120 7828 16172 7880
rect 19432 7828 19484 7880
rect 13452 7692 13504 7744
rect 13636 7803 13688 7812
rect 13636 7769 13645 7803
rect 13645 7769 13679 7803
rect 13679 7769 13688 7803
rect 13636 7760 13688 7769
rect 21364 7760 21416 7812
rect 23204 7828 23256 7880
rect 23388 7871 23440 7880
rect 23388 7837 23397 7871
rect 23397 7837 23431 7871
rect 23431 7837 23440 7871
rect 23388 7828 23440 7837
rect 23940 7828 23992 7880
rect 24032 7871 24084 7880
rect 24032 7837 24041 7871
rect 24041 7837 24075 7871
rect 24075 7837 24084 7871
rect 24032 7828 24084 7837
rect 25596 7896 25648 7948
rect 14188 7692 14240 7744
rect 15660 7692 15712 7744
rect 16856 7692 16908 7744
rect 17316 7692 17368 7744
rect 23664 7735 23716 7744
rect 23664 7701 23673 7735
rect 23673 7701 23707 7735
rect 23707 7701 23716 7735
rect 23664 7692 23716 7701
rect 25412 7692 25464 7744
rect 6814 7590 6866 7642
rect 6878 7590 6930 7642
rect 6942 7590 6994 7642
rect 7006 7590 7058 7642
rect 7070 7590 7122 7642
rect 12679 7590 12731 7642
rect 12743 7590 12795 7642
rect 12807 7590 12859 7642
rect 12871 7590 12923 7642
rect 12935 7590 12987 7642
rect 18544 7590 18596 7642
rect 18608 7590 18660 7642
rect 18672 7590 18724 7642
rect 18736 7590 18788 7642
rect 18800 7590 18852 7642
rect 24409 7590 24461 7642
rect 24473 7590 24525 7642
rect 24537 7590 24589 7642
rect 24601 7590 24653 7642
rect 24665 7590 24717 7642
rect 1768 7488 1820 7540
rect 2688 7488 2740 7540
rect 1400 7352 1452 7404
rect 3148 7420 3200 7472
rect 3516 7352 3568 7404
rect 4068 7488 4120 7540
rect 7380 7488 7432 7540
rect 4160 7420 4212 7472
rect 4528 7420 4580 7472
rect 7472 7420 7524 7472
rect 9588 7420 9640 7472
rect 9680 7420 9732 7472
rect 4252 7352 4304 7404
rect 4988 7352 5040 7404
rect 5448 7352 5500 7404
rect 6368 7352 6420 7404
rect 7564 7352 7616 7404
rect 8668 7395 8720 7404
rect 8668 7361 8677 7395
rect 8677 7361 8711 7395
rect 8711 7361 8720 7395
rect 8668 7352 8720 7361
rect 8944 7395 8996 7404
rect 8944 7361 8953 7395
rect 8953 7361 8987 7395
rect 8987 7361 8996 7395
rect 8944 7352 8996 7361
rect 4068 7216 4120 7268
rect 4344 7148 4396 7200
rect 4712 7191 4764 7200
rect 4712 7157 4721 7191
rect 4721 7157 4755 7191
rect 4755 7157 4764 7191
rect 4712 7148 4764 7157
rect 7932 7327 7984 7336
rect 7932 7293 7941 7327
rect 7941 7293 7975 7327
rect 7975 7293 7984 7327
rect 7932 7284 7984 7293
rect 8300 7284 8352 7336
rect 10140 7395 10192 7404
rect 10140 7361 10149 7395
rect 10149 7361 10183 7395
rect 10183 7361 10192 7395
rect 10140 7352 10192 7361
rect 10232 7395 10284 7404
rect 10232 7361 10241 7395
rect 10241 7361 10275 7395
rect 10275 7361 10284 7395
rect 10232 7352 10284 7361
rect 10324 7352 10376 7404
rect 10784 7420 10836 7472
rect 11796 7420 11848 7472
rect 12072 7463 12124 7472
rect 12072 7429 12081 7463
rect 12081 7429 12115 7463
rect 12115 7429 12124 7463
rect 12072 7420 12124 7429
rect 12164 7420 12216 7472
rect 12348 7420 12400 7472
rect 12440 7463 12492 7472
rect 12440 7429 12449 7463
rect 12449 7429 12483 7463
rect 12483 7429 12492 7463
rect 12440 7420 12492 7429
rect 12992 7420 13044 7472
rect 10048 7284 10100 7336
rect 13084 7352 13136 7404
rect 11888 7284 11940 7336
rect 6276 7148 6328 7200
rect 7564 7148 7616 7200
rect 13452 7488 13504 7540
rect 16580 7488 16632 7540
rect 17776 7488 17828 7540
rect 20628 7488 20680 7540
rect 21180 7488 21232 7540
rect 24032 7488 24084 7540
rect 16396 7420 16448 7472
rect 13636 7216 13688 7268
rect 13268 7148 13320 7200
rect 14280 7352 14332 7404
rect 15660 7395 15712 7404
rect 15660 7361 15669 7395
rect 15669 7361 15703 7395
rect 15703 7361 15712 7395
rect 15660 7352 15712 7361
rect 16488 7352 16540 7404
rect 16948 7352 17000 7404
rect 18144 7352 18196 7404
rect 19432 7352 19484 7404
rect 20352 7420 20404 7472
rect 22100 7420 22152 7472
rect 20076 7395 20128 7404
rect 20076 7361 20083 7395
rect 20083 7361 20117 7395
rect 20117 7361 20128 7395
rect 20076 7352 20128 7361
rect 20168 7352 20220 7404
rect 23020 7352 23072 7404
rect 23296 7399 23348 7404
rect 23296 7365 23305 7399
rect 23305 7365 23339 7399
rect 23339 7365 23348 7399
rect 23296 7352 23348 7365
rect 14832 7284 14884 7336
rect 15016 7284 15068 7336
rect 16028 7284 16080 7336
rect 17224 7327 17276 7336
rect 17224 7293 17233 7327
rect 17233 7293 17267 7327
rect 17267 7293 17276 7327
rect 17224 7284 17276 7293
rect 20812 7284 20864 7336
rect 21364 7284 21416 7336
rect 23848 7352 23900 7404
rect 24032 7395 24084 7404
rect 24032 7361 24041 7395
rect 24041 7361 24075 7395
rect 24075 7361 24084 7395
rect 24032 7352 24084 7361
rect 25044 7352 25096 7404
rect 24860 7284 24912 7336
rect 15200 7216 15252 7268
rect 16212 7216 16264 7268
rect 17132 7148 17184 7200
rect 19892 7148 19944 7200
rect 20812 7191 20864 7200
rect 20812 7157 20821 7191
rect 20821 7157 20855 7191
rect 20855 7157 20864 7191
rect 20812 7148 20864 7157
rect 23572 7148 23624 7200
rect 25136 7148 25188 7200
rect 3882 7046 3934 7098
rect 3946 7046 3998 7098
rect 4010 7046 4062 7098
rect 4074 7046 4126 7098
rect 4138 7046 4190 7098
rect 9747 7046 9799 7098
rect 9811 7046 9863 7098
rect 9875 7046 9927 7098
rect 9939 7046 9991 7098
rect 10003 7046 10055 7098
rect 15612 7046 15664 7098
rect 15676 7046 15728 7098
rect 15740 7046 15792 7098
rect 15804 7046 15856 7098
rect 15868 7046 15920 7098
rect 21477 7046 21529 7098
rect 21541 7046 21593 7098
rect 21605 7046 21657 7098
rect 21669 7046 21721 7098
rect 21733 7046 21785 7098
rect 1584 6987 1636 6996
rect 1584 6953 1593 6987
rect 1593 6953 1627 6987
rect 1627 6953 1636 6987
rect 1584 6944 1636 6953
rect 1676 6944 1728 6996
rect 7380 6944 7432 6996
rect 7472 6987 7524 6996
rect 7472 6953 7481 6987
rect 7481 6953 7515 6987
rect 7515 6953 7524 6987
rect 7472 6944 7524 6953
rect 10232 6944 10284 6996
rect 12072 6944 12124 6996
rect 12440 6944 12492 6996
rect 13360 6944 13412 6996
rect 13544 6944 13596 6996
rect 7288 6876 7340 6928
rect 9496 6876 9548 6928
rect 5632 6851 5684 6860
rect 5632 6817 5641 6851
rect 5641 6817 5675 6851
rect 5675 6817 5684 6851
rect 5632 6808 5684 6817
rect 5908 6808 5960 6860
rect 6276 6851 6328 6860
rect 6276 6817 6285 6851
rect 6285 6817 6319 6851
rect 6319 6817 6328 6851
rect 6276 6808 6328 6817
rect 6644 6851 6696 6860
rect 6644 6817 6678 6851
rect 6678 6817 6696 6851
rect 6644 6808 6696 6817
rect 7380 6808 7432 6860
rect 7932 6808 7984 6860
rect 9772 6808 9824 6860
rect 11060 6808 11112 6860
rect 2596 6783 2648 6792
rect 2596 6749 2605 6783
rect 2605 6749 2648 6783
rect 1492 6715 1544 6724
rect 1492 6681 1501 6715
rect 1501 6681 1535 6715
rect 1535 6681 1544 6715
rect 1492 6672 1544 6681
rect 2596 6740 2648 6749
rect 4252 6783 4304 6792
rect 4252 6749 4261 6783
rect 4261 6749 4295 6783
rect 4295 6749 4304 6783
rect 4252 6740 4304 6749
rect 5540 6740 5592 6792
rect 6552 6783 6604 6792
rect 6552 6749 6561 6783
rect 6561 6749 6595 6783
rect 6595 6749 6604 6783
rect 6552 6740 6604 6749
rect 9312 6740 9364 6792
rect 10048 6740 10100 6792
rect 9220 6672 9272 6724
rect 10232 6672 10284 6724
rect 10600 6740 10652 6792
rect 11336 6672 11388 6724
rect 12072 6740 12124 6792
rect 12348 6740 12400 6792
rect 12808 6740 12860 6792
rect 15200 6987 15252 6996
rect 15200 6953 15209 6987
rect 15209 6953 15243 6987
rect 15243 6953 15252 6987
rect 15200 6944 15252 6953
rect 16396 6944 16448 6996
rect 16948 6944 17000 6996
rect 17132 6944 17184 6996
rect 18236 6876 18288 6928
rect 23020 6944 23072 6996
rect 21824 6876 21876 6928
rect 13912 6672 13964 6724
rect 14096 6740 14148 6792
rect 14648 6672 14700 6724
rect 2228 6604 2280 6656
rect 3240 6604 3292 6656
rect 3332 6647 3384 6656
rect 3332 6613 3341 6647
rect 3341 6613 3375 6647
rect 3375 6613 3384 6647
rect 3332 6604 3384 6613
rect 5632 6604 5684 6656
rect 5724 6604 5776 6656
rect 17776 6740 17828 6792
rect 20720 6808 20772 6860
rect 20812 6851 20864 6860
rect 20812 6817 20821 6851
rect 20821 6817 20855 6851
rect 20855 6817 20864 6851
rect 20812 6808 20864 6817
rect 19248 6783 19300 6792
rect 19248 6749 19257 6783
rect 19257 6749 19291 6783
rect 19291 6749 19300 6783
rect 19248 6740 19300 6749
rect 20628 6740 20680 6792
rect 20996 6783 21048 6792
rect 20996 6749 21005 6783
rect 21005 6749 21039 6783
rect 21039 6749 21048 6783
rect 20996 6740 21048 6749
rect 19616 6604 19668 6656
rect 20628 6604 20680 6656
rect 22284 6783 22336 6792
rect 22284 6749 22293 6783
rect 22293 6749 22327 6783
rect 22327 6749 22336 6783
rect 22284 6740 22336 6749
rect 22560 6783 22612 6792
rect 22560 6749 22569 6783
rect 22569 6749 22603 6783
rect 22603 6749 22612 6783
rect 22560 6740 22612 6749
rect 23112 6783 23164 6792
rect 23112 6749 23121 6783
rect 23121 6749 23155 6783
rect 23155 6749 23164 6783
rect 23112 6740 23164 6749
rect 23480 6783 23532 6792
rect 23480 6749 23489 6783
rect 23489 6749 23523 6783
rect 23523 6749 23532 6783
rect 23480 6740 23532 6749
rect 23848 6783 23900 6792
rect 23848 6749 23857 6783
rect 23857 6749 23891 6783
rect 23891 6749 23900 6783
rect 23848 6740 23900 6749
rect 6814 6502 6866 6554
rect 6878 6502 6930 6554
rect 6942 6502 6994 6554
rect 7006 6502 7058 6554
rect 7070 6502 7122 6554
rect 12679 6502 12731 6554
rect 12743 6502 12795 6554
rect 12807 6502 12859 6554
rect 12871 6502 12923 6554
rect 12935 6502 12987 6554
rect 18544 6502 18596 6554
rect 18608 6502 18660 6554
rect 18672 6502 18724 6554
rect 18736 6502 18788 6554
rect 18800 6502 18852 6554
rect 24409 6502 24461 6554
rect 24473 6502 24525 6554
rect 24537 6502 24589 6554
rect 24601 6502 24653 6554
rect 24665 6502 24717 6554
rect 2136 6400 2188 6452
rect 2780 6400 2832 6452
rect 3240 6400 3292 6452
rect 5724 6400 5776 6452
rect 6276 6400 6328 6452
rect 5540 6332 5592 6384
rect 10048 6400 10100 6452
rect 3792 6307 3844 6316
rect 3792 6273 3826 6307
rect 3826 6273 3844 6307
rect 3792 6264 3844 6273
rect 9680 6332 9732 6384
rect 9772 6332 9824 6384
rect 7472 6264 7524 6316
rect 9128 6264 9180 6316
rect 9312 6264 9364 6316
rect 11428 6264 11480 6316
rect 12348 6332 12400 6384
rect 1400 6239 1452 6248
rect 1400 6205 1409 6239
rect 1409 6205 1443 6239
rect 1443 6205 1452 6239
rect 1400 6196 1452 6205
rect 3332 6196 3384 6248
rect 3240 6128 3292 6180
rect 1308 6060 1360 6112
rect 2412 6060 2464 6112
rect 4344 6196 4396 6248
rect 6184 6196 6236 6248
rect 4344 6060 4396 6112
rect 4620 6103 4672 6112
rect 4620 6069 4629 6103
rect 4629 6069 4663 6103
rect 4663 6069 4672 6103
rect 4620 6060 4672 6069
rect 6368 6128 6420 6180
rect 8944 6196 8996 6248
rect 10600 6196 10652 6248
rect 13728 6332 13780 6384
rect 14188 6443 14240 6452
rect 14188 6409 14197 6443
rect 14197 6409 14231 6443
rect 14231 6409 14240 6443
rect 14188 6400 14240 6409
rect 17224 6400 17276 6452
rect 13360 6264 13412 6316
rect 15476 6264 15528 6316
rect 7656 6103 7708 6112
rect 7656 6069 7665 6103
rect 7665 6069 7699 6103
rect 7699 6069 7708 6103
rect 7656 6060 7708 6069
rect 12072 6128 12124 6180
rect 8852 6060 8904 6112
rect 9128 6060 9180 6112
rect 11612 6060 11664 6112
rect 16304 6196 16356 6248
rect 16672 6239 16724 6248
rect 16672 6205 16681 6239
rect 16681 6205 16715 6239
rect 16715 6205 16724 6239
rect 16672 6196 16724 6205
rect 15476 6128 15528 6180
rect 16028 6128 16080 6180
rect 16212 6128 16264 6180
rect 18144 6443 18196 6452
rect 18144 6409 18153 6443
rect 18153 6409 18187 6443
rect 18187 6409 18196 6443
rect 18144 6400 18196 6409
rect 18236 6400 18288 6452
rect 19248 6400 19300 6452
rect 19340 6400 19392 6452
rect 19984 6400 20036 6452
rect 19892 6332 19944 6384
rect 19432 6264 19484 6316
rect 20628 6400 20680 6452
rect 20996 6443 21048 6452
rect 20996 6409 21005 6443
rect 21005 6409 21039 6443
rect 21039 6409 21048 6443
rect 20996 6400 21048 6409
rect 21088 6400 21140 6452
rect 23020 6400 23072 6452
rect 23112 6443 23164 6452
rect 23112 6409 23121 6443
rect 23121 6409 23155 6443
rect 23155 6409 23164 6443
rect 23112 6400 23164 6409
rect 23480 6400 23532 6452
rect 23664 6400 23716 6452
rect 23848 6443 23900 6452
rect 23848 6409 23857 6443
rect 23857 6409 23891 6443
rect 23891 6409 23900 6443
rect 23848 6400 23900 6409
rect 24308 6400 24360 6452
rect 17776 6196 17828 6248
rect 18604 6239 18656 6248
rect 18604 6205 18613 6239
rect 18613 6205 18647 6239
rect 18647 6205 18656 6239
rect 18604 6196 18656 6205
rect 16396 6060 16448 6112
rect 18512 6128 18564 6180
rect 21272 6264 21324 6316
rect 21364 6307 21416 6316
rect 21364 6273 21373 6307
rect 21373 6273 21407 6307
rect 21407 6273 21416 6307
rect 21364 6264 21416 6273
rect 21824 6264 21876 6316
rect 22100 6307 22152 6316
rect 22100 6273 22109 6307
rect 22109 6273 22143 6307
rect 22143 6273 22152 6307
rect 22100 6264 22152 6273
rect 22836 6264 22888 6316
rect 23572 6264 23624 6316
rect 24032 6307 24084 6316
rect 24032 6273 24041 6307
rect 24041 6273 24075 6307
rect 24075 6273 24084 6307
rect 24032 6264 24084 6273
rect 19524 6060 19576 6112
rect 20168 6103 20220 6112
rect 20168 6069 20177 6103
rect 20177 6069 20211 6103
rect 20211 6069 20220 6103
rect 20168 6060 20220 6069
rect 20536 6060 20588 6112
rect 20720 6060 20772 6112
rect 21548 6060 21600 6112
rect 22376 6060 22428 6112
rect 22560 6060 22612 6112
rect 23112 6060 23164 6112
rect 3882 5958 3934 6010
rect 3946 5958 3998 6010
rect 4010 5958 4062 6010
rect 4074 5958 4126 6010
rect 4138 5958 4190 6010
rect 9747 5958 9799 6010
rect 9811 5958 9863 6010
rect 9875 5958 9927 6010
rect 9939 5958 9991 6010
rect 10003 5958 10055 6010
rect 15612 5958 15664 6010
rect 15676 5958 15728 6010
rect 15740 5958 15792 6010
rect 15804 5958 15856 6010
rect 15868 5958 15920 6010
rect 21477 5958 21529 6010
rect 21541 5958 21593 6010
rect 21605 5958 21657 6010
rect 21669 5958 21721 6010
rect 21733 5958 21785 6010
rect 4436 5856 4488 5908
rect 4896 5856 4948 5908
rect 1676 5763 1728 5772
rect 1676 5729 1685 5763
rect 1685 5729 1719 5763
rect 1719 5729 1728 5763
rect 1676 5720 1728 5729
rect 2136 5763 2188 5772
rect 2136 5729 2145 5763
rect 2145 5729 2179 5763
rect 2179 5729 2188 5763
rect 2136 5720 2188 5729
rect 2412 5763 2464 5772
rect 2412 5729 2421 5763
rect 2421 5729 2455 5763
rect 2455 5729 2464 5763
rect 2412 5720 2464 5729
rect 3792 5720 3844 5772
rect 5080 5763 5132 5772
rect 5080 5729 5089 5763
rect 5089 5729 5123 5763
rect 5123 5729 5132 5763
rect 5080 5720 5132 5729
rect 6460 5856 6512 5908
rect 7380 5899 7432 5908
rect 7380 5865 7389 5899
rect 7389 5865 7423 5899
rect 7423 5865 7432 5899
rect 7380 5856 7432 5865
rect 7656 5856 7708 5908
rect 8300 5856 8352 5908
rect 8760 5856 8812 5908
rect 9312 5856 9364 5908
rect 5632 5763 5684 5772
rect 5632 5729 5641 5763
rect 5641 5729 5675 5763
rect 5675 5729 5684 5763
rect 5632 5720 5684 5729
rect 7472 5720 7524 5772
rect 8668 5720 8720 5772
rect 2688 5695 2740 5704
rect 2688 5661 2697 5695
rect 2697 5661 2731 5695
rect 2731 5661 2740 5695
rect 2688 5652 2740 5661
rect 3424 5695 3476 5704
rect 3424 5661 3433 5695
rect 3433 5661 3467 5695
rect 3467 5661 3476 5695
rect 3424 5652 3476 5661
rect 4068 5695 4120 5704
rect 4068 5661 4077 5695
rect 4077 5661 4111 5695
rect 4111 5661 4120 5695
rect 4068 5652 4120 5661
rect 4528 5652 4580 5704
rect 5356 5695 5408 5704
rect 5356 5661 5365 5695
rect 5365 5661 5399 5695
rect 5399 5661 5408 5695
rect 5356 5652 5408 5661
rect 6368 5695 6420 5704
rect 6368 5661 6377 5695
rect 6377 5661 6411 5695
rect 6411 5661 6420 5695
rect 6368 5652 6420 5661
rect 9312 5652 9364 5704
rect 11060 5856 11112 5908
rect 11612 5856 11664 5908
rect 22100 5856 22152 5908
rect 22284 5856 22336 5908
rect 23940 5856 23992 5908
rect 13912 5788 13964 5840
rect 14740 5788 14792 5840
rect 13820 5720 13872 5772
rect 14280 5720 14332 5772
rect 15016 5720 15068 5772
rect 15108 5763 15160 5772
rect 15108 5729 15117 5763
rect 15117 5729 15151 5763
rect 15151 5729 15160 5763
rect 15108 5720 15160 5729
rect 18512 5788 18564 5840
rect 22468 5831 22520 5840
rect 22468 5797 22477 5831
rect 22477 5797 22511 5831
rect 22511 5797 22520 5831
rect 22468 5788 22520 5797
rect 22652 5788 22704 5840
rect 15476 5763 15528 5772
rect 15476 5729 15510 5763
rect 15510 5729 15528 5763
rect 15476 5720 15528 5729
rect 16028 5720 16080 5772
rect 16672 5720 16724 5772
rect 17408 5720 17460 5772
rect 17776 5763 17828 5772
rect 17776 5729 17785 5763
rect 17785 5729 17819 5763
rect 17819 5729 17828 5763
rect 17776 5720 17828 5729
rect 18604 5720 18656 5772
rect 11704 5652 11756 5704
rect 14832 5652 14884 5704
rect 16304 5652 16356 5704
rect 19248 5652 19300 5704
rect 19432 5695 19484 5704
rect 19432 5661 19441 5695
rect 19441 5661 19475 5695
rect 19475 5661 19484 5695
rect 19432 5652 19484 5661
rect 19616 5695 19668 5704
rect 19616 5661 19625 5695
rect 19625 5661 19659 5695
rect 19659 5661 19668 5695
rect 19616 5652 19668 5661
rect 20168 5695 20220 5704
rect 20168 5661 20177 5695
rect 20177 5661 20211 5695
rect 20211 5661 20220 5695
rect 20168 5652 20220 5661
rect 20444 5652 20496 5704
rect 20536 5695 20588 5704
rect 20536 5661 20545 5695
rect 20545 5661 20579 5695
rect 20579 5661 20588 5695
rect 20536 5652 20588 5661
rect 22192 5720 22244 5772
rect 4988 5516 5040 5568
rect 6276 5559 6328 5568
rect 6276 5525 6285 5559
rect 6285 5525 6319 5559
rect 6319 5525 6328 5559
rect 6276 5516 6328 5525
rect 8024 5516 8076 5568
rect 8576 5516 8628 5568
rect 9404 5516 9456 5568
rect 10140 5516 10192 5568
rect 17684 5584 17736 5636
rect 17776 5516 17828 5568
rect 18052 5516 18104 5568
rect 19524 5584 19576 5636
rect 22284 5695 22336 5704
rect 22284 5661 22293 5695
rect 22293 5661 22327 5695
rect 22327 5661 22336 5695
rect 22284 5652 22336 5661
rect 22744 5695 22796 5704
rect 22744 5661 22753 5695
rect 22753 5661 22787 5695
rect 22787 5661 22796 5695
rect 22744 5652 22796 5661
rect 21180 5584 21232 5636
rect 23296 5584 23348 5636
rect 23664 5584 23716 5636
rect 19984 5516 20036 5568
rect 20536 5516 20588 5568
rect 23480 5516 23532 5568
rect 6814 5414 6866 5466
rect 6878 5414 6930 5466
rect 6942 5414 6994 5466
rect 7006 5414 7058 5466
rect 7070 5414 7122 5466
rect 12679 5414 12731 5466
rect 12743 5414 12795 5466
rect 12807 5414 12859 5466
rect 12871 5414 12923 5466
rect 12935 5414 12987 5466
rect 18544 5414 18596 5466
rect 18608 5414 18660 5466
rect 18672 5414 18724 5466
rect 18736 5414 18788 5466
rect 18800 5414 18852 5466
rect 24409 5414 24461 5466
rect 24473 5414 24525 5466
rect 24537 5414 24589 5466
rect 24601 5414 24653 5466
rect 24665 5414 24717 5466
rect 2688 5312 2740 5364
rect 3240 5355 3292 5364
rect 3240 5321 3249 5355
rect 3249 5321 3283 5355
rect 3283 5321 3292 5355
rect 3240 5312 3292 5321
rect 3516 5312 3568 5364
rect 5080 5312 5132 5364
rect 6552 5312 6604 5364
rect 8576 5312 8628 5364
rect 9128 5312 9180 5364
rect 9680 5312 9732 5364
rect 10324 5312 10376 5364
rect 1676 5249 1728 5296
rect 1400 5219 1452 5228
rect 1400 5185 1409 5219
rect 1409 5185 1443 5219
rect 1443 5185 1452 5219
rect 1400 5176 1452 5185
rect 1676 5244 1701 5249
rect 1701 5244 1728 5249
rect 6276 5244 6328 5296
rect 9404 5244 9456 5296
rect 15200 5312 15252 5364
rect 19340 5312 19392 5364
rect 1216 4972 1268 5024
rect 4160 5219 4212 5228
rect 4160 5185 4169 5219
rect 4169 5185 4203 5219
rect 4203 5185 4212 5219
rect 4160 5176 4212 5185
rect 6736 5176 6788 5228
rect 5908 5108 5960 5160
rect 8576 5219 8628 5228
rect 8576 5185 8585 5219
rect 8585 5185 8619 5219
rect 8619 5185 8628 5219
rect 8576 5176 8628 5185
rect 8852 5219 8904 5228
rect 8852 5185 8861 5219
rect 8861 5185 8895 5219
rect 8895 5185 8904 5219
rect 8852 5176 8904 5185
rect 9496 5219 9548 5228
rect 9496 5185 9505 5219
rect 9505 5185 9539 5219
rect 9539 5185 9548 5219
rect 9496 5176 9548 5185
rect 9680 5176 9732 5228
rect 9956 5176 10008 5228
rect 10140 5219 10192 5228
rect 10140 5185 10149 5219
rect 10149 5185 10183 5219
rect 10183 5185 10192 5219
rect 10140 5176 10192 5185
rect 10784 5244 10836 5296
rect 15108 5244 15160 5296
rect 20904 5312 20956 5364
rect 8208 5108 8260 5160
rect 8300 5151 8352 5160
rect 8300 5117 8309 5151
rect 8309 5117 8343 5151
rect 8343 5117 8352 5151
rect 8300 5108 8352 5117
rect 8668 5108 8720 5160
rect 10232 5108 10284 5160
rect 3516 4972 3568 5024
rect 5540 5040 5592 5092
rect 12532 5176 12584 5228
rect 14004 5219 14056 5228
rect 14004 5185 14013 5219
rect 14013 5185 14047 5219
rect 14047 5185 14056 5219
rect 14004 5176 14056 5185
rect 14648 5176 14700 5228
rect 14740 5219 14792 5228
rect 14740 5185 14749 5219
rect 14749 5185 14783 5219
rect 14783 5185 14792 5219
rect 14740 5176 14792 5185
rect 14924 5176 14976 5228
rect 19248 5176 19300 5228
rect 19524 5186 19576 5238
rect 12440 5108 12492 5160
rect 13084 5108 13136 5160
rect 13728 5151 13780 5160
rect 13728 5117 13737 5151
rect 13737 5117 13771 5151
rect 13771 5117 13780 5151
rect 13728 5108 13780 5117
rect 19800 5176 19852 5228
rect 20904 5219 20956 5228
rect 20904 5185 20913 5219
rect 20913 5185 20947 5219
rect 20947 5185 20956 5219
rect 20904 5176 20956 5185
rect 20996 5176 21048 5228
rect 8024 4972 8076 5024
rect 12624 5040 12676 5092
rect 13452 5083 13504 5092
rect 13452 5049 13461 5083
rect 13461 5049 13495 5083
rect 13495 5049 13504 5083
rect 13452 5040 13504 5049
rect 9404 4972 9456 5024
rect 10968 4972 11020 5024
rect 11796 4972 11848 5024
rect 19156 5015 19208 5024
rect 19156 4981 19165 5015
rect 19165 4981 19199 5015
rect 19199 4981 19208 5015
rect 19156 4972 19208 4981
rect 20168 5108 20220 5160
rect 21916 5176 21968 5228
rect 24124 5244 24176 5296
rect 23020 5219 23072 5228
rect 23020 5185 23029 5219
rect 23029 5185 23063 5219
rect 23063 5185 23072 5219
rect 23020 5176 23072 5185
rect 20260 5040 20312 5092
rect 21364 5040 21416 5092
rect 22100 5040 22152 5092
rect 20352 4972 20404 5024
rect 21180 5015 21232 5024
rect 21180 4981 21189 5015
rect 21189 4981 21223 5015
rect 21223 4981 21232 5015
rect 21180 4972 21232 4981
rect 22008 4972 22060 5024
rect 23388 4972 23440 5024
rect 3882 4870 3934 4922
rect 3946 4870 3998 4922
rect 4010 4870 4062 4922
rect 4074 4870 4126 4922
rect 4138 4870 4190 4922
rect 9747 4870 9799 4922
rect 9811 4870 9863 4922
rect 9875 4870 9927 4922
rect 9939 4870 9991 4922
rect 10003 4870 10055 4922
rect 15612 4870 15664 4922
rect 15676 4870 15728 4922
rect 15740 4870 15792 4922
rect 15804 4870 15856 4922
rect 15868 4870 15920 4922
rect 21477 4870 21529 4922
rect 21541 4870 21593 4922
rect 21605 4870 21657 4922
rect 21669 4870 21721 4922
rect 21733 4870 21785 4922
rect 1308 4768 1360 4820
rect 3700 4768 3752 4820
rect 5080 4811 5132 4820
rect 5080 4777 5089 4811
rect 5089 4777 5123 4811
rect 5123 4777 5132 4811
rect 5080 4768 5132 4777
rect 5540 4811 5592 4820
rect 5540 4777 5549 4811
rect 5549 4777 5583 4811
rect 5583 4777 5592 4811
rect 5540 4768 5592 4777
rect 2136 4700 2188 4752
rect 2596 4700 2648 4752
rect 4436 4700 4488 4752
rect 1400 4675 1452 4684
rect 1400 4641 1409 4675
rect 1409 4641 1443 4675
rect 1443 4641 1452 4675
rect 1400 4632 1452 4641
rect 3148 4632 3200 4684
rect 1676 4607 1728 4616
rect 1676 4573 1683 4607
rect 1683 4573 1717 4607
rect 1717 4573 1728 4607
rect 1676 4564 1728 4573
rect 2596 4564 2648 4616
rect 4620 4564 4672 4616
rect 5080 4564 5132 4616
rect 6368 4768 6420 4820
rect 7104 4768 7156 4820
rect 8300 4743 8352 4752
rect 8300 4709 8309 4743
rect 8309 4709 8343 4743
rect 8343 4709 8352 4743
rect 8300 4700 8352 4709
rect 8668 4700 8720 4752
rect 10232 4768 10284 4820
rect 12624 4811 12676 4820
rect 12624 4777 12633 4811
rect 12633 4777 12667 4811
rect 12667 4777 12676 4811
rect 12624 4768 12676 4777
rect 15200 4768 15252 4820
rect 16028 4768 16080 4820
rect 19156 4768 19208 4820
rect 20168 4768 20220 4820
rect 21916 4768 21968 4820
rect 25504 4768 25556 4820
rect 7104 4564 7156 4616
rect 7288 4607 7340 4616
rect 7288 4573 7297 4607
rect 7297 4573 7331 4607
rect 7331 4573 7340 4607
rect 7288 4564 7340 4573
rect 8024 4564 8076 4616
rect 848 4428 900 4480
rect 3700 4428 3752 4480
rect 4252 4428 4304 4480
rect 4804 4496 4856 4548
rect 8944 4496 8996 4548
rect 11244 4700 11296 4752
rect 11888 4632 11940 4684
rect 14740 4675 14792 4684
rect 14740 4641 14749 4675
rect 14749 4641 14783 4675
rect 14783 4641 14792 4675
rect 14740 4632 14792 4641
rect 9312 4564 9364 4616
rect 11428 4564 11480 4616
rect 11612 4607 11664 4616
rect 11612 4573 11621 4607
rect 11621 4573 11655 4607
rect 11655 4573 11664 4607
rect 11612 4564 11664 4573
rect 12532 4564 12584 4616
rect 15108 4564 15160 4616
rect 10968 4496 11020 4548
rect 11060 4496 11112 4548
rect 17592 4564 17644 4616
rect 18236 4564 18288 4616
rect 18972 4632 19024 4684
rect 5448 4471 5500 4480
rect 5448 4437 5457 4471
rect 5457 4437 5491 4471
rect 5491 4437 5500 4471
rect 5448 4428 5500 4437
rect 7380 4428 7432 4480
rect 7472 4428 7524 4480
rect 10784 4428 10836 4480
rect 11336 4471 11388 4480
rect 11336 4437 11345 4471
rect 11345 4437 11379 4471
rect 11379 4437 11388 4471
rect 11336 4428 11388 4437
rect 11428 4428 11480 4480
rect 17776 4428 17828 4480
rect 18420 4428 18472 4480
rect 19340 4428 19392 4480
rect 19800 4607 19852 4616
rect 19800 4573 19809 4607
rect 19809 4573 19843 4607
rect 19843 4573 19852 4607
rect 19800 4564 19852 4573
rect 20076 4607 20128 4616
rect 20076 4573 20085 4607
rect 20085 4573 20119 4607
rect 20119 4573 20128 4607
rect 20076 4564 20128 4573
rect 20260 4632 20312 4684
rect 20352 4632 20404 4684
rect 20444 4607 20496 4616
rect 20444 4573 20453 4607
rect 20453 4573 20487 4607
rect 20487 4573 20496 4607
rect 20444 4564 20496 4573
rect 22192 4675 22244 4684
rect 22192 4641 22201 4675
rect 22201 4641 22235 4675
rect 22235 4641 22244 4675
rect 22192 4632 22244 4641
rect 21916 4607 21968 4616
rect 21916 4573 21925 4607
rect 21925 4573 21959 4607
rect 21959 4573 21968 4607
rect 21916 4564 21968 4573
rect 22100 4564 22152 4616
rect 22652 4564 22704 4616
rect 22836 4607 22888 4616
rect 22836 4573 22845 4607
rect 22845 4573 22879 4607
rect 22879 4573 22888 4607
rect 22836 4564 22888 4573
rect 19800 4428 19852 4480
rect 20260 4428 20312 4480
rect 25504 4496 25556 4548
rect 6814 4326 6866 4378
rect 6878 4326 6930 4378
rect 6942 4326 6994 4378
rect 7006 4326 7058 4378
rect 7070 4326 7122 4378
rect 12679 4326 12731 4378
rect 12743 4326 12795 4378
rect 12807 4326 12859 4378
rect 12871 4326 12923 4378
rect 12935 4326 12987 4378
rect 18544 4326 18596 4378
rect 18608 4326 18660 4378
rect 18672 4326 18724 4378
rect 18736 4326 18788 4378
rect 18800 4326 18852 4378
rect 24409 4326 24461 4378
rect 24473 4326 24525 4378
rect 24537 4326 24589 4378
rect 24601 4326 24653 4378
rect 24665 4326 24717 4378
rect 2228 4224 2280 4276
rect 3700 4224 3752 4276
rect 4344 4224 4396 4276
rect 4896 4224 4948 4276
rect 5080 4224 5132 4276
rect 1952 4156 2004 4208
rect 2044 4156 2096 4208
rect 1400 4131 1452 4140
rect 1400 4097 1409 4131
rect 1409 4097 1443 4131
rect 1443 4097 1452 4131
rect 1400 4088 1452 4097
rect 2504 4088 2556 4140
rect 2688 4131 2740 4140
rect 2688 4097 2697 4131
rect 2697 4097 2731 4131
rect 2731 4097 2740 4131
rect 2688 4088 2740 4097
rect 3608 4131 3660 4140
rect 3608 4097 3617 4131
rect 3617 4097 3651 4131
rect 3651 4097 3660 4131
rect 3608 4088 3660 4097
rect 6276 4156 6328 4208
rect 8944 4267 8996 4276
rect 8944 4233 8953 4267
rect 8953 4233 8987 4267
rect 8987 4233 8996 4267
rect 8944 4224 8996 4233
rect 11428 4224 11480 4276
rect 12532 4267 12584 4276
rect 12532 4233 12541 4267
rect 12541 4233 12575 4267
rect 12575 4233 12584 4267
rect 12532 4224 12584 4233
rect 14004 4224 14056 4276
rect 14556 4224 14608 4276
rect 18236 4224 18288 4276
rect 18696 4224 18748 4276
rect 19524 4224 19576 4276
rect 10508 4199 10560 4208
rect 10508 4165 10517 4199
rect 10517 4165 10551 4199
rect 10551 4165 10560 4199
rect 10508 4156 10560 4165
rect 11152 4156 11204 4208
rect 11244 4156 11296 4208
rect 14188 4156 14240 4208
rect 5356 4088 5408 4140
rect 5632 4088 5684 4140
rect 6644 4088 6696 4140
rect 7472 4088 7524 4140
rect 8300 4131 8352 4140
rect 8300 4097 8309 4131
rect 8309 4097 8343 4131
rect 8343 4097 8352 4131
rect 8300 4088 8352 4097
rect 8944 4088 8996 4140
rect 10048 4088 10100 4140
rect 10692 4088 10744 4140
rect 13268 4088 13320 4140
rect 17132 4156 17184 4208
rect 19432 4156 19484 4208
rect 17776 4088 17828 4140
rect 17868 4131 17920 4140
rect 17868 4097 17877 4131
rect 17877 4097 17911 4131
rect 17911 4097 17920 4131
rect 17868 4088 17920 4097
rect 18236 4131 18288 4140
rect 18236 4097 18245 4131
rect 18245 4097 18279 4131
rect 18279 4097 18288 4131
rect 18236 4088 18288 4097
rect 18696 4088 18748 4140
rect 19248 4088 19300 4140
rect 20536 4156 20588 4208
rect 20260 4088 20312 4140
rect 20352 4088 20404 4140
rect 23572 4224 23624 4276
rect 21640 4199 21692 4208
rect 21640 4165 21649 4199
rect 21649 4165 21683 4199
rect 21683 4165 21692 4199
rect 21640 4156 21692 4165
rect 21916 4156 21968 4208
rect 2964 3952 3016 4004
rect 3240 3952 3292 4004
rect 3332 3995 3384 4004
rect 3332 3961 3341 3995
rect 3341 3961 3375 3995
rect 3375 3961 3384 3995
rect 3332 3952 3384 3961
rect 1952 3884 2004 3936
rect 3884 4063 3936 4072
rect 3884 4029 3893 4063
rect 3893 4029 3927 4063
rect 3927 4029 3936 4063
rect 3884 4020 3936 4029
rect 7380 4020 7432 4072
rect 8024 4063 8076 4072
rect 8024 4029 8033 4063
rect 8033 4029 8067 4063
rect 8067 4029 8076 4063
rect 8024 4020 8076 4029
rect 8484 4020 8536 4072
rect 7840 3952 7892 4004
rect 4252 3884 4304 3936
rect 4528 3927 4580 3936
rect 4528 3893 4537 3927
rect 4537 3893 4571 3927
rect 4571 3893 4580 3927
rect 4528 3884 4580 3893
rect 4988 3884 5040 3936
rect 11060 4020 11112 4072
rect 11520 4063 11572 4072
rect 11520 4029 11529 4063
rect 11529 4029 11563 4063
rect 11563 4029 11572 4063
rect 11520 4020 11572 4029
rect 9312 3952 9364 4004
rect 10600 3927 10652 3936
rect 10600 3893 10609 3927
rect 10609 3893 10643 3927
rect 10643 3893 10652 3927
rect 10600 3884 10652 3893
rect 11152 3884 11204 3936
rect 12440 3884 12492 3936
rect 12992 3884 13044 3936
rect 14832 3952 14884 4004
rect 18052 3952 18104 4004
rect 18512 3952 18564 4004
rect 13912 3884 13964 3936
rect 14648 3884 14700 3936
rect 18972 3884 19024 3936
rect 21732 4020 21784 4072
rect 22008 4131 22060 4140
rect 22008 4097 22017 4131
rect 22017 4097 22051 4131
rect 22051 4097 22060 4131
rect 22008 4088 22060 4097
rect 22928 4088 22980 4140
rect 22100 4063 22152 4072
rect 22100 4029 22109 4063
rect 22109 4029 22143 4063
rect 22143 4029 22152 4063
rect 22100 4020 22152 4029
rect 24032 4199 24084 4208
rect 24032 4165 24041 4199
rect 24041 4165 24075 4199
rect 24075 4165 24084 4199
rect 24032 4156 24084 4165
rect 23296 4088 23348 4140
rect 23756 4131 23808 4140
rect 23756 4097 23765 4131
rect 23765 4097 23799 4131
rect 23799 4097 23808 4131
rect 23756 4088 23808 4097
rect 24952 4088 25004 4140
rect 21088 3952 21140 4004
rect 21272 3952 21324 4004
rect 21548 3952 21600 4004
rect 22928 3952 22980 4004
rect 23664 3952 23716 4004
rect 19248 3884 19300 3936
rect 19708 3884 19760 3936
rect 20536 3884 20588 3936
rect 23112 3927 23164 3936
rect 23112 3893 23121 3927
rect 23121 3893 23155 3927
rect 23155 3893 23164 3927
rect 23112 3884 23164 3893
rect 23940 3884 23992 3936
rect 3882 3782 3934 3834
rect 3946 3782 3998 3834
rect 4010 3782 4062 3834
rect 4074 3782 4126 3834
rect 4138 3782 4190 3834
rect 9747 3782 9799 3834
rect 9811 3782 9863 3834
rect 9875 3782 9927 3834
rect 9939 3782 9991 3834
rect 10003 3782 10055 3834
rect 15612 3782 15664 3834
rect 15676 3782 15728 3834
rect 15740 3782 15792 3834
rect 15804 3782 15856 3834
rect 15868 3782 15920 3834
rect 21477 3782 21529 3834
rect 21541 3782 21593 3834
rect 21605 3782 21657 3834
rect 21669 3782 21721 3834
rect 21733 3782 21785 3834
rect 1584 3723 1636 3732
rect 1584 3689 1593 3723
rect 1593 3689 1627 3723
rect 1627 3689 1636 3723
rect 1584 3680 1636 3689
rect 3332 3680 3384 3732
rect 4344 3680 4396 3732
rect 3056 3612 3108 3664
rect 4896 3680 4948 3732
rect 5080 3680 5132 3732
rect 1492 3544 1544 3596
rect 3792 3587 3844 3596
rect 3792 3553 3801 3587
rect 3801 3553 3835 3587
rect 3835 3553 3844 3587
rect 3792 3544 3844 3553
rect 664 3476 716 3528
rect 2964 3476 3016 3528
rect 2320 3340 2372 3392
rect 3424 3476 3476 3528
rect 4344 3544 4396 3596
rect 5724 3680 5776 3732
rect 7564 3723 7616 3732
rect 7564 3689 7573 3723
rect 7573 3689 7607 3723
rect 7607 3689 7616 3723
rect 7564 3680 7616 3689
rect 7840 3680 7892 3732
rect 9128 3680 9180 3732
rect 11888 3723 11940 3732
rect 11888 3689 11897 3723
rect 11897 3689 11931 3723
rect 11931 3689 11940 3723
rect 11888 3680 11940 3689
rect 4988 3519 5040 3528
rect 4988 3485 4997 3519
rect 4997 3485 5031 3519
rect 5031 3485 5040 3519
rect 4988 3476 5040 3485
rect 5908 3587 5960 3596
rect 5908 3553 5917 3587
rect 5917 3553 5951 3587
rect 5951 3553 5960 3587
rect 5908 3544 5960 3553
rect 6368 3587 6420 3596
rect 6368 3553 6377 3587
rect 6377 3553 6411 3587
rect 6411 3553 6420 3587
rect 6368 3544 6420 3553
rect 6460 3544 6512 3596
rect 6828 3544 6880 3596
rect 7288 3544 7340 3596
rect 8208 3544 8260 3596
rect 8944 3544 8996 3596
rect 12992 3680 13044 3732
rect 13452 3680 13504 3732
rect 7932 3476 7984 3528
rect 9588 3476 9640 3528
rect 10784 3476 10836 3528
rect 6552 3340 6604 3392
rect 7656 3383 7708 3392
rect 7656 3349 7665 3383
rect 7665 3349 7699 3383
rect 7699 3349 7708 3383
rect 7656 3340 7708 3349
rect 7932 3383 7984 3392
rect 7932 3349 7941 3383
rect 7941 3349 7975 3383
rect 7975 3349 7984 3383
rect 7932 3340 7984 3349
rect 8576 3383 8628 3392
rect 8576 3349 8585 3383
rect 8585 3349 8619 3383
rect 8619 3349 8628 3383
rect 8576 3340 8628 3349
rect 9128 3383 9180 3392
rect 9128 3349 9137 3383
rect 9137 3349 9171 3383
rect 9171 3349 9180 3383
rect 9128 3340 9180 3349
rect 9496 3451 9548 3460
rect 9496 3417 9505 3451
rect 9505 3417 9539 3451
rect 9539 3417 9548 3451
rect 9496 3408 9548 3417
rect 11244 3476 11296 3528
rect 11520 3476 11572 3528
rect 12164 3476 12216 3528
rect 17684 3680 17736 3732
rect 17868 3680 17920 3732
rect 18236 3680 18288 3732
rect 19340 3680 19392 3732
rect 19432 3680 19484 3732
rect 20260 3680 20312 3732
rect 17224 3587 17276 3596
rect 17224 3553 17233 3587
rect 17233 3553 17267 3587
rect 17267 3553 17276 3587
rect 17224 3544 17276 3553
rect 17776 3544 17828 3596
rect 17592 3519 17644 3528
rect 17592 3485 17601 3519
rect 17601 3485 17635 3519
rect 17635 3485 17644 3519
rect 17592 3476 17644 3485
rect 17684 3519 17736 3528
rect 17684 3485 17693 3519
rect 17693 3485 17727 3519
rect 17727 3485 17736 3519
rect 17684 3476 17736 3485
rect 9588 3340 9640 3392
rect 16948 3408 17000 3460
rect 18420 3476 18472 3528
rect 19248 3519 19300 3528
rect 19248 3485 19257 3519
rect 19257 3485 19291 3519
rect 19291 3485 19300 3519
rect 19248 3476 19300 3485
rect 19432 3519 19484 3528
rect 19432 3485 19441 3519
rect 19441 3485 19475 3519
rect 19475 3485 19484 3519
rect 19432 3476 19484 3485
rect 20352 3544 20404 3596
rect 19984 3519 20036 3528
rect 19984 3485 19993 3519
rect 19993 3485 20027 3519
rect 20027 3485 20036 3519
rect 19984 3476 20036 3485
rect 19340 3408 19392 3460
rect 10324 3340 10376 3392
rect 10416 3383 10468 3392
rect 10416 3349 10425 3383
rect 10425 3349 10459 3383
rect 10459 3349 10468 3383
rect 10416 3340 10468 3349
rect 18144 3383 18196 3392
rect 18144 3349 18153 3383
rect 18153 3349 18187 3383
rect 18187 3349 18196 3383
rect 18144 3340 18196 3349
rect 18236 3340 18288 3392
rect 19156 3340 19208 3392
rect 19524 3340 19576 3392
rect 20352 3340 20404 3392
rect 20904 3476 20956 3528
rect 21088 3476 21140 3528
rect 22284 3655 22336 3664
rect 22284 3621 22293 3655
rect 22293 3621 22327 3655
rect 22327 3621 22336 3655
rect 22284 3612 22336 3621
rect 21824 3544 21876 3596
rect 23664 3612 23716 3664
rect 23848 3655 23900 3664
rect 23848 3621 23857 3655
rect 23857 3621 23891 3655
rect 23891 3621 23900 3655
rect 23848 3612 23900 3621
rect 23112 3587 23164 3596
rect 23112 3553 23121 3587
rect 23121 3553 23155 3587
rect 23155 3553 23164 3587
rect 23112 3544 23164 3553
rect 22192 3476 22244 3528
rect 22468 3476 22520 3528
rect 21824 3408 21876 3460
rect 22744 3408 22796 3460
rect 23112 3408 23164 3460
rect 23480 3476 23532 3528
rect 23848 3408 23900 3460
rect 25228 3408 25280 3460
rect 6814 3238 6866 3290
rect 6878 3238 6930 3290
rect 6942 3238 6994 3290
rect 7006 3238 7058 3290
rect 7070 3238 7122 3290
rect 12679 3238 12731 3290
rect 12743 3238 12795 3290
rect 12807 3238 12859 3290
rect 12871 3238 12923 3290
rect 12935 3238 12987 3290
rect 18544 3238 18596 3290
rect 18608 3238 18660 3290
rect 18672 3238 18724 3290
rect 18736 3238 18788 3290
rect 18800 3238 18852 3290
rect 24409 3238 24461 3290
rect 24473 3238 24525 3290
rect 24537 3238 24589 3290
rect 24601 3238 24653 3290
rect 24665 3238 24717 3290
rect 1860 3136 1912 3188
rect 4528 3136 4580 3188
rect 5172 3136 5224 3188
rect 6368 3136 6420 3188
rect 6644 3136 6696 3188
rect 7196 3136 7248 3188
rect 8944 3136 8996 3188
rect 9496 3136 9548 3188
rect 4988 3068 5040 3120
rect 2228 3043 2280 3052
rect 2228 3009 2237 3043
rect 2237 3009 2271 3043
rect 2271 3009 2280 3043
rect 2228 3000 2280 3009
rect 2872 3000 2924 3052
rect 3976 3043 4028 3052
rect 3976 3009 3985 3043
rect 3985 3009 4019 3043
rect 4019 3009 4028 3043
rect 3976 3000 4028 3009
rect 5172 3039 5197 3052
rect 5197 3039 5224 3052
rect 6276 3068 6328 3120
rect 2688 2932 2740 2984
rect 3516 2932 3568 2984
rect 4344 2932 4396 2984
rect 5172 3000 5224 3039
rect 5632 3000 5684 3052
rect 7196 3043 7248 3052
rect 7196 3009 7205 3043
rect 7205 3009 7239 3043
rect 7239 3009 7248 3043
rect 7196 3000 7248 3009
rect 7472 3043 7524 3052
rect 7472 3009 7481 3043
rect 7481 3009 7515 3043
rect 7515 3009 7524 3043
rect 7472 3000 7524 3009
rect 7748 3000 7800 3052
rect 3240 2864 3292 2916
rect 3424 2907 3476 2916
rect 3424 2873 3433 2907
rect 3433 2873 3467 2907
rect 3467 2873 3476 2907
rect 3424 2864 3476 2873
rect 3516 2796 3568 2848
rect 4436 2796 4488 2848
rect 7380 2932 7432 2984
rect 6460 2864 6512 2916
rect 5908 2796 5960 2848
rect 6736 2839 6788 2848
rect 6736 2805 6745 2839
rect 6745 2805 6779 2839
rect 6779 2805 6788 2839
rect 6736 2796 6788 2805
rect 7012 2839 7064 2848
rect 7012 2805 7021 2839
rect 7021 2805 7055 2839
rect 7055 2805 7064 2839
rect 7012 2796 7064 2805
rect 8852 3000 8904 3052
rect 9404 3068 9456 3120
rect 10692 3068 10744 3120
rect 10876 3111 10928 3120
rect 10876 3077 10885 3111
rect 10885 3077 10919 3111
rect 10919 3077 10928 3111
rect 10876 3068 10928 3077
rect 12164 3136 12216 3188
rect 16948 3179 17000 3188
rect 16948 3145 16957 3179
rect 16957 3145 16991 3179
rect 16991 3145 17000 3179
rect 16948 3136 17000 3145
rect 17684 3136 17736 3188
rect 16488 3111 16540 3120
rect 16488 3077 16497 3111
rect 16497 3077 16531 3111
rect 16531 3077 16540 3111
rect 16488 3068 16540 3077
rect 19248 3136 19300 3188
rect 19340 3136 19392 3188
rect 22652 3136 22704 3188
rect 23112 3136 23164 3188
rect 24952 3136 25004 3188
rect 25596 3136 25648 3188
rect 10416 3000 10468 3052
rect 11520 3000 11572 3052
rect 17132 3000 17184 3052
rect 17408 3000 17460 3052
rect 17500 3043 17552 3052
rect 17500 3009 17509 3043
rect 17509 3009 17543 3043
rect 17543 3009 17552 3043
rect 17500 3000 17552 3009
rect 17592 3000 17644 3052
rect 18788 3068 18840 3120
rect 19064 3111 19116 3120
rect 19064 3077 19073 3111
rect 19073 3077 19107 3111
rect 19107 3077 19116 3111
rect 19064 3068 19116 3077
rect 19616 3111 19668 3120
rect 19616 3077 19625 3111
rect 19625 3077 19659 3111
rect 19659 3077 19668 3111
rect 19616 3068 19668 3077
rect 21916 3068 21968 3120
rect 8760 2932 8812 2984
rect 12532 2932 12584 2984
rect 13452 2932 13504 2984
rect 14464 2932 14516 2984
rect 8668 2864 8720 2916
rect 17224 2864 17276 2916
rect 18972 3000 19024 3052
rect 20260 3043 20312 3052
rect 20260 3009 20269 3043
rect 20269 3009 20303 3043
rect 20303 3009 20312 3043
rect 20260 3000 20312 3009
rect 20352 3043 20404 3052
rect 20352 3009 20361 3043
rect 20361 3009 20395 3043
rect 20395 3009 20404 3043
rect 20352 3000 20404 3009
rect 21640 3043 21692 3052
rect 21640 3009 21649 3043
rect 21649 3009 21683 3043
rect 21683 3009 21692 3043
rect 21640 3000 21692 3009
rect 22100 3043 22152 3052
rect 22100 3009 22109 3043
rect 22109 3009 22143 3043
rect 22143 3009 22152 3043
rect 22100 3000 22152 3009
rect 22284 3000 22336 3052
rect 18420 2932 18472 2984
rect 18696 2907 18748 2916
rect 18696 2873 18705 2907
rect 18705 2873 18739 2907
rect 18739 2873 18748 2907
rect 18696 2864 18748 2873
rect 10968 2839 11020 2848
rect 10968 2805 10977 2839
rect 10977 2805 11011 2839
rect 11011 2805 11020 2839
rect 10968 2796 11020 2805
rect 12348 2796 12400 2848
rect 17408 2796 17460 2848
rect 17500 2796 17552 2848
rect 19064 2796 19116 2848
rect 19156 2839 19208 2848
rect 19156 2805 19165 2839
rect 19165 2805 19199 2839
rect 19199 2805 19208 2839
rect 19156 2796 19208 2805
rect 19248 2796 19300 2848
rect 19800 2796 19852 2848
rect 23940 2932 23992 2984
rect 24860 2932 24912 2984
rect 25228 2932 25280 2984
rect 21272 2864 21324 2916
rect 22192 2864 22244 2916
rect 22744 2864 22796 2916
rect 23020 2796 23072 2848
rect 23480 2796 23532 2848
rect 3882 2694 3934 2746
rect 3946 2694 3998 2746
rect 4010 2694 4062 2746
rect 4074 2694 4126 2746
rect 4138 2694 4190 2746
rect 9747 2694 9799 2746
rect 9811 2694 9863 2746
rect 9875 2694 9927 2746
rect 9939 2694 9991 2746
rect 10003 2694 10055 2746
rect 15612 2694 15664 2746
rect 15676 2694 15728 2746
rect 15740 2694 15792 2746
rect 15804 2694 15856 2746
rect 15868 2694 15920 2746
rect 21477 2694 21529 2746
rect 21541 2694 21593 2746
rect 21605 2694 21657 2746
rect 21669 2694 21721 2746
rect 21733 2694 21785 2746
rect 1768 2635 1820 2644
rect 1768 2601 1777 2635
rect 1777 2601 1811 2635
rect 1811 2601 1820 2635
rect 1768 2592 1820 2601
rect 1492 2456 1544 2508
rect 2688 2592 2740 2644
rect 3700 2524 3752 2576
rect 5356 2635 5408 2644
rect 5356 2601 5365 2635
rect 5365 2601 5399 2635
rect 5399 2601 5408 2635
rect 5356 2592 5408 2601
rect 5448 2592 5500 2644
rect 4620 2524 4672 2576
rect 7288 2592 7340 2644
rect 9864 2592 9916 2644
rect 13452 2635 13504 2644
rect 13452 2601 13461 2635
rect 13461 2601 13495 2635
rect 13495 2601 13504 2635
rect 13452 2592 13504 2601
rect 16212 2592 16264 2644
rect 7748 2524 7800 2576
rect 9128 2524 9180 2576
rect 17684 2592 17736 2644
rect 17960 2592 18012 2644
rect 18328 2592 18380 2644
rect 18512 2592 18564 2644
rect 5908 2499 5960 2508
rect 5908 2465 5917 2499
rect 5917 2465 5951 2499
rect 5951 2465 5960 2499
rect 5908 2456 5960 2465
rect 10968 2456 11020 2508
rect 2136 2388 2188 2440
rect 2412 2320 2464 2372
rect 5172 2388 5224 2440
rect 6184 2431 6236 2440
rect 5448 2320 5500 2372
rect 6184 2397 6191 2431
rect 6191 2397 6225 2431
rect 6225 2397 6236 2431
rect 6184 2388 6236 2397
rect 7656 2388 7708 2440
rect 8300 2388 8352 2440
rect 8668 2431 8720 2440
rect 8668 2397 8677 2431
rect 8677 2397 8711 2431
rect 8711 2397 8720 2431
rect 8668 2388 8720 2397
rect 9128 2431 9180 2440
rect 9128 2397 9137 2431
rect 9137 2397 9171 2431
rect 9171 2397 9180 2431
rect 9128 2388 9180 2397
rect 9404 2431 9456 2440
rect 9404 2397 9413 2431
rect 9413 2397 9447 2431
rect 9447 2397 9456 2431
rect 9404 2388 9456 2397
rect 6368 2320 6420 2372
rect 3424 2252 3476 2304
rect 6000 2252 6052 2304
rect 7012 2252 7064 2304
rect 7472 2252 7524 2304
rect 8760 2320 8812 2372
rect 9864 2388 9916 2440
rect 10232 2363 10284 2372
rect 10232 2329 10241 2363
rect 10241 2329 10275 2363
rect 10275 2329 10284 2363
rect 10232 2320 10284 2329
rect 10508 2320 10560 2372
rect 10692 2431 10744 2440
rect 10692 2397 10701 2431
rect 10701 2397 10735 2431
rect 10735 2397 10744 2431
rect 10692 2388 10744 2397
rect 12348 2456 12400 2508
rect 13912 2456 13964 2508
rect 8484 2295 8536 2304
rect 8484 2261 8493 2295
rect 8493 2261 8527 2295
rect 8527 2261 8536 2295
rect 8484 2252 8536 2261
rect 9220 2295 9272 2304
rect 9220 2261 9229 2295
rect 9229 2261 9263 2295
rect 9263 2261 9272 2295
rect 9220 2252 9272 2261
rect 9312 2252 9364 2304
rect 11796 2320 11848 2372
rect 11980 2320 12032 2372
rect 11060 2295 11112 2304
rect 11060 2261 11069 2295
rect 11069 2261 11103 2295
rect 11103 2261 11112 2295
rect 11060 2252 11112 2261
rect 11244 2295 11296 2304
rect 11244 2261 11253 2295
rect 11253 2261 11287 2295
rect 11287 2261 11296 2295
rect 11244 2252 11296 2261
rect 12532 2363 12584 2372
rect 12532 2329 12541 2363
rect 12541 2329 12575 2363
rect 12575 2329 12584 2363
rect 12532 2320 12584 2329
rect 13084 2320 13136 2372
rect 13176 2320 13228 2372
rect 16488 2388 16540 2440
rect 17040 2456 17092 2508
rect 19156 2524 19208 2576
rect 20260 2592 20312 2644
rect 20444 2592 20496 2644
rect 21548 2592 21600 2644
rect 22284 2592 22336 2644
rect 25320 2592 25372 2644
rect 16856 2431 16908 2440
rect 16856 2397 16865 2431
rect 16865 2397 16899 2431
rect 16899 2397 16908 2431
rect 16856 2388 16908 2397
rect 17132 2431 17184 2440
rect 17132 2397 17141 2431
rect 17141 2397 17175 2431
rect 17175 2397 17184 2431
rect 17132 2388 17184 2397
rect 15752 2363 15804 2372
rect 15752 2329 15761 2363
rect 15761 2329 15795 2363
rect 15795 2329 15804 2363
rect 15752 2320 15804 2329
rect 13360 2252 13412 2304
rect 16120 2295 16172 2304
rect 16120 2261 16129 2295
rect 16129 2261 16163 2295
rect 16163 2261 16172 2295
rect 16120 2252 16172 2261
rect 16672 2295 16724 2304
rect 16672 2261 16681 2295
rect 16681 2261 16715 2295
rect 16715 2261 16724 2295
rect 16672 2252 16724 2261
rect 16948 2295 17000 2304
rect 16948 2261 16957 2295
rect 16957 2261 16991 2295
rect 16991 2261 17000 2295
rect 16948 2252 17000 2261
rect 17224 2320 17276 2372
rect 19892 2499 19944 2508
rect 19892 2465 19901 2499
rect 19901 2465 19935 2499
rect 19935 2465 19944 2499
rect 19892 2456 19944 2465
rect 20628 2524 20680 2576
rect 22100 2524 22152 2576
rect 23020 2456 23072 2508
rect 23388 2456 23440 2508
rect 19616 2388 19668 2440
rect 20812 2388 20864 2440
rect 21824 2388 21876 2440
rect 19340 2320 19392 2372
rect 20628 2363 20680 2372
rect 20628 2329 20637 2363
rect 20637 2329 20671 2363
rect 20671 2329 20680 2363
rect 20628 2320 20680 2329
rect 20720 2320 20772 2372
rect 21364 2320 21416 2372
rect 24124 2320 24176 2372
rect 17960 2252 18012 2304
rect 18604 2252 18656 2304
rect 19156 2252 19208 2304
rect 6814 2150 6866 2202
rect 6878 2150 6930 2202
rect 6942 2150 6994 2202
rect 7006 2150 7058 2202
rect 7070 2150 7122 2202
rect 12679 2150 12731 2202
rect 12743 2150 12795 2202
rect 12807 2150 12859 2202
rect 12871 2150 12923 2202
rect 12935 2150 12987 2202
rect 18544 2150 18596 2202
rect 18608 2150 18660 2202
rect 18672 2150 18724 2202
rect 18736 2150 18788 2202
rect 18800 2150 18852 2202
rect 24409 2150 24461 2202
rect 24473 2150 24525 2202
rect 24537 2150 24589 2202
rect 24601 2150 24653 2202
rect 24665 2150 24717 2202
rect 25412 2116 25464 2168
rect 3792 2048 3844 2100
rect 4896 2048 4948 2100
rect 6092 2091 6144 2100
rect 6092 2057 6101 2091
rect 6101 2057 6135 2091
rect 6135 2057 6144 2091
rect 6092 2048 6144 2057
rect 1676 1980 1728 2032
rect 2780 1980 2832 2032
rect 6644 2048 6696 2100
rect 7288 2048 7340 2100
rect 7656 2091 7708 2100
rect 7656 2057 7665 2091
rect 7665 2057 7699 2091
rect 7699 2057 7708 2091
rect 7656 2048 7708 2057
rect 7748 2048 7800 2100
rect 8116 2048 8168 2100
rect 8852 2048 8904 2100
rect 9220 2048 9272 2100
rect 940 1844 992 1896
rect 2688 1912 2740 1964
rect 3976 1912 4028 1964
rect 6460 2023 6512 2032
rect 6460 1989 6469 2023
rect 6469 1989 6503 2023
rect 6503 1989 6512 2023
rect 6460 1980 6512 1989
rect 6736 1980 6788 2032
rect 5356 1912 5408 1964
rect 8024 1912 8076 1964
rect 8392 1912 8444 1964
rect 8484 1912 8536 1964
rect 10048 1980 10100 2032
rect 10784 2048 10836 2100
rect 11336 2048 11388 2100
rect 11612 1980 11664 2032
rect 9496 1844 9548 1896
rect 11520 1912 11572 1964
rect 12532 2048 12584 2100
rect 14464 2091 14516 2100
rect 14464 2057 14473 2091
rect 14473 2057 14507 2091
rect 14507 2057 14516 2091
rect 14464 2048 14516 2057
rect 16672 2048 16724 2100
rect 16948 2048 17000 2100
rect 11888 2023 11940 2032
rect 11888 1989 11897 2023
rect 11897 1989 11931 2023
rect 11931 1989 11940 2023
rect 11888 1980 11940 1989
rect 12256 1912 12308 1964
rect 13268 1980 13320 2032
rect 15384 1980 15436 2032
rect 17132 1980 17184 2032
rect 17408 1980 17460 2032
rect 17960 1980 18012 2032
rect 10048 1887 10100 1896
rect 10048 1853 10057 1887
rect 10057 1853 10091 1887
rect 10091 1853 10100 1887
rect 10048 1844 10100 1853
rect 3608 1708 3660 1760
rect 4988 1708 5040 1760
rect 7932 1776 7984 1828
rect 8392 1819 8444 1828
rect 8392 1785 8401 1819
rect 8401 1785 8435 1819
rect 8435 1785 8444 1819
rect 8392 1776 8444 1785
rect 8484 1776 8536 1828
rect 9680 1776 9732 1828
rect 9956 1776 10008 1828
rect 10784 1776 10836 1828
rect 16028 1955 16080 1964
rect 16028 1921 16037 1955
rect 16037 1921 16071 1955
rect 16071 1921 16080 1955
rect 16028 1912 16080 1921
rect 16304 1912 16356 1964
rect 19064 2091 19116 2100
rect 19064 2057 19073 2091
rect 19073 2057 19107 2091
rect 19107 2057 19116 2091
rect 19064 2048 19116 2057
rect 18236 1844 18288 1896
rect 18328 1844 18380 1896
rect 19892 2048 19944 2100
rect 20076 2048 20128 2100
rect 19340 1912 19392 1964
rect 19984 1980 20036 2032
rect 20168 1980 20220 2032
rect 23664 2048 23716 2100
rect 20904 1980 20956 2032
rect 20720 1844 20772 1896
rect 10508 1708 10560 1760
rect 11796 1708 11848 1760
rect 11980 1751 12032 1760
rect 11980 1717 11989 1751
rect 11989 1717 12023 1751
rect 12023 1717 12032 1751
rect 11980 1708 12032 1717
rect 16672 1776 16724 1828
rect 19064 1776 19116 1828
rect 13728 1751 13780 1760
rect 13728 1717 13737 1751
rect 13737 1717 13771 1751
rect 13771 1717 13780 1751
rect 13728 1708 13780 1717
rect 14188 1708 14240 1760
rect 15292 1708 15344 1760
rect 15936 1708 15988 1760
rect 16396 1708 16448 1760
rect 16948 1708 17000 1760
rect 17684 1708 17736 1760
rect 20168 1708 20220 1760
rect 21088 1887 21140 1896
rect 21088 1853 21097 1887
rect 21097 1853 21131 1887
rect 21131 1853 21140 1887
rect 21088 1844 21140 1853
rect 21548 1844 21600 1896
rect 23756 1955 23808 1964
rect 23756 1921 23765 1955
rect 23765 1921 23799 1955
rect 23799 1921 23808 1955
rect 23756 1912 23808 1921
rect 20904 1776 20956 1828
rect 24676 1708 24728 1760
rect 3882 1606 3934 1658
rect 3946 1606 3998 1658
rect 4010 1606 4062 1658
rect 4074 1606 4126 1658
rect 4138 1606 4190 1658
rect 9747 1606 9799 1658
rect 9811 1606 9863 1658
rect 9875 1606 9927 1658
rect 9939 1606 9991 1658
rect 10003 1606 10055 1658
rect 15612 1606 15664 1658
rect 15676 1606 15728 1658
rect 15740 1606 15792 1658
rect 15804 1606 15856 1658
rect 15868 1606 15920 1658
rect 21477 1606 21529 1658
rect 21541 1606 21593 1658
rect 21605 1606 21657 1658
rect 21669 1606 21721 1658
rect 21733 1606 21785 1658
rect 20 1504 72 1556
rect 6092 1504 6144 1556
rect 8484 1504 8536 1556
rect 1124 1436 1176 1488
rect 4988 1436 5040 1488
rect 6276 1436 6328 1488
rect 572 1300 624 1352
rect 1032 1232 1084 1284
rect 1952 1275 2004 1284
rect 1952 1241 1961 1275
rect 1961 1241 1995 1275
rect 1995 1241 2004 1275
rect 1952 1232 2004 1241
rect 3332 1343 3384 1352
rect 3332 1309 3341 1343
rect 3341 1309 3375 1343
rect 3375 1309 3384 1343
rect 3332 1300 3384 1309
rect 3608 1368 3660 1420
rect 9496 1504 9548 1556
rect 10968 1504 11020 1556
rect 11244 1547 11296 1556
rect 11244 1513 11253 1547
rect 11253 1513 11287 1547
rect 11287 1513 11296 1547
rect 11244 1504 11296 1513
rect 11612 1504 11664 1556
rect 13728 1504 13780 1556
rect 14464 1504 14516 1556
rect 11152 1436 11204 1488
rect 13636 1436 13688 1488
rect 14924 1436 14976 1488
rect 16028 1504 16080 1556
rect 16488 1504 16540 1556
rect 20904 1504 20956 1556
rect 23112 1547 23164 1556
rect 23112 1513 23121 1547
rect 23121 1513 23155 1547
rect 23155 1513 23164 1547
rect 23112 1504 23164 1513
rect 25136 1504 25188 1556
rect 3700 1300 3752 1352
rect 3792 1343 3844 1352
rect 3792 1309 3801 1343
rect 3801 1309 3835 1343
rect 3835 1309 3844 1343
rect 3792 1300 3844 1309
rect 3976 1300 4028 1352
rect 4436 1343 4488 1352
rect 4436 1309 4445 1343
rect 4445 1309 4479 1343
rect 4479 1309 4488 1343
rect 4436 1300 4488 1309
rect 5816 1343 5868 1352
rect 5816 1309 5825 1343
rect 5825 1309 5859 1343
rect 5859 1309 5868 1343
rect 5816 1300 5868 1309
rect 6000 1343 6052 1352
rect 6000 1309 6009 1343
rect 6009 1309 6043 1343
rect 6043 1309 6052 1343
rect 6000 1300 6052 1309
rect 6092 1300 6144 1352
rect 6644 1343 6696 1352
rect 6644 1309 6653 1343
rect 6653 1309 6687 1343
rect 6687 1309 6696 1343
rect 6644 1300 6696 1309
rect 2872 1232 2924 1284
rect 4252 1232 4304 1284
rect 5264 1275 5316 1284
rect 5264 1241 5273 1275
rect 5273 1241 5307 1275
rect 5307 1241 5316 1275
rect 5264 1232 5316 1241
rect 5448 1275 5500 1284
rect 5448 1241 5457 1275
rect 5457 1241 5491 1275
rect 5491 1241 5500 1275
rect 5448 1232 5500 1241
rect 5908 1232 5960 1284
rect 2136 1164 2188 1216
rect 2412 1207 2464 1216
rect 2412 1173 2421 1207
rect 2421 1173 2455 1207
rect 2455 1173 2464 1207
rect 2412 1164 2464 1173
rect 2780 1207 2832 1216
rect 2780 1173 2789 1207
rect 2789 1173 2823 1207
rect 2823 1173 2832 1207
rect 2780 1164 2832 1173
rect 3424 1164 3476 1216
rect 3884 1164 3936 1216
rect 4068 1164 4120 1216
rect 4804 1164 4856 1216
rect 7932 1343 7984 1352
rect 7932 1309 7941 1343
rect 7941 1309 7975 1343
rect 7975 1309 7984 1343
rect 7932 1300 7984 1309
rect 9036 1343 9088 1352
rect 9036 1309 9045 1343
rect 9045 1309 9079 1343
rect 9079 1309 9088 1343
rect 9036 1300 9088 1309
rect 12072 1368 12124 1420
rect 12532 1411 12584 1420
rect 12532 1377 12541 1411
rect 12541 1377 12575 1411
rect 12575 1377 12584 1411
rect 12532 1368 12584 1377
rect 15844 1368 15896 1420
rect 18236 1436 18288 1488
rect 7472 1207 7524 1216
rect 7472 1173 7481 1207
rect 7481 1173 7515 1207
rect 7515 1173 7524 1207
rect 7472 1164 7524 1173
rect 7748 1207 7800 1216
rect 7748 1173 7757 1207
rect 7757 1173 7791 1207
rect 7791 1173 7800 1207
rect 7748 1164 7800 1173
rect 8116 1207 8168 1216
rect 8116 1173 8125 1207
rect 8125 1173 8159 1207
rect 8159 1173 8168 1207
rect 8116 1164 8168 1173
rect 9220 1232 9272 1284
rect 9956 1300 10008 1352
rect 10232 1300 10284 1352
rect 11060 1343 11112 1352
rect 11060 1309 11069 1343
rect 11069 1309 11103 1343
rect 11103 1309 11112 1343
rect 11060 1300 11112 1309
rect 11704 1343 11756 1352
rect 11704 1309 11713 1343
rect 11713 1309 11747 1343
rect 11747 1309 11756 1343
rect 11704 1300 11756 1309
rect 11796 1343 11848 1352
rect 11796 1309 11805 1343
rect 11805 1309 11839 1343
rect 11839 1309 11848 1343
rect 11796 1300 11848 1309
rect 12256 1343 12308 1352
rect 12256 1309 12265 1343
rect 12265 1309 12299 1343
rect 12299 1309 12308 1343
rect 12256 1300 12308 1309
rect 12716 1343 12768 1352
rect 12716 1309 12725 1343
rect 12725 1309 12759 1343
rect 12759 1309 12768 1343
rect 12716 1300 12768 1309
rect 13360 1300 13412 1352
rect 13452 1343 13504 1352
rect 13452 1309 13461 1343
rect 13461 1309 13495 1343
rect 13495 1309 13504 1343
rect 13452 1300 13504 1309
rect 14096 1343 14148 1352
rect 14096 1309 14105 1343
rect 14105 1309 14139 1343
rect 14139 1309 14148 1343
rect 14096 1300 14148 1309
rect 14556 1343 14608 1352
rect 14556 1309 14565 1343
rect 14565 1309 14599 1343
rect 14599 1309 14608 1343
rect 14556 1300 14608 1309
rect 15200 1300 15252 1352
rect 16120 1300 16172 1352
rect 16488 1343 16540 1352
rect 16488 1309 16497 1343
rect 16497 1309 16531 1343
rect 16531 1309 16540 1343
rect 16488 1300 16540 1309
rect 16764 1343 16816 1352
rect 16764 1309 16773 1343
rect 16773 1309 16807 1343
rect 16807 1309 16816 1343
rect 16764 1300 16816 1309
rect 17408 1300 17460 1352
rect 18236 1343 18288 1352
rect 18236 1309 18245 1343
rect 18245 1309 18279 1343
rect 18279 1309 18288 1343
rect 18236 1300 18288 1309
rect 18420 1300 18472 1352
rect 20168 1436 20220 1488
rect 23480 1436 23532 1488
rect 19432 1300 19484 1352
rect 9312 1164 9364 1216
rect 11520 1207 11572 1216
rect 11520 1173 11529 1207
rect 11529 1173 11563 1207
rect 11563 1173 11572 1207
rect 11520 1164 11572 1173
rect 12256 1164 12308 1216
rect 12900 1207 12952 1216
rect 12900 1173 12909 1207
rect 12909 1173 12943 1207
rect 12943 1173 12952 1207
rect 12900 1164 12952 1173
rect 13268 1207 13320 1216
rect 13268 1173 13277 1207
rect 13277 1173 13311 1207
rect 13311 1173 13320 1207
rect 13268 1164 13320 1173
rect 13360 1164 13412 1216
rect 13912 1164 13964 1216
rect 15108 1164 15160 1216
rect 17960 1207 18012 1216
rect 17960 1173 17969 1207
rect 17969 1173 18003 1207
rect 18003 1173 18012 1207
rect 17960 1164 18012 1173
rect 19616 1232 19668 1284
rect 19340 1164 19392 1216
rect 20720 1300 20772 1352
rect 21916 1300 21968 1352
rect 22192 1300 22244 1352
rect 20996 1232 21048 1284
rect 21548 1232 21600 1284
rect 24308 1232 24360 1284
rect 22192 1164 22244 1216
rect 22284 1164 22336 1216
rect 6814 1062 6866 1114
rect 6878 1062 6930 1114
rect 6942 1062 6994 1114
rect 7006 1062 7058 1114
rect 7070 1062 7122 1114
rect 12679 1062 12731 1114
rect 12743 1062 12795 1114
rect 12807 1062 12859 1114
rect 12871 1062 12923 1114
rect 12935 1062 12987 1114
rect 18544 1062 18596 1114
rect 18608 1062 18660 1114
rect 18672 1062 18724 1114
rect 18736 1062 18788 1114
rect 18800 1062 18852 1114
rect 24409 1062 24461 1114
rect 24473 1062 24525 1114
rect 24537 1062 24589 1114
rect 24601 1062 24653 1114
rect 24665 1062 24717 1114
rect 480 620 532 672
rect 6276 960 6328 1012
rect 3424 892 3476 944
rect 5632 892 5684 944
rect 6092 892 6144 944
rect 3332 756 3384 808
rect 5724 756 5776 808
rect 8116 824 8168 876
rect 11428 824 11480 876
rect 5448 688 5500 740
rect 8944 756 8996 808
rect 9864 756 9916 808
rect 9956 756 10008 808
rect 10784 756 10836 808
rect 16580 756 16632 808
rect 19616 960 19668 1012
rect 22100 960 22152 1012
rect 18236 892 18288 944
rect 17132 824 17184 876
rect 6644 688 6696 740
rect 10324 688 10376 740
rect 17132 688 17184 740
rect 17960 756 18012 808
rect 19340 824 19392 876
rect 20536 824 20588 876
rect 22284 824 22336 876
rect 22468 756 22520 808
rect 22928 688 22980 740
rect 2412 552 2464 604
rect 23848 620 23900 672
rect 11244 552 11296 604
rect 11980 552 12032 604
rect 3884 484 3936 536
rect 14372 552 14424 604
rect 14648 552 14700 604
rect 20996 552 21048 604
rect 16488 484 16540 536
rect 25596 484 25648 536
rect 112 416 164 468
rect 5540 416 5592 468
<< metal2 >>
rect 110 44540 166 45000
rect 386 44540 442 45000
rect 662 44540 718 45000
rect 938 44540 994 45000
rect 1214 44540 1270 45000
rect 1490 44540 1546 45000
rect 1766 44540 1822 45000
rect 2042 44540 2098 45000
rect 2318 44540 2374 45000
rect 2594 44540 2650 45000
rect 2870 44540 2926 45000
rect 3146 44540 3202 45000
rect 3422 44540 3478 45000
rect 3698 44540 3754 45000
rect 3974 44540 4030 45000
rect 4250 44540 4306 45000
rect 4526 44540 4582 45000
rect 4802 44540 4858 45000
rect 5078 44540 5134 45000
rect 5354 44540 5410 45000
rect 5630 44540 5686 45000
rect 5906 44540 5962 45000
rect 6182 44540 6238 45000
rect 6458 44540 6514 45000
rect 6734 44540 6790 45000
rect 7010 44540 7066 45000
rect 7286 44540 7342 45000
rect 7562 44540 7618 45000
rect 7838 44540 7894 45000
rect 8114 44540 8170 45000
rect 8390 44540 8446 45000
rect 8666 44540 8722 45000
rect 8942 44540 8998 45000
rect 9218 44540 9274 45000
rect 9494 44540 9550 45000
rect 9770 44540 9826 45000
rect 10046 44540 10102 45000
rect 10322 44540 10378 45000
rect 10598 44540 10654 45000
rect 10874 44540 10930 45000
rect 11150 44540 11206 45000
rect 11426 44540 11482 45000
rect 11702 44540 11758 45000
rect 11978 44540 12034 45000
rect 12254 44540 12310 45000
rect 12530 44540 12586 45000
rect 12806 44540 12862 45000
rect 13082 44540 13138 45000
rect 13358 44540 13414 45000
rect 13634 44540 13690 45000
rect 13910 44540 13966 45000
rect 14186 44540 14242 45000
rect 14462 44540 14518 45000
rect 14738 44540 14794 45000
rect 15014 44540 15070 45000
rect 15290 44540 15346 45000
rect 15566 44540 15622 45000
rect 15842 44540 15898 45000
rect 16118 44540 16174 45000
rect 16394 44540 16450 45000
rect 16670 44540 16726 45000
rect 16946 44540 17002 45000
rect 17222 44540 17278 45000
rect 17498 44540 17554 45000
rect 17774 44540 17830 45000
rect 18050 44540 18106 45000
rect 18326 44540 18382 45000
rect 18602 44540 18658 45000
rect 18878 44540 18934 45000
rect 19154 44540 19210 45000
rect 19430 44540 19486 45000
rect 19706 44540 19762 45000
rect 19982 44540 20038 45000
rect 20258 44540 20314 45000
rect 20534 44540 20590 45000
rect 20810 44540 20866 45000
rect 21086 44540 21142 45000
rect 21362 44540 21418 45000
rect 21638 44540 21694 45000
rect 21914 44540 21970 45000
rect 22190 44540 22246 45000
rect 22466 44540 22522 45000
rect 22742 44540 22798 45000
rect 23018 44540 23074 45000
rect 23294 44540 23350 45000
rect 23570 44540 23626 45000
rect 23846 44540 23902 45000
rect 24122 44540 24178 45000
rect 24398 44540 24454 45000
rect 24674 44540 24730 45000
rect 24950 44540 25006 45000
rect 25226 44540 25282 45000
rect 25502 44540 25558 45000
rect 124 43790 152 44540
rect 112 43784 164 43790
rect 112 43726 164 43732
rect 202 40624 258 40633
rect 202 40559 258 40568
rect 20 38004 72 38010
rect 20 37946 72 37952
rect 32 1562 60 37946
rect 216 3505 244 40559
rect 400 40118 428 44540
rect 676 44334 704 44540
rect 664 44328 716 44334
rect 664 44270 716 44276
rect 952 42702 980 44540
rect 940 42696 992 42702
rect 940 42638 992 42644
rect 1228 42566 1256 44540
rect 1400 43852 1452 43858
rect 1400 43794 1452 43800
rect 1412 43314 1440 43794
rect 1400 43308 1452 43314
rect 1400 43250 1452 43256
rect 1216 42560 1268 42566
rect 1216 42502 1268 42508
rect 1400 41608 1452 41614
rect 1400 41550 1452 41556
rect 1412 41449 1440 41550
rect 1398 41440 1454 41449
rect 1398 41375 1454 41384
rect 1400 41132 1452 41138
rect 1400 41074 1452 41080
rect 848 41064 900 41070
rect 848 41006 900 41012
rect 570 40216 626 40225
rect 570 40151 626 40160
rect 388 40112 440 40118
rect 388 40054 440 40060
rect 386 30424 442 30433
rect 386 30359 442 30368
rect 296 21956 348 21962
rect 296 21898 348 21904
rect 308 14482 336 21898
rect 296 14476 348 14482
rect 296 14418 348 14424
rect 400 11937 428 30359
rect 478 28792 534 28801
rect 478 28727 534 28736
rect 492 18834 520 28727
rect 480 18828 532 18834
rect 480 18770 532 18776
rect 386 11928 442 11937
rect 386 11863 442 11872
rect 202 3496 258 3505
rect 202 3431 258 3440
rect 584 2774 612 40151
rect 756 38276 808 38282
rect 756 38218 808 38224
rect 768 38185 796 38218
rect 754 38176 810 38185
rect 754 38111 810 38120
rect 664 37256 716 37262
rect 664 37198 716 37204
rect 676 36582 704 37198
rect 664 36576 716 36582
rect 664 36518 716 36524
rect 676 20602 704 36518
rect 860 33454 888 41006
rect 1412 39409 1440 41074
rect 1504 39574 1532 44540
rect 1584 43716 1636 43722
rect 1584 43658 1636 43664
rect 1596 43450 1624 43658
rect 1584 43444 1636 43450
rect 1584 43386 1636 43392
rect 1780 43217 1808 44540
rect 1766 43208 1822 43217
rect 1766 43143 1822 43152
rect 1952 42628 2004 42634
rect 1952 42570 2004 42576
rect 1676 42220 1728 42226
rect 1728 42180 1808 42208
rect 1676 42162 1728 42168
rect 1584 42152 1636 42158
rect 1584 42094 1636 42100
rect 1596 40066 1624 42094
rect 1676 40520 1728 40526
rect 1674 40488 1676 40497
rect 1728 40488 1730 40497
rect 1674 40423 1730 40432
rect 1596 40038 1716 40066
rect 1584 39976 1636 39982
rect 1584 39918 1636 39924
rect 1492 39568 1544 39574
rect 1492 39510 1544 39516
rect 1398 39400 1454 39409
rect 1398 39335 1454 39344
rect 1596 38842 1624 39918
rect 1504 38814 1624 38842
rect 1504 38758 1532 38814
rect 1492 38752 1544 38758
rect 1492 38694 1544 38700
rect 1032 38548 1084 38554
rect 1032 38490 1084 38496
rect 938 34776 994 34785
rect 938 34711 994 34720
rect 848 33448 900 33454
rect 848 33390 900 33396
rect 754 29744 810 29753
rect 754 29679 810 29688
rect 768 29646 796 29679
rect 756 29640 808 29646
rect 756 29582 808 29588
rect 756 28484 808 28490
rect 756 28426 808 28432
rect 768 28121 796 28426
rect 754 28112 810 28121
rect 754 28047 810 28056
rect 848 27600 900 27606
rect 848 27542 900 27548
rect 860 27305 888 27542
rect 846 27296 902 27305
rect 846 27231 902 27240
rect 848 25968 900 25974
rect 848 25910 900 25916
rect 860 25401 888 25910
rect 846 25392 902 25401
rect 846 25327 902 25336
rect 848 24812 900 24818
rect 848 24754 900 24760
rect 754 24304 810 24313
rect 754 24239 756 24248
rect 808 24239 810 24248
rect 756 24210 808 24216
rect 860 23769 888 24754
rect 846 23760 902 23769
rect 756 23724 808 23730
rect 846 23695 902 23704
rect 756 23666 808 23672
rect 768 23497 796 23666
rect 754 23488 810 23497
rect 754 23423 810 23432
rect 756 23044 808 23050
rect 756 22986 808 22992
rect 768 22953 796 22986
rect 848 22976 900 22982
rect 754 22944 810 22953
rect 848 22918 900 22924
rect 754 22879 810 22888
rect 860 22681 888 22918
rect 846 22672 902 22681
rect 846 22607 902 22616
rect 952 21962 980 34711
rect 940 21956 992 21962
rect 940 21898 992 21904
rect 938 21856 994 21865
rect 938 21791 994 21800
rect 754 21584 810 21593
rect 754 21519 810 21528
rect 768 20942 796 21519
rect 952 21010 980 21791
rect 940 21004 992 21010
rect 940 20946 992 20952
rect 756 20936 808 20942
rect 756 20878 808 20884
rect 940 20868 992 20874
rect 860 20828 940 20856
rect 664 20596 716 20602
rect 664 20538 716 20544
rect 754 20224 810 20233
rect 754 20159 810 20168
rect 768 19854 796 20159
rect 756 19848 808 19854
rect 756 19790 808 19796
rect 664 19508 716 19514
rect 664 19450 716 19456
rect 676 15094 704 19450
rect 754 19136 810 19145
rect 754 19071 810 19080
rect 768 18290 796 19071
rect 756 18284 808 18290
rect 756 18226 808 18232
rect 756 18012 808 18018
rect 756 17954 808 17960
rect 664 15088 716 15094
rect 664 15030 716 15036
rect 662 13424 718 13433
rect 662 13359 718 13368
rect 676 10810 704 13359
rect 664 10804 716 10810
rect 664 10746 716 10752
rect 768 9654 796 17954
rect 860 17082 888 20828
rect 940 20810 992 20816
rect 940 20528 992 20534
rect 938 20496 940 20505
rect 992 20496 994 20505
rect 938 20431 994 20440
rect 940 18488 992 18494
rect 940 18430 992 18436
rect 952 18018 980 18430
rect 940 18012 992 18018
rect 940 17954 992 17960
rect 860 17054 980 17082
rect 848 16992 900 16998
rect 846 16960 848 16969
rect 900 16960 902 16969
rect 846 16895 902 16904
rect 848 16448 900 16454
rect 848 16390 900 16396
rect 756 9648 808 9654
rect 756 9590 808 9596
rect 860 4486 888 16390
rect 952 15201 980 17054
rect 938 15192 994 15201
rect 938 15127 994 15136
rect 940 14476 992 14482
rect 940 14418 992 14424
rect 848 4480 900 4486
rect 848 4422 900 4428
rect 664 3528 716 3534
rect 664 3470 716 3476
rect 492 2746 612 2774
rect 20 1556 72 1562
rect 20 1498 72 1504
rect 492 678 520 2746
rect 572 1352 624 1358
rect 572 1294 624 1300
rect 480 672 532 678
rect 480 614 532 620
rect 112 468 164 474
rect 112 410 164 416
rect 124 160 152 410
rect 110 -300 166 160
rect 386 82 442 160
rect 584 82 612 1294
rect 676 160 704 3470
rect 952 2774 980 14418
rect 1044 12434 1072 38490
rect 1504 37806 1532 38694
rect 1582 38584 1638 38593
rect 1582 38519 1638 38528
rect 1492 37800 1544 37806
rect 1492 37742 1544 37748
rect 1214 37496 1270 37505
rect 1214 37431 1270 37440
rect 1124 33856 1176 33862
rect 1124 33798 1176 33804
rect 1136 33561 1164 33798
rect 1122 33552 1178 33561
rect 1122 33487 1178 33496
rect 1124 33448 1176 33454
rect 1124 33390 1176 33396
rect 1136 22012 1164 33390
rect 1228 28558 1256 37431
rect 1398 37224 1454 37233
rect 1398 37159 1454 37168
rect 1412 36825 1440 37159
rect 1398 36816 1454 36825
rect 1398 36751 1454 36760
rect 1400 36712 1452 36718
rect 1504 36666 1532 37742
rect 1596 37369 1624 38519
rect 1582 37360 1638 37369
rect 1582 37295 1638 37304
rect 1688 36689 1716 40038
rect 1780 36961 1808 42180
rect 1964 39953 1992 42570
rect 2056 42514 2084 44540
rect 2332 43654 2360 44540
rect 2320 43648 2372 43654
rect 2320 43590 2372 43596
rect 2504 43172 2556 43178
rect 2504 43114 2556 43120
rect 2056 42486 2176 42514
rect 2042 42256 2098 42265
rect 2042 42191 2044 42200
rect 2096 42191 2098 42200
rect 2044 42162 2096 42168
rect 2044 41540 2096 41546
rect 2044 41482 2096 41488
rect 2056 41449 2084 41482
rect 2042 41440 2098 41449
rect 2042 41375 2098 41384
rect 2148 40934 2176 42486
rect 2228 42288 2280 42294
rect 2228 42230 2280 42236
rect 2136 40928 2188 40934
rect 2136 40870 2188 40876
rect 2136 40588 2188 40594
rect 2136 40530 2188 40536
rect 1950 39944 2006 39953
rect 1950 39879 2006 39888
rect 1860 39364 1912 39370
rect 1860 39306 1912 39312
rect 1872 37466 1900 39306
rect 2044 38956 2096 38962
rect 1964 38916 2044 38944
rect 1860 37460 1912 37466
rect 1860 37402 1912 37408
rect 1766 36952 1822 36961
rect 1766 36887 1822 36896
rect 1674 36680 1730 36689
rect 1452 36660 1532 36666
rect 1400 36654 1532 36660
rect 1412 36638 1532 36654
rect 1596 36638 1674 36666
rect 1412 36258 1440 36638
rect 1412 36230 1532 36258
rect 1400 36168 1452 36174
rect 1400 36110 1452 36116
rect 1412 34105 1440 36110
rect 1504 35494 1532 36230
rect 1492 35488 1544 35494
rect 1492 35430 1544 35436
rect 1504 34542 1532 35430
rect 1492 34536 1544 34542
rect 1492 34478 1544 34484
rect 1398 34096 1454 34105
rect 1308 34060 1360 34066
rect 1398 34031 1454 34040
rect 1308 34002 1360 34008
rect 1320 33833 1348 34002
rect 1400 33992 1452 33998
rect 1400 33934 1452 33940
rect 1306 33824 1362 33833
rect 1306 33759 1362 33768
rect 1308 33584 1360 33590
rect 1308 33526 1360 33532
rect 1320 33289 1348 33526
rect 1306 33280 1362 33289
rect 1306 33215 1362 33224
rect 1412 32609 1440 33934
rect 1504 33318 1532 34478
rect 1596 33522 1624 36638
rect 1674 36615 1730 36624
rect 1768 35760 1820 35766
rect 1768 35702 1820 35708
rect 1780 35086 1808 35702
rect 1768 35080 1820 35086
rect 1768 35022 1820 35028
rect 1676 33924 1728 33930
rect 1676 33866 1728 33872
rect 1688 33561 1716 33866
rect 1674 33552 1730 33561
rect 1584 33516 1636 33522
rect 1674 33487 1730 33496
rect 1584 33458 1636 33464
rect 1492 33312 1544 33318
rect 1492 33254 1544 33260
rect 1504 32910 1532 33254
rect 1596 32960 1624 33458
rect 1596 32932 1716 32960
rect 1492 32904 1544 32910
rect 1492 32846 1544 32852
rect 1582 32872 1638 32881
rect 1398 32600 1454 32609
rect 1398 32535 1454 32544
rect 1400 32360 1452 32366
rect 1398 32328 1400 32337
rect 1452 32328 1454 32337
rect 1398 32263 1454 32272
rect 1308 32224 1360 32230
rect 1308 32166 1360 32172
rect 1320 31929 1348 32166
rect 1306 31920 1362 31929
rect 1306 31855 1362 31864
rect 1400 31816 1452 31822
rect 1306 31784 1362 31793
rect 1400 31758 1452 31764
rect 1306 31719 1362 31728
rect 1320 31498 1348 31719
rect 1412 31634 1440 31758
rect 1504 31754 1532 32846
rect 1582 32807 1638 32816
rect 1596 32434 1624 32807
rect 1584 32428 1636 32434
rect 1584 32370 1636 32376
rect 1688 32201 1716 32932
rect 1674 32192 1730 32201
rect 1674 32127 1730 32136
rect 1780 31906 1808 35022
rect 1964 34082 1992 38916
rect 2044 38898 2096 38904
rect 2148 38826 2176 40530
rect 2240 39642 2268 42230
rect 2516 42158 2544 43114
rect 2608 42362 2636 44540
rect 2688 43852 2740 43858
rect 2688 43794 2740 43800
rect 2700 43382 2728 43794
rect 2688 43376 2740 43382
rect 2688 43318 2740 43324
rect 2686 42664 2742 42673
rect 2686 42599 2688 42608
rect 2740 42599 2742 42608
rect 2688 42570 2740 42576
rect 2596 42356 2648 42362
rect 2596 42298 2648 42304
rect 2504 42152 2556 42158
rect 2504 42094 2556 42100
rect 2504 41608 2556 41614
rect 2502 41576 2504 41585
rect 2556 41576 2558 41585
rect 2502 41511 2558 41520
rect 2780 41540 2832 41546
rect 2780 41482 2832 41488
rect 2412 41200 2464 41206
rect 2412 41142 2464 41148
rect 2320 41064 2372 41070
rect 2318 41032 2320 41041
rect 2372 41032 2374 41041
rect 2318 40967 2374 40976
rect 2424 40594 2452 41142
rect 2504 41132 2556 41138
rect 2504 41074 2556 41080
rect 2412 40588 2464 40594
rect 2412 40530 2464 40536
rect 2320 40384 2372 40390
rect 2320 40326 2372 40332
rect 2332 40202 2360 40326
rect 2332 40174 2452 40202
rect 2320 40044 2372 40050
rect 2320 39986 2372 39992
rect 2228 39636 2280 39642
rect 2228 39578 2280 39584
rect 2332 39030 2360 39986
rect 2320 39024 2372 39030
rect 2320 38966 2372 38972
rect 2136 38820 2188 38826
rect 2136 38762 2188 38768
rect 2332 38654 2360 38966
rect 2148 38626 2360 38654
rect 2044 37324 2096 37330
rect 2044 37266 2096 37272
rect 2056 36922 2084 37266
rect 2044 36916 2096 36922
rect 2044 36858 2096 36864
rect 2148 36242 2176 38626
rect 2424 38162 2452 40174
rect 2516 39658 2544 41074
rect 2688 40928 2740 40934
rect 2688 40870 2740 40876
rect 2700 40730 2728 40870
rect 2688 40724 2740 40730
rect 2688 40666 2740 40672
rect 2688 40520 2740 40526
rect 2688 40462 2740 40468
rect 2700 40186 2728 40462
rect 2688 40180 2740 40186
rect 2688 40122 2740 40128
rect 2516 39642 2636 39658
rect 2516 39636 2648 39642
rect 2516 39630 2596 39636
rect 2596 39578 2648 39584
rect 2504 39432 2556 39438
rect 2504 39374 2556 39380
rect 2688 39432 2740 39438
rect 2688 39374 2740 39380
rect 2516 38826 2544 39374
rect 2700 38962 2728 39374
rect 2792 39137 2820 41482
rect 2884 40372 2912 44540
rect 3056 44192 3108 44198
rect 3056 44134 3108 44140
rect 2964 43308 3016 43314
rect 2964 43250 3016 43256
rect 2976 41546 3004 43250
rect 3068 42906 3096 44134
rect 3160 43450 3188 44540
rect 3240 43852 3292 43858
rect 3240 43794 3292 43800
rect 3148 43444 3200 43450
rect 3148 43386 3200 43392
rect 3252 43314 3280 43794
rect 3240 43308 3292 43314
rect 3240 43250 3292 43256
rect 3332 43240 3384 43246
rect 3332 43182 3384 43188
rect 3056 42900 3108 42906
rect 3056 42842 3108 42848
rect 3240 42832 3292 42838
rect 3240 42774 3292 42780
rect 3252 42634 3280 42774
rect 3240 42628 3292 42634
rect 3240 42570 3292 42576
rect 3344 42401 3372 43182
rect 3436 42770 3464 44540
rect 3516 44124 3568 44130
rect 3516 44066 3568 44072
rect 3528 42838 3556 44066
rect 3516 42832 3568 42838
rect 3516 42774 3568 42780
rect 3424 42764 3476 42770
rect 3424 42706 3476 42712
rect 3424 42560 3476 42566
rect 3424 42502 3476 42508
rect 3330 42392 3386 42401
rect 3252 42350 3330 42378
rect 3148 42288 3200 42294
rect 3148 42230 3200 42236
rect 3056 42220 3108 42226
rect 3056 42162 3108 42168
rect 3068 41818 3096 42162
rect 3056 41812 3108 41818
rect 3056 41754 3108 41760
rect 3160 41682 3188 42230
rect 3252 41750 3280 42350
rect 3436 42362 3464 42502
rect 3330 42327 3386 42336
rect 3424 42356 3476 42362
rect 3424 42298 3476 42304
rect 3240 41744 3292 41750
rect 3240 41686 3292 41692
rect 3424 41744 3476 41750
rect 3424 41686 3476 41692
rect 3148 41676 3200 41682
rect 3148 41618 3200 41624
rect 2964 41540 3016 41546
rect 2964 41482 3016 41488
rect 2964 41064 3016 41070
rect 3252 41052 3280 41686
rect 3016 41024 3280 41052
rect 2964 41006 3016 41012
rect 2964 40384 3016 40390
rect 2884 40344 2964 40372
rect 2964 40326 3016 40332
rect 2964 40112 3016 40118
rect 2964 40054 3016 40060
rect 2976 39545 3004 40054
rect 2962 39536 3018 39545
rect 2962 39471 3018 39480
rect 3068 39370 3096 41024
rect 3240 40928 3292 40934
rect 3240 40870 3292 40876
rect 3252 40594 3280 40870
rect 3436 40730 3464 41686
rect 3516 41540 3568 41546
rect 3516 41482 3568 41488
rect 3424 40724 3476 40730
rect 3424 40666 3476 40672
rect 3240 40588 3292 40594
rect 3240 40530 3292 40536
rect 3240 40452 3292 40458
rect 3240 40394 3292 40400
rect 3252 40361 3280 40394
rect 3238 40352 3294 40361
rect 3238 40287 3294 40296
rect 3528 40118 3556 41482
rect 3712 41274 3740 44540
rect 3988 43092 4016 44540
rect 3804 43064 4016 43092
rect 3700 41268 3752 41274
rect 3700 41210 3752 41216
rect 3804 40712 3832 43064
rect 3882 43004 4190 43013
rect 3882 43002 3888 43004
rect 3944 43002 3968 43004
rect 4024 43002 4048 43004
rect 4104 43002 4128 43004
rect 4184 43002 4190 43004
rect 3944 42950 3946 43002
rect 4126 42950 4128 43002
rect 3882 42948 3888 42950
rect 3944 42948 3968 42950
rect 4024 42948 4048 42950
rect 4104 42948 4128 42950
rect 4184 42948 4190 42950
rect 3882 42939 4190 42948
rect 4264 42922 4292 44540
rect 4540 44198 4568 44540
rect 4528 44192 4580 44198
rect 4528 44134 4580 44140
rect 4712 43308 4764 43314
rect 4712 43250 4764 43256
rect 4264 42894 4568 42922
rect 3974 42800 4030 42809
rect 3974 42735 4030 42744
rect 3988 42702 4016 42735
rect 3976 42696 4028 42702
rect 3976 42638 4028 42644
rect 4252 42696 4304 42702
rect 4252 42638 4304 42644
rect 4436 42696 4488 42702
rect 4436 42638 4488 42644
rect 3882 42392 3938 42401
rect 3882 42327 3938 42336
rect 4158 42392 4214 42401
rect 4158 42327 4214 42336
rect 3896 42158 3924 42327
rect 4172 42294 4200 42327
rect 4264 42294 4292 42638
rect 4448 42537 4476 42638
rect 4434 42528 4490 42537
rect 4434 42463 4490 42472
rect 4160 42288 4212 42294
rect 4160 42230 4212 42236
rect 4252 42288 4304 42294
rect 4252 42230 4304 42236
rect 3884 42152 3936 42158
rect 3884 42094 3936 42100
rect 3882 41916 4190 41925
rect 3882 41914 3888 41916
rect 3944 41914 3968 41916
rect 4024 41914 4048 41916
rect 4104 41914 4128 41916
rect 4184 41914 4190 41916
rect 3944 41862 3946 41914
rect 4126 41862 4128 41914
rect 3882 41860 3888 41862
rect 3944 41860 3968 41862
rect 4024 41860 4048 41862
rect 4104 41860 4128 41862
rect 4184 41860 4190 41862
rect 3882 41851 4190 41860
rect 3882 40828 4190 40837
rect 3882 40826 3888 40828
rect 3944 40826 3968 40828
rect 4024 40826 4048 40828
rect 4104 40826 4128 40828
rect 4184 40826 4190 40828
rect 3944 40774 3946 40826
rect 4126 40774 4128 40826
rect 3882 40772 3888 40774
rect 3944 40772 3968 40774
rect 4024 40772 4048 40774
rect 4104 40772 4128 40774
rect 4184 40772 4190 40774
rect 3882 40763 4190 40772
rect 4068 40724 4120 40730
rect 3804 40684 4068 40712
rect 4264 40712 4292 42230
rect 4344 42220 4396 42226
rect 4344 42162 4396 42168
rect 4356 42129 4384 42162
rect 4342 42120 4398 42129
rect 4342 42055 4398 42064
rect 4436 42016 4488 42022
rect 4436 41958 4488 41964
rect 4448 41721 4476 41958
rect 4434 41712 4490 41721
rect 4434 41647 4490 41656
rect 4448 41274 4476 41647
rect 4436 41268 4488 41274
rect 4436 41210 4488 41216
rect 4344 41200 4396 41206
rect 4344 41142 4396 41148
rect 4356 40934 4384 41142
rect 4436 41132 4488 41138
rect 4436 41074 4488 41080
rect 4344 40928 4396 40934
rect 4448 40905 4476 41074
rect 4344 40870 4396 40876
rect 4434 40896 4490 40905
rect 4434 40831 4490 40840
rect 4068 40666 4120 40672
rect 4172 40684 4292 40712
rect 4540 40712 4568 42894
rect 4724 42702 4752 43250
rect 4712 42696 4764 42702
rect 4712 42638 4764 42644
rect 4816 42566 4844 44540
rect 4896 42696 4948 42702
rect 5092 42650 5120 44540
rect 5368 43058 5396 44540
rect 5448 44192 5500 44198
rect 5448 44134 5500 44140
rect 4896 42638 4948 42644
rect 4804 42560 4856 42566
rect 4804 42502 4856 42508
rect 4908 42378 4936 42638
rect 4816 42350 4936 42378
rect 5000 42622 5120 42650
rect 5184 43030 5396 43058
rect 4816 42294 4844 42350
rect 4804 42288 4856 42294
rect 4804 42230 4856 42236
rect 4896 42288 4948 42294
rect 4896 42230 4948 42236
rect 4620 42016 4672 42022
rect 4620 41958 4672 41964
rect 4802 41984 4858 41993
rect 4632 41750 4660 41958
rect 4802 41919 4858 41928
rect 4620 41744 4672 41750
rect 4620 41686 4672 41692
rect 4816 41682 4844 41919
rect 4908 41818 4936 42230
rect 4896 41812 4948 41818
rect 4896 41754 4948 41760
rect 4712 41676 4764 41682
rect 4712 41618 4764 41624
rect 4804 41676 4856 41682
rect 4804 41618 4856 41624
rect 4724 41546 4752 41618
rect 4712 41540 4764 41546
rect 4712 41482 4764 41488
rect 4724 41274 4752 41482
rect 5000 41478 5028 42622
rect 5080 42560 5132 42566
rect 5080 42502 5132 42508
rect 5092 41682 5120 42502
rect 5184 42294 5212 43030
rect 5356 42696 5408 42702
rect 5356 42638 5408 42644
rect 5264 42560 5316 42566
rect 5264 42502 5316 42508
rect 5172 42288 5224 42294
rect 5172 42230 5224 42236
rect 5172 42016 5224 42022
rect 5172 41958 5224 41964
rect 5080 41676 5132 41682
rect 5184 41664 5212 41958
rect 5080 41618 5132 41624
rect 5166 41636 5212 41664
rect 4988 41472 5040 41478
rect 5166 41460 5194 41636
rect 5276 41546 5304 42502
rect 5368 42294 5396 42638
rect 5460 42344 5488 44134
rect 5540 43648 5592 43654
rect 5540 43590 5592 43596
rect 5552 43246 5580 43590
rect 5644 43450 5672 44540
rect 5816 44056 5868 44062
rect 5816 43998 5868 44004
rect 5724 43648 5776 43654
rect 5724 43590 5776 43596
rect 5632 43444 5684 43450
rect 5632 43386 5684 43392
rect 5736 43314 5764 43590
rect 5724 43308 5776 43314
rect 5724 43250 5776 43256
rect 5540 43240 5592 43246
rect 5540 43182 5592 43188
rect 5722 42800 5778 42809
rect 5722 42735 5778 42744
rect 5736 42702 5764 42735
rect 5724 42696 5776 42702
rect 5724 42638 5776 42644
rect 5630 42392 5686 42401
rect 5460 42316 5580 42344
rect 5630 42327 5686 42336
rect 5356 42288 5408 42294
rect 5356 42230 5408 42236
rect 5448 42220 5500 42226
rect 5448 42162 5500 42168
rect 5460 42022 5488 42162
rect 5448 42016 5500 42022
rect 5448 41958 5500 41964
rect 5552 41664 5580 42316
rect 5460 41636 5580 41664
rect 5264 41540 5316 41546
rect 5264 41482 5316 41488
rect 5460 41478 5488 41636
rect 5540 41540 5592 41546
rect 5540 41482 5592 41488
rect 5448 41472 5500 41478
rect 5166 41432 5212 41460
rect 4988 41414 5040 41420
rect 4712 41268 4764 41274
rect 4764 41228 4936 41256
rect 4712 41210 4764 41216
rect 4802 40760 4858 40769
rect 4712 40724 4764 40730
rect 4540 40684 4712 40712
rect 3608 40520 3660 40526
rect 3608 40462 3660 40468
rect 3516 40112 3568 40118
rect 3620 40089 3648 40462
rect 3516 40054 3568 40060
rect 3606 40080 3662 40089
rect 3424 40044 3476 40050
rect 3606 40015 3662 40024
rect 3424 39986 3476 39992
rect 3056 39364 3108 39370
rect 3108 39324 3280 39352
rect 3056 39306 3108 39312
rect 2778 39128 2834 39137
rect 2778 39063 2834 39072
rect 2688 38956 2740 38962
rect 2688 38898 2740 38904
rect 2780 38956 2832 38962
rect 2780 38898 2832 38904
rect 3056 38956 3108 38962
rect 3056 38898 3108 38904
rect 2504 38820 2556 38826
rect 2504 38762 2556 38768
rect 2240 38134 2452 38162
rect 2136 36236 2188 36242
rect 2136 36178 2188 36184
rect 2044 35828 2096 35834
rect 2044 35770 2096 35776
rect 1872 34054 1992 34082
rect 1872 32178 1900 34054
rect 1952 33992 2004 33998
rect 1952 33934 2004 33940
rect 1964 33153 1992 33934
rect 1950 33144 2006 33153
rect 1950 33079 2006 33088
rect 2056 32842 2084 35770
rect 2148 35601 2176 36178
rect 2134 35592 2190 35601
rect 2134 35527 2190 35536
rect 2240 34082 2268 38134
rect 2410 38040 2466 38049
rect 2410 37975 2466 37984
rect 2320 37936 2372 37942
rect 2320 37878 2372 37884
rect 2332 37330 2360 37878
rect 2424 37618 2452 37975
rect 2516 37754 2544 38762
rect 2792 38457 2820 38898
rect 2778 38448 2834 38457
rect 2778 38383 2834 38392
rect 2780 38344 2832 38350
rect 2780 38286 2832 38292
rect 2964 38344 3016 38350
rect 2964 38286 3016 38292
rect 2596 38276 2648 38282
rect 2596 38218 2648 38224
rect 2608 37874 2636 38218
rect 2596 37868 2648 37874
rect 2596 37810 2648 37816
rect 2516 37726 2728 37754
rect 2596 37664 2648 37670
rect 2424 37590 2544 37618
rect 2596 37606 2648 37612
rect 2320 37324 2372 37330
rect 2320 37266 2372 37272
rect 2412 37324 2464 37330
rect 2412 37266 2464 37272
rect 2318 36408 2374 36417
rect 2318 36343 2374 36352
rect 2332 36106 2360 36343
rect 2320 36100 2372 36106
rect 2320 36042 2372 36048
rect 2148 34054 2268 34082
rect 2148 33522 2176 34054
rect 2228 33924 2280 33930
rect 2228 33866 2280 33872
rect 2240 33697 2268 33866
rect 2226 33688 2282 33697
rect 2226 33623 2282 33632
rect 2332 33538 2360 36042
rect 2424 35766 2452 37266
rect 2516 37126 2544 37590
rect 2608 37330 2636 37606
rect 2596 37324 2648 37330
rect 2596 37266 2648 37272
rect 2504 37120 2556 37126
rect 2504 37062 2556 37068
rect 2596 37120 2648 37126
rect 2596 37062 2648 37068
rect 2412 35760 2464 35766
rect 2412 35702 2464 35708
rect 2412 35488 2464 35494
rect 2412 35430 2464 35436
rect 2424 35290 2452 35430
rect 2412 35284 2464 35290
rect 2412 35226 2464 35232
rect 2412 35148 2464 35154
rect 2412 35090 2464 35096
rect 2424 35057 2452 35090
rect 2410 35048 2466 35057
rect 2410 34983 2466 34992
rect 2136 33516 2188 33522
rect 2136 33458 2188 33464
rect 2240 33510 2360 33538
rect 2136 33312 2188 33318
rect 2136 33254 2188 33260
rect 2044 32836 2096 32842
rect 2044 32778 2096 32784
rect 2148 32366 2176 33254
rect 2136 32360 2188 32366
rect 2136 32302 2188 32308
rect 1872 32150 2176 32178
rect 1596 31878 1808 31906
rect 1492 31748 1544 31754
rect 1492 31690 1544 31696
rect 1412 31606 1532 31634
rect 1320 31470 1440 31498
rect 1412 31414 1440 31470
rect 1400 31408 1452 31414
rect 1306 31376 1362 31385
rect 1400 31350 1452 31356
rect 1306 31311 1308 31320
rect 1360 31311 1362 31320
rect 1308 31282 1360 31288
rect 1504 31113 1532 31606
rect 1490 31104 1546 31113
rect 1490 31039 1546 31048
rect 1400 30796 1452 30802
rect 1400 30738 1452 30744
rect 1308 30048 1360 30054
rect 1306 30016 1308 30025
rect 1360 30016 1362 30025
rect 1306 29951 1362 29960
rect 1412 29714 1440 30738
rect 1400 29708 1452 29714
rect 1400 29650 1452 29656
rect 1308 29572 1360 29578
rect 1308 29514 1360 29520
rect 1320 29481 1348 29514
rect 1306 29472 1362 29481
rect 1306 29407 1362 29416
rect 1308 29232 1360 29238
rect 1306 29200 1308 29209
rect 1360 29200 1362 29209
rect 1412 29186 1440 29650
rect 1596 29306 1624 31878
rect 1676 31816 1728 31822
rect 2044 31816 2096 31822
rect 1728 31776 1808 31804
rect 1676 31758 1728 31764
rect 1780 31754 1808 31776
rect 2044 31758 2096 31764
rect 1780 31726 1992 31754
rect 1676 31680 1728 31686
rect 1676 31622 1728 31628
rect 1688 30938 1716 31622
rect 1768 31272 1820 31278
rect 1768 31214 1820 31220
rect 1676 30932 1728 30938
rect 1676 30874 1728 30880
rect 1780 29322 1808 31214
rect 1860 30184 1912 30190
rect 1860 30126 1912 30132
rect 1872 29481 1900 30126
rect 1858 29472 1914 29481
rect 1858 29407 1914 29416
rect 1858 29336 1914 29345
rect 1584 29300 1636 29306
rect 1780 29294 1858 29322
rect 1858 29271 1914 29280
rect 1584 29242 1636 29248
rect 1412 29158 1532 29186
rect 1306 29135 1362 29144
rect 1400 29096 1452 29102
rect 1400 29038 1452 29044
rect 1216 28552 1268 28558
rect 1412 28529 1440 29038
rect 1216 28494 1268 28500
rect 1398 28520 1454 28529
rect 1398 28455 1454 28464
rect 1504 28098 1532 29158
rect 1676 29096 1728 29102
rect 1676 29038 1728 29044
rect 1688 28994 1716 29038
rect 1412 28070 1532 28098
rect 1596 28966 1716 28994
rect 1308 27872 1360 27878
rect 1306 27840 1308 27849
rect 1360 27840 1362 27849
rect 1306 27775 1362 27784
rect 1412 27470 1440 28070
rect 1492 27940 1544 27946
rect 1492 27882 1544 27888
rect 1400 27464 1452 27470
rect 1400 27406 1452 27412
rect 1308 27328 1360 27334
rect 1308 27270 1360 27276
rect 1216 27056 1268 27062
rect 1320 27033 1348 27270
rect 1216 26998 1268 27004
rect 1306 27024 1362 27033
rect 1228 26761 1256 26998
rect 1306 26959 1362 26968
rect 1412 26926 1440 27406
rect 1400 26920 1452 26926
rect 1400 26862 1452 26868
rect 1308 26784 1360 26790
rect 1214 26752 1270 26761
rect 1308 26726 1360 26732
rect 1214 26687 1270 26696
rect 1320 26489 1348 26726
rect 1412 26518 1440 26862
rect 1400 26512 1452 26518
rect 1306 26480 1362 26489
rect 1400 26454 1452 26460
rect 1306 26415 1362 26424
rect 1216 26376 1268 26382
rect 1216 26318 1268 26324
rect 1400 26376 1452 26382
rect 1400 26318 1452 26324
rect 1228 25838 1256 26318
rect 1216 25832 1268 25838
rect 1216 25774 1268 25780
rect 1228 24750 1256 25774
rect 1306 25664 1362 25673
rect 1306 25599 1362 25608
rect 1320 25294 1348 25599
rect 1308 25288 1360 25294
rect 1308 25230 1360 25236
rect 1412 24970 1440 26318
rect 1320 24942 1440 24970
rect 1320 24857 1348 24942
rect 1306 24848 1362 24857
rect 1306 24783 1362 24792
rect 1216 24744 1268 24750
rect 1216 24686 1268 24692
rect 1214 24576 1270 24585
rect 1214 24511 1270 24520
rect 1228 24206 1256 24511
rect 1216 24200 1268 24206
rect 1216 24142 1268 24148
rect 1308 24132 1360 24138
rect 1308 24074 1360 24080
rect 1320 24041 1348 24074
rect 1306 24032 1362 24041
rect 1306 23967 1362 23976
rect 1308 22704 1360 22710
rect 1308 22646 1360 22652
rect 1320 22409 1348 22646
rect 1400 22568 1452 22574
rect 1400 22510 1452 22516
rect 1306 22400 1362 22409
rect 1306 22335 1362 22344
rect 1136 21984 1256 22012
rect 1124 21616 1176 21622
rect 1124 21558 1176 21564
rect 1136 21321 1164 21558
rect 1122 21312 1178 21321
rect 1122 21247 1178 21256
rect 1124 20392 1176 20398
rect 1124 20334 1176 20340
rect 1136 19417 1164 20334
rect 1228 20058 1256 21984
rect 1412 21486 1440 22510
rect 1504 22012 1532 27882
rect 1596 25226 1624 28966
rect 1768 27940 1820 27946
rect 1768 27882 1820 27888
rect 1780 27849 1808 27882
rect 1766 27840 1822 27849
rect 1766 27775 1822 27784
rect 1768 27396 1820 27402
rect 1768 27338 1820 27344
rect 1676 26376 1728 26382
rect 1676 26318 1728 26324
rect 1688 25265 1716 26318
rect 1674 25256 1730 25265
rect 1584 25220 1636 25226
rect 1674 25191 1730 25200
rect 1584 25162 1636 25168
rect 1674 24848 1730 24857
rect 1596 24818 1674 24834
rect 1584 24812 1674 24818
rect 1636 24806 1674 24812
rect 1674 24783 1730 24792
rect 1584 24754 1636 24760
rect 1582 24712 1638 24721
rect 1582 24647 1584 24656
rect 1636 24647 1638 24656
rect 1584 24618 1636 24624
rect 1688 24562 1716 24783
rect 1596 24534 1716 24562
rect 1596 22080 1624 24534
rect 1676 23724 1728 23730
rect 1676 23666 1728 23672
rect 1688 23497 1716 23666
rect 1674 23488 1730 23497
rect 1674 23423 1730 23432
rect 1780 22642 1808 27338
rect 1872 26042 1900 29271
rect 1964 26246 1992 31726
rect 2056 30841 2084 31758
rect 2042 30832 2098 30841
rect 2042 30767 2098 30776
rect 2044 30592 2096 30598
rect 2044 30534 2096 30540
rect 2056 30190 2084 30534
rect 2044 30184 2096 30190
rect 2044 30126 2096 30132
rect 2148 29646 2176 32150
rect 2240 31278 2268 33510
rect 2410 33144 2466 33153
rect 2410 33079 2466 33088
rect 2320 32564 2372 32570
rect 2320 32506 2372 32512
rect 2332 32434 2360 32506
rect 2320 32428 2372 32434
rect 2320 32370 2372 32376
rect 2320 31680 2372 31686
rect 2320 31622 2372 31628
rect 2228 31272 2280 31278
rect 2228 31214 2280 31220
rect 2228 30116 2280 30122
rect 2228 30058 2280 30064
rect 2136 29640 2188 29646
rect 2136 29582 2188 29588
rect 2240 29034 2268 30058
rect 2228 29028 2280 29034
rect 2228 28970 2280 28976
rect 2332 28490 2360 31622
rect 2424 30734 2452 33079
rect 2516 31793 2544 37062
rect 2608 36650 2636 37062
rect 2596 36644 2648 36650
rect 2596 36586 2648 36592
rect 2596 36372 2648 36378
rect 2596 36314 2648 36320
rect 2608 33810 2636 36314
rect 2700 34626 2728 37726
rect 2792 36938 2820 38286
rect 2872 38276 2924 38282
rect 2872 38218 2924 38224
rect 2884 37074 2912 38218
rect 2976 37233 3004 38286
rect 2962 37224 3018 37233
rect 2962 37159 3018 37168
rect 3068 37097 3096 38898
rect 3252 38418 3280 39324
rect 3332 39296 3384 39302
rect 3332 39238 3384 39244
rect 3240 38412 3292 38418
rect 3240 38354 3292 38360
rect 3146 38312 3202 38321
rect 3146 38247 3202 38256
rect 3160 37874 3188 38247
rect 3148 37868 3200 37874
rect 3148 37810 3200 37816
rect 3252 37670 3280 38354
rect 3240 37664 3292 37670
rect 3160 37624 3240 37652
rect 3054 37088 3110 37097
rect 2884 37046 3004 37074
rect 2792 36910 2912 36938
rect 2780 36780 2832 36786
rect 2780 36722 2832 36728
rect 2792 34921 2820 36722
rect 2884 36281 2912 36910
rect 2870 36272 2926 36281
rect 2870 36207 2926 36216
rect 2976 35834 3004 37046
rect 3054 37023 3110 37032
rect 3054 36952 3110 36961
rect 3054 36887 3056 36896
rect 3108 36887 3110 36896
rect 3056 36858 3108 36864
rect 3056 36780 3108 36786
rect 3056 36722 3108 36728
rect 2964 35828 3016 35834
rect 2964 35770 3016 35776
rect 2964 35692 3016 35698
rect 2964 35634 3016 35640
rect 2976 35290 3004 35634
rect 2964 35284 3016 35290
rect 2964 35226 3016 35232
rect 3068 35193 3096 36722
rect 3160 36378 3188 37624
rect 3240 37606 3292 37612
rect 3240 37256 3292 37262
rect 3240 37198 3292 37204
rect 3148 36372 3200 36378
rect 3148 36314 3200 36320
rect 3146 36272 3202 36281
rect 3146 36207 3202 36216
rect 3160 36038 3188 36207
rect 3148 36032 3200 36038
rect 3148 35974 3200 35980
rect 3160 35834 3188 35974
rect 3148 35828 3200 35834
rect 3148 35770 3200 35776
rect 3054 35184 3110 35193
rect 3054 35119 3110 35128
rect 2872 35080 2924 35086
rect 2872 35022 2924 35028
rect 2778 34912 2834 34921
rect 2778 34847 2834 34856
rect 2780 34740 2832 34746
rect 2884 34728 2912 35022
rect 3160 34762 3188 35770
rect 3252 35737 3280 37198
rect 3238 35728 3294 35737
rect 3238 35663 3294 35672
rect 3344 35630 3372 39238
rect 3436 39098 3464 39986
rect 3700 39976 3752 39982
rect 3700 39918 3752 39924
rect 3792 39976 3844 39982
rect 3792 39918 3844 39924
rect 3976 39976 4028 39982
rect 4172 39964 4200 40684
rect 4802 40695 4858 40704
rect 4712 40666 4764 40672
rect 4252 40520 4304 40526
rect 4252 40462 4304 40468
rect 4028 39936 4200 39964
rect 3976 39918 4028 39924
rect 3516 39840 3568 39846
rect 3516 39782 3568 39788
rect 3424 39092 3476 39098
rect 3424 39034 3476 39040
rect 3436 38758 3464 39034
rect 3424 38752 3476 38758
rect 3424 38694 3476 38700
rect 3424 37664 3476 37670
rect 3424 37606 3476 37612
rect 3436 35766 3464 37606
rect 3424 35760 3476 35766
rect 3424 35702 3476 35708
rect 3332 35624 3384 35630
rect 3332 35566 3384 35572
rect 3332 35284 3384 35290
rect 3332 35226 3384 35232
rect 3160 34734 3280 34762
rect 2832 34700 2912 34728
rect 2780 34682 2832 34688
rect 2700 34598 3004 34626
rect 2976 34542 3004 34598
rect 2964 34536 3016 34542
rect 2964 34478 3016 34484
rect 2608 33782 2912 33810
rect 2596 33516 2648 33522
rect 2596 33458 2648 33464
rect 2608 32858 2636 33458
rect 2608 32830 2728 32858
rect 2596 32768 2648 32774
rect 2596 32710 2648 32716
rect 2608 32434 2636 32710
rect 2596 32428 2648 32434
rect 2596 32370 2648 32376
rect 2700 32314 2728 32830
rect 2780 32360 2832 32366
rect 2700 32308 2780 32314
rect 2700 32302 2832 32308
rect 2700 32286 2820 32302
rect 2594 32192 2650 32201
rect 2594 32127 2650 32136
rect 2608 31822 2636 32127
rect 2596 31816 2648 31822
rect 2502 31784 2558 31793
rect 2596 31758 2648 31764
rect 2502 31719 2558 31728
rect 2412 30728 2464 30734
rect 2700 30682 2728 32286
rect 2884 31754 2912 33782
rect 2792 31726 2912 31754
rect 2792 31090 2820 31726
rect 2872 31272 2924 31278
rect 2870 31240 2872 31249
rect 2924 31240 2926 31249
rect 2870 31175 2926 31184
rect 2792 31062 2912 31090
rect 2884 30938 2912 31062
rect 2872 30932 2924 30938
rect 2872 30874 2924 30880
rect 2412 30670 2464 30676
rect 2516 30654 2728 30682
rect 2780 30728 2832 30734
rect 2780 30670 2832 30676
rect 2410 29608 2466 29617
rect 2410 29543 2466 29552
rect 2424 29510 2452 29543
rect 2516 29510 2544 30654
rect 2596 30252 2648 30258
rect 2596 30194 2648 30200
rect 2412 29504 2464 29510
rect 2412 29446 2464 29452
rect 2504 29504 2556 29510
rect 2504 29446 2556 29452
rect 2424 29322 2452 29446
rect 2424 29294 2544 29322
rect 2412 29164 2464 29170
rect 2412 29106 2464 29112
rect 2424 28937 2452 29106
rect 2410 28928 2466 28937
rect 2410 28863 2466 28872
rect 2320 28484 2372 28490
rect 2320 28426 2372 28432
rect 2332 28370 2360 28426
rect 2332 28342 2452 28370
rect 2320 28212 2372 28218
rect 2320 28154 2372 28160
rect 2332 28082 2360 28154
rect 2424 28082 2452 28342
rect 2320 28076 2372 28082
rect 2320 28018 2372 28024
rect 2412 28076 2464 28082
rect 2412 28018 2464 28024
rect 2136 28008 2188 28014
rect 2318 27976 2374 27985
rect 2188 27956 2318 27962
rect 2136 27950 2318 27956
rect 2044 27940 2096 27946
rect 2148 27934 2318 27950
rect 2318 27911 2374 27920
rect 2044 27882 2096 27888
rect 2056 27130 2084 27882
rect 2044 27124 2096 27130
rect 2044 27066 2096 27072
rect 2044 26512 2096 26518
rect 2042 26480 2044 26489
rect 2096 26480 2098 26489
rect 2042 26415 2098 26424
rect 1952 26240 2004 26246
rect 1952 26182 2004 26188
rect 1860 26036 1912 26042
rect 1860 25978 1912 25984
rect 2332 25786 2360 27911
rect 2516 27554 2544 29294
rect 2608 29073 2636 30194
rect 2688 29776 2740 29782
rect 2688 29718 2740 29724
rect 2700 29238 2728 29718
rect 2688 29232 2740 29238
rect 2688 29174 2740 29180
rect 2594 29064 2650 29073
rect 2594 28999 2650 29008
rect 2688 29028 2740 29034
rect 2688 28970 2740 28976
rect 2700 28257 2728 28970
rect 2792 28665 2820 30670
rect 2872 30184 2924 30190
rect 2872 30126 2924 30132
rect 2884 29850 2912 30126
rect 2872 29844 2924 29850
rect 2872 29786 2924 29792
rect 2778 28656 2834 28665
rect 2778 28591 2834 28600
rect 2686 28248 2742 28257
rect 2686 28183 2742 28192
rect 2596 28008 2648 28014
rect 2596 27950 2648 27956
rect 2608 27674 2636 27950
rect 2596 27668 2648 27674
rect 2596 27610 2648 27616
rect 2976 27554 3004 34478
rect 3252 33862 3280 34734
rect 3240 33856 3292 33862
rect 3240 33798 3292 33804
rect 3148 32836 3200 32842
rect 3148 32778 3200 32784
rect 3056 32768 3108 32774
rect 3160 32745 3188 32778
rect 3056 32710 3108 32716
rect 3146 32736 3202 32745
rect 3068 30297 3096 32710
rect 3146 32671 3202 32680
rect 3148 31816 3200 31822
rect 3148 31758 3200 31764
rect 3054 30288 3110 30297
rect 3054 30223 3110 30232
rect 3056 30184 3108 30190
rect 3056 30126 3108 30132
rect 3068 27656 3096 30126
rect 3160 29170 3188 31758
rect 3252 31414 3280 33798
rect 3344 33386 3372 35226
rect 3528 35086 3556 39782
rect 3606 39264 3662 39273
rect 3606 39199 3662 39208
rect 3620 38894 3648 39199
rect 3712 38894 3740 39918
rect 3804 39522 3832 39918
rect 3882 39740 4190 39749
rect 3882 39738 3888 39740
rect 3944 39738 3968 39740
rect 4024 39738 4048 39740
rect 4104 39738 4128 39740
rect 4184 39738 4190 39740
rect 3944 39686 3946 39738
rect 4126 39686 4128 39738
rect 3882 39684 3888 39686
rect 3944 39684 3968 39686
rect 4024 39684 4048 39686
rect 4104 39684 4128 39686
rect 4184 39684 4190 39686
rect 3882 39675 4190 39684
rect 3804 39494 3924 39522
rect 3792 39432 3844 39438
rect 3792 39374 3844 39380
rect 3608 38888 3660 38894
rect 3608 38830 3660 38836
rect 3700 38888 3752 38894
rect 3700 38830 3752 38836
rect 3608 38752 3660 38758
rect 3700 38752 3752 38758
rect 3608 38694 3660 38700
rect 3698 38720 3700 38729
rect 3752 38720 3754 38729
rect 3620 38298 3648 38694
rect 3698 38655 3754 38664
rect 3698 38584 3754 38593
rect 3804 38570 3832 39374
rect 3896 39137 3924 39494
rect 3882 39128 3938 39137
rect 3882 39063 3938 39072
rect 3974 38992 4030 39001
rect 3974 38927 3976 38936
rect 4028 38927 4030 38936
rect 3976 38898 4028 38904
rect 3882 38652 4190 38661
rect 3882 38650 3888 38652
rect 3944 38650 3968 38652
rect 4024 38650 4048 38652
rect 4104 38650 4128 38652
rect 4184 38650 4190 38652
rect 3944 38598 3946 38650
rect 4126 38598 4128 38650
rect 3882 38596 3888 38598
rect 3944 38596 3968 38598
rect 4024 38596 4048 38598
rect 4104 38596 4128 38598
rect 4184 38596 4190 38598
rect 3882 38587 4190 38596
rect 3754 38542 3832 38570
rect 3698 38519 3754 38528
rect 3700 38480 3752 38486
rect 3752 38440 4200 38468
rect 3700 38422 3752 38428
rect 4068 38344 4120 38350
rect 3896 38304 4068 38332
rect 3620 38270 3740 38298
rect 3608 38208 3660 38214
rect 3608 38150 3660 38156
rect 3620 37942 3648 38150
rect 3608 37936 3660 37942
rect 3608 37878 3660 37884
rect 3712 36802 3740 38270
rect 3896 38185 3924 38304
rect 4068 38286 4120 38292
rect 3976 38208 4028 38214
rect 3882 38176 3938 38185
rect 3976 38150 4028 38156
rect 3882 38111 3938 38120
rect 3988 38010 4016 38150
rect 4080 38010 4108 38286
rect 4172 38282 4200 38440
rect 4160 38276 4212 38282
rect 4160 38218 4212 38224
rect 3976 38004 4028 38010
rect 3976 37946 4028 37952
rect 4068 38004 4120 38010
rect 4068 37946 4120 37952
rect 3882 37564 4190 37573
rect 3882 37562 3888 37564
rect 3944 37562 3968 37564
rect 4024 37562 4048 37564
rect 4104 37562 4128 37564
rect 4184 37562 4190 37564
rect 3944 37510 3946 37562
rect 4126 37510 4128 37562
rect 3882 37508 3888 37510
rect 3944 37508 3968 37510
rect 4024 37508 4048 37510
rect 4104 37508 4128 37510
rect 4184 37508 4190 37510
rect 3882 37499 4190 37508
rect 4264 37369 4292 40462
rect 4436 40452 4488 40458
rect 4436 40394 4488 40400
rect 4344 38956 4396 38962
rect 4344 38898 4396 38904
rect 4356 37777 4384 38898
rect 4342 37768 4398 37777
rect 4342 37703 4398 37712
rect 4250 37360 4306 37369
rect 4250 37295 4306 37304
rect 3882 37224 3938 37233
rect 3882 37159 3938 37168
rect 3976 37188 4028 37194
rect 3896 37126 3924 37159
rect 3976 37130 4028 37136
rect 3884 37120 3936 37126
rect 3884 37062 3936 37068
rect 3608 36780 3660 36786
rect 3712 36774 3832 36802
rect 3608 36722 3660 36728
rect 3620 35465 3648 36722
rect 3700 36712 3752 36718
rect 3700 36654 3752 36660
rect 3712 36122 3740 36654
rect 3804 36224 3832 36774
rect 3988 36718 4016 37130
rect 4158 37088 4214 37097
rect 4158 37023 4214 37032
rect 4172 36854 4200 37023
rect 4448 36854 4476 40394
rect 4816 40168 4844 40695
rect 4632 40140 4844 40168
rect 4528 39432 4580 39438
rect 4526 39400 4528 39409
rect 4580 39400 4582 39409
rect 4526 39335 4582 39344
rect 4528 38888 4580 38894
rect 4528 38830 4580 38836
rect 4540 37874 4568 38830
rect 4528 37868 4580 37874
rect 4528 37810 4580 37816
rect 4540 37466 4568 37810
rect 4528 37460 4580 37466
rect 4528 37402 4580 37408
rect 4160 36848 4212 36854
rect 4160 36790 4212 36796
rect 4436 36848 4488 36854
rect 4632 36802 4660 40140
rect 4804 40044 4856 40050
rect 4804 39986 4856 39992
rect 4712 39432 4764 39438
rect 4712 39374 4764 39380
rect 4724 38894 4752 39374
rect 4712 38888 4764 38894
rect 4712 38830 4764 38836
rect 4816 38826 4844 39986
rect 4908 39302 4936 41228
rect 5184 41206 5212 41432
rect 5448 41414 5500 41420
rect 5172 41200 5224 41206
rect 5172 41142 5224 41148
rect 5460 41138 5488 41414
rect 5552 41206 5580 41482
rect 5644 41478 5672 42327
rect 5736 41585 5764 42638
rect 5722 41576 5778 41585
rect 5722 41511 5778 41520
rect 5632 41472 5684 41478
rect 5632 41414 5684 41420
rect 5828 41414 5856 43998
rect 5920 43450 5948 44540
rect 6196 44266 6224 44540
rect 6184 44260 6236 44266
rect 6184 44202 6236 44208
rect 6472 44146 6500 44540
rect 6552 44260 6604 44266
rect 6552 44202 6604 44208
rect 6196 44118 6500 44146
rect 6000 43852 6052 43858
rect 6000 43794 6052 43800
rect 5908 43444 5960 43450
rect 5908 43386 5960 43392
rect 5906 43208 5962 43217
rect 5906 43143 5962 43152
rect 5920 41546 5948 43143
rect 5908 41540 5960 41546
rect 5908 41482 5960 41488
rect 5644 41206 5672 41414
rect 5828 41386 5948 41414
rect 5540 41200 5592 41206
rect 5540 41142 5592 41148
rect 5632 41200 5684 41206
rect 5632 41142 5684 41148
rect 5080 41132 5132 41138
rect 5080 41074 5132 41080
rect 5448 41132 5500 41138
rect 5448 41074 5500 41080
rect 4988 39840 5040 39846
rect 4988 39782 5040 39788
rect 5000 39506 5028 39782
rect 4988 39500 5040 39506
rect 4988 39442 5040 39448
rect 5092 39370 5120 41074
rect 5552 41052 5580 41142
rect 5816 41132 5868 41138
rect 5816 41074 5868 41080
rect 5724 41064 5776 41070
rect 5552 41024 5672 41052
rect 5446 40488 5502 40497
rect 5644 40458 5672 41024
rect 5724 41006 5776 41012
rect 5736 40730 5764 41006
rect 5724 40724 5776 40730
rect 5724 40666 5776 40672
rect 5446 40423 5502 40432
rect 5540 40452 5592 40458
rect 5354 40080 5410 40089
rect 5354 40015 5410 40024
rect 5080 39364 5132 39370
rect 5080 39306 5132 39312
rect 5172 39364 5224 39370
rect 5172 39306 5224 39312
rect 4896 39296 4948 39302
rect 4896 39238 4948 39244
rect 4804 38820 4856 38826
rect 4804 38762 4856 38768
rect 4712 38480 4764 38486
rect 4712 38422 4764 38428
rect 4436 36790 4488 36796
rect 4540 36774 4660 36802
rect 4724 36802 4752 38422
rect 4908 37369 4936 39238
rect 4988 38344 5040 38350
rect 4988 38286 5040 38292
rect 5000 37913 5028 38286
rect 4986 37904 5042 37913
rect 4986 37839 5042 37848
rect 4988 37460 5040 37466
rect 4988 37402 5040 37408
rect 4894 37360 4950 37369
rect 4894 37295 4950 37304
rect 4908 37194 4936 37295
rect 4896 37188 4948 37194
rect 4896 37130 4948 37136
rect 4896 36916 4948 36922
rect 4896 36858 4948 36864
rect 4724 36774 4844 36802
rect 3976 36712 4028 36718
rect 3976 36654 4028 36660
rect 4436 36712 4488 36718
rect 4436 36654 4488 36660
rect 3882 36476 4190 36485
rect 3882 36474 3888 36476
rect 3944 36474 3968 36476
rect 4024 36474 4048 36476
rect 4104 36474 4128 36476
rect 4184 36474 4190 36476
rect 3944 36422 3946 36474
rect 4126 36422 4128 36474
rect 3882 36420 3888 36422
rect 3944 36420 3968 36422
rect 4024 36420 4048 36422
rect 4104 36420 4128 36422
rect 4184 36420 4190 36422
rect 3882 36411 4190 36420
rect 4448 36360 4476 36654
rect 3988 36332 4476 36360
rect 3804 36196 3924 36224
rect 3790 36136 3846 36145
rect 3712 36094 3790 36122
rect 3790 36071 3846 36080
rect 3896 35476 3924 36196
rect 3988 35834 4016 36332
rect 4540 36224 4568 36774
rect 4712 36712 4764 36718
rect 4712 36654 4764 36660
rect 4724 36553 4752 36654
rect 4710 36544 4766 36553
rect 4710 36479 4766 36488
rect 4448 36196 4568 36224
rect 4448 36038 4476 36196
rect 4816 36088 4844 36774
rect 4908 36582 4936 36858
rect 4896 36576 4948 36582
rect 5000 36553 5028 37402
rect 5092 37262 5120 39306
rect 5184 39098 5212 39306
rect 5172 39092 5224 39098
rect 5172 39034 5224 39040
rect 5368 38654 5396 40015
rect 5276 38626 5396 38654
rect 5276 38282 5304 38626
rect 5460 38486 5488 40423
rect 5540 40394 5592 40400
rect 5632 40452 5684 40458
rect 5632 40394 5684 40400
rect 5448 38480 5500 38486
rect 5448 38422 5500 38428
rect 5264 38276 5316 38282
rect 5264 38218 5316 38224
rect 5448 38276 5500 38282
rect 5448 38218 5500 38224
rect 5172 37936 5224 37942
rect 5172 37878 5224 37884
rect 5080 37256 5132 37262
rect 5080 37198 5132 37204
rect 5080 36848 5132 36854
rect 5080 36790 5132 36796
rect 4896 36518 4948 36524
rect 4986 36544 5042 36553
rect 4986 36479 5042 36488
rect 5092 36122 5120 36790
rect 5184 36786 5212 37878
rect 5276 37505 5304 38218
rect 5460 37670 5488 38218
rect 5356 37664 5408 37670
rect 5356 37606 5408 37612
rect 5448 37664 5500 37670
rect 5448 37606 5500 37612
rect 5262 37496 5318 37505
rect 5368 37482 5396 37606
rect 5368 37454 5488 37482
rect 5262 37431 5318 37440
rect 5460 37330 5488 37454
rect 5448 37324 5500 37330
rect 5448 37266 5500 37272
rect 5356 37188 5408 37194
rect 5356 37130 5408 37136
rect 5264 37120 5316 37126
rect 5264 37062 5316 37068
rect 5276 36922 5304 37062
rect 5368 36922 5396 37130
rect 5264 36916 5316 36922
rect 5264 36858 5316 36864
rect 5356 36916 5408 36922
rect 5356 36858 5408 36864
rect 5172 36780 5224 36786
rect 5172 36722 5224 36728
rect 4724 36060 4844 36088
rect 5000 36094 5120 36122
rect 4068 36032 4120 36038
rect 4068 35974 4120 35980
rect 4436 36032 4488 36038
rect 4436 35974 4488 35980
rect 4528 36032 4580 36038
rect 4724 36020 4752 36060
rect 4896 36032 4948 36038
rect 4580 35992 4752 36020
rect 4816 35992 4896 36020
rect 4528 35974 4580 35980
rect 3976 35828 4028 35834
rect 3976 35770 4028 35776
rect 3606 35456 3662 35465
rect 3606 35391 3662 35400
rect 3712 35448 3924 35476
rect 4080 35476 4108 35974
rect 4434 35864 4490 35873
rect 4816 35850 4844 35992
rect 4896 35974 4948 35980
rect 5000 35850 5028 36094
rect 5080 36032 5132 36038
rect 5080 35974 5132 35980
rect 4434 35799 4490 35808
rect 4724 35822 4844 35850
rect 4908 35822 5028 35850
rect 4344 35488 4396 35494
rect 4080 35448 4292 35476
rect 3608 35284 3660 35290
rect 3608 35226 3660 35232
rect 3620 35086 3648 35226
rect 3516 35080 3568 35086
rect 3516 35022 3568 35028
rect 3608 35080 3660 35086
rect 3608 35022 3660 35028
rect 3424 34944 3476 34950
rect 3424 34886 3476 34892
rect 3332 33380 3384 33386
rect 3332 33322 3384 33328
rect 3436 33046 3464 34886
rect 3608 34400 3660 34406
rect 3608 34342 3660 34348
rect 3620 34202 3648 34342
rect 3608 34196 3660 34202
rect 3608 34138 3660 34144
rect 3712 34105 3740 35448
rect 3882 35388 4190 35397
rect 3882 35386 3888 35388
rect 3944 35386 3968 35388
rect 4024 35386 4048 35388
rect 4104 35386 4128 35388
rect 4184 35386 4190 35388
rect 3944 35334 3946 35386
rect 4126 35334 4128 35386
rect 3882 35332 3888 35334
rect 3944 35332 3968 35334
rect 4024 35332 4048 35334
rect 4104 35332 4128 35334
rect 4184 35332 4190 35334
rect 3882 35323 4190 35332
rect 3792 35080 3844 35086
rect 3792 35022 3844 35028
rect 3884 35080 3936 35086
rect 3884 35022 3936 35028
rect 3804 34513 3832 35022
rect 3896 34649 3924 35022
rect 3882 34640 3938 34649
rect 3882 34575 3938 34584
rect 3790 34504 3846 34513
rect 4264 34490 4292 35448
rect 4344 35430 4396 35436
rect 4356 35057 4384 35430
rect 4342 35048 4398 35057
rect 4342 34983 4398 34992
rect 4264 34462 4384 34490
rect 3790 34439 3846 34448
rect 4252 34400 4304 34406
rect 4252 34342 4304 34348
rect 3882 34300 4190 34309
rect 3882 34298 3888 34300
rect 3944 34298 3968 34300
rect 4024 34298 4048 34300
rect 4104 34298 4128 34300
rect 4184 34298 4190 34300
rect 3944 34246 3946 34298
rect 4126 34246 4128 34298
rect 3882 34244 3888 34246
rect 3944 34244 3968 34246
rect 4024 34244 4048 34246
rect 4104 34244 4128 34246
rect 4184 34244 4190 34246
rect 3882 34235 4190 34244
rect 4068 34196 4120 34202
rect 4068 34138 4120 34144
rect 3698 34096 3754 34105
rect 3698 34031 3700 34040
rect 3752 34031 3754 34040
rect 3700 34002 3752 34008
rect 4080 33946 4108 34138
rect 4264 34066 4292 34342
rect 4252 34060 4304 34066
rect 4252 34002 4304 34008
rect 4158 33960 4214 33969
rect 3608 33924 3660 33930
rect 3528 33884 3608 33912
rect 3424 33040 3476 33046
rect 3424 32982 3476 32988
rect 3332 32972 3384 32978
rect 3332 32914 3384 32920
rect 3344 31822 3372 32914
rect 3424 32428 3476 32434
rect 3424 32370 3476 32376
rect 3332 31816 3384 31822
rect 3332 31758 3384 31764
rect 3332 31680 3384 31686
rect 3332 31622 3384 31628
rect 3240 31408 3292 31414
rect 3240 31350 3292 31356
rect 3252 31090 3280 31350
rect 3344 31278 3372 31622
rect 3332 31272 3384 31278
rect 3332 31214 3384 31220
rect 3252 31062 3372 31090
rect 3148 29164 3200 29170
rect 3148 29106 3200 29112
rect 3160 28762 3188 29106
rect 3148 28756 3200 28762
rect 3148 28698 3200 28704
rect 3240 28484 3292 28490
rect 3240 28426 3292 28432
rect 3252 28218 3280 28426
rect 3344 28422 3372 31062
rect 3436 30569 3464 32370
rect 3528 31634 3556 33884
rect 3608 33866 3660 33872
rect 4080 33918 4158 33946
rect 4080 33522 4108 33918
rect 4356 33930 4384 34462
rect 4158 33895 4214 33904
rect 4344 33924 4396 33930
rect 4344 33866 4396 33872
rect 4160 33856 4212 33862
rect 4158 33824 4160 33833
rect 4212 33824 4214 33833
rect 4448 33810 4476 35799
rect 4620 35012 4672 35018
rect 4620 34954 4672 34960
rect 4528 34944 4580 34950
rect 4528 34886 4580 34892
rect 4158 33759 4214 33768
rect 4356 33782 4476 33810
rect 4356 33658 4384 33782
rect 4344 33652 4396 33658
rect 4344 33594 4396 33600
rect 3976 33516 4028 33522
rect 3976 33458 4028 33464
rect 4068 33516 4120 33522
rect 4068 33458 4120 33464
rect 4436 33516 4488 33522
rect 4436 33458 4488 33464
rect 3792 33448 3844 33454
rect 3988 33425 4016 33458
rect 3792 33390 3844 33396
rect 3974 33416 4030 33425
rect 3606 33008 3662 33017
rect 3606 32943 3662 32952
rect 3620 32502 3648 32943
rect 3608 32496 3660 32502
rect 3608 32438 3660 32444
rect 3804 32366 3832 33390
rect 3974 33351 4030 33360
rect 4252 33380 4304 33386
rect 4252 33322 4304 33328
rect 4264 33266 4292 33322
rect 4342 33280 4398 33289
rect 4264 33238 4342 33266
rect 3882 33212 4190 33221
rect 3882 33210 3888 33212
rect 3944 33210 3968 33212
rect 4024 33210 4048 33212
rect 4104 33210 4128 33212
rect 4184 33210 4190 33212
rect 3944 33158 3946 33210
rect 4126 33158 4128 33210
rect 3882 33156 3888 33158
rect 3944 33156 3968 33158
rect 4024 33156 4048 33158
rect 4104 33156 4128 33158
rect 4184 33156 4190 33158
rect 3882 33147 4190 33156
rect 3608 32360 3660 32366
rect 3608 32302 3660 32308
rect 3792 32360 3844 32366
rect 3792 32302 3844 32308
rect 3620 31890 3648 32302
rect 3882 32124 4190 32133
rect 3882 32122 3888 32124
rect 3944 32122 3968 32124
rect 4024 32122 4048 32124
rect 4104 32122 4128 32124
rect 4184 32122 4190 32124
rect 3944 32070 3946 32122
rect 4126 32070 4128 32122
rect 3882 32068 3888 32070
rect 3944 32068 3968 32070
rect 4024 32068 4048 32070
rect 4104 32068 4128 32070
rect 4184 32068 4190 32070
rect 3882 32059 4190 32068
rect 3700 32020 3752 32026
rect 3700 31962 3752 31968
rect 3792 32020 3844 32026
rect 3792 31962 3844 31968
rect 3608 31884 3660 31890
rect 3608 31826 3660 31832
rect 3712 31686 3740 31962
rect 3804 31754 3832 31962
rect 3804 31726 4016 31754
rect 3700 31680 3752 31686
rect 3528 31606 3648 31634
rect 3700 31622 3752 31628
rect 3514 31512 3570 31521
rect 3514 31447 3570 31456
rect 3422 30560 3478 30569
rect 3422 30495 3478 30504
rect 3528 30326 3556 31447
rect 3620 31346 3648 31606
rect 3988 31346 4016 31726
rect 3608 31340 3660 31346
rect 3976 31340 4028 31346
rect 3660 31300 3832 31328
rect 3608 31282 3660 31288
rect 3606 30832 3662 30841
rect 3606 30767 3662 30776
rect 3516 30320 3568 30326
rect 3516 30262 3568 30268
rect 3516 30048 3568 30054
rect 3516 29990 3568 29996
rect 3528 29617 3556 29990
rect 3514 29608 3570 29617
rect 3514 29543 3570 29552
rect 3424 29504 3476 29510
rect 3424 29446 3476 29452
rect 3516 29504 3568 29510
rect 3516 29446 3568 29452
rect 3436 29306 3464 29446
rect 3424 29300 3476 29306
rect 3424 29242 3476 29248
rect 3528 29186 3556 29446
rect 3436 29158 3556 29186
rect 3332 28416 3384 28422
rect 3332 28358 3384 28364
rect 3240 28212 3292 28218
rect 3240 28154 3292 28160
rect 3332 27872 3384 27878
rect 3332 27814 3384 27820
rect 3068 27628 3280 27656
rect 2516 27526 2636 27554
rect 2502 26888 2558 26897
rect 2502 26823 2558 26832
rect 2516 26382 2544 26823
rect 2504 26376 2556 26382
rect 2504 26318 2556 26324
rect 2410 26072 2466 26081
rect 2410 26007 2466 26016
rect 2504 26036 2556 26042
rect 2424 25906 2452 26007
rect 2504 25978 2556 25984
rect 2412 25900 2464 25906
rect 2412 25842 2464 25848
rect 2240 25758 2360 25786
rect 1860 25220 1912 25226
rect 1860 25162 1912 25168
rect 1952 25220 2004 25226
rect 1952 25162 2004 25168
rect 1768 22636 1820 22642
rect 1768 22578 1820 22584
rect 1872 22098 1900 25162
rect 1964 24954 1992 25162
rect 1952 24948 2004 24954
rect 1952 24890 2004 24896
rect 2044 24608 2096 24614
rect 2044 24550 2096 24556
rect 1952 23724 2004 23730
rect 1952 23666 2004 23672
rect 1964 22137 1992 23666
rect 2056 23186 2084 24550
rect 2136 24268 2188 24274
rect 2136 24210 2188 24216
rect 2148 23730 2176 24210
rect 2136 23724 2188 23730
rect 2136 23666 2188 23672
rect 2044 23180 2096 23186
rect 2044 23122 2096 23128
rect 2042 23080 2098 23089
rect 2042 23015 2098 23024
rect 1950 22128 2006 22137
rect 1860 22092 1912 22098
rect 1596 22052 1716 22080
rect 1504 21984 1624 22012
rect 1492 21888 1544 21894
rect 1492 21830 1544 21836
rect 1400 21480 1452 21486
rect 1400 21422 1452 21428
rect 1308 21344 1360 21350
rect 1308 21286 1360 21292
rect 1320 21049 1348 21286
rect 1306 21040 1362 21049
rect 1306 20975 1362 20984
rect 1308 20256 1360 20262
rect 1308 20198 1360 20204
rect 1216 20052 1268 20058
rect 1216 19994 1268 20000
rect 1320 19938 1348 20198
rect 1412 20040 1440 21422
rect 1504 20913 1532 21830
rect 1490 20904 1546 20913
rect 1490 20839 1546 20848
rect 1596 20806 1624 21984
rect 1584 20800 1636 20806
rect 1490 20768 1546 20777
rect 1584 20742 1636 20748
rect 1490 20703 1546 20712
rect 1504 20466 1532 20703
rect 1584 20596 1636 20602
rect 1584 20538 1636 20544
rect 1596 20505 1624 20538
rect 1582 20496 1638 20505
rect 1492 20460 1544 20466
rect 1582 20431 1638 20440
rect 1492 20402 1544 20408
rect 1688 20210 1716 22052
rect 1950 22063 2006 22072
rect 1860 22034 1912 22040
rect 1952 21888 2004 21894
rect 1952 21830 2004 21836
rect 1964 21400 1992 21830
rect 2056 21554 2084 23015
rect 2136 22092 2188 22098
rect 2136 22034 2188 22040
rect 2148 21690 2176 22034
rect 2136 21684 2188 21690
rect 2136 21626 2188 21632
rect 2044 21548 2096 21554
rect 2044 21490 2096 21496
rect 2136 21412 2188 21418
rect 1964 21372 2136 21400
rect 1860 20800 1912 20806
rect 1860 20742 1912 20748
rect 1688 20182 1808 20210
rect 1674 20088 1730 20097
rect 1412 20012 1532 20040
rect 1674 20023 1730 20032
rect 1228 19910 1348 19938
rect 1398 19952 1454 19961
rect 1122 19408 1178 19417
rect 1122 19343 1178 19352
rect 1228 16454 1256 19910
rect 1398 19887 1454 19896
rect 1308 19780 1360 19786
rect 1308 19722 1360 19728
rect 1320 19689 1348 19722
rect 1306 19680 1362 19689
rect 1306 19615 1362 19624
rect 1412 18766 1440 19887
rect 1504 19174 1532 20012
rect 1688 19990 1716 20023
rect 1676 19984 1728 19990
rect 1676 19926 1728 19932
rect 1492 19168 1544 19174
rect 1492 19110 1544 19116
rect 1400 18760 1452 18766
rect 1400 18702 1452 18708
rect 1504 18222 1532 19110
rect 1584 18760 1636 18766
rect 1584 18702 1636 18708
rect 1596 18290 1624 18702
rect 1584 18284 1636 18290
rect 1584 18226 1636 18232
rect 1492 18216 1544 18222
rect 1492 18158 1544 18164
rect 1400 18080 1452 18086
rect 1400 18022 1452 18028
rect 1412 17678 1440 18022
rect 1400 17672 1452 17678
rect 1400 17614 1452 17620
rect 1308 17604 1360 17610
rect 1308 17546 1360 17552
rect 1320 17513 1348 17546
rect 1306 17504 1362 17513
rect 1306 17439 1362 17448
rect 1216 16448 1268 16454
rect 1216 16390 1268 16396
rect 1412 16046 1440 17614
rect 1492 17196 1544 17202
rect 1492 17138 1544 17144
rect 1400 16040 1452 16046
rect 1504 16017 1532 17138
rect 1596 16266 1624 18226
rect 1688 16454 1716 19926
rect 1780 18737 1808 20182
rect 1872 19446 1900 20742
rect 1860 19440 1912 19446
rect 1860 19382 1912 19388
rect 1766 18728 1822 18737
rect 1822 18686 1900 18714
rect 1766 18663 1822 18672
rect 1872 18290 1900 18686
rect 1860 18284 1912 18290
rect 1860 18226 1912 18232
rect 1860 17536 1912 17542
rect 1860 17478 1912 17484
rect 1872 16726 1900 17478
rect 1768 16720 1820 16726
rect 1768 16662 1820 16668
rect 1860 16720 1912 16726
rect 1860 16662 1912 16668
rect 1676 16448 1728 16454
rect 1676 16390 1728 16396
rect 1596 16238 1716 16266
rect 1582 16144 1638 16153
rect 1582 16079 1638 16088
rect 1400 15982 1452 15988
rect 1490 16008 1546 16017
rect 1122 15872 1178 15881
rect 1122 15807 1178 15816
rect 1136 15706 1164 15807
rect 1124 15700 1176 15706
rect 1124 15642 1176 15648
rect 1216 15632 1268 15638
rect 1216 15574 1268 15580
rect 1306 15600 1362 15609
rect 1228 15337 1256 15574
rect 1306 15535 1362 15544
rect 1320 15434 1348 15535
rect 1308 15428 1360 15434
rect 1308 15370 1360 15376
rect 1214 15328 1270 15337
rect 1214 15263 1270 15272
rect 1308 15156 1360 15162
rect 1308 15098 1360 15104
rect 1122 15056 1178 15065
rect 1122 14991 1178 15000
rect 1136 14550 1164 14991
rect 1320 14793 1348 15098
rect 1412 14958 1440 15982
rect 1490 15943 1546 15952
rect 1400 14952 1452 14958
rect 1400 14894 1452 14900
rect 1306 14784 1362 14793
rect 1306 14719 1362 14728
rect 1124 14544 1176 14550
rect 1124 14486 1176 14492
rect 1306 13832 1362 13841
rect 1306 13767 1362 13776
rect 1214 13152 1270 13161
rect 1320 13138 1348 13767
rect 1412 13326 1440 14894
rect 1596 14618 1624 16079
rect 1584 14612 1636 14618
rect 1584 14554 1636 14560
rect 1492 14340 1544 14346
rect 1492 14282 1544 14288
rect 1504 14074 1532 14282
rect 1492 14068 1544 14074
rect 1492 14010 1544 14016
rect 1688 14006 1716 16238
rect 1780 15910 1808 16662
rect 1964 16590 1992 21372
rect 2136 21354 2188 21360
rect 2136 20936 2188 20942
rect 2136 20878 2188 20884
rect 2148 20806 2176 20878
rect 2136 20800 2188 20806
rect 2134 20768 2136 20777
rect 2188 20768 2190 20777
rect 2134 20703 2190 20712
rect 2042 20632 2098 20641
rect 2240 20602 2268 25758
rect 2412 25696 2464 25702
rect 2412 25638 2464 25644
rect 2424 25362 2452 25638
rect 2412 25356 2464 25362
rect 2412 25298 2464 25304
rect 2516 25242 2544 25978
rect 2320 25220 2372 25226
rect 2320 25162 2372 25168
rect 2424 25214 2544 25242
rect 2332 20942 2360 25162
rect 2424 22137 2452 25214
rect 2608 23798 2636 27526
rect 2792 27526 3004 27554
rect 2792 27384 2820 27526
rect 2872 27464 2924 27470
rect 2700 27356 2820 27384
rect 2870 27432 2872 27441
rect 2964 27464 3016 27470
rect 2924 27432 2926 27441
rect 2964 27406 3016 27412
rect 2870 27367 2926 27376
rect 2700 26994 2728 27356
rect 2976 27130 3004 27406
rect 2964 27124 3016 27130
rect 2964 27066 3016 27072
rect 2688 26988 2740 26994
rect 2688 26930 2740 26936
rect 2780 26988 2832 26994
rect 2780 26930 2832 26936
rect 2872 26988 2924 26994
rect 2872 26930 2924 26936
rect 2700 25684 2728 26930
rect 2792 25945 2820 26930
rect 2884 26217 2912 26930
rect 3056 26444 3108 26450
rect 3056 26386 3108 26392
rect 2870 26208 2926 26217
rect 2870 26143 2926 26152
rect 2778 25936 2834 25945
rect 2778 25871 2834 25880
rect 2780 25696 2832 25702
rect 2700 25656 2780 25684
rect 2780 25638 2832 25644
rect 2792 24970 2820 25638
rect 2870 25256 2926 25265
rect 2870 25191 2926 25200
rect 2964 25220 3016 25226
rect 2884 25158 2912 25191
rect 2964 25162 3016 25168
rect 2872 25152 2924 25158
rect 2872 25094 2924 25100
rect 2792 24942 2912 24970
rect 2780 24880 2832 24886
rect 2780 24822 2832 24828
rect 2792 24342 2820 24822
rect 2780 24336 2832 24342
rect 2780 24278 2832 24284
rect 2504 23792 2556 23798
rect 2502 23760 2504 23769
rect 2596 23792 2648 23798
rect 2556 23760 2558 23769
rect 2596 23734 2648 23740
rect 2502 23695 2558 23704
rect 2780 23724 2832 23730
rect 2780 23666 2832 23672
rect 2792 23633 2820 23666
rect 2778 23624 2834 23633
rect 2778 23559 2834 23568
rect 2502 23488 2558 23497
rect 2502 23423 2558 23432
rect 2516 23304 2544 23423
rect 2686 23352 2742 23361
rect 2596 23316 2648 23322
rect 2516 23276 2596 23304
rect 2686 23287 2742 23296
rect 2596 23258 2648 23264
rect 2700 23118 2728 23287
rect 2504 23112 2556 23118
rect 2504 23054 2556 23060
rect 2688 23112 2740 23118
rect 2884 23089 2912 24942
rect 2688 23054 2740 23060
rect 2870 23080 2926 23089
rect 2410 22128 2466 22137
rect 2410 22063 2466 22072
rect 2412 21548 2464 21554
rect 2412 21490 2464 21496
rect 2320 20936 2372 20942
rect 2320 20878 2372 20884
rect 2424 20788 2452 21490
rect 2332 20760 2452 20788
rect 2042 20567 2044 20576
rect 2096 20567 2098 20576
rect 2228 20596 2280 20602
rect 2044 20538 2096 20544
rect 2228 20538 2280 20544
rect 2056 19825 2084 20538
rect 2136 19848 2188 19854
rect 2042 19816 2098 19825
rect 2136 19790 2188 19796
rect 2042 19751 2098 19760
rect 2148 19689 2176 19790
rect 2240 19718 2268 20538
rect 2332 19904 2360 20760
rect 2516 20466 2544 23054
rect 2780 23044 2832 23050
rect 2870 23015 2926 23024
rect 2780 22986 2832 22992
rect 2688 22432 2740 22438
rect 2688 22374 2740 22380
rect 2594 22128 2650 22137
rect 2700 22098 2728 22374
rect 2594 22063 2596 22072
rect 2648 22063 2650 22072
rect 2688 22092 2740 22098
rect 2596 22034 2648 22040
rect 2688 22034 2740 22040
rect 2688 21004 2740 21010
rect 2688 20946 2740 20952
rect 2596 20868 2648 20874
rect 2596 20810 2648 20816
rect 2608 20602 2636 20810
rect 2596 20596 2648 20602
rect 2596 20538 2648 20544
rect 2504 20460 2556 20466
rect 2504 20402 2556 20408
rect 2412 20052 2464 20058
rect 2516 20040 2544 20402
rect 2700 20058 2728 20946
rect 2464 20012 2544 20040
rect 2688 20052 2740 20058
rect 2412 19994 2464 20000
rect 2688 19994 2740 20000
rect 2688 19916 2740 19922
rect 2332 19876 2688 19904
rect 2228 19712 2280 19718
rect 2134 19680 2190 19689
rect 2228 19654 2280 19660
rect 2134 19615 2190 19624
rect 2226 19544 2282 19553
rect 2226 19479 2282 19488
rect 2240 19446 2268 19479
rect 2136 19440 2188 19446
rect 2136 19382 2188 19388
rect 2228 19440 2280 19446
rect 2228 19382 2280 19388
rect 2148 18465 2176 19382
rect 2412 19168 2464 19174
rect 2412 19110 2464 19116
rect 2424 18902 2452 19110
rect 2412 18896 2464 18902
rect 2412 18838 2464 18844
rect 2134 18456 2190 18465
rect 2134 18391 2190 18400
rect 2136 17876 2188 17882
rect 2136 17818 2188 17824
rect 1952 16584 2004 16590
rect 1952 16526 2004 16532
rect 1768 15904 1820 15910
rect 1768 15846 1820 15852
rect 1766 14376 1822 14385
rect 1766 14311 1822 14320
rect 1676 14000 1728 14006
rect 1582 13968 1638 13977
rect 1676 13942 1728 13948
rect 1582 13903 1638 13912
rect 1492 13864 1544 13870
rect 1492 13806 1544 13812
rect 1400 13320 1452 13326
rect 1400 13262 1452 13268
rect 1320 13110 1440 13138
rect 1214 13087 1270 13096
rect 1228 12986 1256 13087
rect 1216 12980 1268 12986
rect 1216 12922 1268 12928
rect 1412 12646 1440 13110
rect 1400 12640 1452 12646
rect 1400 12582 1452 12588
rect 1504 12434 1532 13806
rect 1596 12442 1624 13903
rect 1780 13002 1808 14311
rect 1860 13796 1912 13802
rect 1860 13738 1912 13744
rect 1688 12974 1808 13002
rect 1044 12406 1164 12434
rect 952 2746 1072 2774
rect 940 1896 992 1902
rect 940 1838 992 1844
rect 952 160 980 1838
rect 1044 1290 1072 2746
rect 1136 1494 1164 12406
rect 1412 12406 1532 12434
rect 1584 12436 1636 12442
rect 1306 12064 1362 12073
rect 1412 12050 1440 12406
rect 1584 12378 1636 12384
rect 1492 12232 1544 12238
rect 1490 12200 1492 12209
rect 1544 12200 1546 12209
rect 1490 12135 1546 12144
rect 1412 12022 1532 12050
rect 1306 11999 1362 12008
rect 1320 11354 1348 11999
rect 1504 11694 1532 12022
rect 1492 11688 1544 11694
rect 1492 11630 1544 11636
rect 1582 11520 1638 11529
rect 1582 11455 1638 11464
rect 1308 11348 1360 11354
rect 1308 11290 1360 11296
rect 1308 8424 1360 8430
rect 1492 8424 1544 8430
rect 1308 8366 1360 8372
rect 1490 8392 1492 8401
rect 1544 8392 1546 8401
rect 1320 6118 1348 8366
rect 1490 8327 1546 8336
rect 1400 7404 1452 7410
rect 1400 7346 1452 7352
rect 1412 6254 1440 7346
rect 1596 7002 1624 11455
rect 1688 8498 1716 12974
rect 1766 12608 1822 12617
rect 1766 12543 1822 12552
rect 1780 9722 1808 12543
rect 1872 11898 1900 13738
rect 1964 13734 1992 16526
rect 2044 16244 2096 16250
rect 2044 16186 2096 16192
rect 1952 13728 2004 13734
rect 1952 13670 2004 13676
rect 2056 13258 2084 16186
rect 1952 13252 2004 13258
rect 1952 13194 2004 13200
rect 2044 13252 2096 13258
rect 2044 13194 2096 13200
rect 1860 11892 1912 11898
rect 1860 11834 1912 11840
rect 1860 11688 1912 11694
rect 1860 11630 1912 11636
rect 1872 10033 1900 11630
rect 1964 11014 1992 13194
rect 2148 12918 2176 17818
rect 2226 17368 2282 17377
rect 2226 17303 2282 17312
rect 2240 17202 2268 17303
rect 2228 17196 2280 17202
rect 2228 17138 2280 17144
rect 2516 17082 2544 19876
rect 2688 19858 2740 19864
rect 2792 19530 2820 22986
rect 2872 22432 2924 22438
rect 2872 22374 2924 22380
rect 2884 20754 2912 22374
rect 2976 21434 3004 25162
rect 3068 23662 3096 26386
rect 3148 26240 3200 26246
rect 3148 26182 3200 26188
rect 3160 23866 3188 26182
rect 3148 23860 3200 23866
rect 3148 23802 3200 23808
rect 3148 23724 3200 23730
rect 3148 23666 3200 23672
rect 3056 23656 3108 23662
rect 3056 23598 3108 23604
rect 3160 23322 3188 23666
rect 3148 23316 3200 23322
rect 3148 23258 3200 23264
rect 3252 22778 3280 27628
rect 3344 25498 3372 27814
rect 3332 25492 3384 25498
rect 3332 25434 3384 25440
rect 3240 22772 3292 22778
rect 3240 22714 3292 22720
rect 3252 22438 3280 22714
rect 3240 22432 3292 22438
rect 3240 22374 3292 22380
rect 3344 22094 3372 25434
rect 3436 24954 3464 29158
rect 3514 29064 3570 29073
rect 3514 28999 3570 29008
rect 3528 26790 3556 28999
rect 3620 26994 3648 30767
rect 3700 28960 3752 28966
rect 3700 28902 3752 28908
rect 3712 28558 3740 28902
rect 3700 28552 3752 28558
rect 3700 28494 3752 28500
rect 3712 28393 3740 28494
rect 3804 28490 3832 31300
rect 3976 31282 4028 31288
rect 3882 31036 4190 31045
rect 3882 31034 3888 31036
rect 3944 31034 3968 31036
rect 4024 31034 4048 31036
rect 4104 31034 4128 31036
rect 4184 31034 4190 31036
rect 3944 30982 3946 31034
rect 4126 30982 4128 31034
rect 3882 30980 3888 30982
rect 3944 30980 3968 30982
rect 4024 30980 4048 30982
rect 4104 30980 4128 30982
rect 4184 30980 4190 30982
rect 3882 30971 4190 30980
rect 3976 30932 4028 30938
rect 3976 30874 4028 30880
rect 3988 30190 4016 30874
rect 4160 30592 4212 30598
rect 4160 30534 4212 30540
rect 4172 30433 4200 30534
rect 4158 30424 4214 30433
rect 4158 30359 4214 30368
rect 4264 30258 4292 33238
rect 4342 33215 4398 33224
rect 4448 33153 4476 33458
rect 4434 33144 4490 33153
rect 4434 33079 4490 33088
rect 4344 32428 4396 32434
rect 4344 32370 4396 32376
rect 4356 30977 4384 32370
rect 4540 31736 4568 34886
rect 4632 34678 4660 34954
rect 4620 34672 4672 34678
rect 4620 34614 4672 34620
rect 4632 34406 4660 34614
rect 4620 34400 4672 34406
rect 4620 34342 4672 34348
rect 4724 33930 4752 35822
rect 4804 35624 4856 35630
rect 4804 35566 4856 35572
rect 4816 34678 4844 35566
rect 4908 34950 4936 35822
rect 4988 35760 5040 35766
rect 4988 35702 5040 35708
rect 5000 34950 5028 35702
rect 5092 35698 5120 35974
rect 5080 35692 5132 35698
rect 5080 35634 5132 35640
rect 4896 34944 4948 34950
rect 4896 34886 4948 34892
rect 4988 34944 5040 34950
rect 4988 34886 5040 34892
rect 4988 34740 5040 34746
rect 4988 34682 5040 34688
rect 4804 34672 4856 34678
rect 4804 34614 4856 34620
rect 4896 34604 4948 34610
rect 4896 34546 4948 34552
rect 4802 34504 4858 34513
rect 4802 34439 4858 34448
rect 4712 33924 4764 33930
rect 4712 33866 4764 33872
rect 4620 33856 4672 33862
rect 4620 33798 4672 33804
rect 4448 31708 4568 31736
rect 4448 31482 4476 31708
rect 4632 31634 4660 33798
rect 4540 31606 4660 31634
rect 4540 31482 4568 31606
rect 4436 31476 4488 31482
rect 4436 31418 4488 31424
rect 4528 31476 4580 31482
rect 4528 31418 4580 31424
rect 4434 31104 4490 31113
rect 4434 31039 4490 31048
rect 4342 30968 4398 30977
rect 4448 30938 4476 31039
rect 4342 30903 4398 30912
rect 4436 30932 4488 30938
rect 4252 30252 4304 30258
rect 4252 30194 4304 30200
rect 3976 30184 4028 30190
rect 3976 30126 4028 30132
rect 4066 30152 4122 30161
rect 4066 30087 4122 30096
rect 4080 30054 4108 30087
rect 4068 30048 4120 30054
rect 4068 29990 4120 29996
rect 3882 29948 4190 29957
rect 3882 29946 3888 29948
rect 3944 29946 3968 29948
rect 4024 29946 4048 29948
rect 4104 29946 4128 29948
rect 4184 29946 4190 29948
rect 3944 29894 3946 29946
rect 4126 29894 4128 29946
rect 3882 29892 3888 29894
rect 3944 29892 3968 29894
rect 4024 29892 4048 29894
rect 4104 29892 4128 29894
rect 4184 29892 4190 29894
rect 3882 29883 4190 29892
rect 4264 29186 4292 30194
rect 4172 29158 4292 29186
rect 4172 28966 4200 29158
rect 4252 29096 4304 29102
rect 4252 29038 4304 29044
rect 4160 28960 4212 28966
rect 4160 28902 4212 28908
rect 3882 28860 4190 28869
rect 3882 28858 3888 28860
rect 3944 28858 3968 28860
rect 4024 28858 4048 28860
rect 4104 28858 4128 28860
rect 4184 28858 4190 28860
rect 3944 28806 3946 28858
rect 4126 28806 4128 28858
rect 3882 28804 3888 28806
rect 3944 28804 3968 28806
rect 4024 28804 4048 28806
rect 4104 28804 4128 28806
rect 4184 28804 4190 28806
rect 3882 28795 4190 28804
rect 3792 28484 3844 28490
rect 3792 28426 3844 28432
rect 3698 28384 3754 28393
rect 3698 28319 3754 28328
rect 3700 28076 3752 28082
rect 3700 28018 3752 28024
rect 3712 27577 3740 28018
rect 3698 27568 3754 27577
rect 3698 27503 3754 27512
rect 3608 26988 3660 26994
rect 3608 26930 3660 26936
rect 3516 26784 3568 26790
rect 3516 26726 3568 26732
rect 3620 25786 3648 26930
rect 3804 26450 3832 28426
rect 3882 27772 4190 27781
rect 3882 27770 3888 27772
rect 3944 27770 3968 27772
rect 4024 27770 4048 27772
rect 4104 27770 4128 27772
rect 4184 27770 4190 27772
rect 3944 27718 3946 27770
rect 4126 27718 4128 27770
rect 3882 27716 3888 27718
rect 3944 27716 3968 27718
rect 4024 27716 4048 27718
rect 4104 27716 4128 27718
rect 4184 27716 4190 27718
rect 3882 27707 4190 27716
rect 4066 27568 4122 27577
rect 3896 27526 4066 27554
rect 3896 27441 3924 27526
rect 4066 27503 4122 27512
rect 4068 27464 4120 27470
rect 3882 27432 3938 27441
rect 4068 27406 4120 27412
rect 3882 27367 3938 27376
rect 3896 26994 3924 27367
rect 3976 27328 4028 27334
rect 3976 27270 4028 27276
rect 3988 26994 4016 27270
rect 3884 26988 3936 26994
rect 3884 26930 3936 26936
rect 3976 26988 4028 26994
rect 3976 26930 4028 26936
rect 4080 26790 4108 27406
rect 4068 26784 4120 26790
rect 4068 26726 4120 26732
rect 3882 26684 4190 26693
rect 3882 26682 3888 26684
rect 3944 26682 3968 26684
rect 4024 26682 4048 26684
rect 4104 26682 4128 26684
rect 4184 26682 4190 26684
rect 3944 26630 3946 26682
rect 4126 26630 4128 26682
rect 3882 26628 3888 26630
rect 3944 26628 3968 26630
rect 4024 26628 4048 26630
rect 4104 26628 4128 26630
rect 4184 26628 4190 26630
rect 3882 26619 4190 26628
rect 3792 26444 3844 26450
rect 3792 26386 3844 26392
rect 4158 26344 4214 26353
rect 4158 26279 4214 26288
rect 4172 25906 4200 26279
rect 4160 25900 4212 25906
rect 4160 25842 4212 25848
rect 3528 25758 3648 25786
rect 3528 25702 3556 25758
rect 3516 25696 3568 25702
rect 3516 25638 3568 25644
rect 3608 25696 3660 25702
rect 3608 25638 3660 25644
rect 3698 25664 3754 25673
rect 3424 24948 3476 24954
rect 3424 24890 3476 24896
rect 3422 24712 3478 24721
rect 3422 24647 3478 24656
rect 3436 24313 3464 24647
rect 3422 24304 3478 24313
rect 3422 24239 3478 24248
rect 3528 22778 3556 25638
rect 3620 24410 3648 25638
rect 3698 25599 3754 25608
rect 3608 24404 3660 24410
rect 3608 24346 3660 24352
rect 3712 23882 3740 25599
rect 3882 25596 4190 25605
rect 3882 25594 3888 25596
rect 3944 25594 3968 25596
rect 4024 25594 4048 25596
rect 4104 25594 4128 25596
rect 4184 25594 4190 25596
rect 3944 25542 3946 25594
rect 4126 25542 4128 25594
rect 3882 25540 3888 25542
rect 3944 25540 3968 25542
rect 4024 25540 4048 25542
rect 4104 25540 4128 25542
rect 4184 25540 4190 25542
rect 3882 25531 4190 25540
rect 4264 25158 4292 29038
rect 4356 26738 4384 30903
rect 4436 30874 4488 30880
rect 4436 30592 4488 30598
rect 4436 30534 4488 30540
rect 4448 29782 4476 30534
rect 4436 29776 4488 29782
rect 4436 29718 4488 29724
rect 4448 29102 4476 29718
rect 4436 29096 4488 29102
rect 4436 29038 4488 29044
rect 4436 28960 4488 28966
rect 4436 28902 4488 28908
rect 4448 28558 4476 28902
rect 4540 28558 4568 31418
rect 4620 31340 4672 31346
rect 4724 31328 4752 33866
rect 4816 32366 4844 34439
rect 4908 34241 4936 34546
rect 4894 34232 4950 34241
rect 4894 34167 4950 34176
rect 4894 33824 4950 33833
rect 4894 33759 4950 33768
rect 4908 33658 4936 33759
rect 4896 33652 4948 33658
rect 4896 33594 4948 33600
rect 4804 32360 4856 32366
rect 4804 32302 4856 32308
rect 4896 32360 4948 32366
rect 4896 32302 4948 32308
rect 4908 32042 4936 32302
rect 4816 32014 4936 32042
rect 4816 31414 4844 32014
rect 5000 31940 5028 34682
rect 5092 33862 5120 35634
rect 5184 35068 5212 36722
rect 5448 36168 5500 36174
rect 5368 36128 5448 36156
rect 5368 36009 5396 36128
rect 5448 36110 5500 36116
rect 5448 36032 5500 36038
rect 5354 36000 5410 36009
rect 5448 35974 5500 35980
rect 5354 35935 5410 35944
rect 5262 35728 5318 35737
rect 5262 35663 5264 35672
rect 5316 35663 5318 35672
rect 5264 35634 5316 35640
rect 5184 35040 5396 35068
rect 5172 34944 5224 34950
rect 5172 34886 5224 34892
rect 5264 34944 5316 34950
rect 5264 34886 5316 34892
rect 5080 33856 5132 33862
rect 5080 33798 5132 33804
rect 5184 32960 5212 34886
rect 5276 34202 5304 34886
rect 5264 34196 5316 34202
rect 5264 34138 5316 34144
rect 4908 31912 5028 31940
rect 5092 32932 5212 32960
rect 4804 31408 4856 31414
rect 4804 31350 4856 31356
rect 4672 31300 4752 31328
rect 4620 31282 4672 31288
rect 4618 30696 4674 30705
rect 4618 30631 4674 30640
rect 4632 30598 4660 30631
rect 4620 30592 4672 30598
rect 4620 30534 4672 30540
rect 4436 28552 4488 28558
rect 4436 28494 4488 28500
rect 4528 28552 4580 28558
rect 4528 28494 4580 28500
rect 4724 28490 4752 31300
rect 4804 31204 4856 31210
rect 4804 31146 4856 31152
rect 4816 31113 4844 31146
rect 4802 31104 4858 31113
rect 4802 31039 4858 31048
rect 4908 30954 4936 31912
rect 4988 31816 5040 31822
rect 4988 31758 5040 31764
rect 4816 30926 4936 30954
rect 4816 30841 4844 30926
rect 4802 30832 4858 30841
rect 4802 30767 4858 30776
rect 4896 30796 4948 30802
rect 4896 30738 4948 30744
rect 4804 30592 4856 30598
rect 4804 30534 4856 30540
rect 4816 30433 4844 30534
rect 4802 30424 4858 30433
rect 4908 30394 4936 30738
rect 4802 30359 4858 30368
rect 4896 30388 4948 30394
rect 4896 30330 4948 30336
rect 4804 30252 4856 30258
rect 4804 30194 4856 30200
rect 4816 29238 4844 30194
rect 4804 29232 4856 29238
rect 4804 29174 4856 29180
rect 4712 28484 4764 28490
rect 4712 28426 4764 28432
rect 4620 28416 4672 28422
rect 4620 28358 4672 28364
rect 4528 28144 4580 28150
rect 4528 28086 4580 28092
rect 4540 27849 4568 28086
rect 4526 27840 4582 27849
rect 4526 27775 4582 27784
rect 4356 26710 4568 26738
rect 4342 26616 4398 26625
rect 4342 26551 4398 26560
rect 4356 26450 4384 26551
rect 4436 26512 4488 26518
rect 4436 26454 4488 26460
rect 4344 26444 4396 26450
rect 4344 26386 4396 26392
rect 4252 25152 4304 25158
rect 4252 25094 4304 25100
rect 4250 24984 4306 24993
rect 4250 24919 4306 24928
rect 3792 24744 3844 24750
rect 3792 24686 3844 24692
rect 3804 24324 3832 24686
rect 3882 24508 4190 24517
rect 3882 24506 3888 24508
rect 3944 24506 3968 24508
rect 4024 24506 4048 24508
rect 4104 24506 4128 24508
rect 4184 24506 4190 24508
rect 3944 24454 3946 24506
rect 4126 24454 4128 24506
rect 3882 24452 3888 24454
rect 3944 24452 3968 24454
rect 4024 24452 4048 24454
rect 4104 24452 4128 24454
rect 4184 24452 4190 24454
rect 3882 24443 4190 24452
rect 3804 24296 3924 24324
rect 3620 23854 3740 23882
rect 3620 22982 3648 23854
rect 3700 23792 3752 23798
rect 3700 23734 3752 23740
rect 3608 22976 3660 22982
rect 3608 22918 3660 22924
rect 3516 22772 3568 22778
rect 3516 22714 3568 22720
rect 3528 22522 3556 22714
rect 3608 22636 3660 22642
rect 3608 22578 3660 22584
rect 3436 22494 3556 22522
rect 3436 22234 3464 22494
rect 3620 22386 3648 22578
rect 3528 22358 3648 22386
rect 3424 22228 3476 22234
rect 3424 22170 3476 22176
rect 3344 22066 3464 22094
rect 3332 21888 3384 21894
rect 3160 21848 3332 21876
rect 2976 21406 3096 21434
rect 2964 21344 3016 21350
rect 2964 21286 3016 21292
rect 2976 20942 3004 21286
rect 2964 20936 3016 20942
rect 2964 20878 3016 20884
rect 2884 20726 3004 20754
rect 2700 19502 2820 19530
rect 2594 19272 2650 19281
rect 2594 19207 2650 19216
rect 2608 18766 2636 19207
rect 2596 18760 2648 18766
rect 2596 18702 2648 18708
rect 2608 17513 2636 18702
rect 2594 17504 2650 17513
rect 2594 17439 2650 17448
rect 2596 17332 2648 17338
rect 2596 17274 2648 17280
rect 2240 17054 2544 17082
rect 2240 16250 2268 17054
rect 2608 16658 2636 17274
rect 2320 16652 2372 16658
rect 2596 16652 2648 16658
rect 2372 16612 2452 16640
rect 2320 16594 2372 16600
rect 2228 16244 2280 16250
rect 2228 16186 2280 16192
rect 2320 16108 2372 16114
rect 2320 16050 2372 16056
rect 2228 14816 2280 14822
rect 2228 14758 2280 14764
rect 2240 13870 2268 14758
rect 2332 14385 2360 16050
rect 2318 14376 2374 14385
rect 2318 14311 2374 14320
rect 2320 14272 2372 14278
rect 2320 14214 2372 14220
rect 2228 13864 2280 13870
rect 2228 13806 2280 13812
rect 2228 13184 2280 13190
rect 2228 13126 2280 13132
rect 2240 12918 2268 13126
rect 2136 12912 2188 12918
rect 2136 12854 2188 12860
rect 2228 12912 2280 12918
rect 2228 12854 2280 12860
rect 2332 11744 2360 14214
rect 2424 13938 2452 16612
rect 2596 16594 2648 16600
rect 2608 13938 2636 16594
rect 2700 14414 2728 19502
rect 2780 19372 2832 19378
rect 2780 19314 2832 19320
rect 2792 18873 2820 19314
rect 2778 18864 2834 18873
rect 2778 18799 2834 18808
rect 2872 18760 2924 18766
rect 2872 18702 2924 18708
rect 2884 18426 2912 18702
rect 2872 18420 2924 18426
rect 2872 18362 2924 18368
rect 2976 18329 3004 20726
rect 3068 20058 3096 21406
rect 3056 20052 3108 20058
rect 3056 19994 3108 20000
rect 3056 19304 3108 19310
rect 3056 19246 3108 19252
rect 3068 18834 3096 19246
rect 3056 18828 3108 18834
rect 3056 18770 3108 18776
rect 2778 18320 2834 18329
rect 2778 18255 2834 18264
rect 2962 18320 3018 18329
rect 2962 18255 3018 18264
rect 2792 17678 2820 18255
rect 2780 17672 2832 17678
rect 2780 17614 2832 17620
rect 2976 17082 3004 18255
rect 3068 17270 3096 18770
rect 3056 17264 3108 17270
rect 3056 17206 3108 17212
rect 2976 17054 3096 17082
rect 2964 16652 3016 16658
rect 2964 16594 3016 16600
rect 2780 16584 2832 16590
rect 2780 16526 2832 16532
rect 2792 16250 2820 16526
rect 2780 16244 2832 16250
rect 2780 16186 2832 16192
rect 2976 16182 3004 16594
rect 2964 16176 3016 16182
rect 2964 16118 3016 16124
rect 2780 15904 2832 15910
rect 3068 15892 3096 17054
rect 2780 15846 2832 15852
rect 2884 15864 3096 15892
rect 2688 14408 2740 14414
rect 2688 14350 2740 14356
rect 2412 13932 2464 13938
rect 2412 13874 2464 13880
rect 2596 13932 2648 13938
rect 2596 13874 2648 13880
rect 2424 12850 2452 13874
rect 2608 13376 2636 13874
rect 2688 13864 2740 13870
rect 2688 13806 2740 13812
rect 2700 13530 2728 13806
rect 2688 13524 2740 13530
rect 2688 13466 2740 13472
rect 2516 13348 2728 13376
rect 2412 12844 2464 12850
rect 2412 12786 2464 12792
rect 2424 11762 2452 12786
rect 2516 11762 2544 13348
rect 2700 13258 2728 13348
rect 2596 13252 2648 13258
rect 2596 13194 2648 13200
rect 2688 13252 2740 13258
rect 2688 13194 2740 13200
rect 2608 12238 2636 13194
rect 2688 12844 2740 12850
rect 2792 12832 2820 15846
rect 2884 13870 2912 15864
rect 2964 15428 3016 15434
rect 2964 15370 3016 15376
rect 2976 13977 3004 15370
rect 3054 15328 3110 15337
rect 3054 15263 3110 15272
rect 2962 13968 3018 13977
rect 2962 13903 3018 13912
rect 2872 13864 2924 13870
rect 2872 13806 2924 13812
rect 2872 13728 2924 13734
rect 2872 13670 2924 13676
rect 2884 12850 2912 13670
rect 2740 12804 2820 12832
rect 2872 12844 2924 12850
rect 2688 12786 2740 12792
rect 2872 12786 2924 12792
rect 2884 12646 2912 12786
rect 2872 12640 2924 12646
rect 2872 12582 2924 12588
rect 2596 12232 2648 12238
rect 2596 12174 2648 12180
rect 2240 11716 2360 11744
rect 2412 11756 2464 11762
rect 2136 11620 2188 11626
rect 2136 11562 2188 11568
rect 1952 11008 2004 11014
rect 1952 10950 2004 10956
rect 1858 10024 1914 10033
rect 1964 9994 1992 10950
rect 2148 10266 2176 11562
rect 2240 10674 2268 11716
rect 2412 11698 2464 11704
rect 2504 11756 2556 11762
rect 2504 11698 2556 11704
rect 2318 11656 2374 11665
rect 2318 11591 2374 11600
rect 2332 11150 2360 11591
rect 2516 11218 2544 11698
rect 2688 11688 2740 11694
rect 2688 11630 2740 11636
rect 2700 11354 2728 11630
rect 2780 11552 2832 11558
rect 2780 11494 2832 11500
rect 2688 11348 2740 11354
rect 2688 11290 2740 11296
rect 2504 11212 2556 11218
rect 2504 11154 2556 11160
rect 2320 11144 2372 11150
rect 2594 11112 2650 11121
rect 2320 11086 2372 11092
rect 2516 11070 2594 11098
rect 2412 10736 2464 10742
rect 2412 10678 2464 10684
rect 2228 10668 2280 10674
rect 2228 10610 2280 10616
rect 2136 10260 2188 10266
rect 2136 10202 2188 10208
rect 1858 9959 1914 9968
rect 1952 9988 2004 9994
rect 1952 9930 2004 9936
rect 1768 9716 1820 9722
rect 1964 9674 1992 9930
rect 1768 9658 1820 9664
rect 1872 9646 1992 9674
rect 1872 8974 1900 9646
rect 2136 9580 2188 9586
rect 2136 9522 2188 9528
rect 1860 8968 1912 8974
rect 1860 8910 1912 8916
rect 1676 8492 1728 8498
rect 1676 8434 1728 8440
rect 1688 7002 1716 8434
rect 1872 8090 1900 8910
rect 2044 8832 2096 8838
rect 2044 8774 2096 8780
rect 1950 8528 2006 8537
rect 1950 8463 2006 8472
rect 1964 8090 1992 8463
rect 2056 8430 2084 8774
rect 2148 8673 2176 9522
rect 2240 8974 2268 10610
rect 2320 9512 2372 9518
rect 2320 9454 2372 9460
rect 2228 8968 2280 8974
rect 2228 8910 2280 8916
rect 2332 8820 2360 9454
rect 2240 8792 2360 8820
rect 2134 8664 2190 8673
rect 2134 8599 2190 8608
rect 2044 8424 2096 8430
rect 2044 8366 2096 8372
rect 2136 8356 2188 8362
rect 2136 8298 2188 8304
rect 2044 8288 2096 8294
rect 2044 8230 2096 8236
rect 1860 8084 1912 8090
rect 1780 8044 1860 8072
rect 1780 7546 1808 8044
rect 1860 8026 1912 8032
rect 1952 8084 2004 8090
rect 1952 8026 2004 8032
rect 1858 7984 1914 7993
rect 2056 7970 2084 8230
rect 1858 7919 1914 7928
rect 1964 7942 2084 7970
rect 1768 7540 1820 7546
rect 1768 7482 1820 7488
rect 1584 6996 1636 7002
rect 1584 6938 1636 6944
rect 1676 6996 1728 7002
rect 1676 6938 1728 6944
rect 1490 6760 1546 6769
rect 1490 6695 1492 6704
rect 1544 6695 1546 6704
rect 1492 6666 1544 6672
rect 1400 6248 1452 6254
rect 1400 6190 1452 6196
rect 1308 6112 1360 6118
rect 1308 6054 1360 6060
rect 1412 5234 1440 6190
rect 1688 5778 1716 6938
rect 1676 5772 1728 5778
rect 1676 5714 1728 5720
rect 1674 5536 1730 5545
rect 1674 5471 1730 5480
rect 1688 5302 1716 5471
rect 1766 5400 1822 5409
rect 1766 5335 1822 5344
rect 1676 5296 1728 5302
rect 1676 5238 1728 5244
rect 1400 5228 1452 5234
rect 1400 5170 1452 5176
rect 1216 5024 1268 5030
rect 1216 4966 1268 4972
rect 1306 4992 1362 5001
rect 1124 1488 1176 1494
rect 1124 1430 1176 1436
rect 1032 1284 1084 1290
rect 1032 1226 1084 1232
rect 1228 160 1256 4966
rect 1306 4927 1362 4936
rect 1320 4826 1348 4927
rect 1308 4820 1360 4826
rect 1308 4762 1360 4768
rect 1412 4690 1440 5170
rect 1674 4720 1730 4729
rect 1400 4684 1452 4690
rect 1452 4644 1532 4672
rect 1674 4655 1730 4664
rect 1400 4626 1452 4632
rect 1400 4140 1452 4146
rect 1400 4082 1452 4088
rect 1412 2122 1440 4082
rect 1504 3602 1532 4644
rect 1688 4622 1716 4655
rect 1676 4616 1728 4622
rect 1676 4558 1728 4564
rect 1582 4040 1638 4049
rect 1582 3975 1638 3984
rect 1596 3738 1624 3975
rect 1584 3732 1636 3738
rect 1584 3674 1636 3680
rect 1492 3596 1544 3602
rect 1492 3538 1544 3544
rect 1504 2514 1532 3538
rect 1674 2952 1730 2961
rect 1674 2887 1730 2896
rect 1492 2508 1544 2514
rect 1492 2450 1544 2456
rect 1412 2094 1532 2122
rect 1504 160 1532 2094
rect 1688 2038 1716 2887
rect 1780 2650 1808 5335
rect 1872 3194 1900 7919
rect 1964 4214 1992 7942
rect 2148 6458 2176 8298
rect 2240 6662 2268 8792
rect 2320 8628 2372 8634
rect 2320 8570 2372 8576
rect 2228 6656 2280 6662
rect 2228 6598 2280 6604
rect 2136 6452 2188 6458
rect 2136 6394 2188 6400
rect 2136 5772 2188 5778
rect 2136 5714 2188 5720
rect 2148 4758 2176 5714
rect 2136 4752 2188 4758
rect 2136 4694 2188 4700
rect 2332 4570 2360 8570
rect 2424 8242 2452 10678
rect 2516 8378 2544 11070
rect 2594 11047 2650 11056
rect 2792 10810 2820 11494
rect 2962 11248 3018 11257
rect 2962 11183 3018 11192
rect 2870 10840 2926 10849
rect 2780 10804 2832 10810
rect 2870 10775 2926 10784
rect 2780 10746 2832 10752
rect 2778 10568 2834 10577
rect 2778 10503 2834 10512
rect 2792 9518 2820 10503
rect 2884 10266 2912 10775
rect 2976 10266 3004 11183
rect 2872 10260 2924 10266
rect 2872 10202 2924 10208
rect 2964 10260 3016 10266
rect 2964 10202 3016 10208
rect 2870 9888 2926 9897
rect 3068 9874 3096 15263
rect 3160 11150 3188 21848
rect 3332 21830 3384 21836
rect 3240 21480 3292 21486
rect 3240 21422 3292 21428
rect 3252 20913 3280 21422
rect 3238 20904 3294 20913
rect 3238 20839 3294 20848
rect 3332 20868 3384 20874
rect 3332 20810 3384 20816
rect 3240 19984 3292 19990
rect 3240 19926 3292 19932
rect 3252 19446 3280 19926
rect 3240 19440 3292 19446
rect 3240 19382 3292 19388
rect 3344 18714 3372 20810
rect 3436 20806 3464 22066
rect 3424 20800 3476 20806
rect 3424 20742 3476 20748
rect 3528 20618 3556 22358
rect 3608 22228 3660 22234
rect 3608 22170 3660 22176
rect 3620 22030 3648 22170
rect 3608 22024 3660 22030
rect 3608 21966 3660 21972
rect 3436 20590 3556 20618
rect 3436 20505 3464 20590
rect 3516 20528 3568 20534
rect 3422 20496 3478 20505
rect 3516 20470 3568 20476
rect 3422 20431 3478 20440
rect 3436 19689 3464 20431
rect 3528 19961 3556 20470
rect 3514 19952 3570 19961
rect 3514 19887 3570 19896
rect 3422 19680 3478 19689
rect 3422 19615 3478 19624
rect 3620 18834 3648 21966
rect 3712 21350 3740 23734
rect 3792 23724 3844 23730
rect 3792 23666 3844 23672
rect 3804 23118 3832 23666
rect 3896 23662 3924 24296
rect 4068 24200 4120 24206
rect 4068 24142 4120 24148
rect 4158 24168 4214 24177
rect 4080 23798 4108 24142
rect 4158 24103 4214 24112
rect 4068 23792 4120 23798
rect 4068 23734 4120 23740
rect 4172 23730 4200 24103
rect 4160 23724 4212 23730
rect 4160 23666 4212 23672
rect 3884 23656 3936 23662
rect 3884 23598 3936 23604
rect 3882 23420 4190 23429
rect 3882 23418 3888 23420
rect 3944 23418 3968 23420
rect 4024 23418 4048 23420
rect 4104 23418 4128 23420
rect 4184 23418 4190 23420
rect 3944 23366 3946 23418
rect 4126 23366 4128 23418
rect 3882 23364 3888 23366
rect 3944 23364 3968 23366
rect 4024 23364 4048 23366
rect 4104 23364 4128 23366
rect 4184 23364 4190 23366
rect 3882 23355 4190 23364
rect 3792 23112 3844 23118
rect 3792 23054 3844 23060
rect 3882 22332 4190 22341
rect 3882 22330 3888 22332
rect 3944 22330 3968 22332
rect 4024 22330 4048 22332
rect 4104 22330 4128 22332
rect 4184 22330 4190 22332
rect 3944 22278 3946 22330
rect 4126 22278 4128 22330
rect 3882 22276 3888 22278
rect 3944 22276 3968 22278
rect 4024 22276 4048 22278
rect 4104 22276 4128 22278
rect 4184 22276 4190 22278
rect 3882 22267 4190 22276
rect 4160 21888 4212 21894
rect 4160 21830 4212 21836
rect 3792 21684 3844 21690
rect 3792 21626 3844 21632
rect 3700 21344 3752 21350
rect 3700 21286 3752 21292
rect 3712 21078 3740 21286
rect 3700 21072 3752 21078
rect 3700 21014 3752 21020
rect 3700 20460 3752 20466
rect 3700 20402 3752 20408
rect 3608 18828 3660 18834
rect 3608 18770 3660 18776
rect 3344 18698 3648 18714
rect 3344 18692 3660 18698
rect 3344 18686 3608 18692
rect 3344 18154 3372 18686
rect 3608 18634 3660 18640
rect 3424 18624 3476 18630
rect 3424 18566 3476 18572
rect 3516 18624 3568 18630
rect 3516 18566 3568 18572
rect 3436 18426 3464 18566
rect 3424 18420 3476 18426
rect 3424 18362 3476 18368
rect 3332 18148 3384 18154
rect 3332 18090 3384 18096
rect 3240 18080 3292 18086
rect 3240 18022 3292 18028
rect 3252 17785 3280 18022
rect 3238 17776 3294 17785
rect 3238 17711 3294 17720
rect 3424 17536 3476 17542
rect 3424 17478 3476 17484
rect 3436 17241 3464 17478
rect 3422 17232 3478 17241
rect 3240 17196 3292 17202
rect 3422 17167 3478 17176
rect 3240 17138 3292 17144
rect 3252 15745 3280 17138
rect 3424 16652 3476 16658
rect 3424 16594 3476 16600
rect 3330 16416 3386 16425
rect 3330 16351 3386 16360
rect 3238 15736 3294 15745
rect 3344 15706 3372 16351
rect 3238 15671 3294 15680
rect 3332 15700 3384 15706
rect 3332 15642 3384 15648
rect 3240 13728 3292 13734
rect 3240 13670 3292 13676
rect 3148 11144 3200 11150
rect 3148 11086 3200 11092
rect 3148 11008 3200 11014
rect 3148 10950 3200 10956
rect 3160 10674 3188 10950
rect 3148 10668 3200 10674
rect 3148 10610 3200 10616
rect 3252 10062 3280 13670
rect 3332 12708 3384 12714
rect 3332 12650 3384 12656
rect 3344 12442 3372 12650
rect 3332 12436 3384 12442
rect 3332 12378 3384 12384
rect 3436 12186 3464 16594
rect 3344 12158 3464 12186
rect 3344 11642 3372 12158
rect 3424 12096 3476 12102
rect 3424 12038 3476 12044
rect 3436 11801 3464 12038
rect 3528 11898 3556 18566
rect 3608 18080 3660 18086
rect 3606 18048 3608 18057
rect 3660 18048 3662 18057
rect 3606 17983 3662 17992
rect 3712 17678 3740 20402
rect 3804 19417 3832 21626
rect 3974 21584 4030 21593
rect 3974 21519 4030 21528
rect 3988 21486 4016 21519
rect 3976 21480 4028 21486
rect 4172 21457 4200 21830
rect 3976 21422 4028 21428
rect 4158 21448 4214 21457
rect 4158 21383 4214 21392
rect 4172 21350 4200 21383
rect 4160 21344 4212 21350
rect 4160 21286 4212 21292
rect 3882 21244 4190 21253
rect 3882 21242 3888 21244
rect 3944 21242 3968 21244
rect 4024 21242 4048 21244
rect 4104 21242 4128 21244
rect 4184 21242 4190 21244
rect 3944 21190 3946 21242
rect 4126 21190 4128 21242
rect 3882 21188 3888 21190
rect 3944 21188 3968 21190
rect 4024 21188 4048 21190
rect 4104 21188 4128 21190
rect 4184 21188 4190 21190
rect 3882 21179 4190 21188
rect 4264 21146 4292 24919
rect 4356 23338 4384 26386
rect 4448 26042 4476 26454
rect 4436 26036 4488 26042
rect 4436 25978 4488 25984
rect 4434 25800 4490 25809
rect 4434 25735 4490 25744
rect 4448 23526 4476 25735
rect 4436 23520 4488 23526
rect 4436 23462 4488 23468
rect 4356 23310 4476 23338
rect 4344 22432 4396 22438
rect 4344 22374 4396 22380
rect 4356 21706 4384 22374
rect 4448 22137 4476 23310
rect 4434 22128 4490 22137
rect 4434 22063 4490 22072
rect 4434 21992 4490 22001
rect 4434 21927 4436 21936
rect 4488 21927 4490 21936
rect 4436 21898 4488 21904
rect 4356 21678 4476 21706
rect 4342 21584 4398 21593
rect 4342 21519 4398 21528
rect 4252 21140 4304 21146
rect 4252 21082 4304 21088
rect 4250 21040 4306 21049
rect 4356 21010 4384 21519
rect 4448 21418 4476 21678
rect 4436 21412 4488 21418
rect 4436 21354 4488 21360
rect 4250 20975 4306 20984
rect 4344 21004 4396 21010
rect 3882 20156 4190 20165
rect 3882 20154 3888 20156
rect 3944 20154 3968 20156
rect 4024 20154 4048 20156
rect 4104 20154 4128 20156
rect 4184 20154 4190 20156
rect 3944 20102 3946 20154
rect 4126 20102 4128 20154
rect 3882 20100 3888 20102
rect 3944 20100 3968 20102
rect 4024 20100 4048 20102
rect 4104 20100 4128 20102
rect 4184 20100 4190 20102
rect 3882 20091 4190 20100
rect 4068 20052 4120 20058
rect 4068 19994 4120 20000
rect 4080 19825 4108 19994
rect 4066 19816 4122 19825
rect 4066 19751 4122 19760
rect 3790 19408 3846 19417
rect 3790 19343 3846 19352
rect 4264 19334 4292 20975
rect 4344 20946 4396 20952
rect 4342 20632 4398 20641
rect 4342 20567 4398 20576
rect 4356 20466 4384 20567
rect 4344 20460 4396 20466
rect 4344 20402 4396 20408
rect 4540 19446 4568 26710
rect 4632 26058 4660 28358
rect 4724 26246 4752 28426
rect 4816 28150 4844 29174
rect 4896 28416 4948 28422
rect 4896 28358 4948 28364
rect 4804 28144 4856 28150
rect 4804 28086 4856 28092
rect 4908 27996 4936 28358
rect 4816 27968 4936 27996
rect 4712 26240 4764 26246
rect 4712 26182 4764 26188
rect 4632 26030 4752 26058
rect 4620 24336 4672 24342
rect 4620 24278 4672 24284
rect 4632 20913 4660 24278
rect 4724 23497 4752 26030
rect 4816 24721 4844 27968
rect 5000 27470 5028 31758
rect 5092 30258 5120 32932
rect 5172 32836 5224 32842
rect 5172 32778 5224 32784
rect 5184 32570 5212 32778
rect 5276 32570 5304 34138
rect 5368 32774 5396 35040
rect 5460 35018 5488 35974
rect 5552 35873 5580 40394
rect 5724 40384 5776 40390
rect 5724 40326 5776 40332
rect 5630 39944 5686 39953
rect 5630 39879 5632 39888
rect 5684 39879 5686 39888
rect 5632 39850 5684 39856
rect 5632 39296 5684 39302
rect 5632 39238 5684 39244
rect 5644 38010 5672 39238
rect 5736 38554 5764 40326
rect 5828 40225 5856 41074
rect 5920 40730 5948 41386
rect 6012 41274 6040 43794
rect 6196 43722 6224 44118
rect 6276 43988 6328 43994
rect 6276 43930 6328 43936
rect 6184 43716 6236 43722
rect 6184 43658 6236 43664
rect 6288 42548 6316 43930
rect 6104 42520 6316 42548
rect 6460 42560 6512 42566
rect 6000 41268 6052 41274
rect 6000 41210 6052 41216
rect 6000 40996 6052 41002
rect 6000 40938 6052 40944
rect 5908 40724 5960 40730
rect 5908 40666 5960 40672
rect 5908 40452 5960 40458
rect 5908 40394 5960 40400
rect 5814 40216 5870 40225
rect 5814 40151 5870 40160
rect 5920 39438 5948 40394
rect 5908 39432 5960 39438
rect 5908 39374 5960 39380
rect 5724 38548 5776 38554
rect 5724 38490 5776 38496
rect 5816 38412 5868 38418
rect 5816 38354 5868 38360
rect 5632 38004 5684 38010
rect 5632 37946 5684 37952
rect 5724 37800 5776 37806
rect 5724 37742 5776 37748
rect 5632 37188 5684 37194
rect 5632 37130 5684 37136
rect 5538 35864 5594 35873
rect 5538 35799 5594 35808
rect 5448 35012 5500 35018
rect 5448 34954 5500 34960
rect 5644 34950 5672 37130
rect 5736 36961 5764 37742
rect 5722 36952 5778 36961
rect 5722 36887 5778 36896
rect 5736 36106 5764 36887
rect 5724 36100 5776 36106
rect 5724 36042 5776 36048
rect 5724 35148 5776 35154
rect 5724 35090 5776 35096
rect 5632 34944 5684 34950
rect 5632 34886 5684 34892
rect 5736 34746 5764 35090
rect 5724 34740 5776 34746
rect 5724 34682 5776 34688
rect 5448 34400 5500 34406
rect 5448 34342 5500 34348
rect 5356 32768 5408 32774
rect 5356 32710 5408 32716
rect 5172 32564 5224 32570
rect 5172 32506 5224 32512
rect 5264 32564 5316 32570
rect 5264 32506 5316 32512
rect 5354 32464 5410 32473
rect 5354 32399 5410 32408
rect 5172 32020 5224 32026
rect 5172 31962 5224 31968
rect 5184 31346 5212 31962
rect 5368 31958 5396 32399
rect 5460 32026 5488 34342
rect 5632 33652 5684 33658
rect 5632 33594 5684 33600
rect 5540 33380 5592 33386
rect 5540 33322 5592 33328
rect 5448 32020 5500 32026
rect 5448 31962 5500 31968
rect 5356 31952 5408 31958
rect 5356 31894 5408 31900
rect 5354 31784 5410 31793
rect 5354 31719 5356 31728
rect 5408 31719 5410 31728
rect 5356 31690 5408 31696
rect 5264 31680 5316 31686
rect 5264 31622 5316 31628
rect 5354 31648 5410 31657
rect 5276 31346 5304 31622
rect 5354 31583 5410 31592
rect 5172 31340 5224 31346
rect 5172 31282 5224 31288
rect 5264 31340 5316 31346
rect 5264 31282 5316 31288
rect 5080 30252 5132 30258
rect 5080 30194 5132 30200
rect 5184 29696 5212 31282
rect 5262 30832 5318 30841
rect 5262 30767 5318 30776
rect 5276 30666 5304 30767
rect 5264 30660 5316 30666
rect 5264 30602 5316 30608
rect 5368 30258 5396 31583
rect 5552 31521 5580 33322
rect 5538 31512 5594 31521
rect 5538 31447 5594 31456
rect 5448 31408 5500 31414
rect 5448 31350 5500 31356
rect 5356 30252 5408 30258
rect 5356 30194 5408 30200
rect 5184 29668 5304 29696
rect 5172 29572 5224 29578
rect 5172 29514 5224 29520
rect 5184 29345 5212 29514
rect 5170 29336 5226 29345
rect 5170 29271 5226 29280
rect 5276 29238 5304 29668
rect 5264 29232 5316 29238
rect 5264 29174 5316 29180
rect 5264 28960 5316 28966
rect 5264 28902 5316 28908
rect 5276 28422 5304 28902
rect 5460 28558 5488 31350
rect 5540 30388 5592 30394
rect 5540 30330 5592 30336
rect 5448 28552 5500 28558
rect 5448 28494 5500 28500
rect 5264 28416 5316 28422
rect 5170 28384 5226 28393
rect 5264 28358 5316 28364
rect 5170 28319 5226 28328
rect 4988 27464 5040 27470
rect 4988 27406 5040 27412
rect 5000 27169 5028 27406
rect 5080 27328 5132 27334
rect 5080 27270 5132 27276
rect 4986 27160 5042 27169
rect 4986 27095 5042 27104
rect 4986 27024 5042 27033
rect 4908 26982 4986 27010
rect 4908 26194 4936 26982
rect 4986 26959 5042 26968
rect 4988 26784 5040 26790
rect 4988 26726 5040 26732
rect 5000 26382 5028 26726
rect 4988 26376 5040 26382
rect 4988 26318 5040 26324
rect 4908 26166 5028 26194
rect 4896 25832 4948 25838
rect 4896 25774 4948 25780
rect 4908 25294 4936 25774
rect 4896 25288 4948 25294
rect 4896 25230 4948 25236
rect 4802 24712 4858 24721
rect 4802 24647 4858 24656
rect 4804 24608 4856 24614
rect 4804 24550 4856 24556
rect 4816 24342 4844 24550
rect 4804 24336 4856 24342
rect 4804 24278 4856 24284
rect 4804 23792 4856 23798
rect 4804 23734 4856 23740
rect 4710 23488 4766 23497
rect 4710 23423 4766 23432
rect 4712 22636 4764 22642
rect 4712 22578 4764 22584
rect 4618 20904 4674 20913
rect 4618 20839 4674 20848
rect 4528 19440 4580 19446
rect 4528 19382 4580 19388
rect 4264 19306 4476 19334
rect 4252 19168 4304 19174
rect 4252 19110 4304 19116
rect 3882 19068 4190 19077
rect 3882 19066 3888 19068
rect 3944 19066 3968 19068
rect 4024 19066 4048 19068
rect 4104 19066 4128 19068
rect 4184 19066 4190 19068
rect 3944 19014 3946 19066
rect 4126 19014 4128 19066
rect 3882 19012 3888 19014
rect 3944 19012 3968 19014
rect 4024 19012 4048 19014
rect 4104 19012 4128 19014
rect 4184 19012 4190 19014
rect 3882 19003 4190 19012
rect 3790 18592 3846 18601
rect 3790 18527 3846 18536
rect 3700 17672 3752 17678
rect 3700 17614 3752 17620
rect 3608 16992 3660 16998
rect 3608 16934 3660 16940
rect 3620 16046 3648 16934
rect 3698 16688 3754 16697
rect 3698 16623 3754 16632
rect 3608 16040 3660 16046
rect 3608 15982 3660 15988
rect 3712 15162 3740 16623
rect 3804 16590 3832 18527
rect 4264 18222 4292 19110
rect 4252 18216 4304 18222
rect 4252 18158 4304 18164
rect 4344 18216 4396 18222
rect 4344 18158 4396 18164
rect 4252 18080 4304 18086
rect 4252 18022 4304 18028
rect 3882 17980 4190 17989
rect 3882 17978 3888 17980
rect 3944 17978 3968 17980
rect 4024 17978 4048 17980
rect 4104 17978 4128 17980
rect 4184 17978 4190 17980
rect 3944 17926 3946 17978
rect 4126 17926 4128 17978
rect 3882 17924 3888 17926
rect 3944 17924 3968 17926
rect 4024 17924 4048 17926
rect 4104 17924 4128 17926
rect 4184 17924 4190 17926
rect 3882 17915 4190 17924
rect 4264 17678 4292 18022
rect 4252 17672 4304 17678
rect 4252 17614 4304 17620
rect 4356 17542 4384 18158
rect 4344 17536 4396 17542
rect 4344 17478 4396 17484
rect 4356 17338 4384 17478
rect 4344 17332 4396 17338
rect 4344 17274 4396 17280
rect 4066 17232 4122 17241
rect 4066 17167 4068 17176
rect 4120 17167 4122 17176
rect 4068 17138 4120 17144
rect 4448 17082 4476 19306
rect 4526 19000 4582 19009
rect 4526 18935 4582 18944
rect 4540 18766 4568 18935
rect 4528 18760 4580 18766
rect 4528 18702 4580 18708
rect 4264 17054 4476 17082
rect 3882 16892 4190 16901
rect 3882 16890 3888 16892
rect 3944 16890 3968 16892
rect 4024 16890 4048 16892
rect 4104 16890 4128 16892
rect 4184 16890 4190 16892
rect 3944 16838 3946 16890
rect 4126 16838 4128 16890
rect 3882 16836 3888 16838
rect 3944 16836 3968 16838
rect 4024 16836 4048 16838
rect 4104 16836 4128 16838
rect 4184 16836 4190 16838
rect 3882 16827 4190 16836
rect 4264 16640 4292 17054
rect 4436 16992 4488 16998
rect 4436 16934 4488 16940
rect 4172 16612 4292 16640
rect 3792 16584 3844 16590
rect 3792 16526 3844 16532
rect 3884 16584 3936 16590
rect 3884 16526 3936 16532
rect 3792 15904 3844 15910
rect 3896 15892 3924 16526
rect 4172 16289 4200 16612
rect 4344 16584 4396 16590
rect 4250 16552 4306 16561
rect 4344 16526 4396 16532
rect 4250 16487 4306 16496
rect 4264 16454 4292 16487
rect 4252 16448 4304 16454
rect 4252 16390 4304 16396
rect 4158 16280 4214 16289
rect 4356 16250 4384 16526
rect 4158 16215 4214 16224
rect 4344 16244 4396 16250
rect 4172 16114 4200 16215
rect 4344 16186 4396 16192
rect 4448 16114 4476 16934
rect 4160 16108 4212 16114
rect 4160 16050 4212 16056
rect 4436 16108 4488 16114
rect 4436 16050 4488 16056
rect 3844 15864 3924 15892
rect 4252 15904 4304 15910
rect 3792 15846 3844 15852
rect 4252 15846 4304 15852
rect 3804 15688 3832 15846
rect 3882 15804 4190 15813
rect 3882 15802 3888 15804
rect 3944 15802 3968 15804
rect 4024 15802 4048 15804
rect 4104 15802 4128 15804
rect 4184 15802 4190 15804
rect 3944 15750 3946 15802
rect 4126 15750 4128 15802
rect 3882 15748 3888 15750
rect 3944 15748 3968 15750
rect 4024 15748 4048 15750
rect 4104 15748 4128 15750
rect 4184 15748 4190 15750
rect 3882 15739 4190 15748
rect 3804 15660 3924 15688
rect 3896 15609 3924 15660
rect 3882 15600 3938 15609
rect 3882 15535 3938 15544
rect 3700 15156 3752 15162
rect 3700 15098 3752 15104
rect 3700 15020 3752 15026
rect 3700 14962 3752 14968
rect 3606 13696 3662 13705
rect 3606 13631 3662 13640
rect 3620 12986 3648 13631
rect 3712 13394 3740 14962
rect 4158 14920 4214 14929
rect 3792 14884 3844 14890
rect 4158 14855 4160 14864
rect 3792 14826 3844 14832
rect 4212 14855 4214 14864
rect 4160 14826 4212 14832
rect 3804 13734 3832 14826
rect 3882 14716 4190 14725
rect 3882 14714 3888 14716
rect 3944 14714 3968 14716
rect 4024 14714 4048 14716
rect 4104 14714 4128 14716
rect 4184 14714 4190 14716
rect 3944 14662 3946 14714
rect 4126 14662 4128 14714
rect 3882 14660 3888 14662
rect 3944 14660 3968 14662
rect 4024 14660 4048 14662
rect 4104 14660 4128 14662
rect 4184 14660 4190 14662
rect 3882 14651 4190 14660
rect 3976 14612 4028 14618
rect 3976 14554 4028 14560
rect 3988 14521 4016 14554
rect 4160 14544 4212 14550
rect 3974 14512 4030 14521
rect 4160 14486 4212 14492
rect 3974 14447 4030 14456
rect 4172 14385 4200 14486
rect 4158 14376 4214 14385
rect 4158 14311 4214 14320
rect 3792 13728 3844 13734
rect 3792 13670 3844 13676
rect 3804 13394 3832 13670
rect 3882 13628 4190 13637
rect 3882 13626 3888 13628
rect 3944 13626 3968 13628
rect 4024 13626 4048 13628
rect 4104 13626 4128 13628
rect 4184 13626 4190 13628
rect 3944 13574 3946 13626
rect 4126 13574 4128 13626
rect 3882 13572 3888 13574
rect 3944 13572 3968 13574
rect 4024 13572 4048 13574
rect 4104 13572 4128 13574
rect 4184 13572 4190 13574
rect 3882 13563 4190 13572
rect 3700 13388 3752 13394
rect 3700 13330 3752 13336
rect 3792 13388 3844 13394
rect 3792 13330 3844 13336
rect 3700 13252 3752 13258
rect 3700 13194 3752 13200
rect 3608 12980 3660 12986
rect 3608 12922 3660 12928
rect 3606 12880 3662 12889
rect 3712 12850 3740 13194
rect 3606 12815 3662 12824
rect 3700 12844 3752 12850
rect 3516 11892 3568 11898
rect 3516 11834 3568 11840
rect 3422 11792 3478 11801
rect 3422 11727 3478 11736
rect 3344 11614 3464 11642
rect 3332 11552 3384 11558
rect 3332 11494 3384 11500
rect 3240 10056 3292 10062
rect 3240 9998 3292 10004
rect 2926 9846 3004 9874
rect 3068 9846 3188 9874
rect 2870 9823 2926 9832
rect 2872 9716 2924 9722
rect 2872 9658 2924 9664
rect 2780 9512 2832 9518
rect 2780 9454 2832 9460
rect 2792 8838 2820 9454
rect 2884 9450 2912 9658
rect 2872 9444 2924 9450
rect 2872 9386 2924 9392
rect 2780 8832 2832 8838
rect 2780 8774 2832 8780
rect 2688 8492 2740 8498
rect 2688 8434 2740 8440
rect 2516 8350 2636 8378
rect 2424 8214 2544 8242
rect 2516 7886 2544 8214
rect 2504 7880 2556 7886
rect 2504 7822 2556 7828
rect 2608 7528 2636 8350
rect 2700 7546 2728 8434
rect 2870 7848 2926 7857
rect 2792 7806 2870 7834
rect 2516 7500 2636 7528
rect 2688 7540 2740 7546
rect 2412 6112 2464 6118
rect 2412 6054 2464 6060
rect 2424 5778 2452 6054
rect 2412 5772 2464 5778
rect 2412 5714 2464 5720
rect 2410 5128 2466 5137
rect 2410 5063 2466 5072
rect 2148 4542 2360 4570
rect 1952 4208 2004 4214
rect 1952 4150 2004 4156
rect 2044 4208 2096 4214
rect 2044 4150 2096 4156
rect 1952 3936 2004 3942
rect 1950 3904 1952 3913
rect 2004 3904 2006 3913
rect 1950 3839 2006 3848
rect 1860 3188 1912 3194
rect 1860 3130 1912 3136
rect 1768 2644 1820 2650
rect 1768 2586 1820 2592
rect 1676 2032 1728 2038
rect 1676 1974 1728 1980
rect 1952 1284 2004 1290
rect 1952 1226 2004 1232
rect 1964 626 1992 1226
rect 1780 598 1992 626
rect 1780 160 1808 598
rect 2056 160 2084 4150
rect 2148 2446 2176 4542
rect 2228 4276 2280 4282
rect 2228 4218 2280 4224
rect 2240 3058 2268 4218
rect 2320 3392 2372 3398
rect 2320 3334 2372 3340
rect 2228 3052 2280 3058
rect 2228 2994 2280 3000
rect 2136 2440 2188 2446
rect 2136 2382 2188 2388
rect 2136 1216 2188 1222
rect 2134 1184 2136 1193
rect 2188 1184 2190 1193
rect 2134 1119 2190 1128
rect 2332 160 2360 3334
rect 2424 2378 2452 5063
rect 2516 4146 2544 7500
rect 2688 7482 2740 7488
rect 2596 6792 2648 6798
rect 2596 6734 2648 6740
rect 2608 6497 2636 6734
rect 2594 6488 2650 6497
rect 2792 6458 2820 7806
rect 2870 7783 2926 7792
rect 2870 6624 2926 6633
rect 2870 6559 2926 6568
rect 2594 6423 2650 6432
rect 2780 6452 2832 6458
rect 2780 6394 2832 6400
rect 2594 6352 2650 6361
rect 2594 6287 2650 6296
rect 2608 4758 2636 6287
rect 2778 5808 2834 5817
rect 2778 5743 2834 5752
rect 2688 5704 2740 5710
rect 2688 5646 2740 5652
rect 2700 5370 2728 5646
rect 2688 5364 2740 5370
rect 2688 5306 2740 5312
rect 2596 4752 2648 4758
rect 2596 4694 2648 4700
rect 2596 4616 2648 4622
rect 2596 4558 2648 4564
rect 2504 4140 2556 4146
rect 2504 4082 2556 4088
rect 2412 2372 2464 2378
rect 2412 2314 2464 2320
rect 2412 1216 2464 1222
rect 2412 1158 2464 1164
rect 2424 610 2452 1158
rect 2412 604 2464 610
rect 2412 546 2464 552
rect 2608 160 2636 4558
rect 2686 4312 2742 4321
rect 2686 4247 2742 4256
rect 2700 4146 2728 4247
rect 2688 4140 2740 4146
rect 2688 4082 2740 4088
rect 2700 2990 2728 4082
rect 2688 2984 2740 2990
rect 2688 2926 2740 2932
rect 2688 2644 2740 2650
rect 2688 2586 2740 2592
rect 2700 1970 2728 2586
rect 2792 2038 2820 5743
rect 2884 3058 2912 6559
rect 2976 4010 3004 9846
rect 3056 9444 3108 9450
rect 3056 9386 3108 9392
rect 3068 9178 3096 9386
rect 3056 9172 3108 9178
rect 3056 9114 3108 9120
rect 3056 8900 3108 8906
rect 3056 8842 3108 8848
rect 3068 8430 3096 8842
rect 3056 8424 3108 8430
rect 3056 8366 3108 8372
rect 3054 8256 3110 8265
rect 3054 8191 3110 8200
rect 2964 4004 3016 4010
rect 2964 3946 3016 3952
rect 2962 3904 3018 3913
rect 2962 3839 3018 3848
rect 2976 3534 3004 3839
rect 3068 3670 3096 8191
rect 3160 7478 3188 9846
rect 3240 9716 3292 9722
rect 3240 9658 3292 9664
rect 3252 8786 3280 9658
rect 3344 8974 3372 11494
rect 3332 8968 3384 8974
rect 3436 8945 3464 11614
rect 3620 11354 3648 12815
rect 3700 12786 3752 12792
rect 3700 12436 3752 12442
rect 3700 12378 3752 12384
rect 3712 12345 3740 12378
rect 3698 12336 3754 12345
rect 3804 12306 3832 13330
rect 4264 13274 4292 15846
rect 4436 15156 4488 15162
rect 4436 15098 4488 15104
rect 4344 15088 4396 15094
rect 4344 15030 4396 15036
rect 4356 13326 4384 15030
rect 4448 14414 4476 15098
rect 4540 15094 4568 18702
rect 4724 17678 4752 22578
rect 4816 20534 4844 23734
rect 4908 22574 4936 25230
rect 4896 22568 4948 22574
rect 4896 22510 4948 22516
rect 4908 22234 4936 22510
rect 4896 22228 4948 22234
rect 4896 22170 4948 22176
rect 5000 22030 5028 26166
rect 5092 24886 5120 27270
rect 5184 26790 5212 28319
rect 5276 28082 5304 28358
rect 5264 28076 5316 28082
rect 5264 28018 5316 28024
rect 5172 26784 5224 26790
rect 5172 26726 5224 26732
rect 5170 26208 5226 26217
rect 5170 26143 5226 26152
rect 5184 25906 5212 26143
rect 5172 25900 5224 25906
rect 5172 25842 5224 25848
rect 5172 25152 5224 25158
rect 5172 25094 5224 25100
rect 5080 24880 5132 24886
rect 5080 24822 5132 24828
rect 5184 24410 5212 25094
rect 5172 24404 5224 24410
rect 5172 24346 5224 24352
rect 5172 24200 5224 24206
rect 5172 24142 5224 24148
rect 5080 23724 5132 23730
rect 5080 23666 5132 23672
rect 4988 22024 5040 22030
rect 4988 21966 5040 21972
rect 4896 21956 4948 21962
rect 4896 21898 4948 21904
rect 4804 20528 4856 20534
rect 4804 20470 4856 20476
rect 4816 18970 4844 20470
rect 4908 20040 4936 21898
rect 4988 21888 5040 21894
rect 4988 21830 5040 21836
rect 5000 21554 5028 21830
rect 4988 21548 5040 21554
rect 4988 21490 5040 21496
rect 4908 20012 5028 20040
rect 4896 19916 4948 19922
rect 4896 19858 4948 19864
rect 4908 19378 4936 19858
rect 4896 19372 4948 19378
rect 4896 19314 4948 19320
rect 4804 18964 4856 18970
rect 4804 18906 4856 18912
rect 4804 18624 4856 18630
rect 4804 18566 4856 18572
rect 4816 18290 4844 18566
rect 4804 18284 4856 18290
rect 4804 18226 4856 18232
rect 4712 17672 4764 17678
rect 4712 17614 4764 17620
rect 4724 17354 4752 17614
rect 4620 17332 4672 17338
rect 4724 17326 4936 17354
rect 4620 17274 4672 17280
rect 4632 16726 4660 17274
rect 4712 17128 4764 17134
rect 4712 17070 4764 17076
rect 4620 16720 4672 16726
rect 4618 16688 4620 16697
rect 4672 16688 4674 16697
rect 4618 16623 4674 16632
rect 4724 16504 4752 17070
rect 4678 16476 4752 16504
rect 4678 16402 4706 16476
rect 4678 16374 4752 16402
rect 4724 15502 4752 16374
rect 4908 16266 4936 17326
rect 4816 16238 4936 16266
rect 4816 15502 4844 16238
rect 4712 15496 4764 15502
rect 4712 15438 4764 15444
rect 4804 15496 4856 15502
rect 4804 15438 4856 15444
rect 4528 15088 4580 15094
rect 4528 15030 4580 15036
rect 4528 14952 4580 14958
rect 4580 14912 4660 14940
rect 4528 14894 4580 14900
rect 4436 14408 4488 14414
rect 4436 14350 4488 14356
rect 4528 14340 4580 14346
rect 4528 14282 4580 14288
rect 4436 13728 4488 13734
rect 4436 13670 4488 13676
rect 4080 13246 4292 13274
rect 4344 13320 4396 13326
rect 4344 13262 4396 13268
rect 4080 12866 4108 13246
rect 4080 12838 4292 12866
rect 3882 12540 4190 12549
rect 3882 12538 3888 12540
rect 3944 12538 3968 12540
rect 4024 12538 4048 12540
rect 4104 12538 4128 12540
rect 4184 12538 4190 12540
rect 3944 12486 3946 12538
rect 4126 12486 4128 12538
rect 3882 12484 3888 12486
rect 3944 12484 3968 12486
rect 4024 12484 4048 12486
rect 4104 12484 4128 12486
rect 4184 12484 4190 12486
rect 3882 12475 4190 12484
rect 3698 12271 3754 12280
rect 3792 12300 3844 12306
rect 3792 12242 3844 12248
rect 3700 11688 3752 11694
rect 3700 11630 3752 11636
rect 3608 11348 3660 11354
rect 3608 11290 3660 11296
rect 3712 11234 3740 11630
rect 3620 11218 3740 11234
rect 3608 11212 3740 11218
rect 3660 11206 3740 11212
rect 3608 11154 3660 11160
rect 3620 10690 3648 11154
rect 3528 10662 3648 10690
rect 3698 10704 3754 10713
rect 3528 9722 3556 10662
rect 3698 10639 3754 10648
rect 3606 10432 3662 10441
rect 3606 10367 3662 10376
rect 3620 10266 3648 10367
rect 3608 10260 3660 10266
rect 3608 10202 3660 10208
rect 3712 10198 3740 10639
rect 3804 10248 3832 12242
rect 3882 11452 4190 11461
rect 3882 11450 3888 11452
rect 3944 11450 3968 11452
rect 4024 11450 4048 11452
rect 4104 11450 4128 11452
rect 4184 11450 4190 11452
rect 3944 11398 3946 11450
rect 4126 11398 4128 11450
rect 3882 11396 3888 11398
rect 3944 11396 3968 11398
rect 4024 11396 4048 11398
rect 4104 11396 4128 11398
rect 4184 11396 4190 11398
rect 3882 11387 4190 11396
rect 4264 11082 4292 12838
rect 4448 12782 4476 13670
rect 4540 12782 4568 14282
rect 4632 13734 4660 14912
rect 4620 13728 4672 13734
rect 4620 13670 4672 13676
rect 4436 12776 4488 12782
rect 4436 12718 4488 12724
rect 4528 12776 4580 12782
rect 4528 12718 4580 12724
rect 4344 12708 4396 12714
rect 4344 12650 4396 12656
rect 4252 11076 4304 11082
rect 4252 11018 4304 11024
rect 4356 11014 4384 12650
rect 4528 12640 4580 12646
rect 4434 12608 4490 12617
rect 4580 12600 4660 12628
rect 4528 12582 4580 12588
rect 4434 12543 4490 12552
rect 3884 11008 3936 11014
rect 3976 11008 4028 11014
rect 3884 10950 3936 10956
rect 3974 10976 3976 10985
rect 4344 11008 4396 11014
rect 4028 10976 4030 10985
rect 3896 10742 3924 10950
rect 3974 10911 4030 10920
rect 4158 10976 4214 10985
rect 4344 10950 4396 10956
rect 4158 10911 4214 10920
rect 4172 10810 4200 10911
rect 4160 10804 4212 10810
rect 4160 10746 4212 10752
rect 3884 10736 3936 10742
rect 3884 10678 3936 10684
rect 3882 10364 4190 10373
rect 3882 10362 3888 10364
rect 3944 10362 3968 10364
rect 4024 10362 4048 10364
rect 4104 10362 4128 10364
rect 4184 10362 4190 10364
rect 3944 10310 3946 10362
rect 4126 10310 4128 10362
rect 3882 10308 3888 10310
rect 3944 10308 3968 10310
rect 4024 10308 4048 10310
rect 4104 10308 4128 10310
rect 4184 10308 4190 10310
rect 3882 10299 4190 10308
rect 3804 10220 3924 10248
rect 3700 10192 3752 10198
rect 3700 10134 3752 10140
rect 3792 9988 3844 9994
rect 3792 9930 3844 9936
rect 3698 9888 3754 9897
rect 3698 9823 3754 9832
rect 3516 9716 3568 9722
rect 3516 9658 3568 9664
rect 3608 9580 3660 9586
rect 3608 9522 3660 9528
rect 3516 9512 3568 9518
rect 3516 9454 3568 9460
rect 3332 8910 3384 8916
rect 3422 8936 3478 8945
rect 3528 8906 3556 9454
rect 3422 8871 3478 8880
rect 3516 8900 3568 8906
rect 3516 8842 3568 8848
rect 3514 8800 3570 8809
rect 3252 8758 3464 8786
rect 3240 8560 3292 8566
rect 3238 8528 3240 8537
rect 3292 8528 3294 8537
rect 3238 8463 3294 8472
rect 3148 7472 3200 7478
rect 3148 7414 3200 7420
rect 3146 7304 3202 7313
rect 3146 7239 3202 7248
rect 3160 5250 3188 7239
rect 3240 6656 3292 6662
rect 3240 6598 3292 6604
rect 3332 6656 3384 6662
rect 3332 6598 3384 6604
rect 3252 6458 3280 6598
rect 3240 6452 3292 6458
rect 3240 6394 3292 6400
rect 3344 6254 3372 6598
rect 3332 6248 3384 6254
rect 3238 6216 3294 6225
rect 3436 6225 3464 8758
rect 3514 8735 3570 8744
rect 3528 7410 3556 8735
rect 3620 8090 3648 9522
rect 3712 8498 3740 9823
rect 3804 9194 3832 9930
rect 3896 9364 3924 10220
rect 4066 10160 4122 10169
rect 4066 10095 4122 10104
rect 4344 10124 4396 10130
rect 4080 9722 4108 10095
rect 4344 10066 4396 10072
rect 4160 9920 4212 9926
rect 4160 9862 4212 9868
rect 4068 9716 4120 9722
rect 4068 9658 4120 9664
rect 4066 9616 4122 9625
rect 4172 9602 4200 9862
rect 4356 9625 4384 10066
rect 4122 9574 4200 9602
rect 4342 9616 4398 9625
rect 4066 9551 4122 9560
rect 4342 9551 4398 9560
rect 4344 9376 4396 9382
rect 3896 9336 4292 9364
rect 3882 9276 4190 9285
rect 3882 9274 3888 9276
rect 3944 9274 3968 9276
rect 4024 9274 4048 9276
rect 4104 9274 4128 9276
rect 4184 9274 4190 9276
rect 3944 9222 3946 9274
rect 4126 9222 4128 9274
rect 3882 9220 3888 9222
rect 3944 9220 3968 9222
rect 4024 9220 4048 9222
rect 4104 9220 4128 9222
rect 4184 9220 4190 9222
rect 3882 9211 4190 9220
rect 3804 9178 3857 9194
rect 3792 9172 3857 9178
rect 3844 9132 3857 9172
rect 3792 9114 3844 9120
rect 4068 8968 4120 8974
rect 4068 8910 4120 8916
rect 3700 8492 3752 8498
rect 3700 8434 3752 8440
rect 3792 8424 3844 8430
rect 3792 8366 3844 8372
rect 3882 8392 3938 8401
rect 3608 8084 3660 8090
rect 3608 8026 3660 8032
rect 3606 7984 3662 7993
rect 3606 7919 3608 7928
rect 3660 7919 3662 7928
rect 3608 7890 3660 7896
rect 3516 7404 3568 7410
rect 3516 7346 3568 7352
rect 3514 7168 3570 7177
rect 3514 7103 3570 7112
rect 3332 6190 3384 6196
rect 3422 6216 3478 6225
rect 3238 6151 3240 6160
rect 3292 6151 3294 6160
rect 3422 6151 3478 6160
rect 3240 6122 3292 6128
rect 3238 6080 3294 6089
rect 3238 6015 3294 6024
rect 3252 5370 3280 6015
rect 3424 5704 3476 5710
rect 3424 5646 3476 5652
rect 3240 5364 3292 5370
rect 3240 5306 3292 5312
rect 3160 5222 3280 5250
rect 3148 4684 3200 4690
rect 3148 4626 3200 4632
rect 3056 3664 3108 3670
rect 3056 3606 3108 3612
rect 2964 3528 3016 3534
rect 2964 3470 3016 3476
rect 2872 3052 2924 3058
rect 2872 2994 2924 3000
rect 2780 2032 2832 2038
rect 2780 1974 2832 1980
rect 2688 1964 2740 1970
rect 2688 1906 2740 1912
rect 2872 1284 2924 1290
rect 2872 1226 2924 1232
rect 2780 1216 2832 1222
rect 2780 1158 2832 1164
rect 2792 921 2820 1158
rect 2778 912 2834 921
rect 2778 847 2834 856
rect 2884 160 2912 1226
rect 3160 160 3188 4626
rect 3252 4185 3280 5222
rect 3238 4176 3294 4185
rect 3238 4111 3294 4120
rect 3238 4040 3294 4049
rect 3238 3975 3240 3984
rect 3292 3975 3294 3984
rect 3332 4004 3384 4010
rect 3240 3946 3292 3952
rect 3332 3946 3384 3952
rect 3252 2922 3280 3946
rect 3344 3738 3372 3946
rect 3332 3732 3384 3738
rect 3332 3674 3384 3680
rect 3436 3534 3464 5646
rect 3528 5370 3556 7103
rect 3804 6322 3832 8366
rect 3882 8327 3884 8336
rect 3936 8327 3938 8336
rect 3884 8298 3936 8304
rect 4080 8294 4108 8910
rect 4264 8838 4292 9336
rect 4344 9318 4396 9324
rect 4252 8832 4304 8838
rect 4252 8774 4304 8780
rect 4068 8288 4120 8294
rect 4068 8230 4120 8236
rect 3882 8188 4190 8197
rect 3882 8186 3888 8188
rect 3944 8186 3968 8188
rect 4024 8186 4048 8188
rect 4104 8186 4128 8188
rect 4184 8186 4190 8188
rect 3944 8134 3946 8186
rect 4126 8134 4128 8186
rect 3882 8132 3888 8134
rect 3944 8132 3968 8134
rect 4024 8132 4048 8134
rect 4104 8132 4128 8134
rect 4184 8132 4190 8134
rect 3882 8123 4190 8132
rect 4264 8090 4292 8774
rect 4252 8084 4304 8090
rect 4252 8026 4304 8032
rect 4068 7880 4120 7886
rect 4066 7848 4068 7857
rect 4120 7848 4122 7857
rect 4066 7783 4122 7792
rect 4068 7744 4120 7750
rect 4066 7712 4068 7721
rect 4120 7712 4122 7721
rect 4066 7647 4122 7656
rect 4068 7540 4120 7546
rect 4068 7482 4120 7488
rect 4080 7449 4108 7482
rect 4160 7472 4212 7478
rect 4066 7440 4122 7449
rect 4160 7414 4212 7420
rect 4066 7375 4122 7384
rect 4172 7290 4200 7414
rect 4264 7410 4292 8026
rect 4356 7818 4384 9318
rect 4448 8974 4476 12543
rect 4632 12050 4660 12600
rect 4724 12238 4752 15438
rect 5000 14929 5028 20012
rect 5092 19378 5120 23666
rect 5184 21350 5212 24142
rect 5172 21344 5224 21350
rect 5172 21286 5224 21292
rect 5170 20768 5226 20777
rect 5170 20703 5226 20712
rect 5080 19372 5132 19378
rect 5080 19314 5132 19320
rect 4986 14920 5042 14929
rect 4986 14855 5042 14864
rect 5092 14600 5120 19314
rect 5184 17338 5212 20703
rect 5276 18834 5304 28018
rect 5460 27674 5488 28494
rect 5448 27668 5500 27674
rect 5448 27610 5500 27616
rect 5356 26852 5408 26858
rect 5356 26794 5408 26800
rect 5368 24886 5396 26794
rect 5460 26518 5488 27610
rect 5448 26512 5500 26518
rect 5448 26454 5500 26460
rect 5460 25294 5488 26454
rect 5448 25288 5500 25294
rect 5448 25230 5500 25236
rect 5356 24880 5408 24886
rect 5356 24822 5408 24828
rect 5448 24200 5500 24206
rect 5448 24142 5500 24148
rect 5460 23526 5488 24142
rect 5448 23520 5500 23526
rect 5448 23462 5500 23468
rect 5356 22228 5408 22234
rect 5356 22170 5408 22176
rect 5368 19922 5396 22170
rect 5552 21944 5580 30330
rect 5644 29730 5672 33594
rect 5828 32042 5856 38354
rect 5920 37194 5948 39374
rect 6012 39302 6040 40938
rect 6104 40730 6132 42520
rect 6460 42502 6512 42508
rect 6368 42220 6420 42226
rect 6368 42162 6420 42168
rect 6380 41682 6408 42162
rect 6472 41818 6500 42502
rect 6564 41818 6592 44202
rect 6748 43450 6776 44540
rect 7024 43840 7052 44540
rect 7024 43812 7236 43840
rect 6814 43548 7122 43557
rect 6814 43546 6820 43548
rect 6876 43546 6900 43548
rect 6956 43546 6980 43548
rect 7036 43546 7060 43548
rect 7116 43546 7122 43548
rect 6876 43494 6878 43546
rect 7058 43494 7060 43546
rect 6814 43492 6820 43494
rect 6876 43492 6900 43494
rect 6956 43492 6980 43494
rect 7036 43492 7060 43494
rect 7116 43492 7122 43494
rect 6814 43483 7122 43492
rect 7208 43450 7236 43812
rect 6736 43444 6788 43450
rect 6736 43386 6788 43392
rect 7196 43444 7248 43450
rect 7196 43386 7248 43392
rect 6644 43308 6696 43314
rect 6644 43250 6696 43256
rect 6656 42090 6684 43250
rect 6734 42800 6790 42809
rect 6734 42735 6790 42744
rect 6644 42084 6696 42090
rect 6644 42026 6696 42032
rect 6460 41812 6512 41818
rect 6460 41754 6512 41760
rect 6552 41812 6604 41818
rect 6552 41754 6604 41760
rect 6748 41750 6776 42735
rect 7012 42628 7064 42634
rect 7064 42588 7236 42616
rect 7012 42570 7064 42576
rect 7208 42537 7236 42588
rect 7194 42528 7250 42537
rect 6814 42460 7122 42469
rect 7194 42463 7250 42472
rect 6814 42458 6820 42460
rect 6876 42458 6900 42460
rect 6956 42458 6980 42460
rect 7036 42458 7060 42460
rect 7116 42458 7122 42460
rect 6876 42406 6878 42458
rect 7058 42406 7060 42458
rect 6814 42404 6820 42406
rect 6876 42404 6900 42406
rect 6956 42404 6980 42406
rect 7036 42404 7060 42406
rect 7116 42404 7122 42406
rect 6814 42395 7122 42404
rect 7300 42362 7328 44540
rect 7576 43246 7604 44540
rect 7748 44328 7800 44334
rect 7748 44270 7800 44276
rect 7760 43466 7788 44270
rect 7852 43602 7880 44540
rect 7852 43574 7972 43602
rect 7760 43438 7880 43466
rect 7748 43376 7800 43382
rect 7748 43318 7800 43324
rect 7564 43240 7616 43246
rect 7564 43182 7616 43188
rect 7564 42628 7616 42634
rect 7564 42570 7616 42576
rect 7288 42356 7340 42362
rect 7288 42298 7340 42304
rect 7472 42220 7524 42226
rect 7472 42162 7524 42168
rect 6828 42152 6880 42158
rect 6828 42094 6880 42100
rect 6736 41744 6788 41750
rect 6736 41686 6788 41692
rect 6840 41682 6868 42094
rect 6920 42016 6972 42022
rect 6920 41958 6972 41964
rect 6368 41676 6420 41682
rect 6368 41618 6420 41624
rect 6828 41676 6880 41682
rect 6828 41618 6880 41624
rect 6644 41540 6696 41546
rect 6644 41482 6696 41488
rect 6368 41472 6420 41478
rect 6656 41449 6684 41482
rect 6932 41460 6960 41958
rect 7104 41608 7156 41614
rect 7156 41568 7236 41596
rect 7104 41550 7156 41556
rect 6368 41414 6420 41420
rect 6642 41440 6698 41449
rect 6092 40724 6144 40730
rect 6092 40666 6144 40672
rect 6182 40624 6238 40633
rect 6182 40559 6238 40568
rect 6276 40588 6328 40594
rect 6196 40526 6224 40559
rect 6276 40530 6328 40536
rect 6184 40520 6236 40526
rect 6184 40462 6236 40468
rect 6184 39908 6236 39914
rect 6184 39850 6236 39856
rect 6196 39438 6224 39850
rect 6184 39432 6236 39438
rect 6184 39374 6236 39380
rect 6000 39296 6052 39302
rect 6000 39238 6052 39244
rect 6092 39296 6144 39302
rect 6092 39238 6144 39244
rect 6012 37312 6040 39238
rect 6104 38418 6132 39238
rect 6288 38593 6316 40530
rect 6380 38894 6408 41414
rect 6642 41375 6698 41384
rect 6748 41432 6960 41460
rect 6552 40928 6604 40934
rect 6552 40870 6604 40876
rect 6564 40186 6592 40870
rect 6552 40180 6604 40186
rect 6552 40122 6604 40128
rect 6460 40112 6512 40118
rect 6460 40054 6512 40060
rect 6472 39302 6500 40054
rect 6748 40050 6776 41432
rect 6814 41372 7122 41381
rect 6814 41370 6820 41372
rect 6876 41370 6900 41372
rect 6956 41370 6980 41372
rect 7036 41370 7060 41372
rect 7116 41370 7122 41372
rect 6876 41318 6878 41370
rect 7058 41318 7060 41370
rect 6814 41316 6820 41318
rect 6876 41316 6900 41318
rect 6956 41316 6980 41318
rect 7036 41316 7060 41318
rect 7116 41316 7122 41318
rect 6814 41307 7122 41316
rect 7208 40730 7236 41568
rect 7484 40905 7512 42162
rect 7576 42158 7604 42570
rect 7760 42362 7788 43318
rect 7852 42786 7880 43438
rect 7944 42906 7972 43574
rect 7932 42900 7984 42906
rect 7932 42842 7984 42848
rect 8024 42832 8076 42838
rect 7852 42758 7972 42786
rect 8024 42774 8076 42780
rect 7748 42356 7800 42362
rect 7748 42298 7800 42304
rect 7564 42152 7616 42158
rect 7564 42094 7616 42100
rect 7944 42022 7972 42758
rect 7656 42016 7708 42022
rect 7656 41958 7708 41964
rect 7840 42016 7892 42022
rect 7840 41958 7892 41964
rect 7932 42016 7984 42022
rect 7932 41958 7984 41964
rect 7562 41712 7618 41721
rect 7562 41647 7618 41656
rect 7576 41206 7604 41647
rect 7668 41614 7696 41958
rect 7656 41608 7708 41614
rect 7656 41550 7708 41556
rect 7852 41414 7880 41958
rect 7760 41386 7880 41414
rect 7656 41268 7708 41274
rect 7656 41210 7708 41216
rect 7564 41200 7616 41206
rect 7564 41142 7616 41148
rect 7470 40896 7526 40905
rect 7470 40831 7526 40840
rect 7196 40724 7248 40730
rect 7196 40666 7248 40672
rect 7484 40662 7512 40831
rect 7472 40656 7524 40662
rect 7472 40598 7524 40604
rect 7196 40520 7248 40526
rect 7196 40462 7248 40468
rect 6814 40284 7122 40293
rect 6814 40282 6820 40284
rect 6876 40282 6900 40284
rect 6956 40282 6980 40284
rect 7036 40282 7060 40284
rect 7116 40282 7122 40284
rect 6876 40230 6878 40282
rect 7058 40230 7060 40282
rect 6814 40228 6820 40230
rect 6876 40228 6900 40230
rect 6956 40228 6980 40230
rect 7036 40228 7060 40230
rect 7116 40228 7122 40230
rect 6814 40219 7122 40228
rect 6736 40044 6788 40050
rect 6736 39986 6788 39992
rect 6460 39296 6512 39302
rect 6460 39238 6512 39244
rect 6368 38888 6420 38894
rect 6368 38830 6420 38836
rect 6552 38888 6604 38894
rect 6552 38830 6604 38836
rect 6274 38584 6330 38593
rect 6274 38519 6330 38528
rect 6092 38412 6144 38418
rect 6092 38354 6144 38360
rect 6184 37460 6236 37466
rect 6184 37402 6236 37408
rect 6012 37284 6132 37312
rect 6104 37194 6132 37284
rect 6196 37233 6224 37402
rect 6274 37360 6330 37369
rect 6274 37295 6330 37304
rect 6182 37224 6238 37233
rect 5908 37188 5960 37194
rect 5908 37130 5960 37136
rect 6000 37188 6052 37194
rect 6000 37130 6052 37136
rect 6092 37188 6144 37194
rect 6182 37159 6238 37168
rect 6092 37130 6144 37136
rect 5908 35488 5960 35494
rect 5908 35430 5960 35436
rect 5920 35086 5948 35430
rect 6012 35086 6040 37130
rect 5908 35080 5960 35086
rect 5908 35022 5960 35028
rect 6000 35080 6052 35086
rect 6000 35022 6052 35028
rect 6104 34785 6132 37130
rect 6288 36922 6316 37295
rect 6276 36916 6328 36922
rect 6276 36858 6328 36864
rect 6184 35828 6236 35834
rect 6184 35770 6236 35776
rect 6090 34776 6146 34785
rect 6090 34711 6146 34720
rect 6196 34610 6224 35770
rect 6274 35048 6330 35057
rect 6274 34983 6330 34992
rect 6288 34950 6316 34983
rect 6276 34944 6328 34950
rect 6276 34886 6328 34892
rect 5908 34604 5960 34610
rect 5908 34546 5960 34552
rect 6184 34604 6236 34610
rect 6184 34546 6236 34552
rect 5920 33017 5948 34546
rect 6092 34536 6144 34542
rect 6092 34478 6144 34484
rect 5998 33688 6054 33697
rect 5998 33623 6054 33632
rect 6012 33590 6040 33623
rect 6000 33584 6052 33590
rect 6000 33526 6052 33532
rect 5906 33008 5962 33017
rect 5906 32943 5962 32952
rect 5920 32314 5948 32943
rect 6000 32768 6052 32774
rect 6000 32710 6052 32716
rect 6012 32502 6040 32710
rect 6000 32496 6052 32502
rect 6000 32438 6052 32444
rect 5920 32286 6040 32314
rect 5908 32224 5960 32230
rect 5908 32166 5960 32172
rect 5736 32014 5856 32042
rect 5736 31822 5764 32014
rect 5920 31890 5948 32166
rect 5908 31884 5960 31890
rect 5908 31826 5960 31832
rect 5724 31816 5776 31822
rect 6012 31793 6040 32286
rect 5724 31758 5776 31764
rect 5998 31784 6054 31793
rect 5908 31748 5960 31754
rect 5998 31719 6054 31728
rect 5908 31690 5960 31696
rect 5816 31680 5868 31686
rect 5816 31622 5868 31628
rect 5722 31240 5778 31249
rect 5722 31175 5778 31184
rect 5736 30666 5764 31175
rect 5724 30660 5776 30666
rect 5724 30602 5776 30608
rect 5644 29702 5764 29730
rect 5632 29572 5684 29578
rect 5632 29514 5684 29520
rect 5644 28082 5672 29514
rect 5632 28076 5684 28082
rect 5632 28018 5684 28024
rect 5644 27062 5672 28018
rect 5632 27056 5684 27062
rect 5632 26998 5684 27004
rect 5736 26382 5764 29702
rect 5828 28234 5856 31622
rect 5920 31521 5948 31690
rect 5906 31512 5962 31521
rect 5906 31447 5962 31456
rect 6000 31408 6052 31414
rect 6000 31350 6052 31356
rect 5908 31136 5960 31142
rect 5908 31078 5960 31084
rect 5920 30938 5948 31078
rect 6012 30938 6040 31350
rect 5908 30932 5960 30938
rect 5908 30874 5960 30880
rect 6000 30932 6052 30938
rect 6000 30874 6052 30880
rect 5908 30592 5960 30598
rect 5908 30534 5960 30540
rect 5920 30394 5948 30534
rect 5908 30388 5960 30394
rect 5908 30330 5960 30336
rect 5908 30252 5960 30258
rect 5908 30194 5960 30200
rect 5920 30161 5948 30194
rect 5906 30152 5962 30161
rect 5906 30087 5962 30096
rect 5998 29608 6054 29617
rect 6104 29578 6132 34478
rect 6276 33992 6328 33998
rect 6276 33934 6328 33940
rect 6184 33856 6236 33862
rect 6184 33798 6236 33804
rect 6196 33590 6224 33798
rect 6184 33584 6236 33590
rect 6184 33526 6236 33532
rect 6196 33114 6224 33526
rect 6184 33108 6236 33114
rect 6184 33050 6236 33056
rect 6288 32842 6316 33934
rect 6380 33658 6408 38830
rect 6460 38344 6512 38350
rect 6460 38286 6512 38292
rect 6472 33998 6500 38286
rect 6564 37398 6592 38830
rect 6552 37392 6604 37398
rect 6552 37334 6604 37340
rect 6460 33992 6512 33998
rect 6460 33934 6512 33940
rect 6368 33652 6420 33658
rect 6368 33594 6420 33600
rect 6184 32836 6236 32842
rect 6184 32778 6236 32784
rect 6276 32836 6328 32842
rect 6276 32778 6328 32784
rect 6196 32552 6224 32778
rect 6196 32524 6408 32552
rect 6184 32428 6236 32434
rect 6184 32370 6236 32376
rect 6196 30734 6224 32370
rect 6276 32292 6328 32298
rect 6276 32234 6328 32240
rect 6184 30728 6236 30734
rect 6184 30670 6236 30676
rect 6288 29578 6316 32234
rect 6380 32230 6408 32524
rect 6368 32224 6420 32230
rect 6368 32166 6420 32172
rect 6380 30598 6408 32166
rect 6472 31754 6500 33934
rect 6564 33538 6592 37334
rect 6642 37088 6698 37097
rect 6642 37023 6698 37032
rect 6656 36174 6684 37023
rect 6644 36168 6696 36174
rect 6644 36110 6696 36116
rect 6748 35834 6776 39986
rect 6814 39196 7122 39205
rect 6814 39194 6820 39196
rect 6876 39194 6900 39196
rect 6956 39194 6980 39196
rect 7036 39194 7060 39196
rect 7116 39194 7122 39196
rect 6876 39142 6878 39194
rect 7058 39142 7060 39194
rect 6814 39140 6820 39142
rect 6876 39140 6900 39142
rect 6956 39140 6980 39142
rect 7036 39140 7060 39142
rect 7116 39140 7122 39142
rect 6814 39131 7122 39140
rect 7208 38214 7236 40462
rect 7380 39840 7432 39846
rect 7380 39782 7432 39788
rect 7288 39364 7340 39370
rect 7288 39306 7340 39312
rect 7196 38208 7248 38214
rect 7196 38150 7248 38156
rect 6814 38108 7122 38117
rect 6814 38106 6820 38108
rect 6876 38106 6900 38108
rect 6956 38106 6980 38108
rect 7036 38106 7060 38108
rect 7116 38106 7122 38108
rect 6876 38054 6878 38106
rect 7058 38054 7060 38106
rect 6814 38052 6820 38054
rect 6876 38052 6900 38054
rect 6956 38052 6980 38054
rect 7036 38052 7060 38054
rect 7116 38052 7122 38054
rect 6814 38043 7122 38052
rect 6920 37256 6972 37262
rect 7300 37244 7328 39306
rect 7392 38894 7420 39782
rect 7472 39296 7524 39302
rect 7472 39238 7524 39244
rect 7380 38888 7432 38894
rect 7380 38830 7432 38836
rect 7392 38554 7420 38830
rect 7484 38554 7512 39238
rect 7380 38548 7432 38554
rect 7380 38490 7432 38496
rect 7472 38548 7524 38554
rect 7472 38490 7524 38496
rect 7472 38344 7524 38350
rect 6972 37216 7328 37244
rect 7392 38292 7472 38298
rect 7392 38286 7524 38292
rect 7392 38270 7512 38286
rect 6920 37198 6972 37204
rect 6814 37020 7122 37029
rect 6814 37018 6820 37020
rect 6876 37018 6900 37020
rect 6956 37018 6980 37020
rect 7036 37018 7060 37020
rect 7116 37018 7122 37020
rect 6876 36966 6878 37018
rect 7058 36966 7060 37018
rect 6814 36964 6820 36966
rect 6876 36964 6900 36966
rect 6956 36964 6980 36966
rect 7036 36964 7060 36966
rect 7116 36964 7122 36966
rect 6814 36955 7122 36964
rect 7104 36848 7156 36854
rect 7104 36790 7156 36796
rect 7116 36258 7144 36790
rect 7208 36378 7236 37216
rect 7392 36786 7420 38270
rect 7472 37188 7524 37194
rect 7472 37130 7524 37136
rect 7484 36854 7512 37130
rect 7576 36854 7604 41142
rect 7668 40066 7696 41210
rect 7760 41070 7788 41386
rect 7748 41064 7800 41070
rect 7748 41006 7800 41012
rect 7840 40656 7892 40662
rect 7840 40598 7892 40604
rect 7668 40038 7788 40066
rect 7656 39976 7708 39982
rect 7656 39918 7708 39924
rect 7668 38962 7696 39918
rect 7760 38962 7788 40038
rect 7656 38956 7708 38962
rect 7656 38898 7708 38904
rect 7748 38956 7800 38962
rect 7748 38898 7800 38904
rect 7668 37806 7696 38898
rect 7656 37800 7708 37806
rect 7656 37742 7708 37748
rect 7656 37664 7708 37670
rect 7656 37606 7708 37612
rect 7668 37398 7696 37606
rect 7656 37392 7708 37398
rect 7656 37334 7708 37340
rect 7760 37194 7788 38898
rect 7748 37188 7800 37194
rect 7748 37130 7800 37136
rect 7472 36848 7524 36854
rect 7472 36790 7524 36796
rect 7564 36848 7616 36854
rect 7564 36790 7616 36796
rect 7380 36780 7432 36786
rect 7380 36722 7432 36728
rect 7288 36576 7340 36582
rect 7288 36518 7340 36524
rect 7196 36372 7248 36378
rect 7196 36314 7248 36320
rect 7116 36230 7236 36258
rect 6814 35932 7122 35941
rect 6814 35930 6820 35932
rect 6876 35930 6900 35932
rect 6956 35930 6980 35932
rect 7036 35930 7060 35932
rect 7116 35930 7122 35932
rect 6876 35878 6878 35930
rect 7058 35878 7060 35930
rect 6814 35876 6820 35878
rect 6876 35876 6900 35878
rect 6956 35876 6980 35878
rect 7036 35876 7060 35878
rect 7116 35876 7122 35878
rect 6814 35867 7122 35876
rect 6736 35828 6788 35834
rect 6736 35770 6788 35776
rect 6644 35080 6696 35086
rect 6644 35022 6696 35028
rect 6656 34542 6684 35022
rect 6736 34944 6788 34950
rect 6736 34886 6788 34892
rect 6644 34536 6696 34542
rect 6644 34478 6696 34484
rect 6748 34066 6776 34886
rect 6814 34844 7122 34853
rect 6814 34842 6820 34844
rect 6876 34842 6900 34844
rect 6956 34842 6980 34844
rect 7036 34842 7060 34844
rect 7116 34842 7122 34844
rect 6876 34790 6878 34842
rect 7058 34790 7060 34842
rect 6814 34788 6820 34790
rect 6876 34788 6900 34790
rect 6956 34788 6980 34790
rect 7036 34788 7060 34790
rect 7116 34788 7122 34790
rect 6814 34779 7122 34788
rect 6736 34060 6788 34066
rect 6736 34002 6788 34008
rect 6644 33992 6696 33998
rect 6644 33934 6696 33940
rect 6656 33658 6684 33934
rect 6814 33756 7122 33765
rect 6814 33754 6820 33756
rect 6876 33754 6900 33756
rect 6956 33754 6980 33756
rect 7036 33754 7060 33756
rect 7116 33754 7122 33756
rect 6876 33702 6878 33754
rect 7058 33702 7060 33754
rect 6814 33700 6820 33702
rect 6876 33700 6900 33702
rect 6956 33700 6980 33702
rect 7036 33700 7060 33702
rect 7116 33700 7122 33702
rect 6814 33691 7122 33700
rect 6644 33652 6696 33658
rect 6644 33594 6696 33600
rect 7012 33652 7064 33658
rect 7012 33594 7064 33600
rect 6564 33510 6684 33538
rect 6656 31906 6684 33510
rect 6736 33108 6788 33114
rect 6736 33050 6788 33056
rect 6748 32026 6776 33050
rect 7024 33046 7052 33594
rect 7208 33153 7236 36230
rect 7300 35698 7328 36518
rect 7380 36236 7432 36242
rect 7380 36178 7432 36184
rect 7288 35692 7340 35698
rect 7288 35634 7340 35640
rect 7392 35630 7420 36178
rect 7748 36168 7800 36174
rect 7748 36110 7800 36116
rect 7656 35692 7708 35698
rect 7656 35634 7708 35640
rect 7380 35624 7432 35630
rect 7380 35566 7432 35572
rect 7288 33924 7340 33930
rect 7288 33866 7340 33872
rect 7300 33386 7328 33866
rect 7392 33436 7420 35566
rect 7472 35012 7524 35018
rect 7524 34972 7604 35000
rect 7472 34954 7524 34960
rect 7472 34740 7524 34746
rect 7472 34682 7524 34688
rect 7484 33658 7512 34682
rect 7472 33652 7524 33658
rect 7472 33594 7524 33600
rect 7472 33448 7524 33454
rect 7392 33408 7472 33436
rect 7472 33390 7524 33396
rect 7288 33380 7340 33386
rect 7288 33322 7340 33328
rect 7194 33144 7250 33153
rect 7194 33079 7250 33088
rect 7012 33040 7064 33046
rect 7012 32982 7064 32988
rect 7024 32756 7052 32982
rect 7104 32972 7156 32978
rect 7484 32960 7512 33390
rect 7156 32932 7512 32960
rect 7104 32914 7156 32920
rect 7024 32728 7236 32756
rect 6814 32668 7122 32677
rect 6814 32666 6820 32668
rect 6876 32666 6900 32668
rect 6956 32666 6980 32668
rect 7036 32666 7060 32668
rect 7116 32666 7122 32668
rect 6876 32614 6878 32666
rect 7058 32614 7060 32666
rect 6814 32612 6820 32614
rect 6876 32612 6900 32614
rect 6956 32612 6980 32614
rect 7036 32612 7060 32614
rect 7116 32612 7122 32614
rect 6814 32603 7122 32612
rect 6920 32428 6972 32434
rect 6920 32370 6972 32376
rect 6736 32020 6788 32026
rect 6736 31962 6788 31968
rect 6656 31878 6776 31906
rect 6460 31748 6512 31754
rect 6460 31690 6512 31696
rect 6368 30592 6420 30598
rect 6368 30534 6420 30540
rect 6368 30048 6420 30054
rect 6368 29990 6420 29996
rect 6380 29850 6408 29990
rect 6368 29844 6420 29850
rect 6368 29786 6420 29792
rect 5998 29543 6054 29552
rect 6092 29572 6144 29578
rect 5828 28206 5948 28234
rect 5816 28144 5868 28150
rect 5816 28086 5868 28092
rect 5828 27674 5856 28086
rect 5816 27668 5868 27674
rect 5816 27610 5868 27616
rect 5724 26376 5776 26382
rect 5816 26376 5868 26382
rect 5724 26318 5776 26324
rect 5814 26344 5816 26353
rect 5868 26344 5870 26353
rect 5632 26308 5684 26314
rect 5632 26250 5684 26256
rect 5644 24993 5672 26250
rect 5630 24984 5686 24993
rect 5630 24919 5686 24928
rect 5632 23316 5684 23322
rect 5632 23258 5684 23264
rect 5644 22506 5672 23258
rect 5736 23202 5764 26318
rect 5814 26279 5870 26288
rect 5920 25786 5948 28206
rect 6012 26330 6040 29543
rect 6092 29514 6144 29520
rect 6276 29572 6328 29578
rect 6276 29514 6328 29520
rect 6104 29170 6132 29514
rect 6368 29504 6420 29510
rect 6368 29446 6420 29452
rect 6092 29164 6144 29170
rect 6092 29106 6144 29112
rect 6184 29164 6236 29170
rect 6184 29106 6236 29112
rect 6196 29073 6224 29106
rect 6276 29096 6328 29102
rect 6182 29064 6238 29073
rect 6276 29038 6328 29044
rect 6182 28999 6238 29008
rect 6092 28484 6144 28490
rect 6092 28426 6144 28432
rect 6104 28218 6132 28426
rect 6184 28416 6236 28422
rect 6184 28358 6236 28364
rect 6092 28212 6144 28218
rect 6092 28154 6144 28160
rect 6196 28014 6224 28358
rect 6184 28008 6236 28014
rect 6184 27950 6236 27956
rect 6092 27872 6144 27878
rect 6090 27840 6092 27849
rect 6144 27840 6146 27849
rect 6090 27775 6146 27784
rect 6012 26302 6132 26330
rect 6000 26240 6052 26246
rect 6000 26182 6052 26188
rect 5828 25758 5948 25786
rect 5828 23322 5856 25758
rect 5908 25696 5960 25702
rect 5908 25638 5960 25644
rect 5920 24750 5948 25638
rect 5908 24744 5960 24750
rect 5908 24686 5960 24692
rect 5816 23316 5868 23322
rect 5816 23258 5868 23264
rect 5736 23174 5948 23202
rect 5816 22772 5868 22778
rect 5816 22714 5868 22720
rect 5724 22636 5776 22642
rect 5724 22578 5776 22584
rect 5632 22500 5684 22506
rect 5632 22442 5684 22448
rect 5460 21916 5580 21944
rect 5460 21593 5488 21916
rect 5644 21842 5672 22442
rect 5552 21814 5672 21842
rect 5552 21622 5580 21814
rect 5736 21672 5764 22578
rect 5644 21644 5764 21672
rect 5540 21616 5592 21622
rect 5446 21584 5502 21593
rect 5540 21558 5592 21564
rect 5446 21519 5502 21528
rect 5448 21412 5500 21418
rect 5448 21354 5500 21360
rect 5460 21146 5488 21354
rect 5552 21146 5580 21558
rect 5448 21140 5500 21146
rect 5448 21082 5500 21088
rect 5540 21140 5592 21146
rect 5540 21082 5592 21088
rect 5448 21004 5500 21010
rect 5448 20946 5500 20952
rect 5460 19938 5488 20946
rect 5540 20460 5592 20466
rect 5540 20402 5592 20408
rect 5552 20244 5580 20402
rect 5644 20346 5672 21644
rect 5828 21536 5856 22714
rect 5920 22574 5948 23174
rect 6012 22642 6040 26182
rect 6104 25770 6132 26302
rect 6288 26246 6316 29038
rect 6380 28082 6408 29446
rect 6368 28076 6420 28082
rect 6368 28018 6420 28024
rect 6380 27334 6408 28018
rect 6368 27328 6420 27334
rect 6368 27270 6420 27276
rect 6368 26784 6420 26790
rect 6368 26726 6420 26732
rect 6276 26240 6328 26246
rect 6276 26182 6328 26188
rect 6276 26036 6328 26042
rect 6276 25978 6328 25984
rect 6092 25764 6144 25770
rect 6092 25706 6144 25712
rect 6184 24948 6236 24954
rect 6184 24890 6236 24896
rect 6090 24848 6146 24857
rect 6090 24783 6146 24792
rect 6104 24410 6132 24783
rect 6092 24404 6144 24410
rect 6092 24346 6144 24352
rect 6196 22642 6224 24890
rect 6288 24682 6316 25978
rect 6380 25294 6408 26726
rect 6368 25288 6420 25294
rect 6368 25230 6420 25236
rect 6276 24676 6328 24682
rect 6276 24618 6328 24624
rect 6276 24064 6328 24070
rect 6276 24006 6328 24012
rect 6288 23662 6316 24006
rect 6276 23656 6328 23662
rect 6276 23598 6328 23604
rect 6276 22976 6328 22982
rect 6276 22918 6328 22924
rect 6288 22681 6316 22918
rect 6380 22710 6408 25230
rect 6472 24313 6500 31690
rect 6644 31680 6696 31686
rect 6644 31622 6696 31628
rect 6656 30546 6684 31622
rect 6564 30518 6684 30546
rect 6564 29578 6592 30518
rect 6644 30388 6696 30394
rect 6644 30330 6696 30336
rect 6552 29572 6604 29578
rect 6552 29514 6604 29520
rect 6564 29084 6592 29514
rect 6656 29481 6684 30330
rect 6642 29472 6698 29481
rect 6642 29407 6698 29416
rect 6564 29056 6684 29084
rect 6550 28248 6606 28257
rect 6550 28183 6606 28192
rect 6564 28082 6592 28183
rect 6552 28076 6604 28082
rect 6552 28018 6604 28024
rect 6656 28014 6684 29056
rect 6644 28008 6696 28014
rect 6644 27950 6696 27956
rect 6552 27668 6604 27674
rect 6552 27610 6604 27616
rect 6564 27130 6592 27610
rect 6644 27328 6696 27334
rect 6644 27270 6696 27276
rect 6656 27130 6684 27270
rect 6552 27124 6604 27130
rect 6552 27066 6604 27072
rect 6644 27124 6696 27130
rect 6644 27066 6696 27072
rect 6644 26240 6696 26246
rect 6644 26182 6696 26188
rect 6550 25664 6606 25673
rect 6550 25599 6606 25608
rect 6564 25430 6592 25599
rect 6552 25424 6604 25430
rect 6552 25366 6604 25372
rect 6564 25129 6592 25366
rect 6550 25120 6606 25129
rect 6550 25055 6606 25064
rect 6552 24880 6604 24886
rect 6552 24822 6604 24828
rect 6458 24304 6514 24313
rect 6458 24239 6514 24248
rect 6460 23180 6512 23186
rect 6460 23122 6512 23128
rect 6368 22704 6420 22710
rect 6274 22672 6330 22681
rect 6000 22636 6052 22642
rect 6000 22578 6052 22584
rect 6184 22636 6236 22642
rect 6368 22646 6420 22652
rect 6274 22607 6330 22616
rect 6184 22578 6236 22584
rect 5908 22568 5960 22574
rect 5908 22510 5960 22516
rect 6276 22160 6328 22166
rect 6274 22128 6276 22137
rect 6328 22128 6330 22137
rect 6274 22063 6330 22072
rect 6184 22024 6236 22030
rect 6236 21984 6316 22012
rect 6184 21966 6236 21972
rect 6000 21888 6052 21894
rect 6000 21830 6052 21836
rect 5736 21508 5856 21536
rect 5906 21584 5962 21593
rect 5906 21519 5962 21528
rect 5736 21078 5764 21508
rect 5920 21298 5948 21519
rect 6012 21486 6040 21830
rect 6288 21593 6316 21984
rect 6274 21584 6330 21593
rect 6184 21548 6236 21554
rect 6274 21519 6330 21528
rect 6184 21490 6236 21496
rect 6000 21480 6052 21486
rect 6000 21422 6052 21428
rect 5920 21270 6040 21298
rect 5816 21140 5868 21146
rect 5816 21082 5868 21088
rect 5724 21072 5776 21078
rect 5724 21014 5776 21020
rect 5828 20602 5856 21082
rect 5816 20596 5868 20602
rect 5816 20538 5868 20544
rect 5644 20318 5856 20346
rect 5552 20216 5672 20244
rect 5538 19952 5594 19961
rect 5356 19916 5408 19922
rect 5356 19858 5408 19864
rect 5460 19910 5538 19938
rect 5356 19780 5408 19786
rect 5356 19722 5408 19728
rect 5264 18828 5316 18834
rect 5264 18770 5316 18776
rect 5276 18154 5304 18770
rect 5368 18737 5396 19722
rect 5460 19281 5488 19910
rect 5538 19887 5594 19896
rect 5644 19378 5672 20216
rect 5632 19372 5684 19378
rect 5632 19314 5684 19320
rect 5446 19272 5502 19281
rect 5446 19207 5502 19216
rect 5632 19236 5684 19242
rect 5632 19178 5684 19184
rect 5448 18760 5500 18766
rect 5354 18728 5410 18737
rect 5448 18702 5500 18708
rect 5354 18663 5410 18672
rect 5356 18624 5408 18630
rect 5356 18566 5408 18572
rect 5368 18358 5396 18566
rect 5460 18426 5488 18702
rect 5540 18624 5592 18630
rect 5540 18566 5592 18572
rect 5448 18420 5500 18426
rect 5448 18362 5500 18368
rect 5356 18352 5408 18358
rect 5356 18294 5408 18300
rect 5264 18148 5316 18154
rect 5264 18090 5316 18096
rect 5448 18080 5500 18086
rect 5448 18022 5500 18028
rect 5460 17882 5488 18022
rect 5448 17876 5500 17882
rect 5448 17818 5500 17824
rect 5552 17678 5580 18566
rect 5644 18086 5672 19178
rect 5724 18284 5776 18290
rect 5724 18226 5776 18232
rect 5632 18080 5684 18086
rect 5632 18022 5684 18028
rect 5630 17912 5686 17921
rect 5630 17847 5686 17856
rect 5540 17672 5592 17678
rect 5540 17614 5592 17620
rect 5172 17332 5224 17338
rect 5172 17274 5224 17280
rect 5170 17096 5226 17105
rect 5170 17031 5226 17040
rect 5184 16658 5212 17031
rect 5356 16992 5408 16998
rect 5356 16934 5408 16940
rect 5368 16658 5396 16934
rect 5540 16788 5592 16794
rect 5540 16730 5592 16736
rect 5172 16652 5224 16658
rect 5172 16594 5224 16600
rect 5356 16652 5408 16658
rect 5356 16594 5408 16600
rect 5264 16108 5316 16114
rect 5264 16050 5316 16056
rect 5170 14784 5226 14793
rect 5170 14719 5226 14728
rect 4908 14572 5120 14600
rect 4908 14278 4936 14572
rect 4988 14476 5040 14482
rect 4988 14418 5040 14424
rect 4896 14272 4948 14278
rect 4896 14214 4948 14220
rect 5000 13530 5028 14418
rect 5080 14272 5132 14278
rect 5080 14214 5132 14220
rect 4988 13524 5040 13530
rect 4988 13466 5040 13472
rect 4896 13388 4948 13394
rect 4896 13330 4948 13336
rect 4712 12232 4764 12238
rect 4712 12174 4764 12180
rect 4632 12022 4752 12050
rect 4528 11688 4580 11694
rect 4528 11630 4580 11636
rect 4540 10577 4568 11630
rect 4620 11552 4672 11558
rect 4620 11494 4672 11500
rect 4526 10568 4582 10577
rect 4526 10503 4582 10512
rect 4528 9580 4580 9586
rect 4528 9522 4580 9528
rect 4436 8968 4488 8974
rect 4436 8910 4488 8916
rect 4448 7970 4476 8910
rect 4540 8838 4568 9522
rect 4528 8832 4580 8838
rect 4528 8774 4580 8780
rect 4632 8430 4660 11494
rect 4620 8424 4672 8430
rect 4620 8366 4672 8372
rect 4528 8356 4580 8362
rect 4528 8298 4580 8304
rect 4540 8090 4568 8298
rect 4528 8084 4580 8090
rect 4528 8026 4580 8032
rect 4448 7942 4568 7970
rect 4344 7812 4396 7818
rect 4344 7754 4396 7760
rect 4436 7812 4488 7818
rect 4436 7754 4488 7760
rect 4252 7404 4304 7410
rect 4252 7346 4304 7352
rect 4080 7274 4200 7290
rect 4068 7268 4200 7274
rect 4120 7262 4200 7268
rect 4068 7210 4120 7216
rect 3882 7100 4190 7109
rect 3882 7098 3888 7100
rect 3944 7098 3968 7100
rect 4024 7098 4048 7100
rect 4104 7098 4128 7100
rect 4184 7098 4190 7100
rect 3944 7046 3946 7098
rect 4126 7046 4128 7098
rect 3882 7044 3888 7046
rect 3944 7044 3968 7046
rect 4024 7044 4048 7046
rect 4104 7044 4128 7046
rect 4184 7044 4190 7046
rect 3882 7035 4190 7044
rect 4264 6798 4292 7346
rect 4344 7200 4396 7206
rect 4344 7142 4396 7148
rect 4252 6792 4304 6798
rect 4252 6734 4304 6740
rect 3792 6316 3844 6322
rect 3792 6258 3844 6264
rect 3804 5778 3832 6258
rect 4264 6100 4292 6734
rect 4356 6254 4384 7142
rect 4344 6248 4396 6254
rect 4344 6190 4396 6196
rect 4344 6112 4396 6118
rect 4264 6072 4344 6100
rect 3882 6012 4190 6021
rect 3882 6010 3888 6012
rect 3944 6010 3968 6012
rect 4024 6010 4048 6012
rect 4104 6010 4128 6012
rect 4184 6010 4190 6012
rect 3944 5958 3946 6010
rect 4126 5958 4128 6010
rect 3882 5956 3888 5958
rect 3944 5956 3968 5958
rect 4024 5956 4048 5958
rect 4104 5956 4128 5958
rect 4184 5956 4190 5958
rect 3882 5947 4190 5956
rect 3792 5772 3844 5778
rect 3792 5714 3844 5720
rect 4068 5704 4120 5710
rect 4066 5672 4068 5681
rect 4120 5672 4122 5681
rect 4066 5607 4122 5616
rect 3516 5364 3568 5370
rect 3516 5306 3568 5312
rect 3698 5264 3754 5273
rect 3698 5199 3754 5208
rect 4160 5228 4212 5234
rect 3516 5024 3568 5030
rect 3516 4966 3568 4972
rect 3528 4185 3556 4966
rect 3712 4826 3740 5199
rect 4264 5216 4292 6072
rect 4344 6054 4396 6060
rect 4448 5914 4476 7754
rect 4540 7478 4568 7942
rect 4528 7472 4580 7478
rect 4528 7414 4580 7420
rect 4724 7290 4752 12022
rect 4804 11756 4856 11762
rect 4804 11698 4856 11704
rect 4816 10810 4844 11698
rect 4908 10849 4936 13330
rect 4894 10840 4950 10849
rect 4804 10804 4856 10810
rect 4894 10775 4950 10784
rect 4804 10746 4856 10752
rect 4908 10674 4936 10775
rect 4896 10668 4948 10674
rect 4896 10610 4948 10616
rect 4896 9512 4948 9518
rect 4802 9480 4858 9489
rect 4896 9454 4948 9460
rect 4802 9415 4804 9424
rect 4856 9415 4858 9424
rect 4804 9386 4856 9392
rect 4908 9110 4936 9454
rect 4896 9104 4948 9110
rect 4896 9046 4948 9052
rect 5092 8922 5120 14214
rect 5184 13938 5212 14719
rect 5276 14482 5304 16050
rect 5552 15706 5580 16730
rect 5540 15700 5592 15706
rect 5540 15642 5592 15648
rect 5644 15586 5672 17847
rect 5552 15558 5672 15586
rect 5552 15366 5580 15558
rect 5540 15360 5592 15366
rect 5540 15302 5592 15308
rect 5354 15192 5410 15201
rect 5354 15127 5410 15136
rect 5264 14476 5316 14482
rect 5264 14418 5316 14424
rect 5172 13932 5224 13938
rect 5172 13874 5224 13880
rect 5184 13394 5212 13874
rect 5368 13841 5396 15127
rect 5540 14816 5592 14822
rect 5540 14758 5592 14764
rect 5552 14482 5580 14758
rect 5540 14476 5592 14482
rect 5540 14418 5592 14424
rect 5448 14408 5500 14414
rect 5500 14356 5580 14362
rect 5448 14350 5580 14356
rect 5460 14334 5580 14350
rect 5552 13938 5580 14334
rect 5540 13932 5592 13938
rect 5540 13874 5592 13880
rect 5354 13832 5410 13841
rect 5354 13767 5410 13776
rect 5172 13388 5224 13394
rect 5172 13330 5224 13336
rect 5172 13252 5224 13258
rect 5172 13194 5224 13200
rect 5184 12442 5212 13194
rect 5172 12436 5224 12442
rect 5172 12378 5224 12384
rect 5184 11558 5212 12378
rect 5264 12232 5316 12238
rect 5264 12174 5316 12180
rect 5172 11552 5224 11558
rect 5172 11494 5224 11500
rect 5184 11150 5212 11494
rect 5172 11144 5224 11150
rect 5172 11086 5224 11092
rect 5276 10742 5304 12174
rect 5264 10736 5316 10742
rect 5264 10678 5316 10684
rect 5264 9648 5316 9654
rect 5264 9590 5316 9596
rect 4540 7262 4752 7290
rect 4816 8894 5120 8922
rect 4436 5908 4488 5914
rect 4436 5850 4488 5856
rect 4540 5794 4568 7262
rect 4712 7200 4764 7206
rect 4712 7142 4764 7148
rect 4724 6905 4752 7142
rect 4710 6896 4766 6905
rect 4710 6831 4766 6840
rect 4620 6112 4672 6118
rect 4620 6054 4672 6060
rect 4212 5188 4292 5216
rect 4356 5766 4568 5794
rect 4160 5170 4212 5176
rect 3882 4924 4190 4933
rect 3882 4922 3888 4924
rect 3944 4922 3968 4924
rect 4024 4922 4048 4924
rect 4104 4922 4128 4924
rect 4184 4922 4190 4924
rect 3944 4870 3946 4922
rect 4126 4870 4128 4922
rect 3882 4868 3888 4870
rect 3944 4868 3968 4870
rect 4024 4868 4048 4870
rect 4104 4868 4128 4870
rect 4184 4868 4190 4870
rect 3882 4859 4190 4868
rect 3700 4820 3752 4826
rect 3700 4762 3752 4768
rect 4356 4570 4384 5766
rect 4528 5704 4580 5710
rect 4528 5646 4580 5652
rect 4436 4752 4488 4758
rect 4436 4694 4488 4700
rect 4264 4542 4384 4570
rect 4264 4486 4292 4542
rect 3700 4480 3752 4486
rect 3700 4422 3752 4428
rect 4252 4480 4304 4486
rect 4252 4422 4304 4428
rect 3712 4282 3740 4422
rect 3700 4276 3752 4282
rect 3700 4218 3752 4224
rect 4344 4276 4396 4282
rect 4344 4218 4396 4224
rect 3514 4176 3570 4185
rect 3514 4111 3570 4120
rect 3608 4140 3660 4146
rect 3608 4082 3660 4088
rect 3424 3528 3476 3534
rect 3424 3470 3476 3476
rect 3620 3369 3648 4082
rect 3884 4072 3936 4078
rect 3712 4020 3884 4026
rect 3712 4014 3936 4020
rect 3712 3998 3924 4014
rect 3606 3360 3662 3369
rect 3528 3318 3606 3346
rect 3528 2990 3556 3318
rect 3606 3295 3662 3304
rect 3516 2984 3568 2990
rect 3516 2926 3568 2932
rect 3240 2916 3292 2922
rect 3240 2858 3292 2864
rect 3424 2916 3476 2922
rect 3424 2858 3476 2864
rect 3436 2310 3464 2858
rect 3516 2848 3568 2854
rect 3516 2790 3568 2796
rect 3424 2304 3476 2310
rect 3424 2246 3476 2252
rect 3332 1352 3384 1358
rect 3332 1294 3384 1300
rect 3344 814 3372 1294
rect 3424 1216 3476 1222
rect 3424 1158 3476 1164
rect 3436 950 3464 1158
rect 3424 944 3476 950
rect 3424 886 3476 892
rect 3332 808 3384 814
rect 3528 796 3556 2790
rect 3712 2582 3740 3998
rect 4252 3936 4304 3942
rect 4252 3878 4304 3884
rect 3882 3836 4190 3845
rect 3882 3834 3888 3836
rect 3944 3834 3968 3836
rect 4024 3834 4048 3836
rect 4104 3834 4128 3836
rect 4184 3834 4190 3836
rect 3944 3782 3946 3834
rect 4126 3782 4128 3834
rect 3882 3780 3888 3782
rect 3944 3780 3968 3782
rect 4024 3780 4048 3782
rect 4104 3780 4128 3782
rect 4184 3780 4190 3782
rect 3882 3771 4190 3780
rect 3882 3632 3938 3641
rect 3792 3596 3844 3602
rect 3844 3576 3882 3584
rect 3844 3567 3938 3576
rect 3844 3556 3924 3567
rect 3792 3538 3844 3544
rect 3976 3052 4028 3058
rect 3976 2994 4028 3000
rect 3988 2938 4016 2994
rect 4264 2972 4292 3878
rect 4356 3738 4384 4218
rect 4344 3732 4396 3738
rect 4344 3674 4396 3680
rect 4344 3596 4396 3602
rect 4344 3538 4396 3544
rect 4356 3369 4384 3538
rect 4342 3360 4398 3369
rect 4342 3295 4398 3304
rect 4344 2984 4396 2990
rect 4264 2944 4344 2972
rect 3804 2910 4016 2938
rect 4344 2926 4396 2932
rect 3700 2576 3752 2582
rect 3700 2518 3752 2524
rect 3804 2106 3832 2910
rect 4448 2854 4476 4694
rect 4540 4468 4568 5646
rect 4632 4622 4660 6054
rect 4620 4616 4672 4622
rect 4620 4558 4672 4564
rect 4816 4554 4844 8894
rect 5080 8832 5132 8838
rect 5080 8774 5132 8780
rect 5092 8498 5120 8774
rect 5170 8664 5226 8673
rect 5276 8650 5304 9590
rect 5226 8622 5304 8650
rect 5170 8599 5226 8608
rect 5080 8492 5132 8498
rect 5080 8434 5132 8440
rect 4896 8424 4948 8430
rect 4896 8366 4948 8372
rect 4908 5914 4936 8366
rect 4988 8288 5040 8294
rect 4988 8230 5040 8236
rect 5000 7410 5028 8230
rect 5172 7880 5224 7886
rect 5172 7822 5224 7828
rect 4988 7404 5040 7410
rect 4988 7346 5040 7352
rect 4896 5908 4948 5914
rect 4896 5850 4948 5856
rect 4804 4548 4856 4554
rect 4804 4490 4856 4496
rect 4540 4440 4660 4468
rect 4528 3936 4580 3942
rect 4528 3878 4580 3884
rect 4540 3194 4568 3878
rect 4632 3641 4660 4440
rect 4908 4282 4936 5850
rect 5080 5772 5132 5778
rect 5080 5714 5132 5720
rect 4988 5568 5040 5574
rect 4988 5510 5040 5516
rect 5000 4604 5028 5510
rect 5092 5370 5120 5714
rect 5080 5364 5132 5370
rect 5080 5306 5132 5312
rect 5078 5128 5134 5137
rect 5078 5063 5134 5072
rect 5092 4826 5120 5063
rect 5080 4820 5132 4826
rect 5080 4762 5132 4768
rect 5080 4616 5132 4622
rect 5000 4576 5080 4604
rect 5080 4558 5132 4564
rect 5092 4282 5120 4558
rect 4896 4276 4948 4282
rect 4896 4218 4948 4224
rect 5080 4276 5132 4282
rect 5080 4218 5132 4224
rect 4986 4176 5042 4185
rect 4724 4120 4986 4128
rect 4724 4111 5042 4120
rect 4724 4100 5028 4111
rect 4618 3632 4674 3641
rect 4618 3567 4674 3576
rect 4618 3496 4674 3505
rect 4618 3431 4674 3440
rect 4528 3188 4580 3194
rect 4528 3130 4580 3136
rect 4436 2848 4488 2854
rect 4436 2790 4488 2796
rect 3882 2748 4190 2757
rect 3882 2746 3888 2748
rect 3944 2746 3968 2748
rect 4024 2746 4048 2748
rect 4104 2746 4128 2748
rect 4184 2746 4190 2748
rect 3944 2694 3946 2746
rect 4126 2694 4128 2746
rect 3882 2692 3888 2694
rect 3944 2692 3968 2694
rect 4024 2692 4048 2694
rect 4104 2692 4128 2694
rect 4184 2692 4190 2694
rect 3882 2683 4190 2692
rect 4632 2582 4660 3431
rect 4620 2576 4672 2582
rect 4620 2518 4672 2524
rect 3974 2408 4030 2417
rect 3974 2343 4030 2352
rect 3792 2100 3844 2106
rect 3792 2042 3844 2048
rect 3988 1970 4016 2343
rect 3976 1964 4028 1970
rect 3976 1906 4028 1912
rect 3608 1760 3660 1766
rect 3608 1702 3660 1708
rect 3620 1426 3648 1702
rect 3882 1660 4190 1669
rect 3882 1658 3888 1660
rect 3944 1658 3968 1660
rect 4024 1658 4048 1660
rect 4104 1658 4128 1660
rect 4184 1658 4190 1660
rect 3944 1606 3946 1658
rect 4126 1606 4128 1658
rect 3882 1604 3888 1606
rect 3944 1604 3968 1606
rect 4024 1604 4048 1606
rect 4104 1604 4128 1606
rect 4184 1604 4190 1606
rect 3882 1595 4190 1604
rect 3790 1456 3846 1465
rect 3608 1420 3660 1426
rect 3790 1391 3846 1400
rect 3608 1362 3660 1368
rect 3804 1358 3832 1391
rect 3700 1352 3752 1358
rect 3700 1294 3752 1300
rect 3792 1352 3844 1358
rect 3792 1294 3844 1300
rect 3976 1352 4028 1358
rect 4436 1352 4488 1358
rect 3976 1294 4028 1300
rect 4434 1320 4436 1329
rect 4488 1320 4490 1329
rect 3332 750 3384 756
rect 3436 768 3556 796
rect 3436 160 3464 768
rect 3712 160 3740 1294
rect 3884 1216 3936 1222
rect 3884 1158 3936 1164
rect 3896 542 3924 1158
rect 3884 536 3936 542
rect 3884 478 3936 484
rect 3988 160 4016 1294
rect 4252 1284 4304 1290
rect 4434 1255 4490 1264
rect 4252 1226 4304 1232
rect 4068 1216 4120 1222
rect 4068 1158 4120 1164
rect 4080 785 4108 1158
rect 4066 776 4122 785
rect 4066 711 4122 720
rect 4264 160 4292 1226
rect 386 54 612 82
rect 386 -300 442 54
rect 662 -300 718 160
rect 938 -300 994 160
rect 1214 -300 1270 160
rect 1490 -300 1546 160
rect 1766 -300 1822 160
rect 2042 -300 2098 160
rect 2318 -300 2374 160
rect 2594 -300 2650 160
rect 2870 -300 2926 160
rect 3146 -300 3202 160
rect 3422 -300 3478 160
rect 3698 -300 3754 160
rect 3974 -300 4030 160
rect 4250 -300 4306 160
rect 4526 82 4582 160
rect 4724 82 4752 4100
rect 4988 3936 5040 3942
rect 4988 3878 5040 3884
rect 4802 3768 4858 3777
rect 4802 3703 4858 3712
rect 4896 3732 4948 3738
rect 4816 3369 4844 3703
rect 4896 3674 4948 3680
rect 4802 3360 4858 3369
rect 4802 3295 4858 3304
rect 4908 2106 4936 3674
rect 5000 3534 5028 3878
rect 5080 3732 5132 3738
rect 5080 3674 5132 3680
rect 4988 3528 5040 3534
rect 4988 3470 5040 3476
rect 5092 3210 5120 3674
rect 5000 3182 5120 3210
rect 5184 3194 5212 7822
rect 5368 5710 5396 13767
rect 5736 13326 5764 18226
rect 5724 13320 5776 13326
rect 5724 13262 5776 13268
rect 5540 12096 5592 12102
rect 5540 12038 5592 12044
rect 5448 11552 5500 11558
rect 5448 11494 5500 11500
rect 5460 11218 5488 11494
rect 5552 11354 5580 12038
rect 5632 11892 5684 11898
rect 5632 11834 5684 11840
rect 5540 11348 5592 11354
rect 5540 11290 5592 11296
rect 5448 11212 5500 11218
rect 5448 11154 5500 11160
rect 5644 10062 5672 11834
rect 5736 11694 5764 13262
rect 5724 11688 5776 11694
rect 5724 11630 5776 11636
rect 5724 11212 5776 11218
rect 5724 11154 5776 11160
rect 5736 10810 5764 11154
rect 5724 10804 5776 10810
rect 5724 10746 5776 10752
rect 5632 10056 5684 10062
rect 5632 9998 5684 10004
rect 5540 9716 5592 9722
rect 5540 9658 5592 9664
rect 5446 8936 5502 8945
rect 5446 8871 5502 8880
rect 5460 7410 5488 8871
rect 5552 8090 5580 9658
rect 5632 9512 5684 9518
rect 5632 9454 5684 9460
rect 5644 9042 5672 9454
rect 5724 9104 5776 9110
rect 5724 9046 5776 9052
rect 5632 9036 5684 9042
rect 5632 8978 5684 8984
rect 5540 8084 5592 8090
rect 5540 8026 5592 8032
rect 5448 7404 5500 7410
rect 5448 7346 5500 7352
rect 5644 6866 5672 8978
rect 5736 8362 5764 9046
rect 5724 8356 5776 8362
rect 5724 8298 5776 8304
rect 5736 7993 5764 8298
rect 5722 7984 5778 7993
rect 5722 7919 5778 7928
rect 5632 6860 5684 6866
rect 5632 6802 5684 6808
rect 5540 6792 5592 6798
rect 5540 6734 5592 6740
rect 5552 6390 5580 6734
rect 5632 6656 5684 6662
rect 5632 6598 5684 6604
rect 5724 6656 5776 6662
rect 5724 6598 5776 6604
rect 5540 6384 5592 6390
rect 5540 6326 5592 6332
rect 5644 5778 5672 6598
rect 5736 6458 5764 6598
rect 5724 6452 5776 6458
rect 5724 6394 5776 6400
rect 5632 5772 5684 5778
rect 5632 5714 5684 5720
rect 5356 5704 5408 5710
rect 5356 5646 5408 5652
rect 5368 4842 5396 5646
rect 5540 5092 5592 5098
rect 5540 5034 5592 5040
rect 5276 4814 5396 4842
rect 5552 4826 5580 5034
rect 5540 4820 5592 4826
rect 5276 3777 5304 4814
rect 5540 4762 5592 4768
rect 5448 4480 5500 4486
rect 5448 4422 5500 4428
rect 5356 4140 5408 4146
rect 5356 4082 5408 4088
rect 5262 3768 5318 3777
rect 5262 3703 5318 3712
rect 5172 3188 5224 3194
rect 5000 3126 5028 3182
rect 5172 3130 5224 3136
rect 4988 3120 5040 3126
rect 5368 3097 5396 4082
rect 4988 3062 5040 3068
rect 5354 3088 5410 3097
rect 5172 3052 5224 3058
rect 5354 3023 5410 3032
rect 5172 2994 5224 3000
rect 5184 2446 5212 2994
rect 5354 2680 5410 2689
rect 5460 2650 5488 4422
rect 5722 4312 5778 4321
rect 5722 4247 5778 4256
rect 5630 4176 5686 4185
rect 5630 4111 5632 4120
rect 5684 4111 5686 4120
rect 5632 4082 5684 4088
rect 5736 3738 5764 4247
rect 5724 3732 5776 3738
rect 5724 3674 5776 3680
rect 5632 3052 5684 3058
rect 5632 2994 5684 3000
rect 5354 2615 5356 2624
rect 5408 2615 5410 2624
rect 5448 2644 5500 2650
rect 5356 2586 5408 2592
rect 5448 2586 5500 2592
rect 5172 2440 5224 2446
rect 5172 2382 5224 2388
rect 5460 2378 5488 2586
rect 5448 2372 5500 2378
rect 5448 2314 5500 2320
rect 4896 2100 4948 2106
rect 4896 2042 4948 2048
rect 5356 1964 5408 1970
rect 5356 1906 5408 1912
rect 4988 1760 5040 1766
rect 4988 1702 5040 1708
rect 5000 1494 5028 1702
rect 4988 1488 5040 1494
rect 4988 1430 5040 1436
rect 5264 1284 5316 1290
rect 5264 1226 5316 1232
rect 4804 1216 4856 1222
rect 4804 1158 4856 1164
rect 4816 160 4844 1158
rect 4526 54 4752 82
rect 4526 -300 4582 54
rect 4802 -300 4858 160
rect 5078 82 5134 160
rect 5276 82 5304 1226
rect 5368 160 5396 1906
rect 5448 1284 5500 1290
rect 5448 1226 5500 1232
rect 5460 746 5488 1226
rect 5644 1034 5672 2994
rect 5828 1358 5856 20318
rect 5908 19780 5960 19786
rect 5908 19722 5960 19728
rect 5920 19689 5948 19722
rect 5906 19680 5962 19689
rect 5906 19615 5962 19624
rect 5908 19168 5960 19174
rect 5908 19110 5960 19116
rect 5920 18902 5948 19110
rect 5908 18896 5960 18902
rect 5908 18838 5960 18844
rect 6012 18136 6040 21270
rect 6196 20942 6224 21490
rect 6276 21412 6328 21418
rect 6276 21354 6328 21360
rect 6184 20936 6236 20942
rect 6184 20878 6236 20884
rect 6092 20800 6144 20806
rect 6092 20742 6144 20748
rect 6104 19174 6132 20742
rect 6092 19168 6144 19174
rect 6092 19110 6144 19116
rect 6092 18828 6144 18834
rect 6092 18770 6144 18776
rect 6104 18426 6132 18770
rect 6092 18420 6144 18426
rect 6092 18362 6144 18368
rect 6012 18108 6132 18136
rect 5908 18080 5960 18086
rect 5908 18022 5960 18028
rect 5998 18048 6054 18057
rect 5920 17202 5948 18022
rect 5998 17983 6054 17992
rect 5908 17196 5960 17202
rect 5908 17138 5960 17144
rect 5908 16992 5960 16998
rect 5908 16934 5960 16940
rect 5920 16794 5948 16934
rect 5908 16788 5960 16794
rect 5908 16730 5960 16736
rect 5908 16448 5960 16454
rect 5908 16390 5960 16396
rect 5920 16250 5948 16390
rect 5908 16244 5960 16250
rect 5908 16186 5960 16192
rect 5908 13728 5960 13734
rect 5908 13670 5960 13676
rect 5920 13462 5948 13670
rect 5908 13456 5960 13462
rect 5908 13398 5960 13404
rect 5906 12336 5962 12345
rect 5906 12271 5962 12280
rect 5920 9466 5948 12271
rect 6012 11121 6040 17983
rect 6104 17542 6132 18108
rect 6092 17536 6144 17542
rect 6092 17478 6144 17484
rect 6104 16998 6132 17478
rect 6196 17066 6224 20878
rect 6288 18193 6316 21354
rect 6368 20596 6420 20602
rect 6368 20538 6420 20544
rect 6380 19689 6408 20538
rect 6472 19786 6500 23122
rect 6564 22982 6592 24822
rect 6656 24070 6684 26182
rect 6748 24818 6776 31878
rect 6932 31686 6960 32370
rect 7208 32042 7236 32728
rect 7116 32014 7420 32042
rect 7116 31822 7144 32014
rect 7196 31884 7248 31890
rect 7196 31826 7248 31832
rect 7104 31816 7156 31822
rect 7104 31758 7156 31764
rect 6920 31680 6972 31686
rect 6920 31622 6972 31628
rect 6814 31580 7122 31589
rect 6814 31578 6820 31580
rect 6876 31578 6900 31580
rect 6956 31578 6980 31580
rect 7036 31578 7060 31580
rect 7116 31578 7122 31580
rect 6876 31526 6878 31578
rect 7058 31526 7060 31578
rect 6814 31524 6820 31526
rect 6876 31524 6900 31526
rect 6956 31524 6980 31526
rect 7036 31524 7060 31526
rect 7116 31524 7122 31526
rect 6814 31515 7122 31524
rect 7104 31204 7156 31210
rect 7104 31146 7156 31152
rect 7116 30802 7144 31146
rect 7208 30938 7236 31826
rect 7392 31686 7420 32014
rect 7288 31680 7340 31686
rect 7288 31622 7340 31628
rect 7380 31680 7432 31686
rect 7380 31622 7432 31628
rect 7196 30932 7248 30938
rect 7196 30874 7248 30880
rect 7104 30796 7156 30802
rect 7104 30738 7156 30744
rect 6814 30492 7122 30501
rect 6814 30490 6820 30492
rect 6876 30490 6900 30492
rect 6956 30490 6980 30492
rect 7036 30490 7060 30492
rect 7116 30490 7122 30492
rect 6876 30438 6878 30490
rect 7058 30438 7060 30490
rect 6814 30436 6820 30438
rect 6876 30436 6900 30438
rect 6956 30436 6980 30438
rect 7036 30436 7060 30438
rect 7116 30436 7122 30438
rect 6814 30427 7122 30436
rect 6828 30184 6880 30190
rect 6828 30126 6880 30132
rect 6840 30025 6868 30126
rect 6826 30016 6882 30025
rect 6826 29951 6882 29960
rect 7300 29578 7328 31622
rect 7484 31346 7512 32932
rect 7472 31340 7524 31346
rect 7472 31282 7524 31288
rect 7472 30864 7524 30870
rect 7472 30806 7524 30812
rect 7380 30728 7432 30734
rect 7484 30716 7512 30806
rect 7432 30688 7512 30716
rect 7380 30670 7432 30676
rect 7380 30184 7432 30190
rect 7380 30126 7432 30132
rect 7392 29646 7420 30126
rect 7380 29640 7432 29646
rect 7380 29582 7432 29588
rect 6828 29572 6880 29578
rect 7288 29572 7340 29578
rect 6880 29532 7236 29560
rect 6828 29514 6880 29520
rect 6814 29404 7122 29413
rect 6814 29402 6820 29404
rect 6876 29402 6900 29404
rect 6956 29402 6980 29404
rect 7036 29402 7060 29404
rect 7116 29402 7122 29404
rect 6876 29350 6878 29402
rect 7058 29350 7060 29402
rect 6814 29348 6820 29350
rect 6876 29348 6900 29350
rect 6956 29348 6980 29350
rect 7036 29348 7060 29350
rect 7116 29348 7122 29350
rect 6814 29339 7122 29348
rect 7208 29322 7236 29532
rect 7288 29514 7340 29520
rect 7484 29492 7512 30688
rect 7576 30598 7604 34972
rect 7668 34490 7696 35634
rect 7760 35086 7788 36110
rect 7852 35222 7880 40598
rect 7932 39296 7984 39302
rect 7932 39238 7984 39244
rect 7944 38962 7972 39238
rect 7932 38956 7984 38962
rect 7932 38898 7984 38904
rect 8036 38758 8064 42774
rect 8128 42650 8156 44540
rect 8404 43602 8432 44540
rect 8404 43574 8524 43602
rect 8496 42906 8524 43574
rect 8680 43178 8708 44540
rect 8956 43450 8984 44540
rect 8944 43444 8996 43450
rect 8944 43386 8996 43392
rect 9232 43330 9260 44540
rect 9508 43450 9536 44540
rect 9784 43450 9812 44540
rect 9864 43716 9916 43722
rect 9864 43658 9916 43664
rect 9876 43450 9904 43658
rect 10060 43636 10088 44540
rect 10060 43608 10180 43636
rect 9496 43444 9548 43450
rect 9496 43386 9548 43392
rect 9772 43444 9824 43450
rect 9772 43386 9824 43392
rect 9864 43444 9916 43450
rect 9864 43386 9916 43392
rect 9232 43302 9536 43330
rect 9128 43240 9180 43246
rect 9128 43182 9180 43188
rect 8668 43172 8720 43178
rect 8668 43114 8720 43120
rect 8484 42900 8536 42906
rect 8484 42842 8536 42848
rect 8944 42696 8996 42702
rect 8128 42634 8340 42650
rect 8944 42638 8996 42644
rect 8128 42628 8352 42634
rect 8128 42622 8300 42628
rect 8300 42570 8352 42576
rect 8300 42220 8352 42226
rect 8300 42162 8352 42168
rect 8114 42120 8170 42129
rect 8114 42055 8170 42064
rect 8128 41138 8156 42055
rect 8116 41132 8168 41138
rect 8116 41074 8168 41080
rect 8312 39846 8340 42162
rect 8956 41818 8984 42638
rect 9140 42362 9168 43182
rect 9508 42906 9536 43302
rect 9588 43308 9640 43314
rect 9588 43250 9640 43256
rect 9772 43308 9824 43314
rect 9772 43250 9824 43256
rect 9600 42906 9628 43250
rect 9678 43208 9734 43217
rect 9678 43143 9734 43152
rect 9692 43110 9720 43143
rect 9784 43110 9812 43250
rect 9680 43104 9732 43110
rect 9680 43046 9732 43052
rect 9772 43104 9824 43110
rect 9772 43046 9824 43052
rect 9747 43004 10055 43013
rect 9747 43002 9753 43004
rect 9809 43002 9833 43004
rect 9889 43002 9913 43004
rect 9969 43002 9993 43004
rect 10049 43002 10055 43004
rect 9809 42950 9811 43002
rect 9991 42950 9993 43002
rect 9747 42948 9753 42950
rect 9809 42948 9833 42950
rect 9889 42948 9913 42950
rect 9969 42948 9993 42950
rect 10049 42948 10055 42950
rect 9747 42939 10055 42948
rect 9496 42900 9548 42906
rect 9496 42842 9548 42848
rect 9588 42900 9640 42906
rect 9588 42842 9640 42848
rect 9954 42800 10010 42809
rect 9496 42764 9548 42770
rect 9954 42735 10010 42744
rect 9496 42706 9548 42712
rect 9220 42628 9272 42634
rect 9220 42570 9272 42576
rect 9404 42628 9456 42634
rect 9404 42570 9456 42576
rect 9128 42356 9180 42362
rect 9128 42298 9180 42304
rect 9036 42220 9088 42226
rect 9036 42162 9088 42168
rect 9048 41857 9076 42162
rect 9034 41848 9090 41857
rect 8944 41812 8996 41818
rect 9232 41818 9260 42570
rect 9312 42220 9364 42226
rect 9312 42162 9364 42168
rect 9324 41993 9352 42162
rect 9310 41984 9366 41993
rect 9310 41919 9366 41928
rect 9034 41783 9090 41792
rect 9220 41812 9272 41818
rect 8944 41754 8996 41760
rect 9220 41754 9272 41760
rect 9128 41608 9180 41614
rect 9126 41576 9128 41585
rect 9220 41608 9272 41614
rect 9180 41576 9182 41585
rect 9220 41550 9272 41556
rect 9126 41511 9182 41520
rect 8484 41472 8536 41478
rect 8484 41414 8536 41420
rect 8496 41206 8524 41414
rect 8484 41200 8536 41206
rect 8484 41142 8536 41148
rect 8668 41132 8720 41138
rect 8668 41074 8720 41080
rect 8680 40497 8708 41074
rect 8666 40488 8722 40497
rect 8666 40423 8722 40432
rect 8300 39840 8352 39846
rect 8300 39782 8352 39788
rect 8208 39636 8260 39642
rect 8208 39578 8260 39584
rect 8116 39432 8168 39438
rect 8116 39374 8168 39380
rect 8024 38752 8076 38758
rect 8024 38694 8076 38700
rect 8128 38570 8156 39374
rect 8036 38542 8156 38570
rect 8036 37194 8064 38542
rect 8220 38282 8248 39578
rect 8576 38752 8628 38758
rect 8576 38694 8628 38700
rect 8588 38350 8616 38694
rect 8576 38344 8628 38350
rect 8576 38286 8628 38292
rect 8208 38276 8260 38282
rect 8208 38218 8260 38224
rect 8220 37754 8248 38218
rect 8128 37726 8248 37754
rect 8024 37188 8076 37194
rect 8024 37130 8076 37136
rect 7932 37120 7984 37126
rect 7932 37062 7984 37068
rect 7944 36718 7972 37062
rect 7932 36712 7984 36718
rect 7932 36654 7984 36660
rect 8036 36417 8064 37130
rect 8022 36408 8078 36417
rect 8022 36343 8078 36352
rect 7840 35216 7892 35222
rect 7840 35158 7892 35164
rect 7748 35080 7800 35086
rect 7748 35022 7800 35028
rect 7852 34513 7880 35158
rect 7838 34504 7894 34513
rect 7668 34462 7788 34490
rect 7656 34400 7708 34406
rect 7656 34342 7708 34348
rect 7668 33998 7696 34342
rect 7656 33992 7708 33998
rect 7656 33934 7708 33940
rect 7760 33946 7788 34462
rect 7838 34439 7894 34448
rect 7840 34128 7892 34134
rect 7838 34096 7840 34105
rect 7892 34096 7894 34105
rect 7838 34031 7894 34040
rect 7760 33918 7972 33946
rect 7944 33862 7972 33918
rect 7932 33856 7984 33862
rect 7932 33798 7984 33804
rect 7656 33652 7708 33658
rect 7656 33594 7708 33600
rect 7668 33454 7696 33594
rect 7932 33516 7984 33522
rect 7932 33458 7984 33464
rect 7656 33448 7708 33454
rect 7656 33390 7708 33396
rect 7748 32904 7800 32910
rect 7748 32846 7800 32852
rect 7760 32473 7788 32846
rect 7746 32464 7802 32473
rect 7746 32399 7802 32408
rect 7656 32360 7708 32366
rect 7944 32337 7972 33458
rect 8128 33436 8156 37726
rect 8208 37120 8260 37126
rect 8208 37062 8260 37068
rect 8220 36786 8248 37062
rect 8680 36854 8708 40423
rect 9232 39545 9260 41550
rect 9416 39642 9444 42570
rect 9508 40594 9536 42706
rect 9968 42362 9996 42735
rect 10152 42702 10180 43608
rect 10232 43308 10284 43314
rect 10232 43250 10284 43256
rect 10244 42838 10272 43250
rect 10232 42832 10284 42838
rect 10232 42774 10284 42780
rect 10140 42696 10192 42702
rect 10140 42638 10192 42644
rect 10232 42696 10284 42702
rect 10336 42684 10364 44540
rect 10508 43240 10560 43246
rect 10508 43182 10560 43188
rect 10416 43172 10468 43178
rect 10416 43114 10468 43120
rect 10284 42656 10364 42684
rect 10232 42638 10284 42644
rect 10140 42560 10192 42566
rect 10138 42528 10140 42537
rect 10192 42528 10194 42537
rect 10138 42463 10194 42472
rect 9956 42356 10008 42362
rect 10428 42344 10456 43114
rect 9956 42298 10008 42304
rect 10336 42316 10456 42344
rect 10140 42220 10192 42226
rect 10140 42162 10192 42168
rect 9747 41916 10055 41925
rect 9747 41914 9753 41916
rect 9809 41914 9833 41916
rect 9889 41914 9913 41916
rect 9969 41914 9993 41916
rect 10049 41914 10055 41916
rect 9809 41862 9811 41914
rect 9991 41862 9993 41914
rect 9747 41860 9753 41862
rect 9809 41860 9833 41862
rect 9889 41860 9913 41862
rect 9969 41860 9993 41862
rect 10049 41860 10055 41862
rect 9747 41851 10055 41860
rect 9747 40828 10055 40837
rect 9747 40826 9753 40828
rect 9809 40826 9833 40828
rect 9889 40826 9913 40828
rect 9969 40826 9993 40828
rect 10049 40826 10055 40828
rect 9809 40774 9811 40826
rect 9991 40774 9993 40826
rect 9747 40772 9753 40774
rect 9809 40772 9833 40774
rect 9889 40772 9913 40774
rect 9969 40772 9993 40774
rect 10049 40772 10055 40774
rect 9747 40763 10055 40772
rect 9496 40588 9548 40594
rect 9496 40530 9548 40536
rect 9747 39740 10055 39749
rect 9747 39738 9753 39740
rect 9809 39738 9833 39740
rect 9889 39738 9913 39740
rect 9969 39738 9993 39740
rect 10049 39738 10055 39740
rect 9809 39686 9811 39738
rect 9991 39686 9993 39738
rect 9747 39684 9753 39686
rect 9809 39684 9833 39686
rect 9889 39684 9913 39686
rect 9969 39684 9993 39686
rect 10049 39684 10055 39686
rect 9747 39675 10055 39684
rect 9404 39636 9456 39642
rect 9404 39578 9456 39584
rect 9218 39536 9274 39545
rect 10152 39522 10180 42162
rect 10232 41744 10284 41750
rect 10232 41686 10284 41692
rect 10244 39642 10272 41686
rect 10232 39636 10284 39642
rect 10232 39578 10284 39584
rect 9218 39471 9274 39480
rect 9876 39494 10180 39522
rect 9496 39432 9548 39438
rect 8758 39400 8814 39409
rect 8758 39335 8814 39344
rect 9232 39392 9496 39420
rect 8392 36848 8444 36854
rect 8392 36790 8444 36796
rect 8668 36848 8720 36854
rect 8668 36790 8720 36796
rect 8208 36780 8260 36786
rect 8208 36722 8260 36728
rect 8220 33590 8248 36722
rect 8300 36168 8352 36174
rect 8298 36136 8300 36145
rect 8352 36136 8354 36145
rect 8298 36071 8354 36080
rect 8404 35834 8432 36790
rect 8484 36032 8536 36038
rect 8484 35974 8536 35980
rect 8392 35828 8444 35834
rect 8392 35770 8444 35776
rect 8496 35630 8524 35974
rect 8484 35624 8536 35630
rect 8298 35592 8354 35601
rect 8484 35566 8536 35572
rect 8298 35527 8354 35536
rect 8208 33584 8260 33590
rect 8208 33526 8260 33532
rect 8128 33408 8248 33436
rect 8116 32768 8168 32774
rect 8116 32710 8168 32716
rect 8128 32366 8156 32710
rect 8116 32360 8168 32366
rect 7656 32302 7708 32308
rect 7930 32328 7986 32337
rect 7668 31872 7696 32302
rect 8116 32302 8168 32308
rect 7930 32263 7986 32272
rect 8024 32292 8076 32298
rect 8024 32234 8076 32240
rect 7668 31844 7788 31872
rect 7654 31648 7710 31657
rect 7654 31583 7710 31592
rect 7564 30592 7616 30598
rect 7564 30534 7616 30540
rect 7668 30258 7696 31583
rect 7760 31482 7788 31844
rect 8036 31822 8064 32234
rect 8128 32026 8156 32302
rect 8116 32020 8168 32026
rect 8116 31962 8168 31968
rect 7840 31816 7892 31822
rect 7840 31758 7892 31764
rect 8024 31816 8076 31822
rect 8024 31758 8076 31764
rect 7748 31476 7800 31482
rect 7748 31418 7800 31424
rect 7656 30252 7708 30258
rect 7656 30194 7708 30200
rect 7392 29464 7512 29492
rect 7208 29306 7328 29322
rect 7208 29300 7340 29306
rect 7208 29294 7288 29300
rect 7288 29242 7340 29248
rect 7196 29232 7248 29238
rect 7196 29174 7248 29180
rect 7208 29034 7236 29174
rect 7196 29028 7248 29034
rect 7196 28970 7248 28976
rect 6814 28316 7122 28325
rect 6814 28314 6820 28316
rect 6876 28314 6900 28316
rect 6956 28314 6980 28316
rect 7036 28314 7060 28316
rect 7116 28314 7122 28316
rect 6876 28262 6878 28314
rect 7058 28262 7060 28314
rect 6814 28260 6820 28262
rect 6876 28260 6900 28262
rect 6956 28260 6980 28262
rect 7036 28260 7060 28262
rect 7116 28260 7122 28262
rect 6814 28251 7122 28260
rect 7208 27334 7236 28970
rect 7286 27568 7342 27577
rect 7286 27503 7342 27512
rect 7300 27470 7328 27503
rect 7288 27464 7340 27470
rect 7288 27406 7340 27412
rect 7196 27328 7248 27334
rect 7196 27270 7248 27276
rect 7288 27328 7340 27334
rect 7392 27305 7420 29464
rect 7472 29096 7524 29102
rect 7472 29038 7524 29044
rect 7288 27270 7340 27276
rect 7378 27296 7434 27305
rect 6814 27228 7122 27237
rect 6814 27226 6820 27228
rect 6876 27226 6900 27228
rect 6956 27226 6980 27228
rect 7036 27226 7060 27228
rect 7116 27226 7122 27228
rect 6876 27174 6878 27226
rect 7058 27174 7060 27226
rect 6814 27172 6820 27174
rect 6876 27172 6900 27174
rect 6956 27172 6980 27174
rect 7036 27172 7060 27174
rect 7116 27172 7122 27174
rect 6814 27163 7122 27172
rect 7300 27062 7328 27270
rect 7378 27231 7434 27240
rect 6828 27056 6880 27062
rect 6828 26998 6880 27004
rect 7288 27056 7340 27062
rect 7288 26998 7340 27004
rect 6840 26586 6868 26998
rect 7196 26920 7248 26926
rect 7196 26862 7248 26868
rect 7208 26586 7236 26862
rect 6828 26580 6880 26586
rect 6828 26522 6880 26528
rect 7196 26580 7248 26586
rect 7196 26522 7248 26528
rect 6814 26140 7122 26149
rect 6814 26138 6820 26140
rect 6876 26138 6900 26140
rect 6956 26138 6980 26140
rect 7036 26138 7060 26140
rect 7116 26138 7122 26140
rect 6876 26086 6878 26138
rect 7058 26086 7060 26138
rect 6814 26084 6820 26086
rect 6876 26084 6900 26086
rect 6956 26084 6980 26086
rect 7036 26084 7060 26086
rect 7116 26084 7122 26086
rect 6814 26075 7122 26084
rect 6828 25764 6880 25770
rect 6828 25706 6880 25712
rect 6840 25362 6868 25706
rect 6828 25356 6880 25362
rect 6828 25298 6880 25304
rect 7196 25152 7248 25158
rect 7196 25094 7248 25100
rect 6814 25052 7122 25061
rect 6814 25050 6820 25052
rect 6876 25050 6900 25052
rect 6956 25050 6980 25052
rect 7036 25050 7060 25052
rect 7116 25050 7122 25052
rect 6876 24998 6878 25050
rect 7058 24998 7060 25050
rect 6814 24996 6820 24998
rect 6876 24996 6900 24998
rect 6956 24996 6980 24998
rect 7036 24996 7060 24998
rect 7116 24996 7122 24998
rect 6814 24987 7122 24996
rect 7104 24948 7156 24954
rect 7104 24890 7156 24896
rect 6736 24812 6788 24818
rect 6736 24754 6788 24760
rect 6644 24064 6696 24070
rect 6644 24006 6696 24012
rect 6552 22976 6604 22982
rect 6552 22918 6604 22924
rect 6748 22794 6776 24754
rect 7116 24070 7144 24890
rect 7208 24886 7236 25094
rect 7196 24880 7248 24886
rect 7196 24822 7248 24828
rect 7104 24064 7156 24070
rect 7104 24006 7156 24012
rect 6814 23964 7122 23973
rect 6814 23962 6820 23964
rect 6876 23962 6900 23964
rect 6956 23962 6980 23964
rect 7036 23962 7060 23964
rect 7116 23962 7122 23964
rect 6876 23910 6878 23962
rect 7058 23910 7060 23962
rect 6814 23908 6820 23910
rect 6876 23908 6900 23910
rect 6956 23908 6980 23910
rect 7036 23908 7060 23910
rect 7116 23908 7122 23910
rect 6814 23899 7122 23908
rect 7196 23860 7248 23866
rect 7196 23802 7248 23808
rect 7104 23588 7156 23594
rect 7104 23530 7156 23536
rect 7116 23322 7144 23530
rect 7104 23316 7156 23322
rect 7104 23258 7156 23264
rect 6814 22876 7122 22885
rect 6814 22874 6820 22876
rect 6876 22874 6900 22876
rect 6956 22874 6980 22876
rect 7036 22874 7060 22876
rect 7116 22874 7122 22876
rect 6876 22822 6878 22874
rect 7058 22822 7060 22874
rect 6814 22820 6820 22822
rect 6876 22820 6900 22822
rect 6956 22820 6980 22822
rect 7036 22820 7060 22822
rect 7116 22820 7122 22822
rect 6814 22811 7122 22820
rect 6564 22766 6776 22794
rect 7208 22778 7236 23802
rect 7300 23594 7328 26998
rect 7484 26994 7512 29038
rect 7668 28994 7696 30194
rect 7576 28966 7696 28994
rect 7472 26988 7524 26994
rect 7472 26930 7524 26936
rect 7484 26761 7512 26930
rect 7470 26752 7526 26761
rect 7470 26687 7526 26696
rect 7378 26616 7434 26625
rect 7378 26551 7434 26560
rect 7392 26450 7420 26551
rect 7470 26480 7526 26489
rect 7380 26444 7432 26450
rect 7470 26415 7526 26424
rect 7380 26386 7432 26392
rect 7380 26240 7432 26246
rect 7380 26182 7432 26188
rect 7392 25906 7420 26182
rect 7380 25900 7432 25906
rect 7380 25842 7432 25848
rect 7392 25294 7420 25842
rect 7380 25288 7432 25294
rect 7380 25230 7432 25236
rect 7484 24954 7512 26415
rect 7472 24948 7524 24954
rect 7472 24890 7524 24896
rect 7380 24268 7432 24274
rect 7380 24210 7432 24216
rect 7392 23594 7420 24210
rect 7472 24132 7524 24138
rect 7472 24074 7524 24080
rect 7288 23588 7340 23594
rect 7288 23530 7340 23536
rect 7380 23588 7432 23594
rect 7380 23530 7432 23536
rect 7484 23474 7512 24074
rect 7576 23730 7604 28966
rect 7654 28520 7710 28529
rect 7654 28455 7710 28464
rect 7668 28422 7696 28455
rect 7656 28416 7708 28422
rect 7656 28358 7708 28364
rect 7656 28008 7708 28014
rect 7656 27950 7708 27956
rect 7668 25945 7696 27950
rect 7760 27946 7788 31418
rect 7852 28966 7880 31758
rect 8036 31686 8064 31758
rect 7932 31680 7984 31686
rect 7932 31622 7984 31628
rect 8024 31680 8076 31686
rect 8024 31622 8076 31628
rect 7944 30682 7972 31622
rect 8220 31346 8248 33408
rect 8312 33046 8340 35527
rect 8680 35476 8708 36790
rect 8404 35448 8708 35476
rect 8300 33040 8352 33046
rect 8300 32982 8352 32988
rect 8208 31340 8260 31346
rect 8208 31282 8260 31288
rect 8114 31104 8170 31113
rect 8114 31039 8170 31048
rect 8128 30734 8156 31039
rect 8116 30728 8168 30734
rect 7944 30654 8064 30682
rect 8116 30670 8168 30676
rect 7932 30592 7984 30598
rect 7932 30534 7984 30540
rect 7840 28960 7892 28966
rect 7840 28902 7892 28908
rect 7748 27940 7800 27946
rect 7748 27882 7800 27888
rect 7760 27334 7788 27882
rect 7748 27328 7800 27334
rect 7748 27270 7800 27276
rect 7840 27124 7892 27130
rect 7840 27066 7892 27072
rect 7852 26382 7880 27066
rect 7840 26376 7892 26382
rect 7840 26318 7892 26324
rect 7748 26240 7800 26246
rect 7748 26182 7800 26188
rect 7654 25936 7710 25945
rect 7654 25871 7710 25880
rect 7656 24948 7708 24954
rect 7656 24890 7708 24896
rect 7668 24138 7696 24890
rect 7656 24132 7708 24138
rect 7656 24074 7708 24080
rect 7654 24032 7710 24041
rect 7654 23967 7710 23976
rect 7668 23730 7696 23967
rect 7564 23724 7616 23730
rect 7564 23666 7616 23672
rect 7656 23724 7708 23730
rect 7656 23666 7708 23672
rect 7300 23446 7512 23474
rect 7196 22772 7248 22778
rect 6564 22030 6592 22766
rect 7196 22714 7248 22720
rect 6736 22636 6788 22642
rect 6736 22578 6788 22584
rect 6644 22568 6696 22574
rect 6644 22510 6696 22516
rect 6656 22030 6684 22510
rect 6552 22024 6604 22030
rect 6552 21966 6604 21972
rect 6644 22024 6696 22030
rect 6644 21966 6696 21972
rect 6564 21554 6592 21966
rect 6552 21548 6604 21554
rect 6552 21490 6604 21496
rect 6552 21344 6604 21350
rect 6552 21286 6604 21292
rect 6564 20806 6592 21286
rect 6552 20800 6604 20806
rect 6552 20742 6604 20748
rect 6656 20466 6684 21966
rect 6748 21418 6776 22578
rect 7196 22500 7248 22506
rect 7196 22442 7248 22448
rect 7208 22098 7236 22442
rect 7300 22166 7328 23446
rect 7760 23338 7788 26182
rect 7838 24712 7894 24721
rect 7838 24647 7840 24656
rect 7892 24647 7894 24656
rect 7840 24618 7892 24624
rect 7380 23316 7432 23322
rect 7380 23258 7432 23264
rect 7484 23310 7788 23338
rect 7288 22160 7340 22166
rect 7288 22102 7340 22108
rect 7196 22092 7248 22098
rect 7196 22034 7248 22040
rect 7392 22012 7420 23258
rect 7300 21984 7420 22012
rect 6814 21788 7122 21797
rect 6814 21786 6820 21788
rect 6876 21786 6900 21788
rect 6956 21786 6980 21788
rect 7036 21786 7060 21788
rect 7116 21786 7122 21788
rect 6876 21734 6878 21786
rect 7058 21734 7060 21786
rect 6814 21732 6820 21734
rect 6876 21732 6900 21734
rect 6956 21732 6980 21734
rect 7036 21732 7060 21734
rect 7116 21732 7122 21734
rect 6814 21723 7122 21732
rect 6736 21412 6788 21418
rect 6736 21354 6788 21360
rect 6920 20936 6972 20942
rect 6748 20896 6920 20924
rect 6748 20602 6776 20896
rect 6920 20878 6972 20884
rect 6814 20700 7122 20709
rect 6814 20698 6820 20700
rect 6876 20698 6900 20700
rect 6956 20698 6980 20700
rect 7036 20698 7060 20700
rect 7116 20698 7122 20700
rect 6876 20646 6878 20698
rect 7058 20646 7060 20698
rect 6814 20644 6820 20646
rect 6876 20644 6900 20646
rect 6956 20644 6980 20646
rect 7036 20644 7060 20646
rect 7116 20644 7122 20646
rect 6814 20635 7122 20644
rect 6736 20596 6788 20602
rect 6736 20538 6788 20544
rect 6644 20460 6696 20466
rect 6644 20402 6696 20408
rect 7196 20392 7248 20398
rect 7196 20334 7248 20340
rect 6460 19780 6512 19786
rect 6460 19722 6512 19728
rect 6366 19680 6422 19689
rect 6366 19615 6422 19624
rect 6380 19242 6408 19615
rect 6368 19236 6420 19242
rect 6368 19178 6420 19184
rect 6472 19145 6500 19722
rect 6828 19712 6880 19718
rect 6748 19672 6828 19700
rect 6644 19372 6696 19378
rect 6644 19314 6696 19320
rect 6552 19236 6604 19242
rect 6552 19178 6604 19184
rect 6458 19136 6514 19145
rect 6458 19071 6514 19080
rect 6368 18964 6420 18970
rect 6368 18906 6420 18912
rect 6380 18834 6408 18906
rect 6564 18834 6592 19178
rect 6368 18828 6420 18834
rect 6368 18770 6420 18776
rect 6552 18828 6604 18834
rect 6552 18770 6604 18776
rect 6380 18290 6408 18770
rect 6656 18714 6684 19314
rect 6748 19242 6776 19672
rect 6828 19654 6880 19660
rect 6814 19612 7122 19621
rect 6814 19610 6820 19612
rect 6876 19610 6900 19612
rect 6956 19610 6980 19612
rect 7036 19610 7060 19612
rect 7116 19610 7122 19612
rect 6876 19558 6878 19610
rect 7058 19558 7060 19610
rect 6814 19556 6820 19558
rect 6876 19556 6900 19558
rect 6956 19556 6980 19558
rect 7036 19556 7060 19558
rect 7116 19556 7122 19558
rect 6814 19547 7122 19556
rect 7208 19496 7236 20334
rect 6932 19468 7236 19496
rect 6932 19378 6960 19468
rect 6920 19372 6972 19378
rect 6920 19314 6972 19320
rect 6736 19236 6788 19242
rect 6736 19178 6788 19184
rect 7300 18970 7328 21984
rect 7378 20496 7434 20505
rect 7378 20431 7434 20440
rect 7392 19786 7420 20431
rect 7380 19780 7432 19786
rect 7380 19722 7432 19728
rect 7484 19666 7512 23310
rect 7654 23080 7710 23089
rect 7944 23050 7972 30534
rect 8036 29102 8064 30654
rect 8404 30138 8432 35448
rect 8772 35306 8800 39335
rect 8944 38956 8996 38962
rect 8944 38898 8996 38904
rect 8956 38554 8984 38898
rect 8944 38548 8996 38554
rect 8944 38490 8996 38496
rect 9232 38214 9260 39392
rect 9496 39374 9548 39380
rect 9588 39432 9640 39438
rect 9588 39374 9640 39380
rect 9312 39296 9364 39302
rect 9312 39238 9364 39244
rect 9404 39296 9456 39302
rect 9404 39238 9456 39244
rect 9496 39296 9548 39302
rect 9496 39238 9548 39244
rect 9220 38208 9272 38214
rect 9220 38150 9272 38156
rect 9128 37664 9180 37670
rect 9128 37606 9180 37612
rect 8852 37256 8904 37262
rect 8852 37198 8904 37204
rect 8588 35278 8800 35306
rect 8484 32224 8536 32230
rect 8484 32166 8536 32172
rect 8496 32026 8524 32166
rect 8484 32020 8536 32026
rect 8484 31962 8536 31968
rect 8588 31754 8616 35278
rect 8668 34400 8720 34406
rect 8668 34342 8720 34348
rect 8680 34202 8708 34342
rect 8668 34196 8720 34202
rect 8668 34138 8720 34144
rect 8864 33454 8892 37198
rect 9140 36786 9168 37606
rect 9220 37256 9272 37262
rect 9220 37198 9272 37204
rect 9128 36780 9180 36786
rect 9128 36722 9180 36728
rect 8944 36576 8996 36582
rect 9036 36576 9088 36582
rect 8944 36518 8996 36524
rect 9034 36544 9036 36553
rect 9088 36544 9090 36553
rect 8956 35850 8984 36518
rect 9034 36479 9090 36488
rect 9140 36378 9168 36722
rect 9128 36372 9180 36378
rect 9128 36314 9180 36320
rect 9232 36258 9260 37198
rect 9140 36230 9260 36258
rect 8956 35822 9076 35850
rect 8944 35760 8996 35766
rect 8944 35702 8996 35708
rect 8956 35222 8984 35702
rect 8944 35216 8996 35222
rect 8944 35158 8996 35164
rect 8852 33448 8904 33454
rect 8852 33390 8904 33396
rect 8760 33312 8812 33318
rect 8852 33312 8904 33318
rect 8760 33254 8812 33260
rect 8850 33280 8852 33289
rect 8904 33280 8906 33289
rect 8772 32434 8800 33254
rect 8850 33215 8906 33224
rect 8760 32428 8812 32434
rect 8680 32388 8760 32416
rect 8680 31890 8708 32388
rect 8760 32370 8812 32376
rect 8956 32366 8984 35158
rect 8944 32360 8996 32366
rect 8944 32302 8996 32308
rect 8760 32224 8812 32230
rect 8758 32192 8760 32201
rect 8812 32192 8814 32201
rect 8758 32127 8814 32136
rect 8772 31890 8984 31906
rect 8668 31884 8720 31890
rect 8668 31826 8720 31832
rect 8772 31884 8996 31890
rect 8772 31878 8944 31884
rect 8312 30110 8432 30138
rect 8496 31726 8616 31754
rect 8116 29164 8168 29170
rect 8116 29106 8168 29112
rect 8024 29096 8076 29102
rect 8024 29038 8076 29044
rect 8036 27418 8064 29038
rect 8128 27538 8156 29106
rect 8208 28076 8260 28082
rect 8208 28018 8260 28024
rect 8220 27690 8248 28018
rect 8312 27826 8340 30110
rect 8392 30048 8444 30054
rect 8392 29990 8444 29996
rect 8404 29102 8432 29990
rect 8392 29096 8444 29102
rect 8392 29038 8444 29044
rect 8404 28014 8432 29038
rect 8392 28008 8444 28014
rect 8392 27950 8444 27956
rect 8312 27798 8432 27826
rect 8220 27662 8340 27690
rect 8116 27532 8168 27538
rect 8116 27474 8168 27480
rect 8036 27390 8248 27418
rect 8024 27328 8076 27334
rect 8024 27270 8076 27276
rect 8116 27328 8168 27334
rect 8116 27270 8168 27276
rect 8036 27062 8064 27270
rect 8024 27056 8076 27062
rect 8024 26998 8076 27004
rect 7654 23015 7710 23024
rect 7932 23044 7984 23050
rect 7564 22976 7616 22982
rect 7564 22918 7616 22924
rect 7576 22642 7604 22918
rect 7564 22636 7616 22642
rect 7564 22578 7616 22584
rect 7668 19854 7696 23015
rect 7932 22986 7984 22992
rect 7748 22976 7800 22982
rect 7748 22918 7800 22924
rect 7760 22681 7788 22918
rect 7746 22672 7802 22681
rect 8128 22658 8156 27270
rect 8220 26246 8248 27390
rect 8208 26240 8260 26246
rect 8208 26182 8260 26188
rect 8312 25294 8340 27662
rect 8404 27130 8432 27798
rect 8496 27169 8524 31726
rect 8772 31482 8800 31878
rect 8944 31826 8996 31832
rect 9048 31754 9076 35822
rect 9140 34524 9168 36230
rect 9220 35692 9272 35698
rect 9220 35634 9272 35640
rect 9232 34678 9260 35634
rect 9220 34672 9272 34678
rect 9220 34614 9272 34620
rect 9140 34496 9260 34524
rect 9128 33992 9180 33998
rect 9128 33934 9180 33940
rect 9140 32026 9168 33934
rect 9232 33538 9260 34496
rect 9324 34082 9352 39238
rect 9416 38010 9444 39238
rect 9508 39030 9536 39238
rect 9600 39098 9628 39374
rect 9772 39364 9824 39370
rect 9772 39306 9824 39312
rect 9784 39098 9812 39306
rect 9588 39092 9640 39098
rect 9588 39034 9640 39040
rect 9772 39092 9824 39098
rect 9772 39034 9824 39040
rect 9496 39024 9548 39030
rect 9496 38966 9548 38972
rect 9876 38865 9904 39494
rect 10046 39128 10102 39137
rect 10046 39063 10102 39072
rect 10060 39030 10088 39063
rect 10048 39024 10100 39030
rect 10244 38978 10272 39578
rect 10048 38966 10100 38972
rect 10152 38950 10272 38978
rect 9862 38856 9918 38865
rect 9862 38791 9918 38800
rect 9747 38652 10055 38661
rect 9747 38650 9753 38652
rect 9809 38650 9833 38652
rect 9889 38650 9913 38652
rect 9969 38650 9993 38652
rect 10049 38650 10055 38652
rect 9809 38598 9811 38650
rect 9991 38598 9993 38650
rect 9747 38596 9753 38598
rect 9809 38596 9833 38598
rect 9889 38596 9913 38598
rect 9969 38596 9993 38598
rect 10049 38596 10055 38598
rect 9747 38587 10055 38596
rect 10152 38554 10180 38950
rect 10232 38888 10284 38894
rect 10232 38830 10284 38836
rect 10244 38554 10272 38830
rect 10140 38548 10192 38554
rect 10140 38490 10192 38496
rect 10232 38548 10284 38554
rect 10232 38490 10284 38496
rect 10232 38412 10284 38418
rect 10232 38354 10284 38360
rect 9496 38344 9548 38350
rect 9496 38286 9548 38292
rect 9404 38004 9456 38010
rect 9404 37946 9456 37952
rect 9404 37188 9456 37194
rect 9404 37130 9456 37136
rect 9416 36378 9444 37130
rect 9404 36372 9456 36378
rect 9404 36314 9456 36320
rect 9404 34196 9456 34202
rect 9508 34184 9536 38286
rect 9747 37564 10055 37573
rect 9747 37562 9753 37564
rect 9809 37562 9833 37564
rect 9889 37562 9913 37564
rect 9969 37562 9993 37564
rect 10049 37562 10055 37564
rect 9809 37510 9811 37562
rect 9991 37510 9993 37562
rect 9747 37508 9753 37510
rect 9809 37508 9833 37510
rect 9889 37508 9913 37510
rect 9969 37508 9993 37510
rect 10049 37508 10055 37510
rect 9747 37499 10055 37508
rect 10244 37398 10272 38354
rect 10232 37392 10284 37398
rect 10232 37334 10284 37340
rect 10244 37262 10272 37334
rect 10232 37256 10284 37262
rect 10232 37198 10284 37204
rect 10138 36816 10194 36825
rect 10138 36751 10140 36760
rect 10192 36751 10194 36760
rect 10140 36722 10192 36728
rect 10232 36576 10284 36582
rect 10232 36518 10284 36524
rect 9747 36476 10055 36485
rect 9747 36474 9753 36476
rect 9809 36474 9833 36476
rect 9889 36474 9913 36476
rect 9969 36474 9993 36476
rect 10049 36474 10055 36476
rect 9809 36422 9811 36474
rect 9991 36422 9993 36474
rect 9747 36420 9753 36422
rect 9809 36420 9833 36422
rect 9889 36420 9913 36422
rect 9969 36420 9993 36422
rect 10049 36420 10055 36422
rect 9747 36411 10055 36420
rect 10244 36242 10272 36518
rect 10232 36236 10284 36242
rect 10232 36178 10284 36184
rect 9772 36032 9824 36038
rect 9772 35974 9824 35980
rect 9784 35766 9812 35974
rect 9772 35760 9824 35766
rect 10048 35760 10100 35766
rect 9772 35702 9824 35708
rect 9876 35720 10048 35748
rect 9876 35544 9904 35720
rect 10048 35702 10100 35708
rect 10244 35698 10272 36178
rect 10140 35692 10192 35698
rect 10140 35634 10192 35640
rect 10232 35692 10284 35698
rect 10232 35634 10284 35640
rect 9646 35516 9904 35544
rect 9646 35476 9674 35516
rect 9600 35448 9674 35476
rect 9600 34746 9628 35448
rect 9747 35388 10055 35397
rect 9747 35386 9753 35388
rect 9809 35386 9833 35388
rect 9889 35386 9913 35388
rect 9969 35386 9993 35388
rect 10049 35386 10055 35388
rect 9809 35334 9811 35386
rect 9991 35334 9993 35386
rect 9747 35332 9753 35334
rect 9809 35332 9833 35334
rect 9889 35332 9913 35334
rect 9969 35332 9993 35334
rect 10049 35332 10055 35334
rect 9747 35323 10055 35332
rect 9588 34740 9640 34746
rect 9588 34682 9640 34688
rect 9747 34300 10055 34309
rect 9747 34298 9753 34300
rect 9809 34298 9833 34300
rect 9889 34298 9913 34300
rect 9969 34298 9993 34300
rect 10049 34298 10055 34300
rect 9809 34246 9811 34298
rect 9991 34246 9993 34298
rect 9747 34244 9753 34246
rect 9809 34244 9833 34246
rect 9889 34244 9913 34246
rect 9969 34244 9993 34246
rect 10049 34244 10055 34246
rect 9747 34235 10055 34244
rect 9456 34156 9536 34184
rect 9404 34138 9456 34144
rect 9324 34054 9628 34082
rect 9312 33992 9364 33998
rect 9312 33934 9364 33940
rect 9496 33992 9548 33998
rect 9496 33934 9548 33940
rect 9324 33658 9352 33934
rect 9312 33652 9364 33658
rect 9312 33594 9364 33600
rect 9232 33510 9352 33538
rect 9220 33040 9272 33046
rect 9220 32982 9272 32988
rect 9128 32020 9180 32026
rect 9128 31962 9180 31968
rect 8864 31726 9076 31754
rect 8760 31476 8812 31482
rect 8760 31418 8812 31424
rect 8576 31340 8628 31346
rect 8576 31282 8628 31288
rect 8588 28744 8616 31282
rect 8760 29640 8812 29646
rect 8760 29582 8812 29588
rect 8668 29164 8720 29170
rect 8668 29106 8720 29112
rect 8680 28966 8708 29106
rect 8668 28960 8720 28966
rect 8668 28902 8720 28908
rect 8772 28762 8800 29582
rect 8760 28756 8812 28762
rect 8588 28716 8708 28744
rect 8574 28656 8630 28665
rect 8574 28591 8630 28600
rect 8588 28014 8616 28591
rect 8576 28008 8628 28014
rect 8576 27950 8628 27956
rect 8576 27600 8628 27606
rect 8576 27542 8628 27548
rect 8482 27160 8538 27169
rect 8392 27124 8444 27130
rect 8482 27095 8538 27104
rect 8392 27066 8444 27072
rect 8392 26920 8444 26926
rect 8392 26862 8444 26868
rect 8300 25288 8352 25294
rect 8300 25230 8352 25236
rect 8404 24070 8432 26862
rect 8482 26752 8538 26761
rect 8482 26687 8538 26696
rect 8496 26314 8524 26687
rect 8484 26308 8536 26314
rect 8484 26250 8536 26256
rect 8588 25158 8616 27542
rect 8680 27334 8708 28716
rect 8760 28698 8812 28704
rect 8760 28076 8812 28082
rect 8760 28018 8812 28024
rect 8772 27878 8800 28018
rect 8760 27872 8812 27878
rect 8760 27814 8812 27820
rect 8668 27328 8720 27334
rect 8668 27270 8720 27276
rect 8760 27124 8812 27130
rect 8760 27066 8812 27072
rect 8668 27056 8720 27062
rect 8668 26998 8720 27004
rect 8680 26926 8708 26998
rect 8668 26920 8720 26926
rect 8668 26862 8720 26868
rect 8680 26625 8708 26862
rect 8666 26616 8722 26625
rect 8666 26551 8722 26560
rect 8576 25152 8628 25158
rect 8576 25094 8628 25100
rect 8680 24954 8708 26551
rect 8668 24948 8720 24954
rect 8668 24890 8720 24896
rect 8772 24857 8800 27066
rect 8758 24848 8814 24857
rect 8668 24812 8720 24818
rect 8758 24783 8814 24792
rect 8668 24754 8720 24760
rect 8392 24064 8444 24070
rect 8392 24006 8444 24012
rect 8484 24064 8536 24070
rect 8484 24006 8536 24012
rect 8404 23866 8432 24006
rect 8392 23860 8444 23866
rect 8392 23802 8444 23808
rect 8208 23792 8260 23798
rect 8206 23760 8208 23769
rect 8260 23760 8262 23769
rect 8206 23695 8262 23704
rect 8390 23760 8446 23769
rect 8390 23695 8392 23704
rect 8444 23695 8446 23704
rect 8392 23666 8444 23672
rect 8392 23316 8444 23322
rect 8392 23258 8444 23264
rect 7746 22607 7802 22616
rect 7852 22630 8156 22658
rect 7748 22228 7800 22234
rect 7748 22170 7800 22176
rect 7760 22030 7788 22170
rect 7748 22024 7800 22030
rect 7748 21966 7800 21972
rect 7746 21856 7802 21865
rect 7746 21791 7802 21800
rect 7760 20466 7788 21791
rect 7852 20942 7880 22630
rect 7932 22568 7984 22574
rect 7932 22510 7984 22516
rect 7944 22012 7972 22510
rect 8208 22500 8260 22506
rect 8208 22442 8260 22448
rect 8024 22024 8076 22030
rect 7944 21984 8024 22012
rect 7944 21690 7972 21984
rect 8220 22012 8248 22442
rect 8404 22094 8432 23258
rect 8496 22778 8524 24006
rect 8680 23254 8708 24754
rect 8760 24744 8812 24750
rect 8760 24686 8812 24692
rect 8772 24041 8800 24686
rect 8758 24032 8814 24041
rect 8758 23967 8814 23976
rect 8668 23248 8720 23254
rect 8668 23190 8720 23196
rect 8484 22772 8536 22778
rect 8484 22714 8536 22720
rect 8576 22432 8628 22438
rect 8576 22374 8628 22380
rect 8668 22432 8720 22438
rect 8668 22374 8720 22380
rect 8404 22066 8524 22094
rect 8024 21966 8076 21972
rect 8128 21984 8248 22012
rect 7932 21684 7984 21690
rect 7932 21626 7984 21632
rect 8128 21570 8156 21984
rect 8036 21554 8156 21570
rect 8024 21548 8156 21554
rect 8076 21542 8156 21548
rect 8024 21490 8076 21496
rect 7840 20936 7892 20942
rect 7840 20878 7892 20884
rect 7748 20460 7800 20466
rect 7748 20402 7800 20408
rect 7656 19848 7708 19854
rect 7656 19790 7708 19796
rect 7484 19638 7696 19666
rect 7668 19514 7696 19638
rect 7656 19508 7708 19514
rect 7378 19442 7434 19451
rect 7656 19450 7708 19456
rect 7378 19377 7434 19386
rect 7472 19440 7524 19446
rect 7472 19382 7524 19388
rect 7288 18964 7340 18970
rect 7288 18906 7340 18912
rect 6656 18686 6776 18714
rect 6458 18456 6514 18465
rect 6458 18391 6514 18400
rect 6552 18420 6604 18426
rect 6472 18290 6500 18391
rect 6552 18362 6604 18368
rect 6368 18284 6420 18290
rect 6368 18226 6420 18232
rect 6460 18284 6512 18290
rect 6460 18226 6512 18232
rect 6274 18184 6330 18193
rect 6274 18119 6330 18128
rect 6288 17882 6316 18119
rect 6276 17876 6328 17882
rect 6276 17818 6328 17824
rect 6368 17196 6420 17202
rect 6368 17138 6420 17144
rect 6184 17060 6236 17066
rect 6184 17002 6236 17008
rect 6092 16992 6144 16998
rect 6092 16934 6144 16940
rect 6196 16658 6224 17002
rect 6092 16652 6144 16658
rect 6092 16594 6144 16600
rect 6184 16652 6236 16658
rect 6184 16594 6236 16600
rect 6104 16114 6132 16594
rect 6276 16584 6328 16590
rect 6276 16526 6328 16532
rect 6184 16448 6236 16454
rect 6184 16390 6236 16396
rect 6092 16108 6144 16114
rect 6092 16050 6144 16056
rect 6090 15872 6146 15881
rect 6090 15807 6146 15816
rect 6104 13394 6132 15807
rect 6092 13388 6144 13394
rect 6092 13330 6144 13336
rect 6104 11218 6132 13330
rect 6196 13190 6224 16390
rect 6288 16046 6316 16526
rect 6380 16114 6408 17138
rect 6458 17096 6514 17105
rect 6564 17082 6592 18362
rect 6642 17368 6698 17377
rect 6642 17303 6698 17312
rect 6656 17270 6684 17303
rect 6644 17264 6696 17270
rect 6644 17206 6696 17212
rect 6514 17054 6592 17082
rect 6458 17031 6514 17040
rect 6748 16658 6776 18686
rect 7288 18624 7340 18630
rect 7288 18566 7340 18572
rect 6814 18524 7122 18533
rect 6814 18522 6820 18524
rect 6876 18522 6900 18524
rect 6956 18522 6980 18524
rect 7036 18522 7060 18524
rect 7116 18522 7122 18524
rect 6876 18470 6878 18522
rect 7058 18470 7060 18522
rect 6814 18468 6820 18470
rect 6876 18468 6900 18470
rect 6956 18468 6980 18470
rect 7036 18468 7060 18470
rect 7116 18468 7122 18470
rect 6814 18459 7122 18468
rect 7196 18284 7248 18290
rect 7196 18226 7248 18232
rect 7208 17882 7236 18226
rect 7196 17876 7248 17882
rect 7196 17818 7248 17824
rect 7196 17672 7248 17678
rect 7196 17614 7248 17620
rect 6814 17436 7122 17445
rect 6814 17434 6820 17436
rect 6876 17434 6900 17436
rect 6956 17434 6980 17436
rect 7036 17434 7060 17436
rect 7116 17434 7122 17436
rect 6876 17382 6878 17434
rect 7058 17382 7060 17434
rect 6814 17380 6820 17382
rect 6876 17380 6900 17382
rect 6956 17380 6980 17382
rect 7036 17380 7060 17382
rect 7116 17380 7122 17382
rect 6814 17371 7122 17380
rect 7104 17264 7156 17270
rect 6826 17232 6882 17241
rect 7104 17206 7156 17212
rect 6826 17167 6882 17176
rect 6736 16652 6788 16658
rect 6736 16594 6788 16600
rect 6552 16448 6604 16454
rect 6840 16436 6868 17167
rect 7116 16998 7144 17206
rect 7208 17066 7236 17614
rect 7300 17338 7328 18566
rect 7392 17678 7420 19377
rect 7380 17672 7432 17678
rect 7380 17614 7432 17620
rect 7288 17332 7340 17338
rect 7288 17274 7340 17280
rect 7286 17232 7342 17241
rect 7286 17167 7342 17176
rect 7196 17060 7248 17066
rect 7196 17002 7248 17008
rect 7104 16992 7156 16998
rect 7104 16934 7156 16940
rect 7116 16590 7144 16934
rect 7104 16584 7156 16590
rect 7104 16526 7156 16532
rect 6552 16390 6604 16396
rect 6748 16408 6868 16436
rect 6458 16280 6514 16289
rect 6564 16266 6592 16390
rect 6514 16238 6592 16266
rect 6458 16215 6514 16224
rect 6368 16108 6420 16114
rect 6368 16050 6420 16056
rect 6276 16040 6328 16046
rect 6276 15982 6328 15988
rect 6380 14482 6408 16050
rect 6368 14476 6420 14482
rect 6368 14418 6420 14424
rect 6380 14006 6408 14418
rect 6368 14000 6420 14006
rect 6368 13942 6420 13948
rect 6184 13184 6236 13190
rect 6184 13126 6236 13132
rect 6184 12980 6236 12986
rect 6184 12922 6236 12928
rect 6092 11212 6144 11218
rect 6092 11154 6144 11160
rect 5998 11112 6054 11121
rect 5998 11047 6054 11056
rect 6092 11008 6144 11014
rect 6092 10950 6144 10956
rect 5920 9438 6040 9466
rect 5908 9376 5960 9382
rect 5908 9318 5960 9324
rect 5920 9178 5948 9318
rect 5908 9172 5960 9178
rect 5908 9114 5960 9120
rect 6012 9058 6040 9438
rect 6104 9178 6132 10950
rect 6196 9450 6224 12922
rect 6380 12850 6408 13942
rect 6472 13870 6500 16215
rect 6748 16096 6776 16408
rect 6814 16348 7122 16357
rect 6814 16346 6820 16348
rect 6876 16346 6900 16348
rect 6956 16346 6980 16348
rect 7036 16346 7060 16348
rect 7116 16346 7122 16348
rect 6876 16294 6878 16346
rect 7058 16294 7060 16346
rect 6814 16292 6820 16294
rect 6876 16292 6900 16294
rect 6956 16292 6980 16294
rect 7036 16292 7060 16294
rect 7116 16292 7122 16294
rect 6814 16283 7122 16292
rect 6828 16108 6880 16114
rect 6748 16068 6828 16096
rect 6828 16050 6880 16056
rect 7300 15586 7328 17167
rect 7380 16992 7432 16998
rect 7380 16934 7432 16940
rect 7392 16794 7420 16934
rect 7380 16788 7432 16794
rect 7380 16730 7432 16736
rect 7378 16584 7430 16590
rect 7484 16561 7512 19382
rect 7562 19348 7618 19357
rect 7562 19283 7618 19292
rect 7576 18766 7604 19283
rect 7760 19009 7788 20402
rect 7932 19916 7984 19922
rect 7932 19858 7984 19864
rect 7840 19780 7892 19786
rect 7840 19722 7892 19728
rect 7852 19514 7880 19722
rect 7944 19514 7972 19858
rect 7840 19508 7892 19514
rect 7840 19450 7892 19456
rect 7932 19508 7984 19514
rect 7932 19450 7984 19456
rect 8036 19394 8064 21490
rect 8208 20936 8260 20942
rect 8208 20878 8260 20884
rect 8116 19780 8168 19786
rect 8116 19722 8168 19728
rect 7852 19366 8064 19394
rect 7746 19000 7802 19009
rect 7746 18935 7802 18944
rect 7564 18760 7616 18766
rect 7564 18702 7616 18708
rect 7564 18420 7616 18426
rect 7564 18362 7616 18368
rect 7378 16526 7430 16532
rect 7470 16552 7526 16561
rect 7392 16250 7420 16526
rect 7470 16487 7526 16496
rect 7380 16244 7432 16250
rect 7380 16186 7432 16192
rect 7208 15558 7328 15586
rect 7208 15502 7236 15558
rect 7196 15496 7248 15502
rect 7196 15438 7248 15444
rect 7288 15496 7340 15502
rect 7288 15438 7340 15444
rect 6814 15260 7122 15269
rect 6814 15258 6820 15260
rect 6876 15258 6900 15260
rect 6956 15258 6980 15260
rect 7036 15258 7060 15260
rect 7116 15258 7122 15260
rect 6876 15206 6878 15258
rect 7058 15206 7060 15258
rect 6814 15204 6820 15206
rect 6876 15204 6900 15206
rect 6956 15204 6980 15206
rect 7036 15204 7060 15206
rect 7116 15204 7122 15206
rect 6814 15195 7122 15204
rect 7196 15156 7248 15162
rect 7196 15098 7248 15104
rect 7104 14952 7156 14958
rect 7104 14894 7156 14900
rect 7116 14618 7144 14894
rect 7104 14612 7156 14618
rect 7104 14554 7156 14560
rect 7208 14346 7236 15098
rect 7196 14340 7248 14346
rect 7196 14282 7248 14288
rect 6814 14172 7122 14181
rect 6814 14170 6820 14172
rect 6876 14170 6900 14172
rect 6956 14170 6980 14172
rect 7036 14170 7060 14172
rect 7116 14170 7122 14172
rect 6876 14118 6878 14170
rect 7058 14118 7060 14170
rect 6814 14116 6820 14118
rect 6876 14116 6900 14118
rect 6956 14116 6980 14118
rect 7036 14116 7060 14118
rect 7116 14116 7122 14118
rect 6814 14107 7122 14116
rect 6552 13932 6604 13938
rect 6552 13874 6604 13880
rect 6460 13864 6512 13870
rect 6460 13806 6512 13812
rect 6368 12844 6420 12850
rect 6368 12786 6420 12792
rect 6276 12776 6328 12782
rect 6276 12718 6328 12724
rect 6184 9444 6236 9450
rect 6184 9386 6236 9392
rect 6092 9172 6144 9178
rect 6092 9114 6144 9120
rect 5920 9030 6040 9058
rect 5920 8974 5948 9030
rect 5908 8968 5960 8974
rect 5908 8910 5960 8916
rect 5920 8294 5948 8910
rect 5998 8528 6054 8537
rect 5998 8463 6000 8472
rect 6052 8463 6054 8472
rect 6000 8434 6052 8440
rect 6184 8424 6236 8430
rect 6184 8366 6236 8372
rect 5908 8288 5960 8294
rect 5908 8230 5960 8236
rect 5920 6866 5948 8230
rect 6092 7880 6144 7886
rect 6092 7822 6144 7828
rect 5908 6860 5960 6866
rect 5908 6802 5960 6808
rect 5920 5166 5948 6802
rect 5908 5160 5960 5166
rect 5908 5102 5960 5108
rect 5920 3602 5948 5102
rect 5908 3596 5960 3602
rect 5908 3538 5960 3544
rect 6104 3482 6132 7822
rect 6196 6254 6224 8366
rect 6288 7206 6316 12718
rect 6564 12345 6592 13874
rect 6736 13864 6788 13870
rect 6736 13806 6788 13812
rect 7196 13864 7248 13870
rect 7196 13806 7248 13812
rect 6748 13326 6776 13806
rect 6736 13320 6788 13326
rect 6736 13262 6788 13268
rect 6748 12986 6776 13262
rect 6814 13084 7122 13093
rect 6814 13082 6820 13084
rect 6876 13082 6900 13084
rect 6956 13082 6980 13084
rect 7036 13082 7060 13084
rect 7116 13082 7122 13084
rect 6876 13030 6878 13082
rect 7058 13030 7060 13082
rect 6814 13028 6820 13030
rect 6876 13028 6900 13030
rect 6956 13028 6980 13030
rect 7036 13028 7060 13030
rect 7116 13028 7122 13030
rect 6814 13019 7122 13028
rect 6736 12980 6788 12986
rect 6736 12922 6788 12928
rect 6736 12844 6788 12850
rect 6736 12786 6788 12792
rect 6550 12336 6606 12345
rect 6550 12271 6606 12280
rect 6368 12096 6420 12102
rect 6368 12038 6420 12044
rect 6460 12096 6512 12102
rect 6460 12038 6512 12044
rect 6644 12096 6696 12102
rect 6644 12038 6696 12044
rect 6380 7410 6408 12038
rect 6472 11218 6500 12038
rect 6656 11830 6684 12038
rect 6748 11898 6776 12786
rect 6814 11996 7122 12005
rect 6814 11994 6820 11996
rect 6876 11994 6900 11996
rect 6956 11994 6980 11996
rect 7036 11994 7060 11996
rect 7116 11994 7122 11996
rect 6876 11942 6878 11994
rect 7058 11942 7060 11994
rect 6814 11940 6820 11942
rect 6876 11940 6900 11942
rect 6956 11940 6980 11942
rect 7036 11940 7060 11942
rect 7116 11940 7122 11942
rect 6814 11931 7122 11940
rect 6736 11892 6788 11898
rect 6736 11834 6788 11840
rect 7104 11892 7156 11898
rect 7104 11834 7156 11840
rect 6644 11824 6696 11830
rect 6644 11766 6696 11772
rect 6828 11824 6880 11830
rect 6828 11766 6880 11772
rect 6840 11665 6868 11766
rect 6826 11656 6882 11665
rect 6826 11591 6882 11600
rect 7116 11218 7144 11834
rect 6460 11212 6512 11218
rect 6460 11154 6512 11160
rect 6644 11212 6696 11218
rect 6644 11154 6696 11160
rect 7104 11212 7156 11218
rect 7104 11154 7156 11160
rect 6550 10704 6606 10713
rect 6550 10639 6606 10648
rect 6460 10056 6512 10062
rect 6460 9998 6512 10004
rect 6472 8974 6500 9998
rect 6564 9654 6592 10639
rect 6552 9648 6604 9654
rect 6552 9590 6604 9596
rect 6460 8968 6512 8974
rect 6460 8910 6512 8916
rect 6552 8968 6604 8974
rect 6656 8956 6684 11154
rect 6814 10908 7122 10917
rect 6814 10906 6820 10908
rect 6876 10906 6900 10908
rect 6956 10906 6980 10908
rect 7036 10906 7060 10908
rect 7116 10906 7122 10908
rect 6876 10854 6878 10906
rect 7058 10854 7060 10906
rect 6814 10852 6820 10854
rect 6876 10852 6900 10854
rect 6956 10852 6980 10854
rect 7036 10852 7060 10854
rect 7116 10852 7122 10854
rect 6814 10843 7122 10852
rect 7104 10668 7156 10674
rect 7104 10610 7156 10616
rect 7012 10532 7064 10538
rect 7012 10474 7064 10480
rect 7024 10130 7052 10474
rect 7116 10130 7144 10610
rect 7012 10124 7064 10130
rect 6932 10084 7012 10112
rect 6932 9976 6960 10084
rect 7012 10066 7064 10072
rect 7104 10124 7156 10130
rect 7104 10066 7156 10072
rect 6748 9948 6960 9976
rect 6748 9518 6776 9948
rect 6814 9820 7122 9829
rect 6814 9818 6820 9820
rect 6876 9818 6900 9820
rect 6956 9818 6980 9820
rect 7036 9818 7060 9820
rect 7116 9818 7122 9820
rect 6876 9766 6878 9818
rect 7058 9766 7060 9818
rect 6814 9764 6820 9766
rect 6876 9764 6900 9766
rect 6956 9764 6980 9766
rect 7036 9764 7060 9766
rect 7116 9764 7122 9766
rect 6814 9755 7122 9764
rect 6736 9512 6788 9518
rect 6736 9454 6788 9460
rect 6604 8928 6684 8956
rect 6552 8910 6604 8916
rect 6368 7404 6420 7410
rect 6368 7346 6420 7352
rect 6276 7200 6328 7206
rect 6276 7142 6328 7148
rect 6276 6860 6328 6866
rect 6276 6802 6328 6808
rect 6288 6458 6316 6802
rect 6472 6780 6500 8910
rect 6656 6866 6684 8928
rect 6736 8968 6788 8974
rect 6736 8910 6788 8916
rect 6748 8634 6776 8910
rect 6814 8732 7122 8741
rect 6814 8730 6820 8732
rect 6876 8730 6900 8732
rect 6956 8730 6980 8732
rect 7036 8730 7060 8732
rect 7116 8730 7122 8732
rect 6876 8678 6878 8730
rect 7058 8678 7060 8730
rect 6814 8676 6820 8678
rect 6876 8676 6900 8678
rect 6956 8676 6980 8678
rect 7036 8676 7060 8678
rect 7116 8676 7122 8678
rect 6814 8667 7122 8676
rect 6736 8628 6788 8634
rect 6736 8570 6788 8576
rect 6736 7744 6788 7750
rect 6736 7686 6788 7692
rect 6644 6860 6696 6866
rect 6644 6802 6696 6808
rect 6552 6792 6604 6798
rect 6472 6752 6552 6780
rect 6552 6734 6604 6740
rect 6276 6452 6328 6458
rect 6276 6394 6328 6400
rect 6184 6248 6236 6254
rect 6184 6190 6236 6196
rect 6196 4196 6224 6190
rect 6368 6180 6420 6186
rect 6368 6122 6420 6128
rect 6380 5710 6408 6122
rect 6460 5908 6512 5914
rect 6460 5850 6512 5856
rect 6368 5704 6420 5710
rect 6368 5646 6420 5652
rect 6276 5568 6328 5574
rect 6276 5510 6328 5516
rect 6288 5302 6316 5510
rect 6276 5296 6328 5302
rect 6276 5238 6328 5244
rect 6380 4826 6408 5646
rect 6368 4820 6420 4826
rect 6368 4762 6420 4768
rect 6276 4208 6328 4214
rect 6196 4168 6276 4196
rect 6276 4150 6328 4156
rect 6472 3602 6500 5850
rect 6564 5370 6592 6734
rect 6552 5364 6604 5370
rect 6552 5306 6604 5312
rect 6748 5234 6776 7686
rect 6814 7644 7122 7653
rect 6814 7642 6820 7644
rect 6876 7642 6900 7644
rect 6956 7642 6980 7644
rect 7036 7642 7060 7644
rect 7116 7642 7122 7644
rect 6876 7590 6878 7642
rect 7058 7590 7060 7642
rect 6814 7588 6820 7590
rect 6876 7588 6900 7590
rect 6956 7588 6980 7590
rect 7036 7588 7060 7590
rect 7116 7588 7122 7590
rect 6814 7579 7122 7588
rect 6814 6556 7122 6565
rect 6814 6554 6820 6556
rect 6876 6554 6900 6556
rect 6956 6554 6980 6556
rect 7036 6554 7060 6556
rect 7116 6554 7122 6556
rect 6876 6502 6878 6554
rect 7058 6502 7060 6554
rect 6814 6500 6820 6502
rect 6876 6500 6900 6502
rect 6956 6500 6980 6502
rect 7036 6500 7060 6502
rect 7116 6500 7122 6502
rect 6814 6491 7122 6500
rect 6814 5468 7122 5477
rect 6814 5466 6820 5468
rect 6876 5466 6900 5468
rect 6956 5466 6980 5468
rect 7036 5466 7060 5468
rect 7116 5466 7122 5468
rect 6876 5414 6878 5466
rect 7058 5414 7060 5466
rect 6814 5412 6820 5414
rect 6876 5412 6900 5414
rect 6956 5412 6980 5414
rect 7036 5412 7060 5414
rect 7116 5412 7122 5414
rect 6814 5403 7122 5412
rect 6736 5228 6788 5234
rect 6736 5170 6788 5176
rect 7104 4820 7156 4826
rect 7104 4762 7156 4768
rect 7116 4622 7144 4762
rect 7104 4616 7156 4622
rect 7104 4558 7156 4564
rect 6814 4380 7122 4389
rect 6814 4378 6820 4380
rect 6876 4378 6900 4380
rect 6956 4378 6980 4380
rect 7036 4378 7060 4380
rect 7116 4378 7122 4380
rect 6876 4326 6878 4378
rect 7058 4326 7060 4378
rect 6814 4324 6820 4326
rect 6876 4324 6900 4326
rect 6956 4324 6980 4326
rect 7036 4324 7060 4326
rect 7116 4324 7122 4326
rect 6814 4315 7122 4324
rect 6644 4140 6696 4146
rect 7208 4128 7236 13806
rect 7300 12345 7328 15438
rect 7470 15056 7526 15065
rect 7470 14991 7472 15000
rect 7524 14991 7526 15000
rect 7472 14962 7524 14968
rect 7576 14498 7604 18362
rect 7748 18148 7800 18154
rect 7748 18090 7800 18096
rect 7656 17536 7708 17542
rect 7656 17478 7708 17484
rect 7668 16046 7696 17478
rect 7656 16040 7708 16046
rect 7656 15982 7708 15988
rect 7484 14470 7604 14498
rect 7484 13938 7512 14470
rect 7564 14408 7616 14414
rect 7564 14350 7616 14356
rect 7472 13932 7524 13938
rect 7472 13874 7524 13880
rect 7472 13796 7524 13802
rect 7472 13738 7524 13744
rect 7380 13388 7432 13394
rect 7380 13330 7432 13336
rect 7286 12336 7342 12345
rect 7286 12271 7342 12280
rect 7392 11898 7420 13330
rect 7484 11898 7512 13738
rect 7380 11892 7432 11898
rect 7380 11834 7432 11840
rect 7472 11892 7524 11898
rect 7472 11834 7524 11840
rect 7380 10600 7432 10606
rect 7380 10542 7432 10548
rect 7288 10056 7340 10062
rect 7288 9998 7340 10004
rect 7300 6934 7328 9998
rect 7392 9722 7420 10542
rect 7472 10532 7524 10538
rect 7472 10474 7524 10480
rect 7380 9716 7432 9722
rect 7380 9658 7432 9664
rect 7392 8906 7420 9658
rect 7380 8900 7432 8906
rect 7380 8842 7432 8848
rect 7392 8430 7420 8842
rect 7380 8424 7432 8430
rect 7380 8366 7432 8372
rect 7392 8090 7420 8366
rect 7380 8084 7432 8090
rect 7380 8026 7432 8032
rect 7484 7562 7512 10474
rect 7576 9586 7604 14350
rect 7760 14074 7788 18090
rect 7656 14068 7708 14074
rect 7656 14010 7708 14016
rect 7748 14068 7800 14074
rect 7748 14010 7800 14016
rect 7668 13530 7696 14010
rect 7748 13796 7800 13802
rect 7748 13738 7800 13744
rect 7656 13524 7708 13530
rect 7656 13466 7708 13472
rect 7656 13388 7708 13394
rect 7656 13330 7708 13336
rect 7668 12850 7696 13330
rect 7760 12986 7788 13738
rect 7748 12980 7800 12986
rect 7748 12922 7800 12928
rect 7656 12844 7708 12850
rect 7656 12786 7708 12792
rect 7564 9580 7616 9586
rect 7564 9522 7616 9528
rect 7576 8498 7604 9522
rect 7668 9382 7696 12786
rect 7852 12434 7880 19366
rect 7932 19236 7984 19242
rect 7932 19178 7984 19184
rect 7944 18290 7972 19178
rect 7932 18284 7984 18290
rect 7932 18226 7984 18232
rect 8024 17672 8076 17678
rect 8024 17614 8076 17620
rect 8128 17626 8156 19722
rect 8220 17814 8248 20878
rect 8390 20768 8446 20777
rect 8390 20703 8446 20712
rect 8300 20596 8352 20602
rect 8300 20538 8352 20544
rect 8312 20398 8340 20538
rect 8300 20392 8352 20398
rect 8300 20334 8352 20340
rect 8300 20256 8352 20262
rect 8300 20198 8352 20204
rect 8312 19786 8340 20198
rect 8300 19780 8352 19786
rect 8300 19722 8352 19728
rect 8300 18624 8352 18630
rect 8300 18566 8352 18572
rect 8208 17808 8260 17814
rect 8208 17750 8260 17756
rect 8036 17202 8064 17614
rect 8128 17598 8248 17626
rect 8116 17536 8168 17542
rect 8116 17478 8168 17484
rect 8024 17196 8076 17202
rect 8024 17138 8076 17144
rect 8036 17105 8064 17138
rect 8128 17134 8156 17478
rect 8116 17128 8168 17134
rect 8022 17096 8078 17105
rect 8116 17070 8168 17076
rect 8022 17031 8078 17040
rect 7932 16992 7984 16998
rect 7932 16934 7984 16940
rect 7944 16794 7972 16934
rect 7932 16788 7984 16794
rect 7932 16730 7984 16736
rect 7944 16114 7972 16730
rect 8022 16688 8078 16697
rect 8022 16623 8024 16632
rect 8076 16623 8078 16632
rect 8024 16594 8076 16600
rect 8114 16552 8170 16561
rect 8114 16487 8170 16496
rect 8024 16448 8076 16454
rect 8024 16390 8076 16396
rect 7932 16108 7984 16114
rect 7932 16050 7984 16056
rect 8036 15502 8064 16390
rect 8024 15496 8076 15502
rect 8024 15438 8076 15444
rect 8024 15156 8076 15162
rect 8024 15098 8076 15104
rect 8036 14414 8064 15098
rect 8024 14408 8076 14414
rect 8024 14350 8076 14356
rect 8024 13864 8076 13870
rect 8022 13832 8024 13841
rect 8076 13832 8078 13841
rect 8022 13767 8078 13776
rect 7760 12406 7880 12434
rect 7656 9376 7708 9382
rect 7656 9318 7708 9324
rect 7668 8974 7696 9318
rect 7656 8968 7708 8974
rect 7656 8910 7708 8916
rect 7656 8628 7708 8634
rect 7656 8570 7708 8576
rect 7668 8537 7696 8570
rect 7654 8528 7710 8537
rect 7564 8492 7616 8498
rect 7654 8463 7710 8472
rect 7564 8434 7616 8440
rect 7656 8288 7708 8294
rect 7656 8230 7708 8236
rect 7668 7993 7696 8230
rect 7654 7984 7710 7993
rect 7654 7919 7710 7928
rect 7668 7886 7696 7919
rect 7656 7880 7708 7886
rect 7656 7822 7708 7828
rect 7380 7540 7432 7546
rect 7484 7534 7604 7562
rect 7380 7482 7432 7488
rect 7392 7002 7420 7482
rect 7472 7472 7524 7478
rect 7472 7414 7524 7420
rect 7484 7002 7512 7414
rect 7576 7410 7604 7534
rect 7564 7404 7616 7410
rect 7564 7346 7616 7352
rect 7562 7304 7618 7313
rect 7668 7290 7696 7822
rect 7618 7262 7696 7290
rect 7562 7239 7618 7248
rect 7564 7200 7616 7206
rect 7564 7142 7616 7148
rect 7380 6996 7432 7002
rect 7380 6938 7432 6944
rect 7472 6996 7524 7002
rect 7472 6938 7524 6944
rect 7288 6928 7340 6934
rect 7288 6870 7340 6876
rect 7380 6860 7432 6866
rect 7380 6802 7432 6808
rect 7392 5914 7420 6802
rect 7472 6316 7524 6322
rect 7472 6258 7524 6264
rect 7380 5908 7432 5914
rect 7380 5850 7432 5856
rect 7484 5778 7512 6258
rect 7472 5772 7524 5778
rect 7472 5714 7524 5720
rect 7288 4616 7340 4622
rect 7288 4558 7340 4564
rect 7300 4185 7328 4558
rect 7380 4480 7432 4486
rect 7380 4422 7432 4428
rect 7472 4480 7524 4486
rect 7472 4422 7524 4428
rect 6644 4082 6696 4088
rect 7024 4100 7236 4128
rect 7286 4176 7342 4185
rect 7286 4111 7342 4120
rect 6368 3596 6420 3602
rect 6368 3538 6420 3544
rect 6460 3596 6512 3602
rect 6460 3538 6512 3544
rect 5920 3454 6132 3482
rect 6274 3496 6330 3505
rect 5920 2854 5948 3454
rect 6274 3431 6330 3440
rect 6288 3126 6316 3431
rect 6380 3194 6408 3538
rect 6368 3188 6420 3194
rect 6368 3130 6420 3136
rect 6276 3120 6328 3126
rect 6276 3062 6328 3068
rect 6472 3040 6500 3538
rect 6552 3392 6604 3398
rect 6552 3334 6604 3340
rect 6380 3012 6500 3040
rect 5908 2848 5960 2854
rect 6380 2825 6408 3012
rect 6460 2916 6512 2922
rect 6460 2858 6512 2864
rect 5908 2790 5960 2796
rect 6366 2816 6422 2825
rect 5920 2514 5948 2790
rect 6366 2751 6422 2760
rect 5908 2508 5960 2514
rect 5908 2450 5960 2456
rect 6184 2440 6236 2446
rect 6236 2417 6316 2428
rect 6236 2408 6330 2417
rect 6236 2400 6274 2408
rect 6184 2382 6236 2388
rect 6274 2343 6330 2352
rect 6368 2372 6420 2378
rect 6368 2314 6420 2320
rect 6000 2304 6052 2310
rect 6000 2246 6052 2252
rect 6012 1358 6040 2246
rect 6092 2100 6144 2106
rect 6092 2042 6144 2048
rect 6104 1562 6132 2042
rect 6092 1556 6144 1562
rect 6092 1498 6144 1504
rect 6276 1488 6328 1494
rect 6276 1430 6328 1436
rect 5816 1352 5868 1358
rect 5816 1294 5868 1300
rect 6000 1352 6052 1358
rect 6000 1294 6052 1300
rect 6092 1352 6144 1358
rect 6092 1294 6144 1300
rect 5908 1284 5960 1290
rect 5908 1226 5960 1232
rect 5552 1006 5672 1034
rect 5448 740 5500 746
rect 5448 682 5500 688
rect 5552 474 5580 1006
rect 5632 944 5684 950
rect 5632 886 5684 892
rect 5540 468 5592 474
rect 5540 410 5592 416
rect 5644 160 5672 886
rect 5724 808 5776 814
rect 5724 750 5776 756
rect 5736 490 5764 750
rect 5920 626 5948 1226
rect 6104 950 6132 1294
rect 6288 1018 6316 1430
rect 6380 1204 6408 2314
rect 6472 2038 6500 2858
rect 6460 2032 6512 2038
rect 6460 1974 6512 1980
rect 6380 1176 6500 1204
rect 6276 1012 6328 1018
rect 6276 954 6328 960
rect 6092 944 6144 950
rect 6092 886 6144 892
rect 5920 598 6224 626
rect 5736 462 5948 490
rect 5920 160 5948 462
rect 6196 160 6224 598
rect 6472 160 6500 1176
rect 5078 54 5304 82
rect 5078 -300 5134 54
rect 5354 -300 5410 160
rect 5630 -300 5686 160
rect 5906 -300 5962 160
rect 6182 -300 6238 160
rect 6458 -300 6514 160
rect 6564 82 6592 3334
rect 6656 3194 6684 4082
rect 6828 3596 6880 3602
rect 7024 3584 7052 4100
rect 6880 3556 7052 3584
rect 6828 3538 6880 3544
rect 6814 3292 7122 3301
rect 6814 3290 6820 3292
rect 6876 3290 6900 3292
rect 6956 3290 6980 3292
rect 7036 3290 7060 3292
rect 7116 3290 7122 3292
rect 6876 3238 6878 3290
rect 7058 3238 7060 3290
rect 6814 3236 6820 3238
rect 6876 3236 6900 3238
rect 6956 3236 6980 3238
rect 7036 3236 7060 3238
rect 7116 3236 7122 3238
rect 6814 3227 7122 3236
rect 7208 3194 7236 4100
rect 7392 4078 7420 4422
rect 7484 4146 7512 4422
rect 7472 4140 7524 4146
rect 7472 4082 7524 4088
rect 7380 4072 7432 4078
rect 7380 4014 7432 4020
rect 7378 3768 7434 3777
rect 7576 3738 7604 7142
rect 7656 6112 7708 6118
rect 7656 6054 7708 6060
rect 7668 5914 7696 6054
rect 7656 5908 7708 5914
rect 7656 5850 7708 5856
rect 7378 3703 7434 3712
rect 7564 3732 7616 3738
rect 7288 3596 7340 3602
rect 7288 3538 7340 3544
rect 6644 3188 6696 3194
rect 6644 3130 6696 3136
rect 7196 3188 7248 3194
rect 7196 3130 7248 3136
rect 7196 3052 7248 3058
rect 7196 2994 7248 3000
rect 6736 2848 6788 2854
rect 6642 2816 6698 2825
rect 6736 2790 6788 2796
rect 7012 2848 7064 2854
rect 7012 2790 7064 2796
rect 6642 2751 6698 2760
rect 6656 2106 6684 2751
rect 6644 2100 6696 2106
rect 6644 2042 6696 2048
rect 6748 2038 6776 2790
rect 7024 2310 7052 2790
rect 7012 2304 7064 2310
rect 7012 2246 7064 2252
rect 6814 2204 7122 2213
rect 6814 2202 6820 2204
rect 6876 2202 6900 2204
rect 6956 2202 6980 2204
rect 7036 2202 7060 2204
rect 7116 2202 7122 2204
rect 6876 2150 6878 2202
rect 7058 2150 7060 2202
rect 6814 2148 6820 2150
rect 6876 2148 6900 2150
rect 6956 2148 6980 2150
rect 7036 2148 7060 2150
rect 7116 2148 7122 2150
rect 6814 2139 7122 2148
rect 6736 2032 6788 2038
rect 6736 1974 6788 1980
rect 6644 1352 6696 1358
rect 6644 1294 6696 1300
rect 6656 746 6684 1294
rect 6814 1116 7122 1125
rect 6814 1114 6820 1116
rect 6876 1114 6900 1116
rect 6956 1114 6980 1116
rect 7036 1114 7060 1116
rect 7116 1114 7122 1116
rect 6876 1062 6878 1114
rect 7058 1062 7060 1114
rect 6814 1060 6820 1062
rect 6876 1060 6900 1062
rect 6956 1060 6980 1062
rect 7036 1060 7060 1062
rect 7116 1060 7122 1062
rect 6814 1051 7122 1060
rect 6644 740 6696 746
rect 6644 682 6696 688
rect 6734 82 6790 160
rect 6564 54 6790 82
rect 6734 -300 6790 54
rect 7010 82 7066 160
rect 7208 82 7236 2994
rect 7300 2650 7328 3538
rect 7392 3233 7420 3703
rect 7564 3674 7616 3680
rect 7656 3392 7708 3398
rect 7656 3334 7708 3340
rect 7378 3224 7434 3233
rect 7378 3159 7434 3168
rect 7472 3052 7524 3058
rect 7472 2994 7524 3000
rect 7380 2984 7432 2990
rect 7380 2926 7432 2932
rect 7288 2644 7340 2650
rect 7288 2586 7340 2592
rect 7286 2272 7342 2281
rect 7286 2207 7342 2216
rect 7300 2106 7328 2207
rect 7288 2100 7340 2106
rect 7288 2042 7340 2048
rect 7392 1170 7420 2926
rect 7484 2774 7512 2994
rect 7484 2746 7604 2774
rect 7470 2544 7526 2553
rect 7470 2479 7526 2488
rect 7484 2310 7512 2479
rect 7472 2304 7524 2310
rect 7472 2246 7524 2252
rect 7472 1216 7524 1222
rect 7300 1142 7420 1170
rect 7470 1184 7472 1193
rect 7524 1184 7526 1193
rect 7300 160 7328 1142
rect 7470 1119 7526 1128
rect 7576 160 7604 2746
rect 7668 2446 7696 3334
rect 7760 3058 7788 12406
rect 7932 11552 7984 11558
rect 7932 11494 7984 11500
rect 7838 11384 7894 11393
rect 7838 11319 7894 11328
rect 7852 11150 7880 11319
rect 7840 11144 7892 11150
rect 7840 11086 7892 11092
rect 7852 8294 7880 11086
rect 7944 10674 7972 11494
rect 7932 10668 7984 10674
rect 7932 10610 7984 10616
rect 7840 8288 7892 8294
rect 7840 8230 7892 8236
rect 7944 7342 7972 10610
rect 8024 10056 8076 10062
rect 8024 9998 8076 10004
rect 8036 9722 8064 9998
rect 8024 9716 8076 9722
rect 8024 9658 8076 9664
rect 7932 7336 7984 7342
rect 7932 7278 7984 7284
rect 7944 6866 7972 7278
rect 7932 6860 7984 6866
rect 7932 6802 7984 6808
rect 7944 4060 7972 6802
rect 8024 5568 8076 5574
rect 8024 5510 8076 5516
rect 8036 5030 8064 5510
rect 8024 5024 8076 5030
rect 8024 4966 8076 4972
rect 8024 4616 8076 4622
rect 8022 4584 8024 4593
rect 8076 4584 8078 4593
rect 8022 4519 8078 4528
rect 8024 4072 8076 4078
rect 7944 4049 8024 4060
rect 7930 4040 8024 4049
rect 7840 4004 7892 4010
rect 7986 4032 8024 4040
rect 8024 4014 8076 4020
rect 7930 3975 7986 3984
rect 7840 3946 7892 3952
rect 7852 3738 7880 3946
rect 7840 3732 7892 3738
rect 7840 3674 7892 3680
rect 7932 3528 7984 3534
rect 7852 3476 7932 3482
rect 7852 3470 7984 3476
rect 7852 3454 7972 3470
rect 7748 3052 7800 3058
rect 7748 2994 7800 3000
rect 7760 2825 7788 2994
rect 7746 2816 7802 2825
rect 7746 2751 7802 2760
rect 7748 2576 7800 2582
rect 7748 2518 7800 2524
rect 7656 2440 7708 2446
rect 7656 2382 7708 2388
rect 7760 2106 7788 2518
rect 7656 2100 7708 2106
rect 7656 2042 7708 2048
rect 7748 2100 7800 2106
rect 7748 2042 7800 2048
rect 7668 2009 7696 2042
rect 7654 2000 7710 2009
rect 7654 1935 7710 1944
rect 7748 1216 7800 1222
rect 7748 1158 7800 1164
rect 7760 513 7788 1158
rect 7746 504 7802 513
rect 7746 439 7802 448
rect 7852 160 7880 3454
rect 7932 3392 7984 3398
rect 7932 3334 7984 3340
rect 7944 1834 7972 3334
rect 8128 2774 8156 16487
rect 8220 15201 8248 17598
rect 8312 17338 8340 18566
rect 8300 17332 8352 17338
rect 8300 17274 8352 17280
rect 8298 16144 8354 16153
rect 8298 16079 8300 16088
rect 8352 16079 8354 16088
rect 8300 16050 8352 16056
rect 8312 15473 8340 16050
rect 8298 15464 8354 15473
rect 8298 15399 8354 15408
rect 8206 15192 8262 15201
rect 8206 15127 8262 15136
rect 8300 14952 8352 14958
rect 8298 14920 8300 14929
rect 8352 14920 8354 14929
rect 8298 14855 8354 14864
rect 8300 14272 8352 14278
rect 8300 14214 8352 14220
rect 8312 13938 8340 14214
rect 8300 13932 8352 13938
rect 8300 13874 8352 13880
rect 8208 13864 8260 13870
rect 8208 13806 8260 13812
rect 8220 11762 8248 13806
rect 8208 11756 8260 11762
rect 8208 11698 8260 11704
rect 8220 9722 8248 11698
rect 8300 11552 8352 11558
rect 8300 11494 8352 11500
rect 8312 11354 8340 11494
rect 8300 11348 8352 11354
rect 8300 11290 8352 11296
rect 8404 11121 8432 20703
rect 8496 15026 8524 22066
rect 8588 21049 8616 22374
rect 8574 21040 8630 21049
rect 8574 20975 8630 20984
rect 8680 20942 8708 22374
rect 8760 22160 8812 22166
rect 8760 22102 8812 22108
rect 8668 20936 8720 20942
rect 8668 20878 8720 20884
rect 8668 20528 8720 20534
rect 8668 20470 8720 20476
rect 8576 20256 8628 20262
rect 8576 20198 8628 20204
rect 8588 20058 8616 20198
rect 8576 20052 8628 20058
rect 8576 19994 8628 20000
rect 8576 18760 8628 18766
rect 8576 18702 8628 18708
rect 8588 18601 8616 18702
rect 8574 18592 8630 18601
rect 8574 18527 8630 18536
rect 8588 17202 8616 18527
rect 8576 17196 8628 17202
rect 8576 17138 8628 17144
rect 8574 15600 8630 15609
rect 8574 15535 8630 15544
rect 8484 15020 8536 15026
rect 8484 14962 8536 14968
rect 8588 13258 8616 15535
rect 8680 13394 8708 20470
rect 8772 20058 8800 22102
rect 8760 20052 8812 20058
rect 8760 19994 8812 20000
rect 8758 19136 8814 19145
rect 8758 19071 8814 19080
rect 8772 18970 8800 19071
rect 8760 18964 8812 18970
rect 8760 18906 8812 18912
rect 8758 18864 8814 18873
rect 8758 18799 8814 18808
rect 8772 14521 8800 18799
rect 8864 17338 8892 31726
rect 9128 31408 9180 31414
rect 9128 31350 9180 31356
rect 9036 31340 9088 31346
rect 9036 31282 9088 31288
rect 9048 31142 9076 31282
rect 9036 31136 9088 31142
rect 9036 31078 9088 31084
rect 9048 29889 9076 31078
rect 9140 30977 9168 31350
rect 9126 30968 9182 30977
rect 9126 30903 9182 30912
rect 9034 29880 9090 29889
rect 9034 29815 9090 29824
rect 9232 29646 9260 32982
rect 9324 32774 9352 33510
rect 9404 33516 9456 33522
rect 9404 33458 9456 33464
rect 9312 32768 9364 32774
rect 9312 32710 9364 32716
rect 9416 32570 9444 33458
rect 9508 33386 9536 33934
rect 9496 33380 9548 33386
rect 9496 33322 9548 33328
rect 9404 32564 9456 32570
rect 9404 32506 9456 32512
rect 9508 32450 9536 33322
rect 9324 32422 9536 32450
rect 9220 29640 9272 29646
rect 9220 29582 9272 29588
rect 8944 29504 8996 29510
rect 8944 29446 8996 29452
rect 8956 29170 8984 29446
rect 8944 29164 8996 29170
rect 8996 29124 9076 29152
rect 8944 29106 8996 29112
rect 8944 28552 8996 28558
rect 8944 28494 8996 28500
rect 8956 25906 8984 28494
rect 9048 28082 9076 29124
rect 9232 28994 9260 29582
rect 9140 28966 9260 28994
rect 9036 28076 9088 28082
rect 9036 28018 9088 28024
rect 9036 27328 9088 27334
rect 9036 27270 9088 27276
rect 9048 26042 9076 27270
rect 9036 26036 9088 26042
rect 9036 25978 9088 25984
rect 8944 25900 8996 25906
rect 8944 25842 8996 25848
rect 8944 25356 8996 25362
rect 8944 25298 8996 25304
rect 8956 23254 8984 25298
rect 9140 24886 9168 28966
rect 9220 28008 9272 28014
rect 9220 27950 9272 27956
rect 9232 26314 9260 27950
rect 9324 26489 9352 32422
rect 9404 32360 9456 32366
rect 9404 32302 9456 32308
rect 9416 28014 9444 32302
rect 9496 31748 9548 31754
rect 9496 31690 9548 31696
rect 9508 31482 9536 31690
rect 9496 31476 9548 31482
rect 9496 31418 9548 31424
rect 9600 31385 9628 34054
rect 10152 33538 10180 35634
rect 10230 35592 10286 35601
rect 10230 35527 10232 35536
rect 10284 35527 10286 35536
rect 10232 35498 10284 35504
rect 10336 34746 10364 42316
rect 10416 42220 10468 42226
rect 10416 42162 10468 42168
rect 10428 41585 10456 42162
rect 10414 41576 10470 41585
rect 10414 41511 10470 41520
rect 10520 40526 10548 43182
rect 10612 42702 10640 44540
rect 10692 44124 10744 44130
rect 10692 44066 10744 44072
rect 10600 42696 10652 42702
rect 10600 42638 10652 42644
rect 10704 42548 10732 44066
rect 10888 43874 10916 44540
rect 10888 43846 11008 43874
rect 10980 43314 11008 43846
rect 11060 43648 11112 43654
rect 11060 43590 11112 43596
rect 10968 43308 11020 43314
rect 10968 43250 11020 43256
rect 10876 43104 10928 43110
rect 10876 43046 10928 43052
rect 10784 42628 10836 42634
rect 10784 42570 10836 42576
rect 10612 42520 10732 42548
rect 10508 40520 10560 40526
rect 10508 40462 10560 40468
rect 10520 40050 10548 40462
rect 10508 40044 10560 40050
rect 10508 39986 10560 39992
rect 10416 39296 10468 39302
rect 10416 39238 10468 39244
rect 10428 39098 10456 39238
rect 10416 39092 10468 39098
rect 10416 39034 10468 39040
rect 10416 38480 10468 38486
rect 10416 38422 10468 38428
rect 10324 34740 10376 34746
rect 10324 34682 10376 34688
rect 10324 34604 10376 34610
rect 10324 34546 10376 34552
rect 10336 34202 10364 34546
rect 10324 34196 10376 34202
rect 10324 34138 10376 34144
rect 10336 34066 10364 34138
rect 10428 34066 10456 38422
rect 10508 37460 10560 37466
rect 10508 37402 10560 37408
rect 10520 37126 10548 37402
rect 10508 37120 10560 37126
rect 10508 37062 10560 37068
rect 10508 36916 10560 36922
rect 10508 36858 10560 36864
rect 10324 34060 10376 34066
rect 10324 34002 10376 34008
rect 10416 34060 10468 34066
rect 10416 34002 10468 34008
rect 10322 33960 10378 33969
rect 10322 33895 10324 33904
rect 10376 33895 10378 33904
rect 10324 33866 10376 33872
rect 9968 33510 10180 33538
rect 9968 33300 9996 33510
rect 10048 33448 10100 33454
rect 10428 33402 10456 34002
rect 10100 33396 10456 33402
rect 10048 33390 10456 33396
rect 10060 33374 10456 33390
rect 9968 33272 10180 33300
rect 9747 33212 10055 33221
rect 9747 33210 9753 33212
rect 9809 33210 9833 33212
rect 9889 33210 9913 33212
rect 9969 33210 9993 33212
rect 10049 33210 10055 33212
rect 9809 33158 9811 33210
rect 9991 33158 9993 33210
rect 9747 33156 9753 33158
rect 9809 33156 9833 33158
rect 9889 33156 9913 33158
rect 9969 33156 9993 33158
rect 10049 33156 10055 33158
rect 9747 33147 10055 33156
rect 9680 32768 9732 32774
rect 9680 32710 9732 32716
rect 9692 32178 9720 32710
rect 9674 32150 9720 32178
rect 9674 32042 9702 32150
rect 9747 32124 10055 32133
rect 9747 32122 9753 32124
rect 9809 32122 9833 32124
rect 9889 32122 9913 32124
rect 9969 32122 9993 32124
rect 10049 32122 10055 32124
rect 9809 32070 9811 32122
rect 9991 32070 9993 32122
rect 9747 32068 9753 32070
rect 9809 32068 9833 32070
rect 9889 32068 9913 32070
rect 9969 32068 9993 32070
rect 10049 32068 10055 32070
rect 9747 32059 10055 32068
rect 9674 32014 9720 32042
rect 9586 31376 9642 31385
rect 9692 31346 9720 32014
rect 9862 31920 9918 31929
rect 9862 31855 9918 31864
rect 9876 31822 9904 31855
rect 9864 31816 9916 31822
rect 9864 31758 9916 31764
rect 10152 31686 10180 33272
rect 10230 32872 10286 32881
rect 10230 32807 10286 32816
rect 10244 31686 10272 32807
rect 10140 31680 10192 31686
rect 10140 31622 10192 31628
rect 10232 31680 10284 31686
rect 10232 31622 10284 31628
rect 9772 31476 9824 31482
rect 9956 31476 10008 31482
rect 9824 31436 9956 31464
rect 9772 31418 9824 31424
rect 10336 31464 10364 33374
rect 10520 31754 10548 36858
rect 10612 36632 10640 42520
rect 10796 41414 10824 42570
rect 10704 41386 10824 41414
rect 10704 39409 10732 41386
rect 10784 39840 10836 39846
rect 10784 39782 10836 39788
rect 10690 39400 10746 39409
rect 10690 39335 10746 39344
rect 10690 39264 10746 39273
rect 10690 39199 10746 39208
rect 10704 39030 10732 39199
rect 10692 39024 10744 39030
rect 10692 38966 10744 38972
rect 10796 38486 10824 39782
rect 10784 38480 10836 38486
rect 10784 38422 10836 38428
rect 10796 37194 10824 38422
rect 10784 37188 10836 37194
rect 10784 37130 10836 37136
rect 10692 36644 10744 36650
rect 10612 36604 10692 36632
rect 10692 36586 10744 36592
rect 10796 36530 10824 37130
rect 9956 31418 10008 31424
rect 10244 31436 10364 31464
rect 10428 31726 10548 31754
rect 10612 36502 10824 36530
rect 9586 31311 9642 31320
rect 9680 31340 9732 31346
rect 9680 31282 9732 31288
rect 9747 31036 10055 31045
rect 9747 31034 9753 31036
rect 9809 31034 9833 31036
rect 9889 31034 9913 31036
rect 9969 31034 9993 31036
rect 10049 31034 10055 31036
rect 9809 30982 9811 31034
rect 9991 30982 9993 31034
rect 9747 30980 9753 30982
rect 9809 30980 9833 30982
rect 9889 30980 9913 30982
rect 9969 30980 9993 30982
rect 10049 30980 10055 30982
rect 9747 30971 10055 30980
rect 10244 30870 10272 31436
rect 10324 31340 10376 31346
rect 10324 31282 10376 31288
rect 10232 30864 10284 30870
rect 10232 30806 10284 30812
rect 10048 30728 10100 30734
rect 10048 30670 10100 30676
rect 9588 30592 9640 30598
rect 9588 30534 9640 30540
rect 9496 28960 9548 28966
rect 9496 28902 9548 28908
rect 9508 28626 9536 28902
rect 9496 28620 9548 28626
rect 9496 28562 9548 28568
rect 9404 28008 9456 28014
rect 9404 27950 9456 27956
rect 9404 27532 9456 27538
rect 9404 27474 9456 27480
rect 9416 26994 9444 27474
rect 9404 26988 9456 26994
rect 9404 26930 9456 26936
rect 9496 26784 9548 26790
rect 9496 26726 9548 26732
rect 9310 26480 9366 26489
rect 9310 26415 9366 26424
rect 9508 26314 9536 26726
rect 9220 26308 9272 26314
rect 9220 26250 9272 26256
rect 9496 26308 9548 26314
rect 9496 26250 9548 26256
rect 9600 26194 9628 30534
rect 10060 30258 10088 30670
rect 10048 30252 10100 30258
rect 10232 30252 10284 30258
rect 10100 30212 10180 30240
rect 10048 30194 10100 30200
rect 9747 29948 10055 29957
rect 9747 29946 9753 29948
rect 9809 29946 9833 29948
rect 9889 29946 9913 29948
rect 9969 29946 9993 29948
rect 10049 29946 10055 29948
rect 9809 29894 9811 29946
rect 9991 29894 9993 29946
rect 9747 29892 9753 29894
rect 9809 29892 9833 29894
rect 9889 29892 9913 29894
rect 9969 29892 9993 29894
rect 10049 29892 10055 29894
rect 9747 29883 10055 29892
rect 9956 29844 10008 29850
rect 9956 29786 10008 29792
rect 9968 28948 9996 29786
rect 10152 29209 10180 30212
rect 10232 30194 10284 30200
rect 10244 29850 10272 30194
rect 10232 29844 10284 29850
rect 10232 29786 10284 29792
rect 10232 29572 10284 29578
rect 10232 29514 10284 29520
rect 10244 29306 10272 29514
rect 10232 29300 10284 29306
rect 10232 29242 10284 29248
rect 10138 29200 10194 29209
rect 10138 29135 10194 29144
rect 10140 29096 10192 29102
rect 10336 29050 10364 31282
rect 10140 29038 10192 29044
rect 10048 28960 10100 28966
rect 9968 28920 10048 28948
rect 10048 28902 10100 28908
rect 9747 28860 10055 28869
rect 9747 28858 9753 28860
rect 9809 28858 9833 28860
rect 9889 28858 9913 28860
rect 9969 28858 9993 28860
rect 10049 28858 10055 28860
rect 9809 28806 9811 28858
rect 9991 28806 9993 28858
rect 9747 28804 9753 28806
rect 9809 28804 9833 28806
rect 9889 28804 9913 28806
rect 9969 28804 9993 28806
rect 10049 28804 10055 28806
rect 9747 28795 10055 28804
rect 10152 28218 10180 29038
rect 10244 29022 10364 29050
rect 10140 28212 10192 28218
rect 10140 28154 10192 28160
rect 10140 27872 10192 27878
rect 10138 27840 10140 27849
rect 10192 27840 10194 27849
rect 9747 27772 10055 27781
rect 10138 27775 10194 27784
rect 9747 27770 9753 27772
rect 9809 27770 9833 27772
rect 9889 27770 9913 27772
rect 9969 27770 9993 27772
rect 10049 27770 10055 27772
rect 9809 27718 9811 27770
rect 9991 27718 9993 27770
rect 9747 27716 9753 27718
rect 9809 27716 9833 27718
rect 9889 27716 9913 27718
rect 9969 27716 9993 27718
rect 10049 27716 10055 27718
rect 9747 27707 10055 27716
rect 10140 27532 10192 27538
rect 10140 27474 10192 27480
rect 9747 26684 10055 26693
rect 9747 26682 9753 26684
rect 9809 26682 9833 26684
rect 9889 26682 9913 26684
rect 9969 26682 9993 26684
rect 10049 26682 10055 26684
rect 9809 26630 9811 26682
rect 9991 26630 9993 26682
rect 9747 26628 9753 26630
rect 9809 26628 9833 26630
rect 9889 26628 9913 26630
rect 9969 26628 9993 26630
rect 10049 26628 10055 26630
rect 9747 26619 10055 26628
rect 9324 26166 9628 26194
rect 9862 26208 9918 26217
rect 9324 25838 9352 26166
rect 9862 26143 9918 26152
rect 9680 26036 9732 26042
rect 9680 25978 9732 25984
rect 9692 25922 9720 25978
rect 9416 25894 9720 25922
rect 9876 25906 9904 26143
rect 9864 25900 9916 25906
rect 9312 25832 9364 25838
rect 9312 25774 9364 25780
rect 9128 24880 9180 24886
rect 9128 24822 9180 24828
rect 9036 24608 9088 24614
rect 9036 24550 9088 24556
rect 9312 24608 9364 24614
rect 9312 24550 9364 24556
rect 9048 24410 9076 24550
rect 9036 24404 9088 24410
rect 9036 24346 9088 24352
rect 9324 24274 9352 24550
rect 9312 24268 9364 24274
rect 9232 24228 9312 24256
rect 9128 24200 9180 24206
rect 9128 24142 9180 24148
rect 9140 23866 9168 24142
rect 9128 23860 9180 23866
rect 9128 23802 9180 23808
rect 8944 23248 8996 23254
rect 8944 23190 8996 23196
rect 9036 22432 9088 22438
rect 9036 22374 9088 22380
rect 8944 20052 8996 20058
rect 8944 19994 8996 20000
rect 8956 17678 8984 19994
rect 9048 18426 9076 22374
rect 9126 19000 9182 19009
rect 9126 18935 9182 18944
rect 9036 18420 9088 18426
rect 9036 18362 9088 18368
rect 9140 17746 9168 18935
rect 9128 17740 9180 17746
rect 9128 17682 9180 17688
rect 8944 17672 8996 17678
rect 8944 17614 8996 17620
rect 8852 17332 8904 17338
rect 8852 17274 8904 17280
rect 8852 17196 8904 17202
rect 8852 17138 8904 17144
rect 8864 16250 8892 17138
rect 8852 16244 8904 16250
rect 8852 16186 8904 16192
rect 8956 14940 8984 17614
rect 9128 17264 9180 17270
rect 9128 17206 9180 17212
rect 9140 16522 9168 17206
rect 9232 17082 9260 24228
rect 9312 24210 9364 24216
rect 9312 23656 9364 23662
rect 9312 23598 9364 23604
rect 9324 22098 9352 23598
rect 9416 23050 9444 25894
rect 9864 25842 9916 25848
rect 9496 25832 9548 25838
rect 9496 25774 9548 25780
rect 9588 25832 9640 25838
rect 9588 25774 9640 25780
rect 9508 23186 9536 25774
rect 9600 24886 9628 25774
rect 9747 25596 10055 25605
rect 9747 25594 9753 25596
rect 9809 25594 9833 25596
rect 9889 25594 9913 25596
rect 9969 25594 9993 25596
rect 10049 25594 10055 25596
rect 9809 25542 9811 25594
rect 9991 25542 9993 25594
rect 9747 25540 9753 25542
rect 9809 25540 9833 25542
rect 9889 25540 9913 25542
rect 9969 25540 9993 25542
rect 10049 25540 10055 25542
rect 9747 25531 10055 25540
rect 9956 25356 10008 25362
rect 9956 25298 10008 25304
rect 9588 24880 9640 24886
rect 9588 24822 9640 24828
rect 9968 24818 9996 25298
rect 9956 24812 10008 24818
rect 9956 24754 10008 24760
rect 9747 24508 10055 24517
rect 9747 24506 9753 24508
rect 9809 24506 9833 24508
rect 9889 24506 9913 24508
rect 9969 24506 9993 24508
rect 10049 24506 10055 24508
rect 9809 24454 9811 24506
rect 9991 24454 9993 24506
rect 9747 24452 9753 24454
rect 9809 24452 9833 24454
rect 9889 24452 9913 24454
rect 9969 24452 9993 24454
rect 10049 24452 10055 24454
rect 9747 24443 10055 24452
rect 9588 24336 9640 24342
rect 9588 24278 9640 24284
rect 9600 23633 9628 24278
rect 9680 24268 9732 24274
rect 9680 24210 9732 24216
rect 9772 24268 9824 24274
rect 9772 24210 9824 24216
rect 9692 23905 9720 24210
rect 9678 23896 9734 23905
rect 9678 23831 9734 23840
rect 9586 23624 9642 23633
rect 9784 23594 9812 24210
rect 9864 23656 9916 23662
rect 10048 23656 10100 23662
rect 9864 23598 9916 23604
rect 10046 23624 10048 23633
rect 10100 23624 10102 23633
rect 9586 23559 9642 23568
rect 9772 23588 9824 23594
rect 9772 23530 9824 23536
rect 9876 23526 9904 23598
rect 10046 23559 10102 23568
rect 9588 23520 9640 23526
rect 9588 23462 9640 23468
rect 9864 23520 9916 23526
rect 9864 23462 9916 23468
rect 9496 23180 9548 23186
rect 9496 23122 9548 23128
rect 9404 23044 9456 23050
rect 9404 22986 9456 22992
rect 9600 22574 9628 23462
rect 9747 23420 10055 23429
rect 9747 23418 9753 23420
rect 9809 23418 9833 23420
rect 9889 23418 9913 23420
rect 9969 23418 9993 23420
rect 10049 23418 10055 23420
rect 9809 23366 9811 23418
rect 9991 23366 9993 23418
rect 9747 23364 9753 23366
rect 9809 23364 9833 23366
rect 9889 23364 9913 23366
rect 9969 23364 9993 23366
rect 10049 23364 10055 23366
rect 9747 23355 10055 23364
rect 9588 22568 9640 22574
rect 9588 22510 9640 22516
rect 9312 22092 9364 22098
rect 9600 22094 9628 22510
rect 9747 22332 10055 22341
rect 9747 22330 9753 22332
rect 9809 22330 9833 22332
rect 9889 22330 9913 22332
rect 9969 22330 9993 22332
rect 10049 22330 10055 22332
rect 9809 22278 9811 22330
rect 9991 22278 9993 22330
rect 9747 22276 9753 22278
rect 9809 22276 9833 22278
rect 9889 22276 9913 22278
rect 9969 22276 9993 22278
rect 10049 22276 10055 22278
rect 9747 22267 10055 22276
rect 9600 22066 9720 22094
rect 9312 22034 9364 22040
rect 9404 22024 9456 22030
rect 9404 21966 9456 21972
rect 9416 21350 9444 21966
rect 9588 21888 9640 21894
rect 9588 21830 9640 21836
rect 9404 21344 9456 21350
rect 9404 21286 9456 21292
rect 9416 20942 9444 21286
rect 9600 21146 9628 21830
rect 9692 21486 9720 22066
rect 9680 21480 9732 21486
rect 9680 21422 9732 21428
rect 9747 21244 10055 21253
rect 9747 21242 9753 21244
rect 9809 21242 9833 21244
rect 9889 21242 9913 21244
rect 9969 21242 9993 21244
rect 10049 21242 10055 21244
rect 9809 21190 9811 21242
rect 9991 21190 9993 21242
rect 9747 21188 9753 21190
rect 9809 21188 9833 21190
rect 9889 21188 9913 21190
rect 9969 21188 9993 21190
rect 10049 21188 10055 21190
rect 9747 21179 10055 21188
rect 10152 21146 10180 27474
rect 10244 25401 10272 29022
rect 10322 28928 10378 28937
rect 10322 28863 10378 28872
rect 10336 26042 10364 28863
rect 10428 27538 10456 31726
rect 10508 30796 10560 30802
rect 10508 30738 10560 30744
rect 10520 29628 10548 30738
rect 10612 30433 10640 36502
rect 10784 36100 10836 36106
rect 10784 36042 10836 36048
rect 10692 35692 10744 35698
rect 10692 35634 10744 35640
rect 10704 35154 10732 35634
rect 10692 35148 10744 35154
rect 10692 35090 10744 35096
rect 10796 34746 10824 36042
rect 10784 34740 10836 34746
rect 10784 34682 10836 34688
rect 10784 34536 10836 34542
rect 10784 34478 10836 34484
rect 10796 34202 10824 34478
rect 10784 34196 10836 34202
rect 10784 34138 10836 34144
rect 10784 33992 10836 33998
rect 10784 33934 10836 33940
rect 10796 33658 10824 33934
rect 10784 33652 10836 33658
rect 10784 33594 10836 33600
rect 10692 33040 10744 33046
rect 10692 32982 10744 32988
rect 10598 30424 10654 30433
rect 10598 30359 10654 30368
rect 10704 29646 10732 32982
rect 10784 31748 10836 31754
rect 10784 31690 10836 31696
rect 10796 30938 10824 31690
rect 10784 30932 10836 30938
rect 10784 30874 10836 30880
rect 10782 30560 10838 30569
rect 10782 30495 10838 30504
rect 10796 30326 10824 30495
rect 10784 30320 10836 30326
rect 10784 30262 10836 30268
rect 10784 30048 10836 30054
rect 10784 29990 10836 29996
rect 10600 29640 10652 29646
rect 10520 29600 10600 29628
rect 10600 29582 10652 29588
rect 10692 29640 10744 29646
rect 10692 29582 10744 29588
rect 10796 29170 10824 29990
rect 10784 29164 10836 29170
rect 10784 29106 10836 29112
rect 10508 29096 10560 29102
rect 10560 29044 10732 29050
rect 10508 29038 10732 29044
rect 10520 29022 10732 29038
rect 10508 28960 10560 28966
rect 10508 28902 10560 28908
rect 10520 28150 10548 28902
rect 10704 28762 10732 29022
rect 10784 28960 10836 28966
rect 10784 28902 10836 28908
rect 10692 28756 10744 28762
rect 10692 28698 10744 28704
rect 10600 28552 10652 28558
rect 10600 28494 10652 28500
rect 10508 28144 10560 28150
rect 10508 28086 10560 28092
rect 10612 27826 10640 28494
rect 10704 28014 10732 28698
rect 10796 28082 10824 28902
rect 10784 28076 10836 28082
rect 10784 28018 10836 28024
rect 10692 28008 10744 28014
rect 10692 27950 10744 27956
rect 10520 27798 10640 27826
rect 10784 27872 10836 27878
rect 10784 27814 10836 27820
rect 10520 27538 10548 27798
rect 10690 27704 10746 27713
rect 10612 27662 10690 27690
rect 10416 27532 10468 27538
rect 10416 27474 10468 27480
rect 10508 27532 10560 27538
rect 10508 27474 10560 27480
rect 10416 27396 10468 27402
rect 10416 27338 10468 27344
rect 10428 26586 10456 27338
rect 10416 26580 10468 26586
rect 10416 26522 10468 26528
rect 10324 26036 10376 26042
rect 10324 25978 10376 25984
rect 10324 25900 10376 25906
rect 10324 25842 10376 25848
rect 10230 25392 10286 25401
rect 10230 25327 10286 25336
rect 10230 24576 10286 24585
rect 10230 24511 10286 24520
rect 10244 24274 10272 24511
rect 10336 24426 10364 25842
rect 10612 24857 10640 27662
rect 10690 27639 10746 27648
rect 10692 26308 10744 26314
rect 10692 26250 10744 26256
rect 10704 26042 10732 26250
rect 10692 26036 10744 26042
rect 10692 25978 10744 25984
rect 10796 25945 10824 27814
rect 10888 26246 10916 43046
rect 10968 41540 11020 41546
rect 10968 41482 11020 41488
rect 10980 40050 11008 41482
rect 11072 41414 11100 43590
rect 11164 43314 11192 44540
rect 11152 43308 11204 43314
rect 11152 43250 11204 43256
rect 11440 42702 11468 44540
rect 11428 42696 11480 42702
rect 11716 42684 11744 44540
rect 11992 43874 12020 44540
rect 11992 43846 12112 43874
rect 12084 43314 12112 43846
rect 12164 43444 12216 43450
rect 12164 43386 12216 43392
rect 12072 43308 12124 43314
rect 12072 43250 12124 43256
rect 11888 43172 11940 43178
rect 11888 43114 11940 43120
rect 11796 43104 11848 43110
rect 11796 43046 11848 43052
rect 11808 42945 11836 43046
rect 11794 42936 11850 42945
rect 11794 42871 11850 42880
rect 11796 42696 11848 42702
rect 11716 42656 11796 42684
rect 11428 42638 11480 42644
rect 11796 42638 11848 42644
rect 11520 42560 11572 42566
rect 11520 42502 11572 42508
rect 11612 42560 11664 42566
rect 11612 42502 11664 42508
rect 11072 41386 11192 41414
rect 10968 40044 11020 40050
rect 10968 39986 11020 39992
rect 10966 39536 11022 39545
rect 10966 39471 11022 39480
rect 10980 39030 11008 39471
rect 10968 39024 11020 39030
rect 10968 38966 11020 38972
rect 10968 38752 11020 38758
rect 10968 38694 11020 38700
rect 10980 38486 11008 38694
rect 10968 38480 11020 38486
rect 10968 38422 11020 38428
rect 10968 37324 11020 37330
rect 10968 37266 11020 37272
rect 10980 36922 11008 37266
rect 10968 36916 11020 36922
rect 10968 36858 11020 36864
rect 10968 36644 11020 36650
rect 10968 36586 11020 36592
rect 10980 31346 11008 36586
rect 10968 31340 11020 31346
rect 10968 31282 11020 31288
rect 10966 31240 11022 31249
rect 10966 31175 11022 31184
rect 11060 31204 11112 31210
rect 10980 30734 11008 31175
rect 11060 31146 11112 31152
rect 10968 30728 11020 30734
rect 11072 30705 11100 31146
rect 10968 30670 11020 30676
rect 11058 30696 11114 30705
rect 11058 30631 11114 30640
rect 11164 30598 11192 41386
rect 11532 39137 11560 42502
rect 11518 39128 11574 39137
rect 11518 39063 11574 39072
rect 11336 37868 11388 37874
rect 11336 37810 11388 37816
rect 11242 36680 11298 36689
rect 11242 36615 11298 36624
rect 11152 30592 11204 30598
rect 11152 30534 11204 30540
rect 11058 30424 11114 30433
rect 11114 30382 11192 30410
rect 11058 30359 11114 30368
rect 10968 30320 11020 30326
rect 10966 30288 10968 30297
rect 11020 30288 11022 30297
rect 10966 30223 11022 30232
rect 10968 30116 11020 30122
rect 10968 30058 11020 30064
rect 10980 26625 11008 30058
rect 11060 30048 11112 30054
rect 11060 29990 11112 29996
rect 11072 29714 11100 29990
rect 11060 29708 11112 29714
rect 11060 29650 11112 29656
rect 11060 29572 11112 29578
rect 11060 29514 11112 29520
rect 11072 28966 11100 29514
rect 11060 28960 11112 28966
rect 11060 28902 11112 28908
rect 11060 28212 11112 28218
rect 11060 28154 11112 28160
rect 11072 27033 11100 28154
rect 11058 27024 11114 27033
rect 11058 26959 11114 26968
rect 10966 26616 11022 26625
rect 10966 26551 11022 26560
rect 10968 26376 11020 26382
rect 10968 26318 11020 26324
rect 10876 26240 10928 26246
rect 10876 26182 10928 26188
rect 10782 25936 10838 25945
rect 10782 25871 10838 25880
rect 10876 25900 10928 25906
rect 10876 25842 10928 25848
rect 10692 25288 10744 25294
rect 10692 25230 10744 25236
rect 10598 24848 10654 24857
rect 10598 24783 10654 24792
rect 10508 24608 10560 24614
rect 10508 24550 10560 24556
rect 10414 24440 10470 24449
rect 10336 24398 10414 24426
rect 10414 24375 10470 24384
rect 10520 24274 10548 24550
rect 10232 24268 10284 24274
rect 10508 24268 10560 24274
rect 10284 24228 10456 24256
rect 10232 24210 10284 24216
rect 10232 23656 10284 23662
rect 10232 23598 10284 23604
rect 10244 23254 10272 23598
rect 10232 23248 10284 23254
rect 10232 23190 10284 23196
rect 10232 23044 10284 23050
rect 10232 22986 10284 22992
rect 9588 21140 9640 21146
rect 9588 21082 9640 21088
rect 10140 21140 10192 21146
rect 10140 21082 10192 21088
rect 9862 21040 9918 21049
rect 9600 20998 9862 21026
rect 9404 20936 9456 20942
rect 9404 20878 9456 20884
rect 9494 20632 9550 20641
rect 9600 20618 9628 20998
rect 9862 20975 9918 20984
rect 9550 20590 9628 20618
rect 9494 20567 9550 20576
rect 9312 19848 9364 19854
rect 9312 19790 9364 19796
rect 9324 19446 9352 19790
rect 9508 19446 9536 20567
rect 10244 20534 10272 22986
rect 10324 21956 10376 21962
rect 10324 21898 10376 21904
rect 10232 20528 10284 20534
rect 10232 20470 10284 20476
rect 10138 20360 10194 20369
rect 10138 20295 10194 20304
rect 9747 20156 10055 20165
rect 9747 20154 9753 20156
rect 9809 20154 9833 20156
rect 9889 20154 9913 20156
rect 9969 20154 9993 20156
rect 10049 20154 10055 20156
rect 9809 20102 9811 20154
rect 9991 20102 9993 20154
rect 9747 20100 9753 20102
rect 9809 20100 9833 20102
rect 9889 20100 9913 20102
rect 9969 20100 9993 20102
rect 10049 20100 10055 20102
rect 9747 20091 10055 20100
rect 9588 19848 9640 19854
rect 9588 19790 9640 19796
rect 9600 19718 9628 19790
rect 10152 19786 10180 20295
rect 10140 19780 10192 19786
rect 10140 19722 10192 19728
rect 9588 19712 9640 19718
rect 9588 19654 9640 19660
rect 9600 19446 9628 19654
rect 9312 19440 9364 19446
rect 9312 19382 9364 19388
rect 9496 19440 9548 19446
rect 9496 19382 9548 19388
rect 9588 19440 9640 19446
rect 9588 19382 9640 19388
rect 9324 18222 9352 19382
rect 9404 19304 9456 19310
rect 9404 19246 9456 19252
rect 9416 18766 9444 19246
rect 9680 19168 9732 19174
rect 9680 19110 9732 19116
rect 9690 19094 9720 19110
rect 9690 18986 9718 19094
rect 9747 19068 10055 19077
rect 9747 19066 9753 19068
rect 9809 19066 9833 19068
rect 9889 19066 9913 19068
rect 9969 19066 9993 19068
rect 10049 19066 10055 19068
rect 9809 19014 9811 19066
rect 9991 19014 9993 19066
rect 9747 19012 9753 19014
rect 9809 19012 9833 19014
rect 9889 19012 9913 19014
rect 9969 19012 9993 19014
rect 10049 19012 10055 19014
rect 9747 19003 10055 19012
rect 9690 18958 9720 18986
rect 9692 18834 9720 18958
rect 9954 18864 10010 18873
rect 9680 18828 9732 18834
rect 9954 18799 10010 18808
rect 9680 18770 9732 18776
rect 9968 18766 9996 18799
rect 9404 18760 9456 18766
rect 9404 18702 9456 18708
rect 9496 18760 9548 18766
rect 9956 18760 10008 18766
rect 9548 18708 9628 18714
rect 9496 18702 9628 18708
rect 9956 18702 10008 18708
rect 9508 18686 9628 18702
rect 9600 18680 9628 18686
rect 10232 18692 10284 18698
rect 9600 18652 9720 18680
rect 9402 18456 9458 18465
rect 9692 18426 9720 18652
rect 10232 18634 10284 18640
rect 10244 18601 10272 18634
rect 10230 18592 10286 18601
rect 10230 18527 10286 18536
rect 9402 18391 9458 18400
rect 9680 18420 9732 18426
rect 9312 18216 9364 18222
rect 9312 18158 9364 18164
rect 9324 17678 9352 18158
rect 9312 17672 9364 17678
rect 9312 17614 9364 17620
rect 9310 17232 9366 17241
rect 9310 17167 9312 17176
rect 9364 17167 9366 17176
rect 9312 17138 9364 17144
rect 9232 17054 9352 17082
rect 9220 16992 9272 16998
rect 9220 16934 9272 16940
rect 9128 16516 9180 16522
rect 9128 16458 9180 16464
rect 9128 15904 9180 15910
rect 9128 15846 9180 15852
rect 9036 14952 9088 14958
rect 8956 14912 9036 14940
rect 9036 14894 9088 14900
rect 8758 14512 8814 14521
rect 8758 14447 8814 14456
rect 8772 14414 8800 14447
rect 8760 14408 8812 14414
rect 8760 14350 8812 14356
rect 9036 13728 9088 13734
rect 9036 13670 9088 13676
rect 8668 13388 8720 13394
rect 8668 13330 8720 13336
rect 8576 13252 8628 13258
rect 8576 13194 8628 13200
rect 8680 12306 8708 13330
rect 8758 13152 8814 13161
rect 8758 13087 8814 13096
rect 8668 12300 8720 12306
rect 8668 12242 8720 12248
rect 8484 11620 8536 11626
rect 8484 11562 8536 11568
rect 8496 11354 8524 11562
rect 8484 11348 8536 11354
rect 8484 11290 8536 11296
rect 8576 11144 8628 11150
rect 8390 11112 8446 11121
rect 8390 11047 8446 11056
rect 8496 11104 8576 11132
rect 8496 10996 8524 11104
rect 8576 11086 8628 11092
rect 8404 10968 8524 10996
rect 8300 10124 8352 10130
rect 8300 10066 8352 10072
rect 8312 9722 8340 10066
rect 8208 9716 8260 9722
rect 8208 9658 8260 9664
rect 8300 9716 8352 9722
rect 8300 9658 8352 9664
rect 8404 8498 8432 10968
rect 8484 10260 8536 10266
rect 8484 10202 8536 10208
rect 8496 9178 8524 10202
rect 8484 9172 8536 9178
rect 8484 9114 8536 9120
rect 8484 9036 8536 9042
rect 8484 8978 8536 8984
rect 8392 8492 8444 8498
rect 8392 8434 8444 8440
rect 8300 7744 8352 7750
rect 8300 7686 8352 7692
rect 8312 7342 8340 7686
rect 8300 7336 8352 7342
rect 8300 7278 8352 7284
rect 8300 5908 8352 5914
rect 8300 5850 8352 5856
rect 8312 5166 8340 5850
rect 8208 5160 8260 5166
rect 8208 5102 8260 5108
rect 8300 5160 8352 5166
rect 8300 5102 8352 5108
rect 8220 3602 8248 5102
rect 8300 4752 8352 4758
rect 8300 4694 8352 4700
rect 8312 4146 8340 4694
rect 8300 4140 8352 4146
rect 8300 4082 8352 4088
rect 8496 4078 8524 8978
rect 8680 8090 8708 12242
rect 8772 12170 8800 13087
rect 9048 12434 9076 13670
rect 8956 12406 9076 12434
rect 8760 12164 8812 12170
rect 8760 12106 8812 12112
rect 8772 11150 8800 12106
rect 8760 11144 8812 11150
rect 8760 11086 8812 11092
rect 8760 10464 8812 10470
rect 8760 10406 8812 10412
rect 8772 10266 8800 10406
rect 8760 10260 8812 10266
rect 8760 10202 8812 10208
rect 8760 10056 8812 10062
rect 8956 10044 8984 12406
rect 9036 11756 9088 11762
rect 9036 11698 9088 11704
rect 9048 11354 9076 11698
rect 9036 11348 9088 11354
rect 9036 11290 9088 11296
rect 8812 10016 8984 10044
rect 8760 9998 8812 10004
rect 8772 8974 8800 9998
rect 9140 9674 9168 15846
rect 9232 10266 9260 16934
rect 9324 13938 9352 17054
rect 9416 16522 9444 18391
rect 9680 18362 9732 18368
rect 9588 18284 9640 18290
rect 9640 18244 10180 18272
rect 9588 18226 9640 18232
rect 9494 18184 9550 18193
rect 9494 18119 9550 18128
rect 9508 16998 9536 18119
rect 9747 17980 10055 17989
rect 9747 17978 9753 17980
rect 9809 17978 9833 17980
rect 9889 17978 9913 17980
rect 9969 17978 9993 17980
rect 10049 17978 10055 17980
rect 9809 17926 9811 17978
rect 9991 17926 9993 17978
rect 9747 17924 9753 17926
rect 9809 17924 9833 17926
rect 9889 17924 9913 17926
rect 9969 17924 9993 17926
rect 10049 17924 10055 17926
rect 9747 17915 10055 17924
rect 9680 17808 9732 17814
rect 9680 17750 9732 17756
rect 9864 17808 9916 17814
rect 9864 17750 9916 17756
rect 9496 16992 9548 16998
rect 9496 16934 9548 16940
rect 9588 16992 9640 16998
rect 9692 16946 9720 17750
rect 9876 17202 9904 17750
rect 10152 17678 10180 18244
rect 10140 17672 10192 17678
rect 10140 17614 10192 17620
rect 9864 17196 9916 17202
rect 9864 17138 9916 17144
rect 10336 17082 10364 21898
rect 10428 21894 10456 24228
rect 10508 24210 10560 24216
rect 10598 23896 10654 23905
rect 10598 23831 10654 23840
rect 10506 23624 10562 23633
rect 10506 23559 10562 23568
rect 10520 22794 10548 23559
rect 10612 22982 10640 23831
rect 10704 23322 10732 25230
rect 10888 24410 10916 25842
rect 10980 25498 11008 26318
rect 10968 25492 11020 25498
rect 10968 25434 11020 25440
rect 10968 25288 11020 25294
rect 10968 25230 11020 25236
rect 10876 24404 10928 24410
rect 10876 24346 10928 24352
rect 10782 24304 10838 24313
rect 10782 24239 10838 24248
rect 10876 24268 10928 24274
rect 10692 23316 10744 23322
rect 10692 23258 10744 23264
rect 10692 23180 10744 23186
rect 10692 23122 10744 23128
rect 10600 22976 10652 22982
rect 10600 22918 10652 22924
rect 10520 22766 10640 22794
rect 10508 22704 10560 22710
rect 10612 22681 10640 22766
rect 10508 22646 10560 22652
rect 10598 22672 10654 22681
rect 10416 21888 10468 21894
rect 10416 21830 10468 21836
rect 10416 21684 10468 21690
rect 10416 21626 10468 21632
rect 10428 21593 10456 21626
rect 10414 21584 10470 21593
rect 10520 21570 10548 22646
rect 10598 22607 10654 22616
rect 10612 22506 10640 22607
rect 10600 22500 10652 22506
rect 10600 22442 10652 22448
rect 10704 21978 10732 23122
rect 10796 22710 10824 24239
rect 10876 24210 10928 24216
rect 10888 23662 10916 24210
rect 10980 23866 11008 25230
rect 11060 24200 11112 24206
rect 11060 24142 11112 24148
rect 10968 23860 11020 23866
rect 10968 23802 11020 23808
rect 10876 23656 10928 23662
rect 10876 23598 10928 23604
rect 11072 23526 11100 24142
rect 11060 23520 11112 23526
rect 11060 23462 11112 23468
rect 10968 23316 11020 23322
rect 10968 23258 11020 23264
rect 10784 22704 10836 22710
rect 10784 22646 10836 22652
rect 10980 22438 11008 23258
rect 10784 22432 10836 22438
rect 10784 22374 10836 22380
rect 10968 22432 11020 22438
rect 10968 22374 11020 22380
rect 10796 22098 10824 22374
rect 10784 22092 10836 22098
rect 10784 22034 10836 22040
rect 10980 22030 11008 22374
rect 11164 22094 11192 30382
rect 11256 30122 11284 36615
rect 11348 35086 11376 37810
rect 11426 37768 11482 37777
rect 11426 37703 11482 37712
rect 11440 37194 11468 37703
rect 11520 37664 11572 37670
rect 11520 37606 11572 37612
rect 11428 37188 11480 37194
rect 11428 37130 11480 37136
rect 11532 36854 11560 37606
rect 11520 36848 11572 36854
rect 11520 36790 11572 36796
rect 11428 36236 11480 36242
rect 11428 36178 11480 36184
rect 11336 35080 11388 35086
rect 11336 35022 11388 35028
rect 11336 34400 11388 34406
rect 11336 34342 11388 34348
rect 11348 33590 11376 34342
rect 11336 33584 11388 33590
rect 11336 33526 11388 33532
rect 11336 32224 11388 32230
rect 11336 32166 11388 32172
rect 11348 31822 11376 32166
rect 11336 31816 11388 31822
rect 11336 31758 11388 31764
rect 11336 30592 11388 30598
rect 11336 30534 11388 30540
rect 11244 30116 11296 30122
rect 11244 30058 11296 30064
rect 11244 29572 11296 29578
rect 11244 29514 11296 29520
rect 11256 29209 11284 29514
rect 11242 29200 11298 29209
rect 11242 29135 11298 29144
rect 11242 28656 11298 28665
rect 11242 28591 11298 28600
rect 11256 28558 11284 28591
rect 11244 28552 11296 28558
rect 11244 28494 11296 28500
rect 11348 27130 11376 30534
rect 11440 30054 11468 36178
rect 11520 35284 11572 35290
rect 11520 35226 11572 35232
rect 11532 30682 11560 35226
rect 11624 30841 11652 42502
rect 11704 38752 11756 38758
rect 11702 38720 11704 38729
rect 11756 38720 11758 38729
rect 11702 38655 11758 38664
rect 11796 36032 11848 36038
rect 11796 35974 11848 35980
rect 11808 35630 11836 35974
rect 11796 35624 11848 35630
rect 11796 35566 11848 35572
rect 11796 35080 11848 35086
rect 11796 35022 11848 35028
rect 11702 34640 11758 34649
rect 11702 34575 11758 34584
rect 11716 33658 11744 34575
rect 11704 33652 11756 33658
rect 11704 33594 11756 33600
rect 11716 32910 11744 33594
rect 11704 32904 11756 32910
rect 11704 32846 11756 32852
rect 11704 32768 11756 32774
rect 11704 32710 11756 32716
rect 11716 32337 11744 32710
rect 11702 32328 11758 32337
rect 11702 32263 11758 32272
rect 11704 31476 11756 31482
rect 11704 31418 11756 31424
rect 11716 31346 11744 31418
rect 11704 31340 11756 31346
rect 11704 31282 11756 31288
rect 11610 30832 11666 30841
rect 11610 30767 11666 30776
rect 11532 30654 11652 30682
rect 11520 30592 11572 30598
rect 11520 30534 11572 30540
rect 11532 30258 11560 30534
rect 11520 30252 11572 30258
rect 11520 30194 11572 30200
rect 11518 30152 11574 30161
rect 11518 30087 11574 30096
rect 11428 30048 11480 30054
rect 11428 29990 11480 29996
rect 11532 29617 11560 30087
rect 11624 29714 11652 30654
rect 11704 30592 11756 30598
rect 11704 30534 11756 30540
rect 11612 29708 11664 29714
rect 11612 29650 11664 29656
rect 11716 29646 11744 30534
rect 11808 29782 11836 35022
rect 11900 33046 11928 43114
rect 11980 43104 12032 43110
rect 11980 43046 12032 43052
rect 11992 33590 12020 43046
rect 12072 42628 12124 42634
rect 12072 42570 12124 42576
rect 12084 39302 12112 42570
rect 12072 39296 12124 39302
rect 12072 39238 12124 39244
rect 12084 38962 12112 39238
rect 12072 38956 12124 38962
rect 12072 38898 12124 38904
rect 12176 37482 12204 43386
rect 12268 43382 12296 44540
rect 12544 43432 12572 44540
rect 12820 43874 12848 44540
rect 13096 44010 13124 44540
rect 13096 43982 13216 44010
rect 12820 43846 13124 43874
rect 12679 43548 12987 43557
rect 12679 43546 12685 43548
rect 12741 43546 12765 43548
rect 12821 43546 12845 43548
rect 12901 43546 12925 43548
rect 12981 43546 12987 43548
rect 12741 43494 12743 43546
rect 12923 43494 12925 43546
rect 12679 43492 12685 43494
rect 12741 43492 12765 43494
rect 12821 43492 12845 43494
rect 12901 43492 12925 43494
rect 12981 43492 12987 43494
rect 12679 43483 12987 43492
rect 12544 43404 12664 43432
rect 12256 43376 12308 43382
rect 12256 43318 12308 43324
rect 12348 43308 12400 43314
rect 12348 43250 12400 43256
rect 12084 37454 12204 37482
rect 11980 33584 12032 33590
rect 11980 33526 12032 33532
rect 11888 33040 11940 33046
rect 11888 32982 11940 32988
rect 12084 31482 12112 37454
rect 12164 37392 12216 37398
rect 12162 37360 12164 37369
rect 12216 37360 12218 37369
rect 12162 37295 12218 37304
rect 12256 34740 12308 34746
rect 12256 34682 12308 34688
rect 12268 34610 12296 34682
rect 12256 34604 12308 34610
rect 12256 34546 12308 34552
rect 12164 34128 12216 34134
rect 12164 34070 12216 34076
rect 12072 31476 12124 31482
rect 12072 31418 12124 31424
rect 12072 31272 12124 31278
rect 11978 31240 12034 31249
rect 11888 31204 11940 31210
rect 12072 31214 12124 31220
rect 11978 31175 12034 31184
rect 11888 31146 11940 31152
rect 11900 30433 11928 31146
rect 11886 30424 11942 30433
rect 11886 30359 11942 30368
rect 11888 30252 11940 30258
rect 11888 30194 11940 30200
rect 11796 29776 11848 29782
rect 11796 29718 11848 29724
rect 11704 29640 11756 29646
rect 11518 29608 11574 29617
rect 11704 29582 11756 29588
rect 11518 29543 11574 29552
rect 11532 29510 11560 29543
rect 11520 29504 11572 29510
rect 11520 29446 11572 29452
rect 11796 29504 11848 29510
rect 11796 29446 11848 29452
rect 11428 28960 11480 28966
rect 11428 28902 11480 28908
rect 11518 28928 11574 28937
rect 11440 28558 11468 28902
rect 11518 28863 11574 28872
rect 11532 28762 11560 28863
rect 11520 28756 11572 28762
rect 11520 28698 11572 28704
rect 11428 28552 11480 28558
rect 11428 28494 11480 28500
rect 11336 27124 11388 27130
rect 11336 27066 11388 27072
rect 11440 26926 11468 28494
rect 11612 28416 11664 28422
rect 11612 28358 11664 28364
rect 11624 28150 11652 28358
rect 11612 28144 11664 28150
rect 11612 28086 11664 28092
rect 11704 28144 11756 28150
rect 11704 28086 11756 28092
rect 11612 28008 11664 28014
rect 11716 27985 11744 28086
rect 11808 28082 11836 29446
rect 11796 28076 11848 28082
rect 11796 28018 11848 28024
rect 11612 27950 11664 27956
rect 11702 27976 11758 27985
rect 11624 27606 11652 27950
rect 11702 27911 11758 27920
rect 11612 27600 11664 27606
rect 11612 27542 11664 27548
rect 11796 27464 11848 27470
rect 11702 27432 11758 27441
rect 11796 27406 11848 27412
rect 11702 27367 11758 27376
rect 11428 26920 11480 26926
rect 11348 26880 11428 26908
rect 11348 25362 11376 26880
rect 11428 26862 11480 26868
rect 11612 26852 11664 26858
rect 11612 26794 11664 26800
rect 11428 26376 11480 26382
rect 11428 26318 11480 26324
rect 11440 26042 11468 26318
rect 11520 26308 11572 26314
rect 11520 26250 11572 26256
rect 11428 26036 11480 26042
rect 11428 25978 11480 25984
rect 11532 25906 11560 26250
rect 11624 26042 11652 26794
rect 11612 26036 11664 26042
rect 11612 25978 11664 25984
rect 11520 25900 11572 25906
rect 11520 25842 11572 25848
rect 11336 25356 11388 25362
rect 11256 25316 11336 25344
rect 11256 23866 11284 25316
rect 11336 25298 11388 25304
rect 11520 25356 11572 25362
rect 11520 25298 11572 25304
rect 11428 24880 11480 24886
rect 11334 24848 11390 24857
rect 11428 24822 11480 24828
rect 11334 24783 11390 24792
rect 11244 23860 11296 23866
rect 11244 23802 11296 23808
rect 11072 22066 11192 22094
rect 10968 22024 11020 22030
rect 10600 21956 10652 21962
rect 10704 21950 10916 21978
rect 10968 21966 11020 21972
rect 10600 21898 10652 21904
rect 10612 21690 10640 21898
rect 10692 21888 10744 21894
rect 10692 21830 10744 21836
rect 10600 21684 10652 21690
rect 10600 21626 10652 21632
rect 10520 21542 10640 21570
rect 10414 21519 10470 21528
rect 10506 19952 10562 19961
rect 10506 19887 10562 19896
rect 10520 19718 10548 19887
rect 10508 19712 10560 19718
rect 10508 19654 10560 19660
rect 10508 18760 10560 18766
rect 10508 18702 10560 18708
rect 10520 17660 10548 18702
rect 10612 18290 10640 21542
rect 10600 18284 10652 18290
rect 10600 18226 10652 18232
rect 10600 17672 10652 17678
rect 10520 17632 10600 17660
rect 10600 17614 10652 17620
rect 10416 17332 10468 17338
rect 10416 17274 10468 17280
rect 9588 16934 9640 16940
rect 9600 16794 9628 16934
rect 9690 16918 9720 16946
rect 10152 17054 10364 17082
rect 9690 16810 9718 16918
rect 9747 16892 10055 16901
rect 9747 16890 9753 16892
rect 9809 16890 9833 16892
rect 9889 16890 9913 16892
rect 9969 16890 9993 16892
rect 10049 16890 10055 16892
rect 9809 16838 9811 16890
rect 9991 16838 9993 16890
rect 9747 16836 9753 16838
rect 9809 16836 9833 16838
rect 9889 16836 9913 16838
rect 9969 16836 9993 16838
rect 10049 16836 10055 16838
rect 9747 16827 10055 16836
rect 9588 16788 9640 16794
rect 9690 16782 9720 16810
rect 9588 16730 9640 16736
rect 9692 16658 9720 16782
rect 10046 16688 10102 16697
rect 9680 16652 9732 16658
rect 10046 16623 10102 16632
rect 9680 16594 9732 16600
rect 10060 16590 10088 16623
rect 10048 16584 10100 16590
rect 10048 16526 10100 16532
rect 9404 16516 9456 16522
rect 9404 16458 9456 16464
rect 9496 16448 9548 16454
rect 9496 16390 9548 16396
rect 9508 16114 9536 16390
rect 10152 16130 10180 17054
rect 10232 16992 10284 16998
rect 10232 16934 10284 16940
rect 9496 16108 9548 16114
rect 9496 16050 9548 16056
rect 10060 16102 10180 16130
rect 10060 16046 10088 16102
rect 9588 16040 9640 16046
rect 9588 15982 9640 15988
rect 10048 16040 10100 16046
rect 10048 15982 10100 15988
rect 10140 16040 10192 16046
rect 10244 16028 10272 16934
rect 10322 16824 10378 16833
rect 10322 16759 10378 16768
rect 10192 16000 10272 16028
rect 10140 15982 10192 15988
rect 9600 15638 9628 15982
rect 10060 15892 10088 15982
rect 10060 15864 10180 15892
rect 9747 15804 10055 15813
rect 9747 15802 9753 15804
rect 9809 15802 9833 15804
rect 9889 15802 9913 15804
rect 9969 15802 9993 15804
rect 10049 15802 10055 15804
rect 9809 15750 9811 15802
rect 9991 15750 9993 15802
rect 9747 15748 9753 15750
rect 9809 15748 9833 15750
rect 9889 15748 9913 15750
rect 9969 15748 9993 15750
rect 10049 15748 10055 15750
rect 9747 15739 10055 15748
rect 9588 15632 9640 15638
rect 9588 15574 9640 15580
rect 10152 15502 10180 15864
rect 9404 15496 9456 15502
rect 9404 15438 9456 15444
rect 10140 15496 10192 15502
rect 10140 15438 10192 15444
rect 9416 15026 9444 15438
rect 9404 15020 9456 15026
rect 9404 14962 9456 14968
rect 10232 14952 10284 14958
rect 10232 14894 10284 14900
rect 10140 14884 10192 14890
rect 10140 14826 10192 14832
rect 9747 14716 10055 14725
rect 9747 14714 9753 14716
rect 9809 14714 9833 14716
rect 9889 14714 9913 14716
rect 9969 14714 9993 14716
rect 10049 14714 10055 14716
rect 9809 14662 9811 14714
rect 9991 14662 9993 14714
rect 9747 14660 9753 14662
rect 9809 14660 9833 14662
rect 9889 14660 9913 14662
rect 9969 14660 9993 14662
rect 10049 14660 10055 14662
rect 9747 14651 10055 14660
rect 10152 14618 10180 14826
rect 10140 14612 10192 14618
rect 10140 14554 10192 14560
rect 9312 13932 9364 13938
rect 9312 13874 9364 13880
rect 9747 13628 10055 13637
rect 9747 13626 9753 13628
rect 9809 13626 9833 13628
rect 9889 13626 9913 13628
rect 9969 13626 9993 13628
rect 10049 13626 10055 13628
rect 9809 13574 9811 13626
rect 9991 13574 9993 13626
rect 9747 13572 9753 13574
rect 9809 13572 9833 13574
rect 9889 13572 9913 13574
rect 9969 13572 9993 13574
rect 10049 13572 10055 13574
rect 9747 13563 10055 13572
rect 10244 13326 10272 14894
rect 10336 14385 10364 16759
rect 10322 14376 10378 14385
rect 10322 14311 10378 14320
rect 10232 13320 10284 13326
rect 10284 13280 10364 13308
rect 10232 13262 10284 13268
rect 9956 13184 10008 13190
rect 9956 13126 10008 13132
rect 9496 12912 9548 12918
rect 9494 12880 9496 12889
rect 9548 12880 9550 12889
rect 9494 12815 9550 12824
rect 9508 12434 9536 12815
rect 9968 12782 9996 13126
rect 10140 12844 10192 12850
rect 10140 12786 10192 12792
rect 9956 12776 10008 12782
rect 9956 12718 10008 12724
rect 9747 12540 10055 12549
rect 9747 12538 9753 12540
rect 9809 12538 9833 12540
rect 9889 12538 9913 12540
rect 9969 12538 9993 12540
rect 10049 12538 10055 12540
rect 9809 12486 9811 12538
rect 9991 12486 9993 12538
rect 9747 12484 9753 12486
rect 9809 12484 9833 12486
rect 9889 12484 9913 12486
rect 9969 12484 9993 12486
rect 10049 12484 10055 12486
rect 9747 12475 10055 12484
rect 9324 12406 9536 12434
rect 10048 12436 10100 12442
rect 9220 10260 9272 10266
rect 9220 10202 9272 10208
rect 9324 10112 9352 12406
rect 10152 12424 10180 12786
rect 10100 12396 10180 12424
rect 10048 12378 10100 12384
rect 9588 11688 9640 11694
rect 9588 11630 9640 11636
rect 9496 11552 9548 11558
rect 9496 11494 9548 11500
rect 9048 9646 9168 9674
rect 9232 10084 9352 10112
rect 9232 9654 9260 10084
rect 9508 10010 9536 11494
rect 9324 9982 9536 10010
rect 9220 9648 9272 9654
rect 8760 8968 8812 8974
rect 8760 8910 8812 8916
rect 8668 8084 8720 8090
rect 8668 8026 8720 8032
rect 8772 7886 8800 8910
rect 8852 8492 8904 8498
rect 8852 8434 8904 8440
rect 8760 7880 8812 7886
rect 8760 7822 8812 7828
rect 8668 7744 8720 7750
rect 8668 7686 8720 7692
rect 8680 7410 8708 7686
rect 8668 7404 8720 7410
rect 8668 7346 8720 7352
rect 8680 5778 8708 7346
rect 8772 5914 8800 7822
rect 8864 6236 8892 8434
rect 8944 8288 8996 8294
rect 8944 8230 8996 8236
rect 8956 7410 8984 8230
rect 8944 7404 8996 7410
rect 8944 7346 8996 7352
rect 8944 6248 8996 6254
rect 8864 6208 8944 6236
rect 8944 6190 8996 6196
rect 8852 6112 8904 6118
rect 8852 6054 8904 6060
rect 8760 5908 8812 5914
rect 8760 5850 8812 5856
rect 8668 5772 8720 5778
rect 8668 5714 8720 5720
rect 8576 5568 8628 5574
rect 8576 5510 8628 5516
rect 8588 5370 8616 5510
rect 8576 5364 8628 5370
rect 8576 5306 8628 5312
rect 8588 5234 8616 5306
rect 8576 5228 8628 5234
rect 8576 5170 8628 5176
rect 8668 5160 8720 5166
rect 8668 5102 8720 5108
rect 8680 4758 8708 5102
rect 8668 4752 8720 4758
rect 8668 4694 8720 4700
rect 8484 4072 8536 4078
rect 8484 4014 8536 4020
rect 8208 3596 8260 3602
rect 8208 3538 8260 3544
rect 8220 3505 8248 3538
rect 8206 3496 8262 3505
rect 8206 3431 8262 3440
rect 8576 3392 8628 3398
rect 8576 3334 8628 3340
rect 8588 2774 8616 3334
rect 8772 2990 8800 5850
rect 8864 5234 8892 6054
rect 8956 5273 8984 6190
rect 8942 5264 8998 5273
rect 8852 5228 8904 5234
rect 8942 5199 8998 5208
rect 8852 5170 8904 5176
rect 8944 4548 8996 4554
rect 8944 4490 8996 4496
rect 8956 4282 8984 4490
rect 8944 4276 8996 4282
rect 8944 4218 8996 4224
rect 8944 4140 8996 4146
rect 8864 4100 8944 4128
rect 8864 3097 8892 4100
rect 8944 4082 8996 4088
rect 8944 3596 8996 3602
rect 8944 3538 8996 3544
rect 8956 3194 8984 3538
rect 8944 3188 8996 3194
rect 8944 3130 8996 3136
rect 8850 3088 8906 3097
rect 8850 3023 8852 3032
rect 8904 3023 8906 3032
rect 8852 2994 8904 3000
rect 8760 2984 8812 2990
rect 8760 2926 8812 2932
rect 8668 2916 8720 2922
rect 8668 2858 8720 2864
rect 8036 2746 8156 2774
rect 8404 2746 8616 2774
rect 8036 1970 8064 2746
rect 8300 2440 8352 2446
rect 8220 2400 8300 2428
rect 8114 2272 8170 2281
rect 8114 2207 8170 2216
rect 8128 2106 8156 2207
rect 8116 2100 8168 2106
rect 8116 2042 8168 2048
rect 8024 1964 8076 1970
rect 8024 1906 8076 1912
rect 7932 1828 7984 1834
rect 7932 1770 7984 1776
rect 7932 1352 7984 1358
rect 7930 1320 7932 1329
rect 7984 1320 7986 1329
rect 7930 1255 7986 1264
rect 8116 1216 8168 1222
rect 8116 1158 8168 1164
rect 8128 882 8156 1158
rect 8116 876 8168 882
rect 8116 818 8168 824
rect 7010 54 7236 82
rect 7010 -300 7066 54
rect 7286 -300 7342 160
rect 7562 -300 7618 160
rect 7838 -300 7894 160
rect 8114 82 8170 160
rect 8220 82 8248 2400
rect 8300 2382 8352 2388
rect 8404 1970 8432 2746
rect 8680 2666 8708 2858
rect 8680 2638 8984 2666
rect 8668 2440 8720 2446
rect 8588 2400 8668 2428
rect 8484 2304 8536 2310
rect 8484 2246 8536 2252
rect 8496 1970 8524 2246
rect 8392 1964 8444 1970
rect 8392 1906 8444 1912
rect 8484 1964 8536 1970
rect 8484 1906 8536 1912
rect 8390 1864 8446 1873
rect 8390 1799 8392 1808
rect 8444 1799 8446 1808
rect 8484 1828 8536 1834
rect 8392 1770 8444 1776
rect 8484 1770 8536 1776
rect 8496 1562 8524 1770
rect 8484 1556 8536 1562
rect 8484 1498 8536 1504
rect 8588 1204 8616 2400
rect 8668 2382 8720 2388
rect 8760 2372 8812 2378
rect 8760 2314 8812 2320
rect 8772 1204 8800 2314
rect 8850 2272 8906 2281
rect 8850 2207 8906 2216
rect 8864 2106 8892 2207
rect 8852 2100 8904 2106
rect 8852 2042 8904 2048
rect 8404 1176 8616 1204
rect 8680 1176 8800 1204
rect 8404 160 8432 1176
rect 8680 160 8708 1176
rect 8956 814 8984 2638
rect 9048 1358 9076 9646
rect 9220 9590 9272 9596
rect 9324 7750 9352 9982
rect 9496 9920 9548 9926
rect 9496 9862 9548 9868
rect 9404 9648 9456 9654
rect 9404 9590 9456 9596
rect 9416 7750 9444 9590
rect 9508 9518 9536 9862
rect 9496 9512 9548 9518
rect 9496 9454 9548 9460
rect 9312 7744 9364 7750
rect 9312 7686 9364 7692
rect 9404 7744 9456 7750
rect 9404 7686 9456 7692
rect 9600 7478 9628 11630
rect 9747 11452 10055 11461
rect 9747 11450 9753 11452
rect 9809 11450 9833 11452
rect 9889 11450 9913 11452
rect 9969 11450 9993 11452
rect 10049 11450 10055 11452
rect 9809 11398 9811 11450
rect 9991 11398 9993 11450
rect 9747 11396 9753 11398
rect 9809 11396 9833 11398
rect 9889 11396 9913 11398
rect 9969 11396 9993 11398
rect 10049 11396 10055 11398
rect 9747 11387 10055 11396
rect 10232 11212 10284 11218
rect 10232 11154 10284 11160
rect 10140 11144 10192 11150
rect 10140 11086 10192 11092
rect 9747 10364 10055 10373
rect 9747 10362 9753 10364
rect 9809 10362 9833 10364
rect 9889 10362 9913 10364
rect 9969 10362 9993 10364
rect 10049 10362 10055 10364
rect 9809 10310 9811 10362
rect 9991 10310 9993 10362
rect 9747 10308 9753 10310
rect 9809 10308 9833 10310
rect 9889 10308 9913 10310
rect 9969 10308 9993 10310
rect 10049 10308 10055 10310
rect 9747 10299 10055 10308
rect 10152 9586 10180 11086
rect 10244 9586 10272 11154
rect 10336 10674 10364 13280
rect 10324 10668 10376 10674
rect 10324 10610 10376 10616
rect 10324 9648 10376 9654
rect 10324 9590 10376 9596
rect 10140 9580 10192 9586
rect 10140 9522 10192 9528
rect 10232 9580 10284 9586
rect 10232 9522 10284 9528
rect 9747 9276 10055 9285
rect 9747 9274 9753 9276
rect 9809 9274 9833 9276
rect 9889 9274 9913 9276
rect 9969 9274 9993 9276
rect 10049 9274 10055 9276
rect 9809 9222 9811 9274
rect 9991 9222 9993 9274
rect 9747 9220 9753 9222
rect 9809 9220 9833 9222
rect 9889 9220 9913 9222
rect 9969 9220 9993 9222
rect 10049 9220 10055 9222
rect 9747 9211 10055 9220
rect 10048 9172 10100 9178
rect 10048 9114 10100 9120
rect 10060 8566 10088 9114
rect 10048 8560 10100 8566
rect 10048 8502 10100 8508
rect 9747 8188 10055 8197
rect 9747 8186 9753 8188
rect 9809 8186 9833 8188
rect 9889 8186 9913 8188
rect 9969 8186 9993 8188
rect 10049 8186 10055 8188
rect 9809 8134 9811 8186
rect 9991 8134 9993 8186
rect 9747 8132 9753 8134
rect 9809 8132 9833 8134
rect 9889 8132 9913 8134
rect 9969 8132 9993 8134
rect 10049 8132 10055 8134
rect 9747 8123 10055 8132
rect 9770 7984 9826 7993
rect 9826 7954 9904 7970
rect 9826 7948 9916 7954
rect 9826 7942 9864 7948
rect 9770 7919 9826 7928
rect 9864 7890 9916 7896
rect 9680 7744 9732 7750
rect 9680 7686 9732 7692
rect 10048 7744 10100 7750
rect 10048 7686 10100 7692
rect 9692 7478 9720 7686
rect 9588 7472 9640 7478
rect 9588 7414 9640 7420
rect 9680 7472 9732 7478
rect 9680 7414 9732 7420
rect 9692 7154 9720 7414
rect 10060 7342 10088 7686
rect 10152 7410 10180 9522
rect 10244 7698 10272 9522
rect 10336 9178 10364 9590
rect 10324 9172 10376 9178
rect 10324 9114 10376 9120
rect 10324 8832 10376 8838
rect 10324 8774 10376 8780
rect 10336 7818 10364 8774
rect 10324 7812 10376 7818
rect 10324 7754 10376 7760
rect 10244 7670 10364 7698
rect 10336 7410 10364 7670
rect 10140 7404 10192 7410
rect 10140 7346 10192 7352
rect 10232 7404 10284 7410
rect 10232 7346 10284 7352
rect 10324 7404 10376 7410
rect 10324 7346 10376 7352
rect 10048 7336 10100 7342
rect 10048 7278 10100 7284
rect 9600 7126 9720 7154
rect 9496 6928 9548 6934
rect 9496 6870 9548 6876
rect 9312 6792 9364 6798
rect 9312 6734 9364 6740
rect 9220 6724 9272 6730
rect 9220 6666 9272 6672
rect 9126 6352 9182 6361
rect 9126 6287 9128 6296
rect 9180 6287 9182 6296
rect 9128 6258 9180 6264
rect 9126 6216 9182 6225
rect 9126 6151 9182 6160
rect 9140 6118 9168 6151
rect 9128 6112 9180 6118
rect 9128 6054 9180 6060
rect 9128 5364 9180 5370
rect 9128 5306 9180 5312
rect 9140 3738 9168 5306
rect 9128 3732 9180 3738
rect 9128 3674 9180 3680
rect 9140 3398 9168 3674
rect 9128 3392 9180 3398
rect 9128 3334 9180 3340
rect 9232 2774 9260 6666
rect 9324 6322 9352 6734
rect 9312 6316 9364 6322
rect 9312 6258 9364 6264
rect 9324 5914 9352 6258
rect 9312 5908 9364 5914
rect 9312 5850 9364 5856
rect 9312 5704 9364 5710
rect 9312 5646 9364 5652
rect 9324 4622 9352 5646
rect 9404 5568 9456 5574
rect 9404 5510 9456 5516
rect 9416 5302 9444 5510
rect 9404 5296 9456 5302
rect 9404 5238 9456 5244
rect 9508 5234 9536 6870
rect 9600 5930 9628 7126
rect 9747 7100 10055 7109
rect 9747 7098 9753 7100
rect 9809 7098 9833 7100
rect 9889 7098 9913 7100
rect 9969 7098 9993 7100
rect 10049 7098 10055 7100
rect 9809 7046 9811 7098
rect 9991 7046 9993 7098
rect 9747 7044 9753 7046
rect 9809 7044 9833 7046
rect 9889 7044 9913 7046
rect 9969 7044 9993 7046
rect 10049 7044 10055 7046
rect 9747 7035 10055 7044
rect 9772 6860 9824 6866
rect 9772 6802 9824 6808
rect 9678 6760 9734 6769
rect 9678 6695 9734 6704
rect 9692 6390 9720 6695
rect 9784 6390 9812 6802
rect 10048 6792 10100 6798
rect 10048 6734 10100 6740
rect 10060 6458 10088 6734
rect 10048 6452 10100 6458
rect 10048 6394 10100 6400
rect 9680 6384 9732 6390
rect 9680 6326 9732 6332
rect 9772 6384 9824 6390
rect 9772 6326 9824 6332
rect 9747 6012 10055 6021
rect 9747 6010 9753 6012
rect 9809 6010 9833 6012
rect 9889 6010 9913 6012
rect 9969 6010 9993 6012
rect 10049 6010 10055 6012
rect 9809 5958 9811 6010
rect 9991 5958 9993 6010
rect 9747 5956 9753 5958
rect 9809 5956 9833 5958
rect 9889 5956 9913 5958
rect 9969 5956 9993 5958
rect 10049 5956 10055 5958
rect 9747 5947 10055 5956
rect 9600 5902 9720 5930
rect 9692 5370 9720 5902
rect 10152 5794 10180 7346
rect 10244 7002 10272 7346
rect 10232 6996 10284 7002
rect 10232 6938 10284 6944
rect 10232 6724 10284 6730
rect 10232 6666 10284 6672
rect 10244 6633 10272 6666
rect 10230 6624 10286 6633
rect 10230 6559 10286 6568
rect 9968 5766 10180 5794
rect 9680 5364 9732 5370
rect 9680 5306 9732 5312
rect 9968 5234 9996 5766
rect 10140 5568 10192 5574
rect 10140 5510 10192 5516
rect 10152 5234 10180 5510
rect 10336 5370 10364 7346
rect 10428 6440 10456 17274
rect 10612 17134 10640 17614
rect 10600 17128 10652 17134
rect 10600 17070 10652 17076
rect 10554 16040 10606 16046
rect 10704 16028 10732 21830
rect 10784 21140 10836 21146
rect 10784 21082 10836 21088
rect 10606 16000 10732 16028
rect 10554 15982 10606 15988
rect 10508 15496 10560 15502
rect 10508 15438 10560 15444
rect 10520 13433 10548 15438
rect 10600 14816 10652 14822
rect 10600 14758 10652 14764
rect 10506 13424 10562 13433
rect 10506 13359 10562 13368
rect 10508 13320 10560 13326
rect 10508 13262 10560 13268
rect 10520 12918 10548 13262
rect 10612 13002 10640 14758
rect 10704 13841 10732 16000
rect 10796 15586 10824 21082
rect 10888 16833 10916 21950
rect 10968 21548 11020 21554
rect 10968 21490 11020 21496
rect 10980 21457 11008 21490
rect 10966 21448 11022 21457
rect 10966 21383 11022 21392
rect 10968 20868 11020 20874
rect 10968 20810 11020 20816
rect 10980 19174 11008 20810
rect 10968 19168 11020 19174
rect 10968 19110 11020 19116
rect 10968 18420 11020 18426
rect 10968 18362 11020 18368
rect 10874 16824 10930 16833
rect 10874 16759 10930 16768
rect 10876 16720 10928 16726
rect 10876 16662 10928 16668
rect 10888 16046 10916 16662
rect 10876 16040 10928 16046
rect 10876 15982 10928 15988
rect 10796 15558 10916 15586
rect 10888 14482 10916 15558
rect 10876 14476 10928 14482
rect 10876 14418 10928 14424
rect 10690 13832 10746 13841
rect 10690 13767 10746 13776
rect 10704 13240 10732 13767
rect 10876 13728 10928 13734
rect 10876 13670 10928 13676
rect 10888 13394 10916 13670
rect 10876 13388 10928 13394
rect 10876 13330 10928 13336
rect 10704 13212 10916 13240
rect 10782 13152 10838 13161
rect 10782 13087 10838 13096
rect 10612 12974 10732 13002
rect 10508 12912 10560 12918
rect 10508 12854 10560 12860
rect 10600 12912 10652 12918
rect 10600 12854 10652 12860
rect 10508 9988 10560 9994
rect 10508 9930 10560 9936
rect 10520 9110 10548 9930
rect 10612 9654 10640 12854
rect 10704 11354 10732 12974
rect 10796 12782 10824 13087
rect 10784 12776 10836 12782
rect 10784 12718 10836 12724
rect 10692 11348 10744 11354
rect 10692 11290 10744 11296
rect 10600 9648 10652 9654
rect 10652 9608 10824 9636
rect 10600 9590 10652 9596
rect 10692 9376 10744 9382
rect 10692 9318 10744 9324
rect 10508 9104 10560 9110
rect 10508 9046 10560 9052
rect 10600 8492 10652 8498
rect 10600 8434 10652 8440
rect 10612 7886 10640 8434
rect 10600 7880 10652 7886
rect 10600 7822 10652 7828
rect 10600 6792 10652 6798
rect 10600 6734 10652 6740
rect 10428 6412 10548 6440
rect 10324 5364 10376 5370
rect 10324 5306 10376 5312
rect 9496 5228 9548 5234
rect 9496 5170 9548 5176
rect 9680 5228 9732 5234
rect 9680 5170 9732 5176
rect 9956 5228 10008 5234
rect 9956 5170 10008 5176
rect 10140 5228 10192 5234
rect 10140 5170 10192 5176
rect 9404 5024 9456 5030
rect 9692 4978 9720 5170
rect 10232 5160 10284 5166
rect 10232 5102 10284 5108
rect 9404 4966 9456 4972
rect 9312 4616 9364 4622
rect 9312 4558 9364 4564
rect 9324 4010 9352 4558
rect 9312 4004 9364 4010
rect 9312 3946 9364 3952
rect 9416 3126 9444 4966
rect 9600 4950 9720 4978
rect 9600 4842 9628 4950
rect 9747 4924 10055 4933
rect 9747 4922 9753 4924
rect 9809 4922 9833 4924
rect 9889 4922 9913 4924
rect 9969 4922 9993 4924
rect 10049 4922 10055 4924
rect 9809 4870 9811 4922
rect 9991 4870 9993 4922
rect 9747 4868 9753 4870
rect 9809 4868 9833 4870
rect 9889 4868 9913 4870
rect 9969 4868 9993 4870
rect 10049 4868 10055 4870
rect 9747 4859 10055 4868
rect 9600 4814 9720 4842
rect 10244 4826 10272 5102
rect 9692 4128 9720 4814
rect 10232 4820 10284 4826
rect 10232 4762 10284 4768
rect 9600 4100 9720 4128
rect 10048 4140 10100 4146
rect 9600 3534 9628 4100
rect 10100 4100 10180 4128
rect 10048 4082 10100 4088
rect 9747 3836 10055 3845
rect 9747 3834 9753 3836
rect 9809 3834 9833 3836
rect 9889 3834 9913 3836
rect 9969 3834 9993 3836
rect 10049 3834 10055 3836
rect 9809 3782 9811 3834
rect 9991 3782 9993 3834
rect 9747 3780 9753 3782
rect 9809 3780 9833 3782
rect 9889 3780 9913 3782
rect 9969 3780 9993 3782
rect 10049 3780 10055 3782
rect 9747 3771 10055 3780
rect 9588 3528 9640 3534
rect 9588 3470 9640 3476
rect 9496 3460 9548 3466
rect 9496 3402 9548 3408
rect 9508 3194 9536 3402
rect 9588 3392 9640 3398
rect 9588 3334 9640 3340
rect 9496 3188 9548 3194
rect 9496 3130 9548 3136
rect 9404 3120 9456 3126
rect 9404 3062 9456 3068
rect 9140 2746 9260 2774
rect 9140 2582 9168 2746
rect 9128 2576 9180 2582
rect 9128 2518 9180 2524
rect 9128 2440 9180 2446
rect 9128 2382 9180 2388
rect 9404 2440 9456 2446
rect 9404 2382 9456 2388
rect 9036 1352 9088 1358
rect 9036 1294 9088 1300
rect 8944 808 8996 814
rect 8944 750 8996 756
rect 8114 54 8248 82
rect 8114 -300 8170 54
rect 8390 -300 8446 160
rect 8666 -300 8722 160
rect 8942 82 8998 160
rect 9140 82 9168 2382
rect 9220 2304 9272 2310
rect 9220 2246 9272 2252
rect 9312 2304 9364 2310
rect 9312 2246 9364 2252
rect 9232 2106 9260 2246
rect 9220 2100 9272 2106
rect 9220 2042 9272 2048
rect 9220 1284 9272 1290
rect 9220 1226 9272 1232
rect 9232 1193 9260 1226
rect 9324 1222 9352 2246
rect 9312 1216 9364 1222
rect 9218 1184 9274 1193
rect 9312 1158 9364 1164
rect 9218 1119 9274 1128
rect 8942 54 9168 82
rect 9218 82 9274 160
rect 9416 82 9444 2382
rect 9494 2000 9550 2009
rect 9494 1935 9550 1944
rect 9508 1902 9536 1935
rect 9496 1896 9548 1902
rect 9496 1838 9548 1844
rect 9600 1578 9628 3334
rect 9747 2748 10055 2757
rect 9747 2746 9753 2748
rect 9809 2746 9833 2748
rect 9889 2746 9913 2748
rect 9969 2746 9993 2748
rect 10049 2746 10055 2748
rect 9809 2694 9811 2746
rect 9991 2694 9993 2746
rect 9747 2692 9753 2694
rect 9809 2692 9833 2694
rect 9889 2692 9913 2694
rect 9969 2692 9993 2694
rect 10049 2692 10055 2694
rect 9747 2683 10055 2692
rect 9864 2644 9916 2650
rect 9864 2586 9916 2592
rect 9876 2446 9904 2586
rect 9864 2440 9916 2446
rect 9864 2382 9916 2388
rect 9678 2272 9734 2281
rect 9678 2207 9734 2216
rect 9692 1834 9720 2207
rect 10048 2032 10100 2038
rect 10152 2020 10180 4100
rect 10336 3398 10364 5306
rect 10520 4214 10548 6412
rect 10612 6254 10640 6734
rect 10600 6248 10652 6254
rect 10600 6190 10652 6196
rect 10508 4208 10560 4214
rect 10508 4150 10560 4156
rect 10704 4146 10732 9318
rect 10796 7478 10824 9608
rect 10784 7472 10836 7478
rect 10784 7414 10836 7420
rect 10796 5302 10824 7414
rect 10888 5794 10916 13212
rect 10980 11218 11008 18362
rect 11072 12434 11100 22066
rect 11242 21040 11298 21049
rect 11242 20975 11298 20984
rect 11256 20942 11284 20975
rect 11244 20936 11296 20942
rect 11150 20904 11206 20913
rect 11244 20878 11296 20884
rect 11150 20839 11206 20848
rect 11164 20534 11192 20839
rect 11152 20528 11204 20534
rect 11152 20470 11204 20476
rect 11152 20256 11204 20262
rect 11152 20198 11204 20204
rect 11164 19854 11192 20198
rect 11152 19848 11204 19854
rect 11152 19790 11204 19796
rect 11244 19780 11296 19786
rect 11244 19722 11296 19728
rect 11256 18970 11284 19722
rect 11244 18964 11296 18970
rect 11244 18906 11296 18912
rect 11244 18760 11296 18766
rect 11150 18728 11206 18737
rect 11244 18702 11296 18708
rect 11150 18663 11206 18672
rect 11164 17678 11192 18663
rect 11256 18329 11284 18702
rect 11242 18320 11298 18329
rect 11242 18255 11298 18264
rect 11152 17672 11204 17678
rect 11152 17614 11204 17620
rect 11152 17536 11204 17542
rect 11152 17478 11204 17484
rect 11164 17270 11192 17478
rect 11152 17264 11204 17270
rect 11152 17206 11204 17212
rect 11164 12782 11192 17206
rect 11348 16266 11376 24783
rect 11440 21978 11468 24822
rect 11532 24274 11560 25298
rect 11624 24750 11652 25978
rect 11716 25906 11744 27367
rect 11704 25900 11756 25906
rect 11704 25842 11756 25848
rect 11704 25288 11756 25294
rect 11704 25230 11756 25236
rect 11612 24744 11664 24750
rect 11612 24686 11664 24692
rect 11520 24268 11572 24274
rect 11520 24210 11572 24216
rect 11624 23730 11652 24686
rect 11716 24206 11744 25230
rect 11808 24562 11836 27406
rect 11900 24886 11928 30194
rect 11992 26897 12020 31175
rect 12084 30734 12112 31214
rect 12072 30728 12124 30734
rect 12072 30670 12124 30676
rect 12072 30592 12124 30598
rect 12072 30534 12124 30540
rect 12084 29510 12112 30534
rect 12072 29504 12124 29510
rect 12072 29446 12124 29452
rect 12084 29345 12112 29446
rect 12070 29336 12126 29345
rect 12070 29271 12126 29280
rect 12072 28688 12124 28694
rect 12072 28630 12124 28636
rect 12084 28082 12112 28630
rect 12072 28076 12124 28082
rect 12072 28018 12124 28024
rect 11978 26888 12034 26897
rect 11978 26823 12034 26832
rect 11978 26480 12034 26489
rect 11978 26415 12034 26424
rect 11888 24880 11940 24886
rect 11888 24822 11940 24828
rect 11992 24750 12020 26415
rect 12072 25424 12124 25430
rect 12070 25392 12072 25401
rect 12124 25392 12126 25401
rect 12070 25327 12126 25336
rect 11980 24744 12032 24750
rect 11980 24686 12032 24692
rect 11808 24534 11928 24562
rect 11704 24200 11756 24206
rect 11704 24142 11756 24148
rect 11704 23860 11756 23866
rect 11704 23802 11756 23808
rect 11612 23724 11664 23730
rect 11612 23666 11664 23672
rect 11520 23316 11572 23322
rect 11520 23258 11572 23264
rect 11532 22710 11560 23258
rect 11612 23044 11664 23050
rect 11716 23032 11744 23802
rect 11900 23769 11928 24534
rect 11886 23760 11942 23769
rect 11886 23695 11888 23704
rect 11940 23695 11942 23704
rect 11888 23666 11940 23672
rect 11900 23100 11928 23666
rect 11900 23072 12020 23100
rect 11716 23004 11928 23032
rect 11612 22986 11664 22992
rect 11520 22704 11572 22710
rect 11520 22646 11572 22652
rect 11520 22500 11572 22506
rect 11520 22442 11572 22448
rect 11532 22234 11560 22442
rect 11520 22228 11572 22234
rect 11520 22170 11572 22176
rect 11440 21950 11560 21978
rect 11428 21888 11480 21894
rect 11428 21830 11480 21836
rect 11440 16454 11468 21830
rect 11532 21554 11560 21950
rect 11520 21548 11572 21554
rect 11520 21490 11572 21496
rect 11532 21146 11560 21490
rect 11520 21140 11572 21146
rect 11520 21082 11572 21088
rect 11520 20392 11572 20398
rect 11518 20360 11520 20369
rect 11572 20360 11574 20369
rect 11518 20295 11574 20304
rect 11624 19854 11652 22986
rect 11796 22636 11848 22642
rect 11796 22578 11848 22584
rect 11702 21992 11758 22001
rect 11702 21927 11758 21936
rect 11716 21622 11744 21927
rect 11808 21894 11836 22578
rect 11796 21888 11848 21894
rect 11796 21830 11848 21836
rect 11794 21720 11850 21729
rect 11794 21655 11850 21664
rect 11704 21616 11756 21622
rect 11704 21558 11756 21564
rect 11612 19848 11664 19854
rect 11612 19790 11664 19796
rect 11716 18358 11744 21558
rect 11704 18352 11756 18358
rect 11704 18294 11756 18300
rect 11520 18284 11572 18290
rect 11520 18226 11572 18232
rect 11428 16448 11480 16454
rect 11428 16390 11480 16396
rect 11348 16238 11468 16266
rect 11336 15700 11388 15706
rect 11336 15642 11388 15648
rect 11244 15428 11296 15434
rect 11244 15370 11296 15376
rect 11152 12776 11204 12782
rect 11152 12718 11204 12724
rect 11072 12406 11192 12434
rect 10968 11212 11020 11218
rect 10968 11154 11020 11160
rect 11060 11212 11112 11218
rect 11060 11154 11112 11160
rect 11072 10810 11100 11154
rect 11060 10804 11112 10810
rect 11060 10746 11112 10752
rect 10968 10668 11020 10674
rect 10968 10610 11020 10616
rect 10980 8498 11008 10610
rect 11058 9480 11114 9489
rect 11058 9415 11114 9424
rect 10968 8492 11020 8498
rect 10968 8434 11020 8440
rect 11072 8362 11100 9415
rect 11164 8945 11192 12406
rect 11256 12238 11284 15370
rect 11348 14618 11376 15642
rect 11440 15366 11468 16238
rect 11428 15360 11480 15366
rect 11428 15302 11480 15308
rect 11532 14929 11560 18226
rect 11704 18216 11756 18222
rect 11704 18158 11756 18164
rect 11610 16688 11666 16697
rect 11610 16623 11612 16632
rect 11664 16623 11666 16632
rect 11612 16594 11664 16600
rect 11612 15632 11664 15638
rect 11612 15574 11664 15580
rect 11518 14920 11574 14929
rect 11518 14855 11574 14864
rect 11336 14612 11388 14618
rect 11336 14554 11388 14560
rect 11624 13870 11652 15574
rect 11612 13864 11664 13870
rect 11612 13806 11664 13812
rect 11336 13796 11388 13802
rect 11336 13738 11388 13744
rect 11348 12918 11376 13738
rect 11612 13728 11664 13734
rect 11612 13670 11664 13676
rect 11624 13433 11652 13670
rect 11610 13424 11666 13433
rect 11610 13359 11666 13368
rect 11716 13326 11744 18158
rect 11808 13802 11836 21655
rect 11900 18222 11928 23004
rect 11992 18714 12020 23072
rect 12084 22094 12112 25327
rect 12176 22506 12204 34070
rect 12268 33946 12296 34546
rect 12360 34134 12388 43250
rect 12532 43104 12584 43110
rect 12530 43072 12532 43081
rect 12584 43072 12586 43081
rect 12530 43007 12586 43016
rect 12636 42702 12664 43404
rect 13096 43314 13124 43846
rect 13188 43382 13216 43982
rect 13176 43376 13228 43382
rect 13372 43364 13400 44540
rect 13648 43602 13676 44540
rect 13648 43574 13768 43602
rect 13544 43376 13596 43382
rect 13372 43336 13544 43364
rect 13176 43318 13228 43324
rect 13544 43318 13596 43324
rect 13084 43308 13136 43314
rect 13084 43250 13136 43256
rect 13176 43240 13228 43246
rect 13176 43182 13228 43188
rect 13084 42764 13136 42770
rect 13084 42706 13136 42712
rect 12624 42696 12676 42702
rect 12624 42638 12676 42644
rect 12440 42560 12492 42566
rect 12440 42502 12492 42508
rect 12452 41449 12480 42502
rect 12679 42460 12987 42469
rect 12679 42458 12685 42460
rect 12741 42458 12765 42460
rect 12821 42458 12845 42460
rect 12901 42458 12925 42460
rect 12981 42458 12987 42460
rect 12741 42406 12743 42458
rect 12923 42406 12925 42458
rect 12679 42404 12685 42406
rect 12741 42404 12765 42406
rect 12821 42404 12845 42406
rect 12901 42404 12925 42406
rect 12981 42404 12987 42406
rect 12679 42395 12987 42404
rect 12438 41440 12494 41449
rect 12438 41375 12494 41384
rect 12679 41372 12987 41381
rect 12679 41370 12685 41372
rect 12741 41370 12765 41372
rect 12821 41370 12845 41372
rect 12901 41370 12925 41372
rect 12981 41370 12987 41372
rect 12741 41318 12743 41370
rect 12923 41318 12925 41370
rect 12679 41316 12685 41318
rect 12741 41316 12765 41318
rect 12821 41316 12845 41318
rect 12901 41316 12925 41318
rect 12981 41316 12987 41318
rect 12679 41307 12987 41316
rect 12679 40284 12987 40293
rect 12679 40282 12685 40284
rect 12741 40282 12765 40284
rect 12821 40282 12845 40284
rect 12901 40282 12925 40284
rect 12981 40282 12987 40284
rect 12741 40230 12743 40282
rect 12923 40230 12925 40282
rect 12679 40228 12685 40230
rect 12741 40228 12765 40230
rect 12821 40228 12845 40230
rect 12901 40228 12925 40230
rect 12981 40228 12987 40230
rect 12679 40219 12987 40228
rect 12440 39432 12492 39438
rect 12440 39374 12492 39380
rect 12452 36038 12480 39374
rect 12679 39196 12987 39205
rect 12679 39194 12685 39196
rect 12741 39194 12765 39196
rect 12821 39194 12845 39196
rect 12901 39194 12925 39196
rect 12981 39194 12987 39196
rect 12741 39142 12743 39194
rect 12923 39142 12925 39194
rect 12679 39140 12685 39142
rect 12741 39140 12765 39142
rect 12821 39140 12845 39142
rect 12901 39140 12925 39142
rect 12981 39140 12987 39142
rect 12679 39131 12987 39140
rect 12679 38108 12987 38117
rect 12679 38106 12685 38108
rect 12741 38106 12765 38108
rect 12821 38106 12845 38108
rect 12901 38106 12925 38108
rect 12981 38106 12987 38108
rect 12741 38054 12743 38106
rect 12923 38054 12925 38106
rect 12679 38052 12685 38054
rect 12741 38052 12765 38054
rect 12821 38052 12845 38054
rect 12901 38052 12925 38054
rect 12981 38052 12987 38054
rect 12679 38043 12987 38052
rect 12532 37664 12584 37670
rect 12532 37606 12584 37612
rect 12544 37262 12572 37606
rect 12532 37256 12584 37262
rect 12532 37198 12584 37204
rect 12679 37020 12987 37029
rect 12679 37018 12685 37020
rect 12741 37018 12765 37020
rect 12821 37018 12845 37020
rect 12901 37018 12925 37020
rect 12981 37018 12987 37020
rect 12741 36966 12743 37018
rect 12923 36966 12925 37018
rect 12679 36964 12685 36966
rect 12741 36964 12765 36966
rect 12821 36964 12845 36966
rect 12901 36964 12925 36966
rect 12981 36964 12987 36966
rect 12679 36955 12987 36964
rect 12440 36032 12492 36038
rect 12440 35974 12492 35980
rect 12679 35932 12987 35941
rect 12679 35930 12685 35932
rect 12741 35930 12765 35932
rect 12821 35930 12845 35932
rect 12901 35930 12925 35932
rect 12981 35930 12987 35932
rect 12741 35878 12743 35930
rect 12923 35878 12925 35930
rect 12679 35876 12685 35878
rect 12741 35876 12765 35878
rect 12821 35876 12845 35878
rect 12901 35876 12925 35878
rect 12981 35876 12987 35878
rect 12679 35867 12987 35876
rect 12532 35624 12584 35630
rect 12532 35566 12584 35572
rect 12716 35624 12768 35630
rect 12716 35566 12768 35572
rect 12544 34746 12572 35566
rect 12728 35290 12756 35566
rect 12716 35284 12768 35290
rect 12716 35226 12768 35232
rect 12679 34844 12987 34853
rect 12679 34842 12685 34844
rect 12741 34842 12765 34844
rect 12821 34842 12845 34844
rect 12901 34842 12925 34844
rect 12981 34842 12987 34844
rect 12741 34790 12743 34842
rect 12923 34790 12925 34842
rect 12679 34788 12685 34790
rect 12741 34788 12765 34790
rect 12821 34788 12845 34790
rect 12901 34788 12925 34790
rect 12981 34788 12987 34790
rect 12679 34779 12987 34788
rect 12532 34740 12584 34746
rect 12532 34682 12584 34688
rect 13096 34649 13124 42706
rect 13188 36564 13216 43182
rect 13360 43172 13412 43178
rect 13360 43114 13412 43120
rect 13268 36576 13320 36582
rect 13188 36536 13268 36564
rect 13268 36518 13320 36524
rect 13176 36100 13228 36106
rect 13176 36042 13228 36048
rect 13082 34640 13138 34649
rect 13082 34575 13138 34584
rect 12348 34128 12400 34134
rect 12348 34070 12400 34076
rect 12268 33918 12388 33946
rect 12256 33856 12308 33862
rect 12256 33798 12308 33804
rect 12268 33658 12296 33798
rect 12256 33652 12308 33658
rect 12256 33594 12308 33600
rect 12254 33416 12310 33425
rect 12254 33351 12310 33360
rect 12268 31249 12296 33351
rect 12360 32994 12388 33918
rect 13084 33924 13136 33930
rect 13084 33866 13136 33872
rect 12679 33756 12987 33765
rect 12679 33754 12685 33756
rect 12741 33754 12765 33756
rect 12821 33754 12845 33756
rect 12901 33754 12925 33756
rect 12981 33754 12987 33756
rect 12741 33702 12743 33754
rect 12923 33702 12925 33754
rect 12679 33700 12685 33702
rect 12741 33700 12765 33702
rect 12821 33700 12845 33702
rect 12901 33700 12925 33702
rect 12981 33700 12987 33702
rect 12679 33691 12987 33700
rect 13096 33658 13124 33866
rect 13084 33652 13136 33658
rect 13084 33594 13136 33600
rect 12808 33584 12860 33590
rect 12438 33552 12494 33561
rect 12808 33526 12860 33532
rect 12438 33487 12440 33496
rect 12492 33487 12494 33496
rect 12532 33516 12584 33522
rect 12440 33458 12492 33464
rect 12532 33458 12584 33464
rect 12360 32966 12480 32994
rect 12544 32978 12572 33458
rect 12820 33289 12848 33526
rect 13084 33312 13136 33318
rect 12806 33280 12862 33289
rect 13084 33254 13136 33260
rect 12806 33215 12862 33224
rect 12348 32904 12400 32910
rect 12348 32846 12400 32852
rect 12360 31890 12388 32846
rect 12348 31884 12400 31890
rect 12348 31826 12400 31832
rect 12360 31346 12388 31826
rect 12348 31340 12400 31346
rect 12348 31282 12400 31288
rect 12254 31240 12310 31249
rect 12254 31175 12310 31184
rect 12256 31136 12308 31142
rect 12452 31090 12480 32966
rect 12532 32972 12584 32978
rect 12532 32914 12584 32920
rect 13096 32842 13124 33254
rect 13084 32836 13136 32842
rect 13084 32778 13136 32784
rect 12679 32668 12987 32677
rect 12679 32666 12685 32668
rect 12741 32666 12765 32668
rect 12821 32666 12845 32668
rect 12901 32666 12925 32668
rect 12981 32666 12987 32668
rect 12741 32614 12743 32666
rect 12923 32614 12925 32666
rect 12679 32612 12685 32614
rect 12741 32612 12765 32614
rect 12821 32612 12845 32614
rect 12901 32612 12925 32614
rect 12981 32612 12987 32614
rect 12679 32603 12987 32612
rect 12624 32020 12676 32026
rect 12256 31078 12308 31084
rect 12268 30666 12296 31078
rect 12360 31062 12480 31090
rect 12544 31980 12624 32008
rect 12256 30660 12308 30666
rect 12256 30602 12308 30608
rect 12360 30546 12388 31062
rect 12544 30682 12572 31980
rect 12624 31962 12676 31968
rect 12679 31580 12987 31589
rect 12679 31578 12685 31580
rect 12741 31578 12765 31580
rect 12821 31578 12845 31580
rect 12901 31578 12925 31580
rect 12981 31578 12987 31580
rect 12741 31526 12743 31578
rect 12923 31526 12925 31578
rect 12679 31524 12685 31526
rect 12741 31524 12765 31526
rect 12821 31524 12845 31526
rect 12901 31524 12925 31526
rect 12981 31524 12987 31526
rect 12679 31515 12987 31524
rect 13096 31464 13124 32778
rect 13188 31822 13216 36042
rect 13268 34196 13320 34202
rect 13268 34138 13320 34144
rect 13280 33590 13308 34138
rect 13268 33584 13320 33590
rect 13268 33526 13320 33532
rect 13268 33312 13320 33318
rect 13268 33254 13320 33260
rect 13280 32434 13308 33254
rect 13268 32428 13320 32434
rect 13268 32370 13320 32376
rect 13176 31816 13228 31822
rect 13176 31758 13228 31764
rect 13176 31680 13228 31686
rect 13176 31622 13228 31628
rect 13004 31436 13124 31464
rect 12808 31272 12860 31278
rect 12806 31240 12808 31249
rect 12860 31240 12862 31249
rect 12806 31175 12862 31184
rect 12268 30518 12388 30546
rect 12452 30654 12572 30682
rect 13004 30666 13032 31436
rect 13084 30796 13136 30802
rect 13084 30738 13136 30744
rect 12992 30660 13044 30666
rect 12268 26382 12296 30518
rect 12452 30326 12480 30654
rect 12992 30602 13044 30608
rect 12532 30592 12584 30598
rect 12530 30560 12532 30569
rect 12584 30560 12586 30569
rect 12530 30495 12586 30504
rect 12679 30492 12987 30501
rect 12679 30490 12685 30492
rect 12741 30490 12765 30492
rect 12821 30490 12845 30492
rect 12901 30490 12925 30492
rect 12981 30490 12987 30492
rect 12741 30438 12743 30490
rect 12923 30438 12925 30490
rect 12679 30436 12685 30438
rect 12741 30436 12765 30438
rect 12821 30436 12845 30438
rect 12901 30436 12925 30438
rect 12981 30436 12987 30438
rect 12679 30427 12987 30436
rect 12440 30320 12492 30326
rect 12440 30262 12492 30268
rect 13096 30122 13124 30738
rect 13188 30734 13216 31622
rect 13268 31476 13320 31482
rect 13268 31418 13320 31424
rect 13176 30728 13228 30734
rect 13176 30670 13228 30676
rect 13280 30326 13308 31418
rect 13176 30320 13228 30326
rect 13176 30262 13228 30268
rect 13268 30320 13320 30326
rect 13268 30262 13320 30268
rect 13084 30116 13136 30122
rect 13084 30058 13136 30064
rect 12348 30048 12400 30054
rect 12400 29996 12572 30002
rect 12348 29990 12572 29996
rect 12360 29974 12572 29990
rect 12452 28234 12480 29974
rect 12544 29850 12572 29974
rect 12532 29844 12584 29850
rect 12532 29786 12584 29792
rect 12532 29708 12584 29714
rect 12532 29650 12584 29656
rect 12360 28206 12480 28234
rect 12360 27962 12388 28206
rect 12438 28112 12494 28121
rect 12438 28047 12440 28056
rect 12492 28047 12494 28056
rect 12440 28018 12492 28024
rect 12360 27934 12480 27962
rect 12256 26376 12308 26382
rect 12254 26344 12256 26353
rect 12308 26344 12310 26353
rect 12254 26279 12310 26288
rect 12348 25900 12400 25906
rect 12348 25842 12400 25848
rect 12256 25356 12308 25362
rect 12256 25298 12308 25304
rect 12268 24886 12296 25298
rect 12256 24880 12308 24886
rect 12256 24822 12308 24828
rect 12360 24410 12388 25842
rect 12452 25242 12480 27934
rect 12544 26024 12572 29650
rect 12679 29404 12987 29413
rect 12679 29402 12685 29404
rect 12741 29402 12765 29404
rect 12821 29402 12845 29404
rect 12901 29402 12925 29404
rect 12981 29402 12987 29404
rect 12741 29350 12743 29402
rect 12923 29350 12925 29402
rect 12679 29348 12685 29350
rect 12741 29348 12765 29350
rect 12821 29348 12845 29350
rect 12901 29348 12925 29350
rect 12981 29348 12987 29350
rect 12679 29339 12987 29348
rect 13084 29096 13136 29102
rect 13084 29038 13136 29044
rect 12679 28316 12987 28325
rect 12679 28314 12685 28316
rect 12741 28314 12765 28316
rect 12821 28314 12845 28316
rect 12901 28314 12925 28316
rect 12981 28314 12987 28316
rect 12741 28262 12743 28314
rect 12923 28262 12925 28314
rect 12679 28260 12685 28262
rect 12741 28260 12765 28262
rect 12821 28260 12845 28262
rect 12901 28260 12925 28262
rect 12981 28260 12987 28262
rect 12679 28251 12987 28260
rect 12900 28144 12952 28150
rect 12900 28086 12952 28092
rect 12912 27418 12940 28086
rect 12990 27976 13046 27985
rect 12990 27911 12992 27920
rect 13044 27911 13046 27920
rect 12992 27882 13044 27888
rect 13096 27713 13124 29038
rect 13188 28994 13216 30262
rect 13280 29578 13308 30262
rect 13268 29572 13320 29578
rect 13268 29514 13320 29520
rect 13188 28966 13308 28994
rect 13176 28484 13228 28490
rect 13176 28426 13228 28432
rect 13188 28082 13216 28426
rect 13176 28076 13228 28082
rect 13176 28018 13228 28024
rect 13082 27704 13138 27713
rect 13082 27639 13138 27648
rect 12912 27390 13124 27418
rect 12679 27228 12987 27237
rect 12679 27226 12685 27228
rect 12741 27226 12765 27228
rect 12821 27226 12845 27228
rect 12901 27226 12925 27228
rect 12981 27226 12987 27228
rect 12741 27174 12743 27226
rect 12923 27174 12925 27226
rect 12679 27172 12685 27174
rect 12741 27172 12765 27174
rect 12821 27172 12845 27174
rect 12901 27172 12925 27174
rect 12981 27172 12987 27174
rect 12679 27163 12987 27172
rect 13096 26586 13124 27390
rect 13176 26784 13228 26790
rect 13176 26726 13228 26732
rect 13084 26580 13136 26586
rect 13084 26522 13136 26528
rect 13084 26240 13136 26246
rect 13084 26182 13136 26188
rect 12679 26140 12987 26149
rect 12679 26138 12685 26140
rect 12741 26138 12765 26140
rect 12821 26138 12845 26140
rect 12901 26138 12925 26140
rect 12981 26138 12987 26140
rect 12741 26086 12743 26138
rect 12923 26086 12925 26138
rect 12679 26084 12685 26086
rect 12741 26084 12765 26086
rect 12821 26084 12845 26086
rect 12901 26084 12925 26086
rect 12981 26084 12987 26086
rect 12679 26075 12987 26084
rect 12544 25996 12756 26024
rect 12532 25696 12584 25702
rect 12532 25638 12584 25644
rect 12544 25498 12572 25638
rect 12532 25492 12584 25498
rect 12532 25434 12584 25440
rect 12530 25392 12586 25401
rect 12530 25327 12532 25336
rect 12584 25327 12586 25336
rect 12532 25298 12584 25304
rect 12728 25242 12756 25996
rect 13096 25362 13124 26182
rect 13084 25356 13136 25362
rect 13084 25298 13136 25304
rect 12452 25214 12572 25242
rect 12728 25214 13124 25242
rect 12348 24404 12400 24410
rect 12348 24346 12400 24352
rect 12348 24268 12400 24274
rect 12348 24210 12400 24216
rect 12440 24268 12492 24274
rect 12440 24210 12492 24216
rect 12360 23254 12388 24210
rect 12452 23866 12480 24210
rect 12440 23860 12492 23866
rect 12440 23802 12492 23808
rect 12544 23780 12572 25214
rect 12679 25052 12987 25061
rect 12679 25050 12685 25052
rect 12741 25050 12765 25052
rect 12821 25050 12845 25052
rect 12901 25050 12925 25052
rect 12981 25050 12987 25052
rect 12741 24998 12743 25050
rect 12923 24998 12925 25050
rect 12679 24996 12685 24998
rect 12741 24996 12765 24998
rect 12821 24996 12845 24998
rect 12901 24996 12925 24998
rect 12981 24996 12987 24998
rect 12679 24987 12987 24996
rect 12716 24200 12768 24206
rect 12768 24160 12848 24188
rect 12716 24142 12768 24148
rect 12820 24052 12848 24160
rect 13096 24154 13124 25214
rect 13188 24274 13216 26726
rect 13176 24268 13228 24274
rect 13176 24210 13228 24216
rect 13096 24126 13216 24154
rect 12820 24024 13124 24052
rect 12679 23964 12987 23973
rect 12679 23962 12685 23964
rect 12741 23962 12765 23964
rect 12821 23962 12845 23964
rect 12901 23962 12925 23964
rect 12981 23962 12987 23964
rect 12741 23910 12743 23962
rect 12923 23910 12925 23962
rect 12679 23908 12685 23910
rect 12741 23908 12765 23910
rect 12821 23908 12845 23910
rect 12901 23908 12925 23910
rect 12981 23908 12987 23910
rect 12679 23899 12987 23908
rect 13096 23866 13124 24024
rect 13084 23860 13136 23866
rect 13084 23802 13136 23808
rect 12544 23752 12664 23780
rect 12348 23248 12400 23254
rect 12348 23190 12400 23196
rect 12256 22976 12308 22982
rect 12256 22918 12308 22924
rect 12164 22500 12216 22506
rect 12164 22442 12216 22448
rect 12084 22066 12204 22094
rect 12072 21888 12124 21894
rect 12176 21865 12204 22066
rect 12268 22030 12296 22918
rect 12360 22642 12388 23190
rect 12532 23112 12584 23118
rect 12532 23054 12584 23060
rect 12440 22976 12492 22982
rect 12440 22918 12492 22924
rect 12452 22642 12480 22918
rect 12348 22636 12400 22642
rect 12348 22578 12400 22584
rect 12440 22636 12492 22642
rect 12440 22578 12492 22584
rect 12440 22092 12492 22098
rect 12440 22034 12492 22040
rect 12256 22024 12308 22030
rect 12256 21966 12308 21972
rect 12348 21956 12400 21962
rect 12348 21898 12400 21904
rect 12072 21830 12124 21836
rect 12162 21856 12218 21865
rect 12084 21690 12112 21830
rect 12162 21791 12218 21800
rect 12360 21690 12388 21898
rect 12072 21684 12124 21690
rect 12348 21684 12400 21690
rect 12124 21644 12204 21672
rect 12072 21626 12124 21632
rect 12072 21548 12124 21554
rect 12072 21490 12124 21496
rect 12084 19922 12112 21490
rect 12176 21434 12204 21644
rect 12348 21626 12400 21632
rect 12176 21406 12296 21434
rect 12164 21344 12216 21350
rect 12164 21286 12216 21292
rect 12176 21078 12204 21286
rect 12164 21072 12216 21078
rect 12164 21014 12216 21020
rect 12268 20924 12296 21406
rect 12452 21146 12480 22034
rect 12544 21962 12572 23054
rect 12636 22964 12664 23752
rect 12602 22936 12664 22964
rect 12602 22692 12630 22936
rect 12679 22876 12987 22885
rect 12679 22874 12685 22876
rect 12741 22874 12765 22876
rect 12821 22874 12845 22876
rect 12901 22874 12925 22876
rect 12981 22874 12987 22876
rect 12741 22822 12743 22874
rect 12923 22822 12925 22874
rect 12679 22820 12685 22822
rect 12741 22820 12765 22822
rect 12821 22820 12845 22822
rect 12901 22820 12925 22822
rect 12981 22820 12987 22822
rect 12679 22811 12987 22820
rect 12716 22704 12768 22710
rect 12602 22664 12716 22692
rect 12716 22646 12768 22652
rect 13096 22098 13124 23802
rect 13188 23338 13216 24126
rect 13280 23497 13308 28966
rect 13266 23488 13322 23497
rect 13266 23423 13322 23432
rect 13188 23310 13308 23338
rect 13280 22250 13308 23310
rect 13188 22222 13308 22250
rect 13084 22092 13136 22098
rect 13084 22034 13136 22040
rect 13188 21978 13216 22222
rect 13268 22160 13320 22166
rect 13266 22128 13268 22137
rect 13320 22128 13322 22137
rect 13266 22063 13322 22072
rect 12532 21956 12584 21962
rect 12532 21898 12584 21904
rect 13096 21950 13216 21978
rect 12440 21140 12492 21146
rect 12440 21082 12492 21088
rect 12544 20942 12572 21898
rect 12679 21788 12987 21797
rect 12679 21786 12685 21788
rect 12741 21786 12765 21788
rect 12821 21786 12845 21788
rect 12901 21786 12925 21788
rect 12981 21786 12987 21788
rect 12741 21734 12743 21786
rect 12923 21734 12925 21786
rect 12679 21732 12685 21734
rect 12741 21732 12765 21734
rect 12821 21732 12845 21734
rect 12901 21732 12925 21734
rect 12981 21732 12987 21734
rect 12679 21723 12987 21732
rect 12900 21412 12952 21418
rect 12900 21354 12952 21360
rect 12912 21078 12940 21354
rect 12900 21072 12952 21078
rect 12900 21014 12952 21020
rect 12176 20896 12296 20924
rect 12532 20936 12584 20942
rect 12072 19916 12124 19922
rect 12072 19858 12124 19864
rect 12084 19417 12112 19858
rect 12070 19408 12126 19417
rect 12070 19343 12072 19352
rect 12124 19343 12126 19352
rect 12072 19314 12124 19320
rect 11992 18686 12112 18714
rect 11980 18624 12032 18630
rect 11980 18566 12032 18572
rect 11992 18290 12020 18566
rect 11980 18284 12032 18290
rect 11980 18226 12032 18232
rect 11888 18216 11940 18222
rect 11888 18158 11940 18164
rect 11888 18080 11940 18086
rect 11888 18022 11940 18028
rect 11900 17882 11928 18022
rect 11888 17876 11940 17882
rect 11888 17818 11940 17824
rect 11888 17536 11940 17542
rect 11888 17478 11940 17484
rect 11900 14550 11928 17478
rect 11980 16516 12032 16522
rect 11980 16458 12032 16464
rect 11992 14958 12020 16458
rect 11980 14952 12032 14958
rect 11980 14894 12032 14900
rect 11888 14544 11940 14550
rect 11888 14486 11940 14492
rect 11980 14544 12032 14550
rect 11980 14486 12032 14492
rect 11796 13796 11848 13802
rect 11796 13738 11848 13744
rect 11900 13530 11928 14486
rect 11888 13524 11940 13530
rect 11888 13466 11940 13472
rect 11992 13394 12020 14486
rect 12084 14074 12112 18686
rect 12176 15638 12204 20896
rect 12532 20878 12584 20884
rect 12440 20868 12492 20874
rect 12440 20810 12492 20816
rect 12256 20528 12308 20534
rect 12256 20470 12308 20476
rect 12346 20496 12402 20505
rect 12268 20058 12296 20470
rect 12346 20431 12348 20440
rect 12400 20431 12402 20440
rect 12348 20402 12400 20408
rect 12256 20052 12308 20058
rect 12256 19994 12308 20000
rect 12256 19780 12308 19786
rect 12256 19722 12308 19728
rect 12268 18766 12296 19722
rect 12452 19334 12480 20810
rect 12679 20700 12987 20709
rect 12679 20698 12685 20700
rect 12741 20698 12765 20700
rect 12821 20698 12845 20700
rect 12901 20698 12925 20700
rect 12981 20698 12987 20700
rect 12741 20646 12743 20698
rect 12923 20646 12925 20698
rect 12679 20644 12685 20646
rect 12741 20644 12765 20646
rect 12821 20644 12845 20646
rect 12901 20644 12925 20646
rect 12981 20644 12987 20646
rect 12679 20635 12987 20644
rect 12532 20256 12584 20262
rect 12532 20198 12584 20204
rect 12360 19306 12480 19334
rect 12256 18760 12308 18766
rect 12256 18702 12308 18708
rect 12256 17672 12308 17678
rect 12256 17614 12308 17620
rect 12268 17338 12296 17614
rect 12256 17332 12308 17338
rect 12256 17274 12308 17280
rect 12256 16992 12308 16998
rect 12256 16934 12308 16940
rect 12268 16794 12296 16934
rect 12256 16788 12308 16794
rect 12256 16730 12308 16736
rect 12268 15706 12296 16730
rect 12360 15978 12388 19306
rect 12440 19168 12492 19174
rect 12440 19110 12492 19116
rect 12452 18970 12480 19110
rect 12440 18964 12492 18970
rect 12440 18906 12492 18912
rect 12440 17672 12492 17678
rect 12440 17614 12492 17620
rect 12452 17338 12480 17614
rect 12440 17332 12492 17338
rect 12440 17274 12492 17280
rect 12440 16448 12492 16454
rect 12440 16390 12492 16396
rect 12452 16046 12480 16390
rect 12440 16040 12492 16046
rect 12440 15982 12492 15988
rect 12348 15972 12400 15978
rect 12348 15914 12400 15920
rect 12256 15700 12308 15706
rect 12256 15642 12308 15648
rect 12164 15632 12216 15638
rect 12164 15574 12216 15580
rect 12544 15552 12572 20198
rect 12679 19612 12987 19621
rect 12679 19610 12685 19612
rect 12741 19610 12765 19612
rect 12821 19610 12845 19612
rect 12901 19610 12925 19612
rect 12981 19610 12987 19612
rect 12741 19558 12743 19610
rect 12923 19558 12925 19610
rect 12679 19556 12685 19558
rect 12741 19556 12765 19558
rect 12821 19556 12845 19558
rect 12901 19556 12925 19558
rect 12981 19556 12987 19558
rect 12679 19547 12987 19556
rect 13096 19334 13124 21950
rect 13176 21888 13228 21894
rect 13176 21830 13228 21836
rect 13188 20874 13216 21830
rect 13176 20868 13228 20874
rect 13176 20810 13228 20816
rect 13188 20466 13216 20810
rect 13372 20618 13400 43114
rect 13636 43104 13688 43110
rect 13636 43046 13688 43052
rect 13648 41414 13676 43046
rect 13740 42702 13768 43574
rect 13924 43296 13952 44540
rect 14200 43602 14228 44540
rect 14200 43574 14320 43602
rect 14096 43308 14148 43314
rect 13924 43268 14096 43296
rect 14096 43250 14148 43256
rect 14188 43172 14240 43178
rect 14188 43114 14240 43120
rect 13728 42696 13780 42702
rect 13728 42638 13780 42644
rect 14096 42560 14148 42566
rect 13464 41386 13676 41414
rect 13740 42520 14096 42548
rect 13464 30682 13492 41386
rect 13544 40452 13596 40458
rect 13544 40394 13596 40400
rect 13556 37806 13584 40394
rect 13636 39908 13688 39914
rect 13636 39850 13688 39856
rect 13648 38321 13676 39850
rect 13634 38312 13690 38321
rect 13634 38247 13690 38256
rect 13544 37800 13596 37806
rect 13596 37760 13676 37788
rect 13544 37742 13596 37748
rect 13544 36576 13596 36582
rect 13544 36518 13596 36524
rect 13556 31226 13584 36518
rect 13648 35834 13676 37760
rect 13636 35828 13688 35834
rect 13636 35770 13688 35776
rect 13648 33658 13676 35770
rect 13636 33652 13688 33658
rect 13636 33594 13688 33600
rect 13636 33040 13688 33046
rect 13636 32982 13688 32988
rect 13648 32842 13676 32982
rect 13636 32836 13688 32842
rect 13636 32778 13688 32784
rect 13636 32292 13688 32298
rect 13636 32234 13688 32240
rect 13648 32026 13676 32234
rect 13636 32020 13688 32026
rect 13636 31962 13688 31968
rect 13636 31816 13688 31822
rect 13636 31758 13688 31764
rect 13648 31414 13676 31758
rect 13740 31482 13768 42520
rect 14096 42502 14148 42508
rect 14200 42378 14228 43114
rect 14292 42702 14320 43574
rect 14476 43314 14504 44540
rect 14464 43308 14516 43314
rect 14752 43296 14780 44540
rect 15028 43602 15056 44540
rect 15028 43574 15148 43602
rect 14832 43308 14884 43314
rect 14752 43268 14832 43296
rect 14464 43250 14516 43256
rect 14832 43250 14884 43256
rect 15016 43240 15068 43246
rect 15016 43182 15068 43188
rect 14648 43104 14700 43110
rect 14648 43046 14700 43052
rect 14280 42696 14332 42702
rect 14280 42638 14332 42644
rect 14016 42350 14228 42378
rect 13912 41676 13964 41682
rect 13912 41618 13964 41624
rect 13820 41608 13872 41614
rect 13820 41550 13872 41556
rect 13832 41177 13860 41550
rect 13924 41206 13952 41618
rect 13912 41200 13964 41206
rect 13818 41168 13874 41177
rect 13912 41142 13964 41148
rect 13818 41103 13874 41112
rect 14016 41041 14044 42350
rect 14094 42256 14150 42265
rect 14094 42191 14150 42200
rect 14002 41032 14058 41041
rect 14002 40967 14058 40976
rect 13820 37800 13872 37806
rect 13820 37742 13872 37748
rect 13832 36854 13860 37742
rect 13820 36848 13872 36854
rect 13820 36790 13872 36796
rect 13820 36032 13872 36038
rect 14108 35986 14136 42191
rect 14660 38826 14688 43046
rect 15028 42945 15056 43182
rect 15014 42936 15070 42945
rect 14924 42900 14976 42906
rect 15014 42871 15070 42880
rect 14924 42842 14976 42848
rect 14648 38820 14700 38826
rect 14648 38762 14700 38768
rect 14188 36780 14240 36786
rect 14188 36722 14240 36728
rect 13820 35974 13872 35980
rect 13832 35766 13860 35974
rect 13924 35958 14136 35986
rect 13820 35760 13872 35766
rect 13820 35702 13872 35708
rect 13832 34610 13860 35702
rect 13820 34604 13872 34610
rect 13820 34546 13872 34552
rect 13820 33108 13872 33114
rect 13820 33050 13872 33056
rect 13832 32366 13860 33050
rect 13820 32360 13872 32366
rect 13820 32302 13872 32308
rect 13924 31754 13952 35958
rect 14004 32768 14056 32774
rect 14004 32710 14056 32716
rect 14016 31890 14044 32710
rect 14200 32450 14228 36722
rect 14556 36168 14608 36174
rect 14556 36110 14608 36116
rect 14568 35834 14596 36110
rect 14740 36032 14792 36038
rect 14740 35974 14792 35980
rect 14556 35828 14608 35834
rect 14556 35770 14608 35776
rect 14752 35630 14780 35974
rect 14936 35834 14964 42842
rect 15120 42702 15148 43574
rect 15304 43382 15332 44540
rect 15292 43376 15344 43382
rect 15292 43318 15344 43324
rect 15580 43314 15608 44540
rect 15856 43364 15884 44540
rect 16132 43450 16160 44540
rect 16120 43444 16172 43450
rect 16120 43386 16172 43392
rect 16028 43376 16080 43382
rect 15856 43336 16028 43364
rect 16028 43318 16080 43324
rect 16408 43314 16436 44540
rect 15568 43308 15620 43314
rect 15568 43250 15620 43256
rect 16396 43308 16448 43314
rect 16396 43250 16448 43256
rect 16684 43246 16712 44540
rect 16856 43648 16908 43654
rect 16856 43590 16908 43596
rect 16868 43382 16896 43590
rect 16856 43376 16908 43382
rect 16960 43364 16988 44540
rect 17236 43874 17264 44540
rect 17512 44010 17540 44540
rect 17788 44146 17816 44540
rect 17788 44118 18000 44146
rect 18064 44130 18092 44540
rect 17972 44062 18000 44118
rect 18052 44124 18104 44130
rect 18052 44066 18104 44072
rect 17960 44056 18012 44062
rect 17512 43994 17816 44010
rect 17960 43998 18012 44004
rect 17512 43988 17828 43994
rect 17512 43982 17776 43988
rect 17776 43930 17828 43936
rect 17236 43846 18092 43874
rect 17316 43444 17368 43450
rect 17316 43386 17368 43392
rect 17224 43376 17276 43382
rect 16960 43336 17224 43364
rect 16856 43318 16908 43324
rect 17224 43318 17276 43324
rect 16672 43240 16724 43246
rect 16672 43182 16724 43188
rect 15476 43104 15528 43110
rect 15476 43046 15528 43052
rect 16304 43104 16356 43110
rect 16304 43046 16356 43052
rect 15488 42945 15516 43046
rect 15612 43004 15920 43013
rect 15612 43002 15618 43004
rect 15674 43002 15698 43004
rect 15754 43002 15778 43004
rect 15834 43002 15858 43004
rect 15914 43002 15920 43004
rect 15674 42950 15676 43002
rect 15856 42950 15858 43002
rect 15612 42948 15618 42950
rect 15674 42948 15698 42950
rect 15754 42948 15778 42950
rect 15834 42948 15858 42950
rect 15914 42948 15920 42950
rect 15474 42936 15530 42945
rect 15612 42939 15920 42948
rect 15474 42871 15530 42880
rect 15108 42696 15160 42702
rect 15108 42638 15160 42644
rect 15612 41916 15920 41925
rect 15612 41914 15618 41916
rect 15674 41914 15698 41916
rect 15754 41914 15778 41916
rect 15834 41914 15858 41916
rect 15914 41914 15920 41916
rect 15674 41862 15676 41914
rect 15856 41862 15858 41914
rect 15612 41860 15618 41862
rect 15674 41860 15698 41862
rect 15754 41860 15778 41862
rect 15834 41860 15858 41862
rect 15914 41860 15920 41862
rect 15612 41851 15920 41860
rect 15200 41812 15252 41818
rect 15200 41754 15252 41760
rect 15212 39001 15240 41754
rect 16212 41064 16264 41070
rect 16212 41006 16264 41012
rect 15612 40828 15920 40837
rect 15612 40826 15618 40828
rect 15674 40826 15698 40828
rect 15754 40826 15778 40828
rect 15834 40826 15858 40828
rect 15914 40826 15920 40828
rect 15674 40774 15676 40826
rect 15856 40774 15858 40826
rect 15612 40772 15618 40774
rect 15674 40772 15698 40774
rect 15754 40772 15778 40774
rect 15834 40772 15858 40774
rect 15914 40772 15920 40774
rect 15612 40763 15920 40772
rect 15612 39740 15920 39749
rect 15612 39738 15618 39740
rect 15674 39738 15698 39740
rect 15754 39738 15778 39740
rect 15834 39738 15858 39740
rect 15914 39738 15920 39740
rect 15674 39686 15676 39738
rect 15856 39686 15858 39738
rect 15612 39684 15618 39686
rect 15674 39684 15698 39686
rect 15754 39684 15778 39686
rect 15834 39684 15858 39686
rect 15914 39684 15920 39686
rect 15612 39675 15920 39684
rect 15198 38992 15254 39001
rect 15198 38927 15254 38936
rect 15612 38652 15920 38661
rect 15612 38650 15618 38652
rect 15674 38650 15698 38652
rect 15754 38650 15778 38652
rect 15834 38650 15858 38652
rect 15914 38650 15920 38652
rect 15674 38598 15676 38650
rect 15856 38598 15858 38650
rect 15612 38596 15618 38598
rect 15674 38596 15698 38598
rect 15754 38596 15778 38598
rect 15834 38596 15858 38598
rect 15914 38596 15920 38598
rect 15612 38587 15920 38596
rect 15476 38276 15528 38282
rect 15476 38218 15528 38224
rect 15488 37874 15516 38218
rect 15476 37868 15528 37874
rect 15476 37810 15528 37816
rect 15016 36168 15068 36174
rect 15016 36110 15068 36116
rect 14924 35828 14976 35834
rect 14924 35770 14976 35776
rect 14924 35692 14976 35698
rect 14924 35634 14976 35640
rect 14740 35624 14792 35630
rect 14740 35566 14792 35572
rect 14936 35290 14964 35634
rect 15028 35290 15056 36110
rect 14924 35284 14976 35290
rect 14924 35226 14976 35232
rect 15016 35284 15068 35290
rect 15016 35226 15068 35232
rect 14924 35080 14976 35086
rect 14924 35022 14976 35028
rect 15200 35080 15252 35086
rect 15200 35022 15252 35028
rect 14648 33448 14700 33454
rect 14648 33390 14700 33396
rect 14832 33448 14884 33454
rect 14832 33390 14884 33396
rect 14372 33312 14424 33318
rect 14372 33254 14424 33260
rect 14280 32904 14332 32910
rect 14384 32881 14412 33254
rect 14464 32904 14516 32910
rect 14280 32846 14332 32852
rect 14370 32872 14426 32881
rect 14108 32422 14228 32450
rect 14004 31884 14056 31890
rect 14004 31826 14056 31832
rect 14108 31754 14136 32422
rect 14188 32360 14240 32366
rect 14292 32337 14320 32846
rect 14464 32846 14516 32852
rect 14370 32807 14426 32816
rect 14384 32434 14412 32807
rect 14372 32428 14424 32434
rect 14372 32370 14424 32376
rect 14188 32302 14240 32308
rect 14278 32328 14334 32337
rect 14200 31958 14228 32302
rect 14278 32263 14334 32272
rect 14280 32224 14332 32230
rect 14280 32166 14332 32172
rect 14188 31952 14240 31958
rect 14188 31894 14240 31900
rect 13924 31726 14044 31754
rect 14108 31726 14253 31754
rect 13728 31476 13780 31482
rect 13728 31418 13780 31424
rect 13636 31408 13688 31414
rect 13636 31350 13688 31356
rect 13556 31198 13952 31226
rect 13636 31136 13688 31142
rect 13636 31078 13688 31084
rect 13820 31136 13872 31142
rect 13820 31078 13872 31084
rect 13648 30734 13676 31078
rect 13636 30728 13688 30734
rect 13464 30654 13584 30682
rect 13636 30670 13688 30676
rect 13452 30592 13504 30598
rect 13452 30534 13504 30540
rect 13464 30394 13492 30534
rect 13556 30410 13584 30654
rect 13636 30592 13688 30598
rect 13688 30552 13768 30580
rect 13636 30534 13688 30540
rect 13452 30388 13504 30394
rect 13556 30382 13676 30410
rect 13452 30330 13504 30336
rect 13452 30048 13504 30054
rect 13452 29990 13504 29996
rect 13464 29073 13492 29990
rect 13450 29064 13506 29073
rect 13450 28999 13506 29008
rect 13544 29028 13596 29034
rect 13544 28970 13596 28976
rect 13556 28762 13584 28970
rect 13544 28756 13596 28762
rect 13544 28698 13596 28704
rect 13648 28642 13676 30382
rect 13556 28614 13676 28642
rect 13452 27396 13504 27402
rect 13452 27338 13504 27344
rect 13464 26586 13492 27338
rect 13452 26580 13504 26586
rect 13452 26522 13504 26528
rect 13452 24880 13504 24886
rect 13452 24822 13504 24828
rect 13464 22681 13492 24822
rect 13450 22672 13506 22681
rect 13450 22607 13452 22616
rect 13504 22607 13506 22616
rect 13452 22578 13504 22584
rect 13452 22092 13504 22098
rect 13452 22034 13504 22040
rect 13280 20590 13400 20618
rect 13464 20618 13492 22034
rect 13556 20777 13584 28614
rect 13636 28552 13688 28558
rect 13636 28494 13688 28500
rect 13542 20768 13598 20777
rect 13542 20703 13598 20712
rect 13464 20590 13584 20618
rect 13176 20460 13228 20466
rect 13176 20402 13228 20408
rect 13174 19680 13230 19689
rect 13174 19615 13230 19624
rect 13188 19446 13216 19615
rect 13176 19440 13228 19446
rect 13176 19382 13228 19388
rect 13096 19306 13216 19334
rect 12679 18524 12987 18533
rect 12679 18522 12685 18524
rect 12741 18522 12765 18524
rect 12821 18522 12845 18524
rect 12901 18522 12925 18524
rect 12981 18522 12987 18524
rect 12741 18470 12743 18522
rect 12923 18470 12925 18522
rect 12679 18468 12685 18470
rect 12741 18468 12765 18470
rect 12821 18468 12845 18470
rect 12901 18468 12925 18470
rect 12981 18468 12987 18470
rect 12679 18459 12987 18468
rect 12679 17436 12987 17445
rect 12679 17434 12685 17436
rect 12741 17434 12765 17436
rect 12821 17434 12845 17436
rect 12901 17434 12925 17436
rect 12981 17434 12987 17436
rect 12741 17382 12743 17434
rect 12923 17382 12925 17434
rect 12679 17380 12685 17382
rect 12741 17380 12765 17382
rect 12821 17380 12845 17382
rect 12901 17380 12925 17382
rect 12981 17380 12987 17382
rect 12679 17371 12987 17380
rect 13084 16448 13136 16454
rect 13084 16390 13136 16396
rect 12679 16348 12987 16357
rect 12679 16346 12685 16348
rect 12741 16346 12765 16348
rect 12821 16346 12845 16348
rect 12901 16346 12925 16348
rect 12981 16346 12987 16348
rect 12741 16294 12743 16346
rect 12923 16294 12925 16346
rect 12679 16292 12685 16294
rect 12741 16292 12765 16294
rect 12821 16292 12845 16294
rect 12901 16292 12925 16294
rect 12981 16292 12987 16294
rect 12679 16283 12987 16292
rect 12992 16244 13044 16250
rect 12992 16186 13044 16192
rect 12268 15524 12572 15552
rect 12072 14068 12124 14074
rect 12072 14010 12124 14016
rect 12164 14068 12216 14074
rect 12164 14010 12216 14016
rect 11980 13388 12032 13394
rect 11980 13330 12032 13336
rect 11704 13320 11756 13326
rect 11756 13280 11836 13308
rect 11704 13262 11756 13268
rect 11612 13184 11664 13190
rect 11612 13126 11664 13132
rect 11624 12918 11652 13126
rect 11336 12912 11388 12918
rect 11336 12854 11388 12860
rect 11612 12912 11664 12918
rect 11612 12854 11664 12860
rect 11808 12832 11836 13280
rect 12084 13258 12112 14010
rect 12072 13252 12124 13258
rect 12072 13194 12124 13200
rect 11980 13184 12032 13190
rect 11980 13126 12032 13132
rect 11888 12844 11940 12850
rect 11808 12804 11888 12832
rect 11520 12776 11572 12782
rect 11520 12718 11572 12724
rect 11244 12232 11296 12238
rect 11244 12174 11296 12180
rect 11256 10674 11284 12174
rect 11532 11694 11560 12718
rect 11520 11688 11572 11694
rect 11520 11630 11572 11636
rect 11336 11144 11388 11150
rect 11336 11086 11388 11092
rect 11244 10668 11296 10674
rect 11244 10610 11296 10616
rect 11242 9072 11298 9081
rect 11242 9007 11298 9016
rect 11150 8936 11206 8945
rect 11150 8871 11206 8880
rect 11152 8832 11204 8838
rect 11152 8774 11204 8780
rect 11060 8356 11112 8362
rect 11060 8298 11112 8304
rect 10968 7948 11020 7954
rect 11020 7908 11100 7936
rect 10968 7890 11020 7896
rect 11072 6866 11100 7908
rect 11060 6860 11112 6866
rect 11060 6802 11112 6808
rect 11072 5914 11100 6802
rect 11060 5908 11112 5914
rect 11060 5850 11112 5856
rect 10888 5766 11008 5794
rect 10784 5296 10836 5302
rect 10784 5238 10836 5244
rect 10796 4486 10824 5238
rect 10980 5030 11008 5766
rect 10968 5024 11020 5030
rect 10968 4966 11020 4972
rect 10980 4554 11008 4966
rect 11164 4593 11192 8774
rect 11256 8634 11284 9007
rect 11348 8634 11376 11086
rect 11532 10742 11560 11630
rect 11612 11144 11664 11150
rect 11612 11086 11664 11092
rect 11624 10810 11652 11086
rect 11612 10804 11664 10810
rect 11612 10746 11664 10752
rect 11520 10736 11572 10742
rect 11520 10678 11572 10684
rect 11808 9897 11836 12804
rect 11888 12786 11940 12792
rect 11888 12436 11940 12442
rect 11888 12378 11940 12384
rect 11900 9994 11928 12378
rect 11992 12288 12020 13126
rect 12176 12442 12204 14010
rect 12164 12436 12216 12442
rect 12164 12378 12216 12384
rect 12164 12300 12216 12306
rect 11992 12260 12164 12288
rect 12164 12242 12216 12248
rect 11980 12164 12032 12170
rect 11980 12106 12032 12112
rect 11992 11937 12020 12106
rect 11978 11928 12034 11937
rect 11978 11863 12034 11872
rect 12268 11642 12296 15524
rect 12530 15464 12586 15473
rect 12530 15399 12586 15408
rect 12440 14272 12492 14278
rect 12440 14214 12492 14220
rect 12346 13968 12402 13977
rect 12452 13938 12480 14214
rect 12346 13903 12402 13912
rect 12440 13932 12492 13938
rect 12360 12458 12388 13903
rect 12440 13874 12492 13880
rect 12438 13832 12494 13841
rect 12438 13767 12494 13776
rect 12452 12782 12480 13767
rect 12440 12776 12492 12782
rect 12440 12718 12492 12724
rect 12544 12730 12572 15399
rect 13004 15348 13032 16186
rect 13096 16046 13124 16390
rect 13188 16250 13216 19306
rect 13176 16244 13228 16250
rect 13176 16186 13228 16192
rect 13084 16040 13136 16046
rect 13084 15982 13136 15988
rect 13174 16008 13230 16017
rect 13174 15943 13230 15952
rect 13004 15320 13124 15348
rect 12679 15260 12987 15269
rect 12679 15258 12685 15260
rect 12741 15258 12765 15260
rect 12821 15258 12845 15260
rect 12901 15258 12925 15260
rect 12981 15258 12987 15260
rect 12741 15206 12743 15258
rect 12923 15206 12925 15258
rect 12679 15204 12685 15206
rect 12741 15204 12765 15206
rect 12821 15204 12845 15206
rect 12901 15204 12925 15206
rect 12981 15204 12987 15206
rect 12679 15195 12987 15204
rect 13096 14618 13124 15320
rect 13188 14958 13216 15943
rect 13176 14952 13228 14958
rect 13176 14894 13228 14900
rect 13084 14612 13136 14618
rect 13084 14554 13136 14560
rect 13084 14272 13136 14278
rect 13084 14214 13136 14220
rect 12679 14172 12987 14181
rect 12679 14170 12685 14172
rect 12741 14170 12765 14172
rect 12821 14170 12845 14172
rect 12901 14170 12925 14172
rect 12981 14170 12987 14172
rect 12741 14118 12743 14170
rect 12923 14118 12925 14170
rect 12679 14116 12685 14118
rect 12741 14116 12765 14118
rect 12821 14116 12845 14118
rect 12901 14116 12925 14118
rect 12981 14116 12987 14118
rect 12679 14107 12987 14116
rect 12716 13932 12768 13938
rect 12716 13874 12768 13880
rect 12728 13530 12756 13874
rect 13096 13870 13124 14214
rect 13084 13864 13136 13870
rect 13084 13806 13136 13812
rect 13084 13728 13136 13734
rect 13084 13670 13136 13676
rect 12716 13524 12768 13530
rect 12716 13466 12768 13472
rect 12679 13084 12987 13093
rect 12679 13082 12685 13084
rect 12741 13082 12765 13084
rect 12821 13082 12845 13084
rect 12901 13082 12925 13084
rect 12981 13082 12987 13084
rect 12741 13030 12743 13082
rect 12923 13030 12925 13082
rect 12679 13028 12685 13030
rect 12741 13028 12765 13030
rect 12821 13028 12845 13030
rect 12901 13028 12925 13030
rect 12981 13028 12987 13030
rect 12679 13019 12987 13028
rect 12992 12776 13044 12782
rect 12544 12702 12664 12730
rect 12992 12718 13044 12724
rect 12532 12640 12584 12646
rect 12532 12582 12584 12588
rect 12360 12442 12480 12458
rect 12360 12436 12492 12442
rect 12360 12430 12440 12436
rect 12440 12378 12492 12384
rect 12544 12374 12572 12582
rect 12348 12368 12400 12374
rect 12532 12368 12584 12374
rect 12400 12316 12480 12322
rect 12348 12310 12480 12316
rect 12532 12310 12584 12316
rect 12360 12294 12480 12310
rect 12452 11898 12480 12294
rect 12636 12084 12664 12702
rect 13004 12306 13032 12718
rect 12992 12300 13044 12306
rect 12992 12242 13044 12248
rect 13096 12238 13124 13670
rect 13280 12434 13308 20590
rect 13360 20460 13412 20466
rect 13360 20402 13412 20408
rect 13372 20058 13400 20402
rect 13452 20392 13504 20398
rect 13452 20334 13504 20340
rect 13360 20052 13412 20058
rect 13360 19994 13412 20000
rect 13464 19514 13492 20334
rect 13452 19508 13504 19514
rect 13452 19450 13504 19456
rect 13358 19408 13414 19417
rect 13358 19343 13414 19352
rect 13452 19372 13504 19378
rect 13372 18698 13400 19343
rect 13452 19314 13504 19320
rect 13360 18692 13412 18698
rect 13360 18634 13412 18640
rect 13372 16697 13400 18634
rect 13464 18358 13492 19314
rect 13452 18352 13504 18358
rect 13452 18294 13504 18300
rect 13452 18216 13504 18222
rect 13452 18158 13504 18164
rect 13464 17202 13492 18158
rect 13452 17196 13504 17202
rect 13452 17138 13504 17144
rect 13358 16688 13414 16697
rect 13358 16623 13414 16632
rect 13360 16584 13412 16590
rect 13360 16526 13412 16532
rect 13372 16114 13400 16526
rect 13452 16244 13504 16250
rect 13452 16186 13504 16192
rect 13360 16108 13412 16114
rect 13360 16050 13412 16056
rect 13464 15450 13492 16186
rect 13372 15422 13492 15450
rect 13372 14074 13400 15422
rect 13452 15360 13504 15366
rect 13452 15302 13504 15308
rect 13464 14278 13492 15302
rect 13452 14272 13504 14278
rect 13452 14214 13504 14220
rect 13360 14068 13412 14074
rect 13360 14010 13412 14016
rect 13360 13184 13412 13190
rect 13360 13126 13412 13132
rect 13188 12406 13308 12434
rect 13084 12232 13136 12238
rect 13084 12174 13136 12180
rect 12544 12056 12664 12084
rect 12440 11892 12492 11898
rect 12440 11834 12492 11840
rect 12438 11792 12494 11801
rect 12438 11727 12494 11736
rect 12544 11744 12572 12056
rect 12679 11996 12987 12005
rect 12679 11994 12685 11996
rect 12741 11994 12765 11996
rect 12821 11994 12845 11996
rect 12901 11994 12925 11996
rect 12981 11994 12987 11996
rect 12741 11942 12743 11994
rect 12923 11942 12925 11994
rect 12679 11940 12685 11942
rect 12741 11940 12765 11942
rect 12821 11940 12845 11942
rect 12901 11940 12925 11942
rect 12981 11940 12987 11942
rect 12679 11931 12987 11940
rect 12716 11892 12768 11898
rect 12716 11834 12768 11840
rect 12624 11756 12676 11762
rect 12176 11614 12296 11642
rect 11980 11552 12032 11558
rect 12032 11500 12112 11506
rect 11980 11494 12112 11500
rect 11992 11478 12112 11494
rect 12084 11286 12112 11478
rect 12072 11280 12124 11286
rect 12072 11222 12124 11228
rect 12176 11098 12204 11614
rect 12452 11354 12480 11727
rect 12544 11716 12624 11744
rect 12624 11698 12676 11704
rect 12440 11348 12492 11354
rect 12440 11290 12492 11296
rect 12346 11248 12402 11257
rect 12346 11183 12402 11192
rect 12360 11150 12388 11183
rect 12348 11144 12400 11150
rect 12176 11070 12296 11098
rect 12348 11086 12400 11092
rect 12164 10668 12216 10674
rect 12164 10610 12216 10616
rect 11980 10260 12032 10266
rect 11980 10202 12032 10208
rect 11888 9988 11940 9994
rect 11888 9930 11940 9936
rect 11794 9888 11850 9897
rect 11794 9823 11850 9832
rect 11808 9674 11836 9823
rect 11716 9646 11836 9674
rect 11428 9512 11480 9518
rect 11428 9454 11480 9460
rect 11440 9042 11468 9454
rect 11428 9036 11480 9042
rect 11428 8978 11480 8984
rect 11244 8628 11296 8634
rect 11244 8570 11296 8576
rect 11336 8628 11388 8634
rect 11336 8570 11388 8576
rect 11336 8084 11388 8090
rect 11336 8026 11388 8032
rect 11348 6730 11376 8026
rect 11336 6724 11388 6730
rect 11336 6666 11388 6672
rect 11440 6322 11468 8978
rect 11428 6316 11480 6322
rect 11428 6258 11480 6264
rect 11612 6112 11664 6118
rect 11612 6054 11664 6060
rect 11624 5914 11652 6054
rect 11612 5908 11664 5914
rect 11612 5850 11664 5856
rect 11716 5710 11744 9646
rect 11796 7812 11848 7818
rect 11796 7754 11848 7760
rect 11808 7478 11836 7754
rect 11888 7744 11940 7750
rect 11888 7686 11940 7692
rect 11796 7472 11848 7478
rect 11796 7414 11848 7420
rect 11900 7342 11928 7686
rect 11888 7336 11940 7342
rect 11888 7278 11940 7284
rect 11704 5704 11756 5710
rect 11704 5646 11756 5652
rect 11610 5536 11666 5545
rect 11610 5471 11666 5480
rect 11426 4992 11482 5001
rect 11426 4927 11482 4936
rect 11244 4752 11296 4758
rect 11244 4694 11296 4700
rect 11150 4584 11206 4593
rect 10968 4548 11020 4554
rect 10968 4490 11020 4496
rect 11060 4548 11112 4554
rect 11150 4519 11206 4528
rect 11060 4490 11112 4496
rect 10784 4480 10836 4486
rect 10784 4422 10836 4428
rect 10692 4140 10744 4146
rect 10692 4082 10744 4088
rect 10600 3936 10652 3942
rect 10600 3878 10652 3884
rect 10324 3392 10376 3398
rect 10324 3334 10376 3340
rect 10416 3392 10468 3398
rect 10416 3334 10468 3340
rect 10230 2544 10286 2553
rect 10230 2479 10286 2488
rect 10244 2378 10272 2479
rect 10232 2372 10284 2378
rect 10232 2314 10284 2320
rect 10100 1992 10180 2020
rect 10048 1974 10100 1980
rect 10048 1896 10100 1902
rect 9954 1864 10010 1873
rect 9680 1828 9732 1834
rect 10100 1856 10272 1884
rect 10048 1838 10100 1844
rect 9954 1799 9956 1808
rect 9680 1770 9732 1776
rect 10008 1799 10010 1808
rect 9956 1770 10008 1776
rect 10244 1737 10272 1856
rect 10230 1728 10286 1737
rect 9747 1660 10055 1669
rect 10230 1663 10286 1672
rect 9747 1658 9753 1660
rect 9809 1658 9833 1660
rect 9889 1658 9913 1660
rect 9969 1658 9993 1660
rect 10049 1658 10055 1660
rect 9809 1606 9811 1658
rect 9991 1606 9993 1658
rect 9747 1604 9753 1606
rect 9809 1604 9833 1606
rect 9889 1604 9913 1606
rect 9969 1604 9993 1606
rect 10049 1604 10055 1606
rect 9747 1595 10055 1604
rect 9496 1556 9548 1562
rect 9600 1550 9720 1578
rect 9496 1498 9548 1504
rect 9508 1306 9536 1498
rect 9692 1408 9720 1550
rect 9692 1380 9870 1408
rect 9632 1320 9688 1329
rect 9508 1278 9632 1306
rect 9632 1255 9688 1264
rect 9842 1204 9870 1380
rect 10244 1358 10272 1663
rect 9956 1352 10008 1358
rect 10232 1352 10284 1358
rect 9956 1294 10008 1300
rect 10046 1320 10102 1329
rect 9600 1176 9870 1204
rect 9218 54 9444 82
rect 9494 82 9550 160
rect 9600 82 9628 1176
rect 9968 898 9996 1294
rect 10232 1294 10284 1300
rect 10046 1255 10102 1264
rect 9876 870 9996 898
rect 9876 814 9904 870
rect 9864 808 9916 814
rect 9864 750 9916 756
rect 9956 808 10008 814
rect 9956 750 10008 756
rect 9494 54 9628 82
rect 9770 82 9826 160
rect 9968 82 9996 750
rect 10060 160 10088 1255
rect 10336 746 10364 3334
rect 10428 3058 10456 3334
rect 10416 3052 10468 3058
rect 10416 2994 10468 3000
rect 10612 2774 10640 3878
rect 10796 3534 10824 4422
rect 11072 4078 11100 4490
rect 11164 4214 11192 4519
rect 11256 4214 11284 4694
rect 11440 4622 11468 4927
rect 11624 4622 11652 5471
rect 11796 5024 11848 5030
rect 11796 4966 11848 4972
rect 11428 4616 11480 4622
rect 11334 4584 11390 4593
rect 11428 4558 11480 4564
rect 11612 4616 11664 4622
rect 11612 4558 11664 4564
rect 11334 4519 11390 4528
rect 11348 4486 11376 4519
rect 11336 4480 11388 4486
rect 11336 4422 11388 4428
rect 11428 4480 11480 4486
rect 11428 4422 11480 4428
rect 11152 4208 11204 4214
rect 11152 4150 11204 4156
rect 11244 4208 11296 4214
rect 11244 4150 11296 4156
rect 11060 4072 11112 4078
rect 10874 4040 10930 4049
rect 11060 4014 11112 4020
rect 10874 3975 10930 3984
rect 10784 3528 10836 3534
rect 10784 3470 10836 3476
rect 10888 3126 10916 3975
rect 11152 3936 11204 3942
rect 11152 3878 11204 3884
rect 10692 3120 10744 3126
rect 10692 3062 10744 3068
rect 10876 3120 10928 3126
rect 10876 3062 10928 3068
rect 10520 2746 10640 2774
rect 10520 2530 10548 2746
rect 10428 2502 10548 2530
rect 10324 740 10376 746
rect 10324 682 10376 688
rect 9770 54 9996 82
rect 8942 -300 8998 54
rect 9218 -300 9274 54
rect 9494 -300 9550 54
rect 9770 -300 9826 54
rect 10046 -300 10102 160
rect 10322 82 10378 160
rect 10428 82 10456 2502
rect 10704 2446 10732 3062
rect 10968 2848 11020 2854
rect 10888 2796 10968 2802
rect 10888 2790 11020 2796
rect 10888 2774 11008 2790
rect 10692 2440 10744 2446
rect 10692 2382 10744 2388
rect 10508 2372 10560 2378
rect 10508 2314 10560 2320
rect 10520 2122 10548 2314
rect 10520 2106 10824 2122
rect 10520 2100 10836 2106
rect 10520 2094 10784 2100
rect 10784 2042 10836 2048
rect 10784 1828 10836 1834
rect 10784 1770 10836 1776
rect 10508 1760 10560 1766
rect 10508 1702 10560 1708
rect 10520 898 10548 1702
rect 10520 870 10640 898
rect 10612 160 10640 870
rect 10796 814 10824 1770
rect 10784 808 10836 814
rect 10784 750 10836 756
rect 10888 160 10916 2774
rect 10968 2508 11020 2514
rect 10968 2450 11020 2456
rect 10980 1562 11008 2450
rect 11060 2304 11112 2310
rect 11164 2281 11192 3878
rect 11256 3534 11284 4150
rect 11244 3528 11296 3534
rect 11244 3470 11296 3476
rect 11242 2408 11298 2417
rect 11242 2343 11298 2352
rect 11256 2310 11284 2343
rect 11244 2304 11296 2310
rect 11060 2246 11112 2252
rect 11150 2272 11206 2281
rect 10968 1556 11020 1562
rect 10968 1498 11020 1504
rect 11072 1465 11100 2246
rect 11244 2246 11296 2252
rect 11150 2207 11206 2216
rect 11348 2106 11376 4422
rect 11440 4282 11468 4422
rect 11428 4276 11480 4282
rect 11428 4218 11480 4224
rect 11520 4072 11572 4078
rect 11572 4049 11652 4060
rect 11572 4040 11666 4049
rect 11572 4032 11610 4040
rect 11520 4014 11572 4020
rect 11532 3534 11560 4014
rect 11610 3975 11666 3984
rect 11520 3528 11572 3534
rect 11520 3470 11572 3476
rect 11532 3058 11560 3470
rect 11520 3052 11572 3058
rect 11520 2994 11572 3000
rect 11336 2100 11388 2106
rect 11336 2042 11388 2048
rect 11532 1970 11560 2994
rect 11808 2961 11836 4966
rect 11888 4684 11940 4690
rect 11888 4626 11940 4632
rect 11900 3738 11928 4626
rect 11888 3732 11940 3738
rect 11888 3674 11940 3680
rect 11794 2952 11850 2961
rect 11794 2887 11850 2896
rect 11992 2774 12020 10202
rect 12072 9988 12124 9994
rect 12072 9930 12124 9936
rect 12084 7750 12112 9930
rect 12176 9625 12204 10610
rect 12162 9616 12218 9625
rect 12162 9551 12218 9560
rect 12176 8090 12204 9551
rect 12164 8084 12216 8090
rect 12164 8026 12216 8032
rect 12072 7744 12124 7750
rect 12072 7686 12124 7692
rect 12072 7472 12124 7478
rect 12072 7414 12124 7420
rect 12164 7472 12216 7478
rect 12164 7414 12216 7420
rect 12084 7002 12112 7414
rect 12072 6996 12124 7002
rect 12072 6938 12124 6944
rect 12072 6792 12124 6798
rect 12072 6734 12124 6740
rect 12084 6186 12112 6734
rect 12072 6180 12124 6186
rect 12072 6122 12124 6128
rect 12176 3534 12204 7414
rect 12164 3528 12216 3534
rect 12164 3470 12216 3476
rect 12176 3369 12204 3470
rect 12162 3360 12218 3369
rect 12162 3295 12218 3304
rect 12176 3194 12204 3295
rect 12164 3188 12216 3194
rect 12164 3130 12216 3136
rect 12268 2774 12296 11070
rect 12728 11064 12756 11834
rect 13096 11830 13124 12174
rect 13084 11824 13136 11830
rect 13084 11766 13136 11772
rect 12900 11552 12952 11558
rect 12900 11494 12952 11500
rect 12912 11150 12940 11494
rect 12900 11144 12952 11150
rect 12900 11086 12952 11092
rect 12544 11036 12756 11064
rect 12544 10146 12572 11036
rect 12679 10908 12987 10917
rect 12679 10906 12685 10908
rect 12741 10906 12765 10908
rect 12821 10906 12845 10908
rect 12901 10906 12925 10908
rect 12981 10906 12987 10908
rect 12741 10854 12743 10906
rect 12923 10854 12925 10906
rect 12679 10852 12685 10854
rect 12741 10852 12765 10854
rect 12821 10852 12845 10854
rect 12901 10852 12925 10854
rect 12981 10852 12987 10854
rect 12679 10843 12987 10852
rect 12440 10124 12492 10130
rect 12544 10118 12664 10146
rect 12440 10066 12492 10072
rect 12452 9178 12480 10066
rect 12636 10062 12664 10118
rect 12624 10056 12676 10062
rect 12624 9998 12676 10004
rect 12532 9988 12584 9994
rect 12532 9930 12584 9936
rect 13084 9988 13136 9994
rect 13084 9930 13136 9936
rect 12544 9722 12572 9930
rect 12679 9820 12987 9829
rect 12679 9818 12685 9820
rect 12741 9818 12765 9820
rect 12821 9818 12845 9820
rect 12901 9818 12925 9820
rect 12981 9818 12987 9820
rect 12741 9766 12743 9818
rect 12923 9766 12925 9818
rect 12679 9764 12685 9766
rect 12741 9764 12765 9766
rect 12821 9764 12845 9766
rect 12901 9764 12925 9766
rect 12981 9764 12987 9766
rect 12679 9755 12987 9764
rect 12532 9716 12584 9722
rect 12532 9658 12584 9664
rect 12440 9172 12492 9178
rect 12440 9114 12492 9120
rect 12348 8968 12400 8974
rect 12348 8910 12400 8916
rect 12360 7478 12388 8910
rect 12679 8732 12987 8741
rect 12679 8730 12685 8732
rect 12741 8730 12765 8732
rect 12821 8730 12845 8732
rect 12901 8730 12925 8732
rect 12981 8730 12987 8732
rect 12741 8678 12743 8730
rect 12923 8678 12925 8730
rect 12679 8676 12685 8678
rect 12741 8676 12765 8678
rect 12821 8676 12845 8678
rect 12901 8676 12925 8678
rect 12981 8676 12987 8678
rect 12679 8667 12987 8676
rect 13096 7818 13124 9930
rect 13084 7812 13136 7818
rect 13084 7754 13136 7760
rect 12532 7744 12584 7750
rect 12532 7686 12584 7692
rect 12348 7472 12400 7478
rect 12348 7414 12400 7420
rect 12440 7472 12492 7478
rect 12440 7414 12492 7420
rect 12452 7002 12480 7414
rect 12440 6996 12492 7002
rect 12440 6938 12492 6944
rect 12348 6792 12400 6798
rect 12348 6734 12400 6740
rect 12360 6390 12388 6734
rect 12452 6633 12480 6938
rect 12438 6624 12494 6633
rect 12438 6559 12494 6568
rect 12348 6384 12400 6390
rect 12348 6326 12400 6332
rect 12544 5234 12572 7686
rect 12679 7644 12987 7653
rect 12679 7642 12685 7644
rect 12741 7642 12765 7644
rect 12821 7642 12845 7644
rect 12901 7642 12925 7644
rect 12981 7642 12987 7644
rect 12741 7590 12743 7642
rect 12923 7590 12925 7642
rect 12679 7588 12685 7590
rect 12741 7588 12765 7590
rect 12821 7588 12845 7590
rect 12901 7588 12925 7590
rect 12981 7588 12987 7590
rect 12679 7579 12987 7588
rect 12992 7472 13044 7478
rect 12992 7414 13044 7420
rect 13004 7290 13032 7414
rect 13096 7410 13124 7754
rect 13084 7404 13136 7410
rect 13084 7346 13136 7352
rect 13004 7262 13124 7290
rect 12808 6792 12860 6798
rect 12806 6760 12808 6769
rect 12860 6760 12862 6769
rect 12806 6695 12862 6704
rect 12679 6556 12987 6565
rect 12679 6554 12685 6556
rect 12741 6554 12765 6556
rect 12821 6554 12845 6556
rect 12901 6554 12925 6556
rect 12981 6554 12987 6556
rect 12741 6502 12743 6554
rect 12923 6502 12925 6554
rect 12679 6500 12685 6502
rect 12741 6500 12765 6502
rect 12821 6500 12845 6502
rect 12901 6500 12925 6502
rect 12981 6500 12987 6502
rect 12679 6491 12987 6500
rect 12679 5468 12987 5477
rect 12679 5466 12685 5468
rect 12741 5466 12765 5468
rect 12821 5466 12845 5468
rect 12901 5466 12925 5468
rect 12981 5466 12987 5468
rect 12741 5414 12743 5466
rect 12923 5414 12925 5466
rect 12679 5412 12685 5414
rect 12741 5412 12765 5414
rect 12821 5412 12845 5414
rect 12901 5412 12925 5414
rect 12981 5412 12987 5414
rect 12679 5403 12987 5412
rect 12532 5228 12584 5234
rect 12532 5170 12584 5176
rect 13096 5166 13124 7262
rect 12440 5160 12492 5166
rect 12440 5102 12492 5108
rect 13084 5160 13136 5166
rect 13084 5102 13136 5108
rect 12452 3942 12480 5102
rect 12624 5092 12676 5098
rect 12624 5034 12676 5040
rect 12636 4826 12664 5034
rect 12624 4820 12676 4826
rect 12624 4762 12676 4768
rect 12532 4616 12584 4622
rect 12532 4558 12584 4564
rect 12544 4282 12572 4558
rect 12679 4380 12987 4389
rect 12679 4378 12685 4380
rect 12741 4378 12765 4380
rect 12821 4378 12845 4380
rect 12901 4378 12925 4380
rect 12981 4378 12987 4380
rect 12741 4326 12743 4378
rect 12923 4326 12925 4378
rect 12679 4324 12685 4326
rect 12741 4324 12765 4326
rect 12821 4324 12845 4326
rect 12901 4324 12925 4326
rect 12981 4324 12987 4326
rect 12679 4315 12987 4324
rect 12532 4276 12584 4282
rect 12532 4218 12584 4224
rect 12990 4176 13046 4185
rect 12990 4111 13046 4120
rect 13004 3942 13032 4111
rect 12440 3936 12492 3942
rect 12440 3878 12492 3884
rect 12992 3936 13044 3942
rect 12992 3878 13044 3884
rect 13004 3738 13032 3878
rect 12992 3732 13044 3738
rect 12992 3674 13044 3680
rect 12679 3292 12987 3301
rect 12679 3290 12685 3292
rect 12741 3290 12765 3292
rect 12821 3290 12845 3292
rect 12901 3290 12925 3292
rect 12981 3290 12987 3292
rect 12741 3238 12743 3290
rect 12923 3238 12925 3290
rect 12679 3236 12685 3238
rect 12741 3236 12765 3238
rect 12821 3236 12845 3238
rect 12901 3236 12925 3238
rect 12981 3236 12987 3238
rect 12530 3224 12586 3233
rect 12679 3227 12987 3236
rect 12530 3159 12586 3168
rect 12544 2990 12572 3159
rect 12532 2984 12584 2990
rect 12532 2926 12584 2932
rect 12348 2848 12400 2854
rect 12348 2790 12400 2796
rect 11992 2746 12112 2774
rect 11794 2680 11850 2689
rect 11794 2615 11850 2624
rect 11808 2378 11836 2615
rect 11886 2408 11942 2417
rect 11796 2372 11848 2378
rect 11886 2343 11942 2352
rect 11980 2372 12032 2378
rect 11796 2314 11848 2320
rect 11612 2032 11664 2038
rect 11612 1974 11664 1980
rect 11520 1964 11572 1970
rect 11520 1906 11572 1912
rect 11532 1737 11560 1906
rect 11518 1728 11574 1737
rect 11518 1663 11574 1672
rect 11624 1562 11652 1974
rect 11808 1850 11836 2314
rect 11900 2038 11928 2343
rect 11980 2314 12032 2320
rect 11992 2281 12020 2314
rect 11978 2272 12034 2281
rect 11978 2207 12034 2216
rect 11888 2032 11940 2038
rect 11888 1974 11940 1980
rect 11716 1822 11836 1850
rect 11244 1556 11296 1562
rect 11244 1498 11296 1504
rect 11612 1556 11664 1562
rect 11612 1498 11664 1504
rect 11152 1488 11204 1494
rect 11058 1456 11114 1465
rect 11152 1430 11204 1436
rect 11058 1391 11114 1400
rect 11060 1352 11112 1358
rect 11058 1320 11060 1329
rect 11112 1320 11114 1329
rect 11058 1255 11114 1264
rect 11164 160 11192 1430
rect 11256 610 11284 1498
rect 11716 1358 11744 1822
rect 11796 1760 11848 1766
rect 11796 1702 11848 1708
rect 11980 1760 12032 1766
rect 11980 1702 12032 1708
rect 11808 1358 11836 1702
rect 11704 1352 11756 1358
rect 11704 1294 11756 1300
rect 11796 1352 11848 1358
rect 11796 1294 11848 1300
rect 11520 1216 11572 1222
rect 11518 1184 11520 1193
rect 11572 1184 11574 1193
rect 11518 1119 11574 1128
rect 11992 898 12020 1702
rect 12084 1426 12112 2746
rect 12176 2746 12296 2774
rect 12072 1420 12124 1426
rect 12072 1362 12124 1368
rect 12176 1340 12204 2746
rect 12360 2514 12388 2790
rect 12348 2508 12400 2514
rect 12348 2450 12400 2456
rect 13188 2378 13216 12406
rect 13268 12232 13320 12238
rect 13268 12174 13320 12180
rect 13280 11898 13308 12174
rect 13268 11892 13320 11898
rect 13268 11834 13320 11840
rect 13268 11688 13320 11694
rect 13268 11630 13320 11636
rect 13280 11014 13308 11630
rect 13268 11008 13320 11014
rect 13268 10950 13320 10956
rect 13268 10532 13320 10538
rect 13268 10474 13320 10480
rect 13280 9926 13308 10474
rect 13372 10062 13400 13126
rect 13464 10538 13492 14214
rect 13556 13734 13584 20590
rect 13648 16250 13676 28494
rect 13636 16244 13688 16250
rect 13636 16186 13688 16192
rect 13636 16108 13688 16114
rect 13636 16050 13688 16056
rect 13648 15706 13676 16050
rect 13636 15700 13688 15706
rect 13636 15642 13688 15648
rect 13544 13728 13596 13734
rect 13544 13670 13596 13676
rect 13544 12640 13596 12646
rect 13544 12582 13596 12588
rect 13556 12209 13584 12582
rect 13740 12434 13768 30552
rect 13832 30190 13860 31078
rect 13820 30184 13872 30190
rect 13820 30126 13872 30132
rect 13924 29102 13952 31198
rect 13820 29096 13872 29102
rect 13820 29038 13872 29044
rect 13912 29096 13964 29102
rect 13912 29038 13964 29044
rect 13832 28762 13860 29038
rect 13820 28756 13872 28762
rect 13820 28698 13872 28704
rect 13924 28558 13952 29038
rect 13912 28552 13964 28558
rect 13912 28494 13964 28500
rect 13820 28484 13872 28490
rect 13820 28426 13872 28432
rect 13832 27062 13860 28426
rect 13912 28008 13964 28014
rect 13912 27950 13964 27956
rect 13820 27056 13872 27062
rect 13820 26998 13872 27004
rect 13820 26240 13872 26246
rect 13820 26182 13872 26188
rect 13832 26042 13860 26182
rect 13820 26036 13872 26042
rect 13820 25978 13872 25984
rect 13832 25906 13860 25978
rect 13820 25900 13872 25906
rect 13820 25842 13872 25848
rect 13820 25764 13872 25770
rect 13924 25752 13952 27950
rect 13872 25724 13952 25752
rect 13820 25706 13872 25712
rect 13820 25288 13872 25294
rect 14016 25265 14044 31726
rect 14225 31498 14253 31726
rect 14200 31470 14253 31498
rect 14096 31272 14148 31278
rect 14094 31240 14096 31249
rect 14148 31240 14150 31249
rect 14094 31175 14150 31184
rect 14096 29096 14148 29102
rect 14096 29038 14148 29044
rect 14108 28218 14136 29038
rect 14200 28558 14228 31470
rect 14292 30598 14320 32166
rect 14372 31816 14424 31822
rect 14372 31758 14424 31764
rect 14280 30592 14332 30598
rect 14280 30534 14332 30540
rect 14280 30320 14332 30326
rect 14280 30262 14332 30268
rect 14292 29102 14320 30262
rect 14280 29096 14332 29102
rect 14280 29038 14332 29044
rect 14384 28994 14412 31758
rect 14476 31754 14504 32846
rect 14476 31726 14596 31754
rect 14464 31680 14516 31686
rect 14464 31622 14516 31628
rect 14476 31482 14504 31622
rect 14464 31476 14516 31482
rect 14464 31418 14516 31424
rect 14568 31414 14596 31726
rect 14556 31408 14608 31414
rect 14556 31350 14608 31356
rect 14464 31136 14516 31142
rect 14464 31078 14516 31084
rect 14476 30326 14504 31078
rect 14464 30320 14516 30326
rect 14464 30262 14516 30268
rect 14660 29753 14688 33390
rect 14740 32224 14792 32230
rect 14740 32166 14792 32172
rect 14752 31890 14780 32166
rect 14740 31884 14792 31890
rect 14740 31826 14792 31832
rect 14646 29744 14702 29753
rect 14646 29679 14702 29688
rect 14660 29073 14688 29679
rect 14646 29064 14702 29073
rect 14646 28999 14702 29008
rect 14292 28966 14412 28994
rect 14188 28552 14240 28558
rect 14188 28494 14240 28500
rect 14096 28212 14148 28218
rect 14096 28154 14148 28160
rect 14096 27464 14148 27470
rect 14094 27432 14096 27441
rect 14148 27432 14150 27441
rect 14094 27367 14150 27376
rect 14188 27396 14240 27402
rect 14188 27338 14240 27344
rect 14096 27328 14148 27334
rect 14096 27270 14148 27276
rect 13820 25230 13872 25236
rect 14002 25256 14058 25265
rect 13832 24886 13860 25230
rect 14002 25191 14058 25200
rect 14004 25152 14056 25158
rect 14004 25094 14056 25100
rect 13820 24880 13872 24886
rect 13820 24822 13872 24828
rect 13832 24070 13860 24822
rect 13912 24744 13964 24750
rect 13912 24686 13964 24692
rect 13820 24064 13872 24070
rect 13820 24006 13872 24012
rect 13820 23112 13872 23118
rect 13820 23054 13872 23060
rect 13832 22574 13860 23054
rect 13924 22574 13952 24686
rect 14016 23118 14044 25094
rect 14004 23112 14056 23118
rect 14004 23054 14056 23060
rect 14004 22976 14056 22982
rect 14004 22918 14056 22924
rect 13820 22568 13872 22574
rect 13820 22510 13872 22516
rect 13912 22568 13964 22574
rect 13912 22510 13964 22516
rect 13924 21690 13952 22510
rect 13912 21684 13964 21690
rect 13912 21626 13964 21632
rect 13924 20534 13952 21626
rect 13912 20528 13964 20534
rect 13912 20470 13964 20476
rect 13820 20460 13872 20466
rect 13820 20402 13872 20408
rect 13832 20369 13860 20402
rect 13818 20360 13874 20369
rect 13818 20295 13874 20304
rect 13832 20058 13860 20295
rect 13820 20052 13872 20058
rect 13820 19994 13872 20000
rect 13910 19816 13966 19825
rect 14016 19802 14044 22918
rect 13966 19774 14044 19802
rect 13910 19751 13966 19760
rect 13924 19334 13952 19751
rect 13832 19306 13952 19334
rect 13832 18630 13860 19306
rect 13820 18624 13872 18630
rect 13820 18566 13872 18572
rect 13912 18624 13964 18630
rect 13912 18566 13964 18572
rect 13832 17678 13860 18566
rect 13820 17672 13872 17678
rect 13820 17614 13872 17620
rect 13832 17241 13860 17614
rect 13818 17232 13874 17241
rect 13818 17167 13874 17176
rect 13832 12646 13860 17167
rect 13924 15366 13952 18566
rect 14108 16590 14136 27270
rect 14200 27130 14228 27338
rect 14188 27124 14240 27130
rect 14188 27066 14240 27072
rect 14186 26616 14242 26625
rect 14186 26551 14242 26560
rect 14200 26382 14228 26551
rect 14188 26376 14240 26382
rect 14188 26318 14240 26324
rect 14188 26240 14240 26246
rect 14292 26228 14320 28966
rect 14556 28960 14608 28966
rect 14556 28902 14608 28908
rect 14568 28558 14596 28902
rect 14556 28552 14608 28558
rect 14556 28494 14608 28500
rect 14372 28484 14424 28490
rect 14372 28426 14424 28432
rect 14240 26200 14320 26228
rect 14188 26182 14240 26188
rect 14280 24948 14332 24954
rect 14280 24890 14332 24896
rect 14188 24608 14240 24614
rect 14188 24550 14240 24556
rect 14200 22098 14228 24550
rect 14292 24274 14320 24890
rect 14280 24268 14332 24274
rect 14280 24210 14332 24216
rect 14280 24132 14332 24138
rect 14280 24074 14332 24080
rect 14188 22092 14240 22098
rect 14188 22034 14240 22040
rect 14188 21956 14240 21962
rect 14188 21898 14240 21904
rect 14200 21593 14228 21898
rect 14186 21584 14242 21593
rect 14186 21519 14242 21528
rect 14200 21010 14228 21519
rect 14188 21004 14240 21010
rect 14188 20946 14240 20952
rect 14186 20632 14242 20641
rect 14186 20567 14242 20576
rect 14096 16584 14148 16590
rect 14096 16526 14148 16532
rect 14108 16250 14136 16526
rect 14096 16244 14148 16250
rect 14096 16186 14148 16192
rect 14096 15496 14148 15502
rect 14096 15438 14148 15444
rect 13912 15360 13964 15366
rect 13912 15302 13964 15308
rect 13910 15192 13966 15201
rect 13910 15127 13966 15136
rect 13924 13938 13952 15127
rect 14108 14414 14136 15438
rect 14096 14408 14148 14414
rect 14096 14350 14148 14356
rect 13912 13932 13964 13938
rect 13912 13874 13964 13880
rect 14004 13932 14056 13938
rect 14004 13874 14056 13880
rect 13820 12640 13872 12646
rect 13820 12582 13872 12588
rect 13648 12406 13768 12434
rect 13542 12200 13598 12209
rect 13542 12135 13598 12144
rect 13544 11756 13596 11762
rect 13544 11698 13596 11704
rect 13556 10996 13584 11698
rect 13648 11098 13676 12406
rect 13924 11830 13952 13874
rect 14016 13530 14044 13874
rect 14004 13524 14056 13530
rect 14004 13466 14056 13472
rect 14004 13252 14056 13258
rect 14004 13194 14056 13200
rect 14016 12442 14044 13194
rect 14108 12764 14136 14350
rect 14200 14346 14228 20567
rect 14292 20398 14320 24074
rect 14384 20602 14412 28426
rect 14568 27441 14596 28494
rect 14554 27432 14610 27441
rect 14554 27367 14610 27376
rect 14568 27334 14596 27367
rect 14556 27328 14608 27334
rect 14556 27270 14608 27276
rect 14568 26450 14596 27270
rect 14556 26444 14608 26450
rect 14556 26386 14608 26392
rect 14464 25968 14516 25974
rect 14464 25910 14516 25916
rect 14476 24392 14504 25910
rect 14568 25906 14596 26386
rect 14752 25974 14780 31826
rect 14844 30870 14872 33390
rect 14936 32570 14964 35022
rect 15108 34944 15160 34950
rect 15108 34886 15160 34892
rect 15120 34406 15148 34886
rect 15108 34400 15160 34406
rect 15108 34342 15160 34348
rect 15120 33998 15148 34342
rect 15016 33992 15068 33998
rect 15016 33934 15068 33940
rect 15108 33992 15160 33998
rect 15108 33934 15160 33940
rect 15028 33017 15056 33934
rect 15108 33312 15160 33318
rect 15108 33254 15160 33260
rect 15014 33008 15070 33017
rect 15120 32978 15148 33254
rect 15212 33114 15240 35022
rect 15384 33856 15436 33862
rect 15384 33798 15436 33804
rect 15396 33538 15424 33798
rect 15304 33510 15424 33538
rect 15304 33454 15332 33510
rect 15292 33448 15344 33454
rect 15488 33436 15516 37810
rect 15612 37564 15920 37573
rect 15612 37562 15618 37564
rect 15674 37562 15698 37564
rect 15754 37562 15778 37564
rect 15834 37562 15858 37564
rect 15914 37562 15920 37564
rect 15674 37510 15676 37562
rect 15856 37510 15858 37562
rect 15612 37508 15618 37510
rect 15674 37508 15698 37510
rect 15754 37508 15778 37510
rect 15834 37508 15858 37510
rect 15914 37508 15920 37510
rect 15612 37499 15920 37508
rect 15612 36476 15920 36485
rect 15612 36474 15618 36476
rect 15674 36474 15698 36476
rect 15754 36474 15778 36476
rect 15834 36474 15858 36476
rect 15914 36474 15920 36476
rect 15674 36422 15676 36474
rect 15856 36422 15858 36474
rect 15612 36420 15618 36422
rect 15674 36420 15698 36422
rect 15754 36420 15778 36422
rect 15834 36420 15858 36422
rect 15914 36420 15920 36422
rect 15612 36411 15920 36420
rect 15612 35388 15920 35397
rect 15612 35386 15618 35388
rect 15674 35386 15698 35388
rect 15754 35386 15778 35388
rect 15834 35386 15858 35388
rect 15914 35386 15920 35388
rect 15674 35334 15676 35386
rect 15856 35334 15858 35386
rect 15612 35332 15618 35334
rect 15674 35332 15698 35334
rect 15754 35332 15778 35334
rect 15834 35332 15858 35334
rect 15914 35332 15920 35334
rect 15612 35323 15920 35332
rect 15612 34300 15920 34309
rect 15612 34298 15618 34300
rect 15674 34298 15698 34300
rect 15754 34298 15778 34300
rect 15834 34298 15858 34300
rect 15914 34298 15920 34300
rect 15674 34246 15676 34298
rect 15856 34246 15858 34298
rect 15612 34244 15618 34246
rect 15674 34244 15698 34246
rect 15754 34244 15778 34246
rect 15834 34244 15858 34246
rect 15914 34244 15920 34246
rect 15612 34235 15920 34244
rect 15936 34060 15988 34066
rect 15936 34002 15988 34008
rect 15568 33516 15620 33522
rect 15568 33458 15620 33464
rect 15292 33390 15344 33396
rect 15396 33408 15516 33436
rect 15200 33108 15252 33114
rect 15200 33050 15252 33056
rect 15014 32943 15070 32952
rect 15108 32972 15160 32978
rect 15108 32914 15160 32920
rect 15118 32858 15146 32914
rect 15292 32904 15344 32910
rect 15028 32830 15146 32858
rect 15290 32872 15292 32881
rect 15344 32872 15346 32881
rect 14924 32564 14976 32570
rect 14924 32506 14976 32512
rect 14924 31952 14976 31958
rect 14924 31894 14976 31900
rect 14832 30864 14884 30870
rect 14832 30806 14884 30812
rect 14936 30734 14964 31894
rect 14924 30728 14976 30734
rect 14924 30670 14976 30676
rect 14832 30592 14884 30598
rect 14832 30534 14884 30540
rect 14844 28014 14872 30534
rect 14936 30258 14964 30670
rect 15028 30394 15056 32830
rect 15290 32807 15346 32816
rect 15396 32756 15424 33408
rect 15580 33368 15608 33458
rect 15304 32728 15424 32756
rect 15488 33340 15608 33368
rect 15106 32464 15162 32473
rect 15162 32422 15240 32450
rect 15106 32399 15162 32408
rect 15212 31822 15240 32422
rect 15200 31816 15252 31822
rect 15200 31758 15252 31764
rect 15212 30870 15240 31758
rect 15108 30864 15160 30870
rect 15108 30806 15160 30812
rect 15200 30864 15252 30870
rect 15200 30806 15252 30812
rect 15120 30394 15148 30806
rect 15200 30728 15252 30734
rect 15200 30670 15252 30676
rect 15016 30388 15068 30394
rect 15016 30330 15068 30336
rect 15108 30388 15160 30394
rect 15108 30330 15160 30336
rect 14924 30252 14976 30258
rect 14924 30194 14976 30200
rect 14924 29776 14976 29782
rect 14924 29718 14976 29724
rect 14832 28008 14884 28014
rect 14832 27950 14884 27956
rect 14832 27872 14884 27878
rect 14832 27814 14884 27820
rect 14844 25974 14872 27814
rect 14740 25968 14792 25974
rect 14740 25910 14792 25916
rect 14832 25968 14884 25974
rect 14832 25910 14884 25916
rect 14556 25900 14608 25906
rect 14556 25842 14608 25848
rect 14936 25786 14964 29718
rect 15014 29064 15070 29073
rect 15014 28999 15070 29008
rect 15028 26790 15056 28999
rect 15212 28218 15240 30670
rect 15200 28212 15252 28218
rect 15200 28154 15252 28160
rect 15212 27674 15240 28154
rect 15200 27668 15252 27674
rect 15200 27610 15252 27616
rect 15304 27402 15332 32728
rect 15384 30252 15436 30258
rect 15488 30240 15516 33340
rect 15612 33212 15920 33221
rect 15612 33210 15618 33212
rect 15674 33210 15698 33212
rect 15754 33210 15778 33212
rect 15834 33210 15858 33212
rect 15914 33210 15920 33212
rect 15674 33158 15676 33210
rect 15856 33158 15858 33210
rect 15612 33156 15618 33158
rect 15674 33156 15698 33158
rect 15754 33156 15778 33158
rect 15834 33156 15858 33158
rect 15914 33156 15920 33158
rect 15612 33147 15920 33156
rect 15842 33008 15898 33017
rect 15842 32943 15844 32952
rect 15896 32943 15898 32952
rect 15844 32914 15896 32920
rect 15948 32910 15976 34002
rect 15936 32904 15988 32910
rect 15936 32846 15988 32852
rect 16120 32768 16172 32774
rect 16120 32710 16172 32716
rect 15612 32124 15920 32133
rect 15612 32122 15618 32124
rect 15674 32122 15698 32124
rect 15754 32122 15778 32124
rect 15834 32122 15858 32124
rect 15914 32122 15920 32124
rect 15674 32070 15676 32122
rect 15856 32070 15858 32122
rect 15612 32068 15618 32070
rect 15674 32068 15698 32070
rect 15754 32068 15778 32070
rect 15834 32068 15858 32070
rect 15914 32068 15920 32070
rect 15612 32059 15920 32068
rect 16028 32020 16080 32026
rect 16028 31962 16080 31968
rect 15936 31680 15988 31686
rect 15936 31622 15988 31628
rect 15612 31036 15920 31045
rect 15612 31034 15618 31036
rect 15674 31034 15698 31036
rect 15754 31034 15778 31036
rect 15834 31034 15858 31036
rect 15914 31034 15920 31036
rect 15674 30982 15676 31034
rect 15856 30982 15858 31034
rect 15612 30980 15618 30982
rect 15674 30980 15698 30982
rect 15754 30980 15778 30982
rect 15834 30980 15858 30982
rect 15914 30980 15920 30982
rect 15612 30971 15920 30980
rect 15948 30870 15976 31622
rect 15568 30864 15620 30870
rect 15568 30806 15620 30812
rect 15936 30864 15988 30870
rect 15936 30806 15988 30812
rect 15436 30212 15516 30240
rect 15384 30194 15436 30200
rect 15396 29238 15424 30194
rect 15580 30036 15608 30806
rect 15936 30184 15988 30190
rect 15936 30126 15988 30132
rect 15488 30008 15608 30036
rect 15488 29594 15516 30008
rect 15612 29948 15920 29957
rect 15612 29946 15618 29948
rect 15674 29946 15698 29948
rect 15754 29946 15778 29948
rect 15834 29946 15858 29948
rect 15914 29946 15920 29948
rect 15674 29894 15676 29946
rect 15856 29894 15858 29946
rect 15612 29892 15618 29894
rect 15674 29892 15698 29894
rect 15754 29892 15778 29894
rect 15834 29892 15858 29894
rect 15914 29892 15920 29894
rect 15612 29883 15920 29892
rect 15752 29776 15804 29782
rect 15658 29744 15714 29753
rect 15948 29730 15976 30126
rect 15804 29724 15976 29730
rect 15752 29718 15976 29724
rect 15764 29702 15976 29718
rect 15658 29679 15714 29688
rect 15672 29646 15700 29679
rect 15660 29640 15712 29646
rect 15488 29578 15608 29594
rect 15660 29582 15712 29588
rect 15488 29572 15620 29578
rect 15488 29566 15568 29572
rect 15568 29514 15620 29520
rect 15476 29504 15528 29510
rect 15476 29446 15528 29452
rect 15384 29232 15436 29238
rect 15384 29174 15436 29180
rect 15384 28416 15436 28422
rect 15384 28358 15436 28364
rect 15396 28014 15424 28358
rect 15384 28008 15436 28014
rect 15384 27950 15436 27956
rect 15488 27826 15516 29446
rect 15934 29336 15990 29345
rect 15934 29271 15990 29280
rect 15948 29034 15976 29271
rect 15936 29028 15988 29034
rect 15936 28970 15988 28976
rect 15612 28860 15920 28869
rect 15612 28858 15618 28860
rect 15674 28858 15698 28860
rect 15754 28858 15778 28860
rect 15834 28858 15858 28860
rect 15914 28858 15920 28860
rect 15674 28806 15676 28858
rect 15856 28806 15858 28858
rect 15612 28804 15618 28806
rect 15674 28804 15698 28806
rect 15754 28804 15778 28806
rect 15834 28804 15858 28806
rect 15914 28804 15920 28806
rect 15612 28795 15920 28804
rect 15948 28098 15976 28970
rect 15764 28082 15976 28098
rect 15752 28076 15976 28082
rect 15804 28070 15976 28076
rect 15752 28018 15804 28024
rect 15568 28008 15620 28014
rect 15568 27950 15620 27956
rect 15580 27878 15608 27950
rect 16040 27878 16068 31962
rect 16132 30734 16160 32710
rect 16120 30728 16172 30734
rect 16120 30670 16172 30676
rect 15396 27798 15516 27826
rect 15568 27872 15620 27878
rect 15568 27814 15620 27820
rect 16028 27872 16080 27878
rect 16028 27814 16080 27820
rect 15292 27396 15344 27402
rect 15292 27338 15344 27344
rect 15108 27328 15160 27334
rect 15108 27270 15160 27276
rect 15016 26784 15068 26790
rect 15016 26726 15068 26732
rect 14648 25764 14700 25770
rect 14648 25706 14700 25712
rect 14752 25758 14964 25786
rect 14660 25498 14688 25706
rect 14648 25492 14700 25498
rect 14648 25434 14700 25440
rect 14648 25152 14700 25158
rect 14648 25094 14700 25100
rect 14660 24818 14688 25094
rect 14648 24812 14700 24818
rect 14648 24754 14700 24760
rect 14556 24744 14608 24750
rect 14556 24686 14608 24692
rect 14752 24698 14780 25758
rect 14832 25696 14884 25702
rect 14832 25638 14884 25644
rect 14844 24818 14872 25638
rect 15120 25498 15148 27270
rect 15198 27024 15254 27033
rect 15254 26982 15332 27010
rect 15198 26959 15254 26968
rect 15304 26382 15332 26982
rect 15200 26376 15252 26382
rect 15200 26318 15252 26324
rect 15292 26376 15344 26382
rect 15292 26318 15344 26324
rect 15212 26042 15240 26318
rect 15200 26036 15252 26042
rect 15200 25978 15252 25984
rect 15108 25492 15160 25498
rect 15108 25434 15160 25440
rect 15016 25288 15068 25294
rect 14936 25248 15016 25276
rect 14832 24812 14884 24818
rect 14832 24754 14884 24760
rect 14568 24585 14596 24686
rect 14752 24670 14872 24698
rect 14554 24576 14610 24585
rect 14554 24511 14610 24520
rect 14476 24364 14596 24392
rect 14464 24268 14516 24274
rect 14464 24210 14516 24216
rect 14476 24070 14504 24210
rect 14464 24064 14516 24070
rect 14464 24006 14516 24012
rect 14476 23322 14504 24006
rect 14464 23316 14516 23322
rect 14464 23258 14516 23264
rect 14476 22681 14504 23258
rect 14462 22672 14518 22681
rect 14462 22607 14518 22616
rect 14464 22500 14516 22506
rect 14464 22442 14516 22448
rect 14476 22166 14504 22442
rect 14464 22160 14516 22166
rect 14464 22102 14516 22108
rect 14464 21548 14516 21554
rect 14464 21490 14516 21496
rect 14372 20596 14424 20602
rect 14372 20538 14424 20544
rect 14476 20466 14504 21490
rect 14568 21457 14596 24364
rect 14648 23520 14700 23526
rect 14648 23462 14700 23468
rect 14660 21554 14688 23462
rect 14844 23118 14872 24670
rect 14936 24614 14964 25248
rect 15016 25230 15068 25236
rect 15108 25288 15160 25294
rect 15108 25230 15160 25236
rect 15396 25242 15424 27798
rect 15612 27772 15920 27781
rect 15612 27770 15618 27772
rect 15674 27770 15698 27772
rect 15754 27770 15778 27772
rect 15834 27770 15858 27772
rect 15914 27770 15920 27772
rect 15674 27718 15676 27770
rect 15856 27718 15858 27770
rect 15612 27716 15618 27718
rect 15674 27716 15698 27718
rect 15754 27716 15778 27718
rect 15834 27716 15858 27718
rect 15914 27716 15920 27718
rect 15612 27707 15920 27716
rect 16028 27396 16080 27402
rect 16028 27338 16080 27344
rect 15936 27056 15988 27062
rect 15936 26998 15988 27004
rect 15612 26684 15920 26693
rect 15612 26682 15618 26684
rect 15674 26682 15698 26684
rect 15754 26682 15778 26684
rect 15834 26682 15858 26684
rect 15914 26682 15920 26684
rect 15674 26630 15676 26682
rect 15856 26630 15858 26682
rect 15612 26628 15618 26630
rect 15674 26628 15698 26630
rect 15754 26628 15778 26630
rect 15834 26628 15858 26630
rect 15914 26628 15920 26630
rect 15612 26619 15920 26628
rect 15476 26240 15528 26246
rect 15476 26182 15528 26188
rect 15488 25362 15516 26182
rect 15612 25596 15920 25605
rect 15612 25594 15618 25596
rect 15674 25594 15698 25596
rect 15754 25594 15778 25596
rect 15834 25594 15858 25596
rect 15914 25594 15920 25596
rect 15674 25542 15676 25594
rect 15856 25542 15858 25594
rect 15612 25540 15618 25542
rect 15674 25540 15698 25542
rect 15754 25540 15778 25542
rect 15834 25540 15858 25542
rect 15914 25540 15920 25542
rect 15612 25531 15920 25540
rect 15476 25356 15528 25362
rect 15476 25298 15528 25304
rect 15844 25356 15896 25362
rect 15844 25298 15896 25304
rect 15016 24744 15068 24750
rect 15016 24686 15068 24692
rect 14924 24608 14976 24614
rect 14924 24550 14976 24556
rect 14832 23112 14884 23118
rect 14832 23054 14884 23060
rect 14740 22772 14792 22778
rect 14740 22714 14792 22720
rect 14832 22772 14884 22778
rect 14832 22714 14884 22720
rect 14752 22250 14780 22714
rect 14844 22642 14872 22714
rect 14832 22636 14884 22642
rect 14832 22578 14884 22584
rect 14844 22438 14872 22578
rect 14832 22432 14884 22438
rect 14832 22374 14884 22380
rect 14752 22234 14872 22250
rect 14752 22228 14884 22234
rect 14752 22222 14832 22228
rect 14832 22170 14884 22176
rect 14832 22092 14884 22098
rect 15028 22094 15056 24686
rect 15120 22778 15148 25230
rect 15396 25214 15516 25242
rect 15384 25152 15436 25158
rect 15384 25094 15436 25100
rect 15200 23520 15252 23526
rect 15200 23462 15252 23468
rect 15212 23186 15240 23462
rect 15200 23180 15252 23186
rect 15200 23122 15252 23128
rect 15200 22976 15252 22982
rect 15200 22918 15252 22924
rect 15108 22772 15160 22778
rect 15108 22714 15160 22720
rect 15212 22574 15240 22918
rect 15200 22568 15252 22574
rect 15200 22510 15252 22516
rect 15108 22094 15160 22098
rect 15028 22092 15160 22094
rect 14884 22052 14964 22080
rect 15028 22066 15108 22092
rect 14832 22034 14884 22040
rect 14648 21548 14700 21554
rect 14648 21490 14700 21496
rect 14554 21448 14610 21457
rect 14554 21383 14610 21392
rect 14464 20460 14516 20466
rect 14384 20420 14464 20448
rect 14280 20392 14332 20398
rect 14280 20334 14332 20340
rect 14280 20256 14332 20262
rect 14280 20198 14332 20204
rect 14292 19417 14320 20198
rect 14278 19408 14334 19417
rect 14278 19343 14334 19352
rect 14384 19258 14412 20420
rect 14464 20402 14516 20408
rect 14464 20324 14516 20330
rect 14464 20266 14516 20272
rect 14292 19242 14412 19258
rect 14280 19236 14412 19242
rect 14332 19230 14412 19236
rect 14280 19178 14332 19184
rect 14292 16436 14320 19178
rect 14372 19168 14424 19174
rect 14372 19110 14424 19116
rect 14384 18290 14412 19110
rect 14372 18284 14424 18290
rect 14372 18226 14424 18232
rect 14384 17134 14412 18226
rect 14372 17128 14424 17134
rect 14372 17070 14424 17076
rect 14476 16504 14504 20266
rect 14568 19334 14596 21383
rect 14936 19334 14964 22052
rect 15212 22094 15240 22510
rect 15292 22094 15344 22098
rect 15212 22092 15344 22094
rect 15212 22066 15292 22092
rect 15108 22034 15160 22040
rect 15292 22034 15344 22040
rect 15016 22024 15068 22030
rect 15016 21966 15068 21972
rect 15028 21894 15056 21966
rect 15016 21888 15068 21894
rect 15016 21830 15068 21836
rect 15396 21690 15424 25094
rect 15384 21684 15436 21690
rect 15304 21644 15384 21672
rect 15200 21344 15252 21350
rect 15200 21286 15252 21292
rect 15108 20460 15160 20466
rect 15108 20402 15160 20408
rect 14568 19306 14872 19334
rect 14936 19306 15056 19334
rect 14556 18284 14608 18290
rect 14556 18226 14608 18232
rect 14568 17882 14596 18226
rect 14556 17876 14608 17882
rect 14556 17818 14608 17824
rect 14738 17776 14794 17785
rect 14738 17711 14794 17720
rect 14752 17678 14780 17711
rect 14740 17672 14792 17678
rect 14740 17614 14792 17620
rect 14740 17128 14792 17134
rect 14740 17070 14792 17076
rect 14752 16810 14780 17070
rect 14660 16782 14780 16810
rect 14556 16516 14608 16522
rect 14476 16476 14556 16504
rect 14556 16458 14608 16464
rect 14372 16448 14424 16454
rect 14292 16408 14372 16436
rect 14372 16390 14424 16396
rect 14384 15570 14412 16390
rect 14372 15564 14424 15570
rect 14372 15506 14424 15512
rect 14280 15360 14332 15366
rect 14280 15302 14332 15308
rect 14292 14890 14320 15302
rect 14464 14952 14516 14958
rect 14464 14894 14516 14900
rect 14280 14884 14332 14890
rect 14280 14826 14332 14832
rect 14188 14340 14240 14346
rect 14188 14282 14240 14288
rect 14188 13932 14240 13938
rect 14188 13874 14240 13880
rect 14200 13190 14228 13874
rect 14292 13326 14320 14826
rect 14372 13524 14424 13530
rect 14372 13466 14424 13472
rect 14280 13320 14332 13326
rect 14280 13262 14332 13268
rect 14188 13184 14240 13190
rect 14188 13126 14240 13132
rect 14280 12776 14332 12782
rect 14108 12736 14280 12764
rect 14280 12718 14332 12724
rect 14096 12640 14148 12646
rect 14096 12582 14148 12588
rect 14004 12436 14056 12442
rect 14004 12378 14056 12384
rect 14004 12096 14056 12102
rect 14004 12038 14056 12044
rect 13912 11824 13964 11830
rect 13912 11766 13964 11772
rect 13820 11756 13872 11762
rect 13820 11698 13872 11704
rect 13726 11112 13782 11121
rect 13648 11070 13726 11098
rect 13726 11047 13782 11056
rect 13556 10968 13768 10996
rect 13452 10532 13504 10538
rect 13504 10492 13676 10520
rect 13452 10474 13504 10480
rect 13360 10056 13412 10062
rect 13360 9998 13412 10004
rect 13268 9920 13320 9926
rect 13268 9862 13320 9868
rect 13268 8628 13320 8634
rect 13268 8570 13320 8576
rect 13280 7206 13308 8570
rect 13372 7818 13400 9998
rect 13544 7948 13596 7954
rect 13544 7890 13596 7896
rect 13360 7812 13412 7818
rect 13360 7754 13412 7760
rect 13268 7200 13320 7206
rect 13268 7142 13320 7148
rect 13372 7002 13400 7754
rect 13452 7744 13504 7750
rect 13452 7686 13504 7692
rect 13464 7546 13492 7686
rect 13452 7540 13504 7546
rect 13452 7482 13504 7488
rect 13556 7002 13584 7890
rect 13648 7818 13676 10492
rect 13636 7812 13688 7818
rect 13636 7754 13688 7760
rect 13648 7274 13676 7754
rect 13636 7268 13688 7274
rect 13636 7210 13688 7216
rect 13360 6996 13412 7002
rect 13360 6938 13412 6944
rect 13544 6996 13596 7002
rect 13544 6938 13596 6944
rect 13740 6390 13768 10968
rect 13832 10674 13860 11698
rect 14016 11257 14044 12038
rect 14002 11248 14058 11257
rect 14002 11183 14058 11192
rect 13912 10736 13964 10742
rect 13912 10678 13964 10684
rect 13820 10668 13872 10674
rect 13820 10610 13872 10616
rect 13728 6384 13780 6390
rect 13358 6352 13414 6361
rect 13728 6326 13780 6332
rect 13358 6287 13360 6296
rect 13412 6287 13414 6296
rect 13360 6258 13412 6264
rect 13832 5896 13860 10610
rect 13924 9586 13952 10678
rect 14016 9722 14044 11183
rect 14004 9716 14056 9722
rect 14004 9658 14056 9664
rect 13912 9580 13964 9586
rect 13912 9522 13964 9528
rect 14016 8090 14044 9658
rect 14004 8084 14056 8090
rect 14004 8026 14056 8032
rect 14108 7936 14136 12582
rect 14188 12436 14240 12442
rect 14188 12378 14240 12384
rect 14200 11898 14228 12378
rect 14188 11892 14240 11898
rect 14188 11834 14240 11840
rect 14292 11801 14320 12718
rect 14384 12102 14412 13466
rect 14476 13394 14504 14894
rect 14568 13938 14596 16458
rect 14556 13932 14608 13938
rect 14556 13874 14608 13880
rect 14464 13388 14516 13394
rect 14464 13330 14516 13336
rect 14568 13274 14596 13874
rect 14476 13246 14596 13274
rect 14372 12096 14424 12102
rect 14372 12038 14424 12044
rect 14278 11792 14334 11801
rect 14278 11727 14334 11736
rect 14292 11558 14320 11727
rect 14280 11552 14332 11558
rect 14280 11494 14332 11500
rect 14476 11370 14504 13246
rect 14556 12164 14608 12170
rect 14660 12152 14688 16782
rect 14844 15502 14872 19306
rect 15028 17202 15056 19306
rect 15016 17196 15068 17202
rect 15016 17138 15068 17144
rect 15120 16538 15148 20402
rect 15212 20398 15240 21286
rect 15200 20392 15252 20398
rect 15200 20334 15252 20340
rect 15198 19544 15254 19553
rect 15198 19479 15254 19488
rect 15212 18630 15240 19479
rect 15200 18624 15252 18630
rect 15200 18566 15252 18572
rect 15200 18080 15252 18086
rect 15200 18022 15252 18028
rect 15212 17184 15240 18022
rect 15304 17338 15332 21644
rect 15384 21626 15436 21632
rect 15384 20256 15436 20262
rect 15384 20198 15436 20204
rect 15396 19990 15424 20198
rect 15384 19984 15436 19990
rect 15384 19926 15436 19932
rect 15488 19938 15516 25214
rect 15856 25140 15884 25298
rect 15948 25294 15976 26998
rect 15936 25288 15988 25294
rect 15936 25230 15988 25236
rect 15856 25112 15976 25140
rect 15612 24508 15920 24517
rect 15612 24506 15618 24508
rect 15674 24506 15698 24508
rect 15754 24506 15778 24508
rect 15834 24506 15858 24508
rect 15914 24506 15920 24508
rect 15674 24454 15676 24506
rect 15856 24454 15858 24506
rect 15612 24452 15618 24454
rect 15674 24452 15698 24454
rect 15754 24452 15778 24454
rect 15834 24452 15858 24454
rect 15914 24452 15920 24454
rect 15612 24443 15920 24452
rect 15612 23420 15920 23429
rect 15612 23418 15618 23420
rect 15674 23418 15698 23420
rect 15754 23418 15778 23420
rect 15834 23418 15858 23420
rect 15914 23418 15920 23420
rect 15674 23366 15676 23418
rect 15856 23366 15858 23418
rect 15612 23364 15618 23366
rect 15674 23364 15698 23366
rect 15754 23364 15778 23366
rect 15834 23364 15858 23366
rect 15914 23364 15920 23366
rect 15612 23355 15920 23364
rect 15612 22332 15920 22341
rect 15612 22330 15618 22332
rect 15674 22330 15698 22332
rect 15754 22330 15778 22332
rect 15834 22330 15858 22332
rect 15914 22330 15920 22332
rect 15674 22278 15676 22330
rect 15856 22278 15858 22330
rect 15612 22276 15618 22278
rect 15674 22276 15698 22278
rect 15754 22276 15778 22278
rect 15834 22276 15858 22278
rect 15914 22276 15920 22278
rect 15612 22267 15920 22276
rect 15612 21244 15920 21253
rect 15612 21242 15618 21244
rect 15674 21242 15698 21244
rect 15754 21242 15778 21244
rect 15834 21242 15858 21244
rect 15914 21242 15920 21244
rect 15674 21190 15676 21242
rect 15856 21190 15858 21242
rect 15612 21188 15618 21190
rect 15674 21188 15698 21190
rect 15754 21188 15778 21190
rect 15834 21188 15858 21190
rect 15914 21188 15920 21190
rect 15612 21179 15920 21188
rect 15612 20156 15920 20165
rect 15612 20154 15618 20156
rect 15674 20154 15698 20156
rect 15754 20154 15778 20156
rect 15834 20154 15858 20156
rect 15914 20154 15920 20156
rect 15674 20102 15676 20154
rect 15856 20102 15858 20154
rect 15612 20100 15618 20102
rect 15674 20100 15698 20102
rect 15754 20100 15778 20102
rect 15834 20100 15858 20102
rect 15914 20100 15920 20102
rect 15612 20091 15920 20100
rect 15488 19910 15700 19938
rect 15672 19854 15700 19910
rect 15660 19848 15712 19854
rect 15660 19790 15712 19796
rect 15844 19848 15896 19854
rect 15844 19790 15896 19796
rect 15672 19378 15700 19790
rect 15856 19514 15884 19790
rect 15844 19508 15896 19514
rect 15844 19450 15896 19456
rect 15660 19372 15712 19378
rect 15660 19314 15712 19320
rect 15612 19068 15920 19077
rect 15612 19066 15618 19068
rect 15674 19066 15698 19068
rect 15754 19066 15778 19068
rect 15834 19066 15858 19068
rect 15914 19066 15920 19068
rect 15674 19014 15676 19066
rect 15856 19014 15858 19066
rect 15612 19012 15618 19014
rect 15674 19012 15698 19014
rect 15754 19012 15778 19014
rect 15834 19012 15858 19014
rect 15914 19012 15920 19014
rect 15612 19003 15920 19012
rect 15612 17980 15920 17989
rect 15612 17978 15618 17980
rect 15674 17978 15698 17980
rect 15754 17978 15778 17980
rect 15834 17978 15858 17980
rect 15914 17978 15920 17980
rect 15674 17926 15676 17978
rect 15856 17926 15858 17978
rect 15612 17924 15618 17926
rect 15674 17924 15698 17926
rect 15754 17924 15778 17926
rect 15834 17924 15858 17926
rect 15914 17924 15920 17926
rect 15612 17915 15920 17924
rect 15568 17672 15620 17678
rect 15568 17614 15620 17620
rect 15292 17332 15344 17338
rect 15292 17274 15344 17280
rect 15580 17202 15608 17614
rect 15568 17196 15620 17202
rect 15212 17156 15424 17184
rect 15292 17060 15344 17066
rect 15292 17002 15344 17008
rect 15304 16794 15332 17002
rect 15292 16788 15344 16794
rect 15292 16730 15344 16736
rect 15028 16510 15148 16538
rect 14832 15496 14884 15502
rect 14738 15464 14794 15473
rect 14884 15456 14964 15484
rect 14832 15438 14884 15444
rect 14738 15399 14740 15408
rect 14792 15399 14794 15408
rect 14740 15370 14792 15376
rect 14832 15360 14884 15366
rect 14832 15302 14884 15308
rect 14844 15042 14872 15302
rect 14936 15178 14964 15456
rect 15028 15366 15056 16510
rect 15108 16448 15160 16454
rect 15108 16390 15160 16396
rect 15120 16046 15148 16390
rect 15200 16176 15252 16182
rect 15200 16118 15252 16124
rect 15290 16144 15346 16153
rect 15108 16040 15160 16046
rect 15108 15982 15160 15988
rect 15120 15434 15148 15982
rect 15108 15428 15160 15434
rect 15108 15370 15160 15376
rect 15016 15360 15068 15366
rect 15016 15302 15068 15308
rect 14936 15150 15148 15178
rect 14844 15014 15056 15042
rect 14832 14952 14884 14958
rect 14832 14894 14884 14900
rect 14740 14272 14792 14278
rect 14740 14214 14792 14220
rect 14752 14006 14780 14214
rect 14740 14000 14792 14006
rect 14740 13942 14792 13948
rect 14844 13734 14872 14894
rect 14924 14884 14976 14890
rect 14924 14826 14976 14832
rect 14936 14618 14964 14826
rect 14924 14612 14976 14618
rect 14924 14554 14976 14560
rect 15028 14362 15056 15014
rect 14936 14334 15056 14362
rect 14832 13728 14884 13734
rect 14832 13670 14884 13676
rect 14832 12640 14884 12646
rect 14752 12600 14832 12628
rect 14752 12238 14780 12600
rect 14832 12582 14884 12588
rect 14936 12458 14964 14334
rect 15016 14272 15068 14278
rect 15016 14214 15068 14220
rect 15028 13870 15056 14214
rect 15016 13864 15068 13870
rect 15016 13806 15068 13812
rect 14844 12430 14964 12458
rect 14740 12232 14792 12238
rect 14740 12174 14792 12180
rect 14608 12124 14688 12152
rect 14556 12106 14608 12112
rect 14200 11342 14504 11370
rect 14200 9994 14228 11342
rect 14568 11286 14596 12106
rect 14556 11280 14608 11286
rect 14556 11222 14608 11228
rect 14648 11280 14700 11286
rect 14648 11222 14700 11228
rect 14280 11212 14332 11218
rect 14280 11154 14332 11160
rect 14292 10130 14320 11154
rect 14464 10464 14516 10470
rect 14464 10406 14516 10412
rect 14476 10266 14504 10406
rect 14464 10260 14516 10266
rect 14464 10202 14516 10208
rect 14556 10192 14608 10198
rect 14660 10180 14688 11222
rect 14740 10464 14792 10470
rect 14740 10406 14792 10412
rect 14752 10266 14780 10406
rect 14740 10260 14792 10266
rect 14740 10202 14792 10208
rect 14608 10152 14688 10180
rect 14738 10160 14794 10169
rect 14556 10134 14608 10140
rect 14280 10124 14332 10130
rect 14738 10095 14794 10104
rect 14280 10066 14332 10072
rect 14188 9988 14240 9994
rect 14188 9930 14240 9936
rect 14016 7908 14136 7936
rect 13912 7880 13964 7886
rect 13912 7822 13964 7828
rect 13924 6730 13952 7822
rect 13912 6724 13964 6730
rect 13912 6666 13964 6672
rect 13740 5868 13860 5896
rect 13740 5250 13768 5868
rect 13924 5846 13952 6666
rect 13912 5840 13964 5846
rect 13912 5782 13964 5788
rect 13820 5772 13872 5778
rect 13820 5714 13872 5720
rect 13648 5222 13768 5250
rect 13452 5092 13504 5098
rect 13452 5034 13504 5040
rect 13268 4140 13320 4146
rect 13268 4082 13320 4088
rect 12532 2372 12584 2378
rect 12532 2314 12584 2320
rect 13084 2372 13136 2378
rect 13084 2314 13136 2320
rect 13176 2372 13228 2378
rect 13176 2314 13228 2320
rect 12254 2136 12310 2145
rect 12544 2106 12572 2314
rect 12679 2204 12987 2213
rect 12679 2202 12685 2204
rect 12741 2202 12765 2204
rect 12821 2202 12845 2204
rect 12901 2202 12925 2204
rect 12981 2202 12987 2204
rect 12741 2150 12743 2202
rect 12923 2150 12925 2202
rect 12679 2148 12685 2150
rect 12741 2148 12765 2150
rect 12821 2148 12845 2150
rect 12901 2148 12925 2150
rect 12981 2148 12987 2150
rect 12679 2139 12987 2148
rect 12254 2071 12310 2080
rect 12532 2100 12584 2106
rect 12268 1970 12296 2071
rect 12532 2042 12584 2048
rect 12256 1964 12308 1970
rect 12256 1906 12308 1912
rect 13096 1873 13124 2314
rect 13280 2038 13308 4082
rect 13464 3738 13492 5034
rect 13648 5001 13676 5222
rect 13728 5160 13780 5166
rect 13832 5148 13860 5714
rect 14016 5692 14044 7908
rect 14200 7834 14228 9930
rect 14108 7806 14228 7834
rect 14108 6798 14136 7806
rect 14188 7744 14240 7750
rect 14188 7686 14240 7692
rect 14096 6792 14148 6798
rect 14096 6734 14148 6740
rect 13780 5120 13860 5148
rect 13924 5664 14044 5692
rect 13728 5102 13780 5108
rect 13634 4992 13690 5001
rect 13634 4927 13690 4936
rect 13924 3942 13952 5664
rect 14004 5228 14056 5234
rect 14004 5170 14056 5176
rect 14016 4282 14044 5170
rect 14004 4276 14056 4282
rect 14004 4218 14056 4224
rect 14108 4196 14136 6734
rect 14200 6458 14228 7686
rect 14292 7410 14320 10066
rect 14464 10056 14516 10062
rect 14370 10024 14426 10033
rect 14464 9998 14516 10004
rect 14646 10024 14702 10033
rect 14370 9959 14426 9968
rect 14384 9586 14412 9959
rect 14476 9738 14504 9998
rect 14646 9959 14702 9968
rect 14554 9752 14610 9761
rect 14476 9710 14554 9738
rect 14554 9687 14610 9696
rect 14556 9648 14608 9654
rect 14556 9590 14608 9596
rect 14372 9580 14424 9586
rect 14372 9522 14424 9528
rect 14464 8832 14516 8838
rect 14464 8774 14516 8780
rect 14370 8392 14426 8401
rect 14370 8327 14426 8336
rect 14280 7404 14332 7410
rect 14280 7346 14332 7352
rect 14188 6452 14240 6458
rect 14188 6394 14240 6400
rect 14292 5778 14320 7346
rect 14280 5772 14332 5778
rect 14280 5714 14332 5720
rect 14188 4208 14240 4214
rect 14108 4168 14188 4196
rect 14188 4150 14240 4156
rect 13912 3936 13964 3942
rect 13912 3878 13964 3884
rect 13452 3732 13504 3738
rect 13452 3674 13504 3680
rect 13452 2984 13504 2990
rect 13452 2926 13504 2932
rect 13464 2650 13492 2926
rect 13452 2644 13504 2650
rect 13452 2586 13504 2592
rect 13910 2544 13966 2553
rect 13910 2479 13912 2488
rect 13964 2479 13966 2488
rect 13912 2450 13964 2456
rect 13360 2304 13412 2310
rect 13360 2246 13412 2252
rect 13268 2032 13320 2038
rect 13268 1974 13320 1980
rect 13082 1864 13138 1873
rect 13082 1799 13138 1808
rect 12532 1420 12584 1426
rect 12532 1362 12584 1368
rect 12256 1352 12308 1358
rect 12176 1312 12256 1340
rect 12256 1294 12308 1300
rect 12256 1216 12308 1222
rect 12256 1158 12308 1164
rect 11428 876 11480 882
rect 11428 818 11480 824
rect 11716 870 12020 898
rect 11244 604 11296 610
rect 11244 546 11296 552
rect 11440 160 11468 818
rect 11716 160 11744 870
rect 11980 604 12032 610
rect 11980 546 12032 552
rect 11992 160 12020 546
rect 12268 160 12296 1158
rect 12544 160 12572 1362
rect 13372 1358 13400 2246
rect 13728 1760 13780 1766
rect 13728 1702 13780 1708
rect 14188 1760 14240 1766
rect 14188 1702 14240 1708
rect 13740 1562 13768 1702
rect 13728 1556 13780 1562
rect 13728 1498 13780 1504
rect 13636 1488 13688 1494
rect 13636 1430 13688 1436
rect 12716 1352 12768 1358
rect 12714 1320 12716 1329
rect 13360 1352 13412 1358
rect 12768 1320 12770 1329
rect 13452 1352 13504 1358
rect 13360 1294 13412 1300
rect 13450 1320 13452 1329
rect 13504 1320 13506 1329
rect 12714 1255 12770 1264
rect 13450 1255 13506 1264
rect 12900 1216 12952 1222
rect 13268 1216 13320 1222
rect 12952 1176 13124 1204
rect 12900 1158 12952 1164
rect 12679 1116 12987 1125
rect 12679 1114 12685 1116
rect 12741 1114 12765 1116
rect 12821 1114 12845 1116
rect 12901 1114 12925 1116
rect 12981 1114 12987 1116
rect 12741 1062 12743 1114
rect 12923 1062 12925 1114
rect 12679 1060 12685 1062
rect 12741 1060 12765 1062
rect 12821 1060 12845 1062
rect 12901 1060 12925 1062
rect 12981 1060 12987 1062
rect 12679 1051 12987 1060
rect 13096 490 13124 1176
rect 13004 462 13124 490
rect 13188 1176 13268 1204
rect 10322 54 10456 82
rect 10322 -300 10378 54
rect 10598 -300 10654 160
rect 10874 -300 10930 160
rect 11150 -300 11206 160
rect 11426 -300 11482 160
rect 11702 -300 11758 160
rect 11978 -300 12034 160
rect 12254 -300 12310 160
rect 12530 -300 12586 160
rect 12806 82 12862 160
rect 13004 82 13032 462
rect 13188 218 13216 1176
rect 13268 1158 13320 1164
rect 13360 1216 13412 1222
rect 13360 1158 13412 1164
rect 13096 190 13216 218
rect 13096 160 13124 190
rect 13372 160 13400 1158
rect 13648 160 13676 1430
rect 14096 1352 14148 1358
rect 14094 1320 14096 1329
rect 14148 1320 14150 1329
rect 14094 1255 14150 1264
rect 13912 1216 13964 1222
rect 13912 1158 13964 1164
rect 13924 160 13952 1158
rect 14200 160 14228 1702
rect 14384 610 14412 8327
rect 14476 2990 14504 8774
rect 14568 4282 14596 9590
rect 14660 6730 14688 9959
rect 14752 8820 14780 10095
rect 14844 8974 14872 12430
rect 14924 12300 14976 12306
rect 14924 12242 14976 12248
rect 14936 11898 14964 12242
rect 15016 12096 15068 12102
rect 15016 12038 15068 12044
rect 15028 11898 15056 12038
rect 14924 11892 14976 11898
rect 14924 11834 14976 11840
rect 15016 11892 15068 11898
rect 15016 11834 15068 11840
rect 14924 11552 14976 11558
rect 14924 11494 14976 11500
rect 14936 11354 14964 11494
rect 14924 11348 14976 11354
rect 14924 11290 14976 11296
rect 15120 11234 15148 15150
rect 15212 14958 15240 16118
rect 15290 16079 15292 16088
rect 15344 16079 15346 16088
rect 15292 16050 15344 16056
rect 15200 14952 15252 14958
rect 15200 14894 15252 14900
rect 15212 14618 15240 14894
rect 15200 14612 15252 14618
rect 15200 14554 15252 14560
rect 15200 14408 15252 14414
rect 15200 14350 15252 14356
rect 14936 11206 15148 11234
rect 14936 10538 14964 11206
rect 15016 11144 15068 11150
rect 15016 11086 15068 11092
rect 14924 10532 14976 10538
rect 14924 10474 14976 10480
rect 14936 9382 14964 10474
rect 15028 10062 15056 11086
rect 15212 10742 15240 14350
rect 15304 14006 15332 16050
rect 15292 14000 15344 14006
rect 15292 13942 15344 13948
rect 15292 13320 15344 13326
rect 15292 13262 15344 13268
rect 15200 10736 15252 10742
rect 15200 10678 15252 10684
rect 15198 10160 15254 10169
rect 15304 10146 15332 13262
rect 15254 10118 15332 10146
rect 15198 10095 15254 10104
rect 15016 10056 15068 10062
rect 15016 9998 15068 10004
rect 15200 10056 15252 10062
rect 15200 9998 15252 10004
rect 15292 10056 15344 10062
rect 15292 9998 15344 10004
rect 15028 9926 15056 9998
rect 15016 9920 15068 9926
rect 15016 9862 15068 9868
rect 15016 9716 15068 9722
rect 15212 9704 15240 9998
rect 15304 9722 15332 9998
rect 15068 9676 15240 9704
rect 15292 9716 15344 9722
rect 15016 9658 15068 9664
rect 15292 9658 15344 9664
rect 15396 9602 15424 17156
rect 15568 17138 15620 17144
rect 15612 16892 15920 16901
rect 15612 16890 15618 16892
rect 15674 16890 15698 16892
rect 15754 16890 15778 16892
rect 15834 16890 15858 16892
rect 15914 16890 15920 16892
rect 15674 16838 15676 16890
rect 15856 16838 15858 16890
rect 15612 16836 15618 16838
rect 15674 16836 15698 16838
rect 15754 16836 15778 16838
rect 15834 16836 15858 16838
rect 15914 16836 15920 16838
rect 15612 16827 15920 16836
rect 15612 15804 15920 15813
rect 15612 15802 15618 15804
rect 15674 15802 15698 15804
rect 15754 15802 15778 15804
rect 15834 15802 15858 15804
rect 15914 15802 15920 15804
rect 15674 15750 15676 15802
rect 15856 15750 15858 15802
rect 15612 15748 15618 15750
rect 15674 15748 15698 15750
rect 15754 15748 15778 15750
rect 15834 15748 15858 15750
rect 15914 15748 15920 15750
rect 15612 15739 15920 15748
rect 15948 15706 15976 25112
rect 16040 21622 16068 27338
rect 16132 23050 16160 30670
rect 16224 28966 16252 41006
rect 16212 28960 16264 28966
rect 16212 28902 16264 28908
rect 16212 27328 16264 27334
rect 16212 27270 16264 27276
rect 16224 27062 16252 27270
rect 16212 27056 16264 27062
rect 16212 26998 16264 27004
rect 16316 26568 16344 43046
rect 17328 42702 17356 43386
rect 18064 43246 18092 43846
rect 18052 43240 18104 43246
rect 18052 43182 18104 43188
rect 18340 43194 18368 44540
rect 18420 43988 18472 43994
rect 18420 43930 18472 43936
rect 18432 43382 18460 43930
rect 18616 43874 18644 44540
rect 18892 44010 18920 44540
rect 19168 44282 19196 44540
rect 19168 44254 19288 44282
rect 19156 44124 19208 44130
rect 19156 44066 19208 44072
rect 19064 44056 19116 44062
rect 18892 43982 19012 44010
rect 19064 43998 19116 44004
rect 18616 43846 18920 43874
rect 18544 43548 18852 43557
rect 18544 43546 18550 43548
rect 18606 43546 18630 43548
rect 18686 43546 18710 43548
rect 18766 43546 18790 43548
rect 18846 43546 18852 43548
rect 18606 43494 18608 43546
rect 18788 43494 18790 43546
rect 18544 43492 18550 43494
rect 18606 43492 18630 43494
rect 18686 43492 18710 43494
rect 18766 43492 18790 43494
rect 18846 43492 18852 43494
rect 18544 43483 18852 43492
rect 18892 43382 18920 43846
rect 18420 43376 18472 43382
rect 18420 43318 18472 43324
rect 18880 43376 18932 43382
rect 18880 43318 18932 43324
rect 18696 43240 18748 43246
rect 18340 43188 18696 43194
rect 18340 43182 18748 43188
rect 18984 43194 19012 43982
rect 19076 43314 19104 43998
rect 19168 43314 19196 44066
rect 19064 43308 19116 43314
rect 19064 43250 19116 43256
rect 19156 43308 19208 43314
rect 19156 43250 19208 43256
rect 19260 43194 19288 44254
rect 19444 43602 19472 44540
rect 19444 43574 19656 43602
rect 17868 43172 17920 43178
rect 18340 43166 18736 43182
rect 18984 43166 19104 43194
rect 17868 43114 17920 43120
rect 17592 43104 17644 43110
rect 17592 43046 17644 43052
rect 17776 43104 17828 43110
rect 17776 43046 17828 43052
rect 17604 42945 17632 43046
rect 17590 42936 17646 42945
rect 17590 42871 17646 42880
rect 17788 42838 17816 43046
rect 17776 42832 17828 42838
rect 17776 42774 17828 42780
rect 17880 42702 17908 43114
rect 18052 43104 18104 43110
rect 18052 43046 18104 43052
rect 18604 43104 18656 43110
rect 18604 43046 18656 43052
rect 18064 42702 18092 43046
rect 18616 42906 18644 43046
rect 18604 42900 18656 42906
rect 18604 42842 18656 42848
rect 17316 42696 17368 42702
rect 17316 42638 17368 42644
rect 17868 42696 17920 42702
rect 17868 42638 17920 42644
rect 18052 42696 18104 42702
rect 18328 42696 18380 42702
rect 18052 42638 18104 42644
rect 18326 42664 18328 42673
rect 18380 42664 18382 42673
rect 16488 42628 16540 42634
rect 16488 42570 16540 42576
rect 17960 42628 18012 42634
rect 18326 42599 18382 42608
rect 17960 42570 18012 42576
rect 16500 42362 16528 42570
rect 16764 42560 16816 42566
rect 16764 42502 16816 42508
rect 17132 42560 17184 42566
rect 17132 42502 17184 42508
rect 17500 42560 17552 42566
rect 17500 42502 17552 42508
rect 16776 42362 16804 42502
rect 16488 42356 16540 42362
rect 16488 42298 16540 42304
rect 16764 42356 16816 42362
rect 16764 42298 16816 42304
rect 16396 42288 16448 42294
rect 16396 42230 16448 42236
rect 16408 33658 16436 42230
rect 17040 40928 17092 40934
rect 17040 40870 17092 40876
rect 16580 40044 16632 40050
rect 16580 39986 16632 39992
rect 16488 34944 16540 34950
rect 16488 34886 16540 34892
rect 16396 33652 16448 33658
rect 16396 33594 16448 33600
rect 16500 33538 16528 34886
rect 16408 33510 16528 33538
rect 16408 28218 16436 33510
rect 16488 33448 16540 33454
rect 16488 33390 16540 33396
rect 16500 33114 16528 33390
rect 16488 33108 16540 33114
rect 16488 33050 16540 33056
rect 16592 32042 16620 39986
rect 16672 34604 16724 34610
rect 16672 34546 16724 34552
rect 16684 32774 16712 34546
rect 16762 33960 16818 33969
rect 16762 33895 16818 33904
rect 16776 33590 16804 33895
rect 16764 33584 16816 33590
rect 16764 33526 16816 33532
rect 16856 33516 16908 33522
rect 16856 33458 16908 33464
rect 16672 32768 16724 32774
rect 16672 32710 16724 32716
rect 16762 32328 16818 32337
rect 16762 32263 16818 32272
rect 16500 32014 16620 32042
rect 16500 31770 16528 32014
rect 16578 31920 16634 31929
rect 16634 31878 16712 31906
rect 16578 31855 16634 31864
rect 16684 31822 16712 31878
rect 16672 31816 16724 31822
rect 16500 31742 16620 31770
rect 16672 31758 16724 31764
rect 16488 30048 16540 30054
rect 16488 29990 16540 29996
rect 16500 29073 16528 29990
rect 16486 29064 16542 29073
rect 16486 28999 16542 29008
rect 16488 28416 16540 28422
rect 16488 28358 16540 28364
rect 16396 28212 16448 28218
rect 16396 28154 16448 28160
rect 16500 28121 16528 28358
rect 16486 28112 16542 28121
rect 16486 28047 16542 28056
rect 16488 28008 16540 28014
rect 16488 27950 16540 27956
rect 16396 27872 16448 27878
rect 16396 27814 16448 27820
rect 16224 26540 16344 26568
rect 16120 23044 16172 23050
rect 16120 22986 16172 22992
rect 16224 21842 16252 26540
rect 16304 26444 16356 26450
rect 16304 26386 16356 26392
rect 16316 23730 16344 26386
rect 16304 23724 16356 23730
rect 16304 23666 16356 23672
rect 16304 23044 16356 23050
rect 16304 22986 16356 22992
rect 16132 21814 16252 21842
rect 16028 21616 16080 21622
rect 16028 21558 16080 21564
rect 16040 20874 16068 21558
rect 16028 20868 16080 20874
rect 16028 20810 16080 20816
rect 16028 20256 16080 20262
rect 16028 20198 16080 20204
rect 16040 19922 16068 20198
rect 16028 19916 16080 19922
rect 16028 19858 16080 19864
rect 16132 18426 16160 21814
rect 16212 21344 16264 21350
rect 16212 21286 16264 21292
rect 16224 21146 16252 21286
rect 16212 21140 16264 21146
rect 16212 21082 16264 21088
rect 16212 20868 16264 20874
rect 16212 20810 16264 20816
rect 16224 19310 16252 20810
rect 16212 19304 16264 19310
rect 16212 19246 16264 19252
rect 16120 18420 16172 18426
rect 16120 18362 16172 18368
rect 16120 18284 16172 18290
rect 16120 18226 16172 18232
rect 16028 17128 16080 17134
rect 16028 17070 16080 17076
rect 16040 16250 16068 17070
rect 16028 16244 16080 16250
rect 16028 16186 16080 16192
rect 16132 16096 16160 18226
rect 16040 16068 16160 16096
rect 15936 15700 15988 15706
rect 15936 15642 15988 15648
rect 15476 15360 15528 15366
rect 15476 15302 15528 15308
rect 15488 15026 15516 15302
rect 15476 15020 15528 15026
rect 15476 14962 15528 14968
rect 15612 14716 15920 14725
rect 15612 14714 15618 14716
rect 15674 14714 15698 14716
rect 15754 14714 15778 14716
rect 15834 14714 15858 14716
rect 15914 14714 15920 14716
rect 15674 14662 15676 14714
rect 15856 14662 15858 14714
rect 15612 14660 15618 14662
rect 15674 14660 15698 14662
rect 15754 14660 15778 14662
rect 15834 14660 15858 14662
rect 15914 14660 15920 14662
rect 15612 14651 15920 14660
rect 15936 14612 15988 14618
rect 15936 14554 15988 14560
rect 15568 14000 15620 14006
rect 15016 9580 15068 9586
rect 15016 9522 15068 9528
rect 15304 9574 15424 9602
rect 15488 13960 15568 13988
rect 14924 9376 14976 9382
rect 14924 9318 14976 9324
rect 14832 8968 14884 8974
rect 14832 8910 14884 8916
rect 14924 8968 14976 8974
rect 14924 8910 14976 8916
rect 14936 8820 14964 8910
rect 14752 8792 14964 8820
rect 14740 8424 14792 8430
rect 14740 8366 14792 8372
rect 14752 7886 14780 8366
rect 14740 7880 14792 7886
rect 14740 7822 14792 7828
rect 14844 7342 14872 8792
rect 15028 8650 15056 9522
rect 15108 9512 15160 9518
rect 15108 9454 15160 9460
rect 15120 9194 15148 9454
rect 15120 9166 15240 9194
rect 15108 9104 15160 9110
rect 15106 9072 15108 9081
rect 15160 9072 15162 9081
rect 15106 9007 15162 9016
rect 15212 8906 15240 9166
rect 15200 8900 15252 8906
rect 15200 8842 15252 8848
rect 14936 8622 15056 8650
rect 14832 7336 14884 7342
rect 14832 7278 14884 7284
rect 14648 6724 14700 6730
rect 14648 6666 14700 6672
rect 14660 5234 14688 6666
rect 14740 5840 14792 5846
rect 14740 5782 14792 5788
rect 14752 5234 14780 5782
rect 14844 5710 14872 7278
rect 14832 5704 14884 5710
rect 14832 5646 14884 5652
rect 14648 5228 14700 5234
rect 14648 5170 14700 5176
rect 14740 5228 14792 5234
rect 14740 5170 14792 5176
rect 14752 4690 14780 5170
rect 14740 4684 14792 4690
rect 14740 4626 14792 4632
rect 14556 4276 14608 4282
rect 14556 4218 14608 4224
rect 14844 4010 14872 5646
rect 14936 5522 14964 8622
rect 15212 7970 15240 8842
rect 15120 7942 15240 7970
rect 15120 7886 15148 7942
rect 15108 7880 15160 7886
rect 15108 7822 15160 7828
rect 15200 7880 15252 7886
rect 15200 7822 15252 7828
rect 15212 7426 15240 7822
rect 15304 7528 15332 9574
rect 15384 9512 15436 9518
rect 15488 9500 15516 13960
rect 15568 13942 15620 13948
rect 15612 13628 15920 13637
rect 15612 13626 15618 13628
rect 15674 13626 15698 13628
rect 15754 13626 15778 13628
rect 15834 13626 15858 13628
rect 15914 13626 15920 13628
rect 15674 13574 15676 13626
rect 15856 13574 15858 13626
rect 15612 13572 15618 13574
rect 15674 13572 15698 13574
rect 15754 13572 15778 13574
rect 15834 13572 15858 13574
rect 15914 13572 15920 13574
rect 15612 13563 15920 13572
rect 15948 12850 15976 14554
rect 16040 13530 16068 16068
rect 16224 16028 16252 19246
rect 16316 18290 16344 22986
rect 16408 19496 16436 27814
rect 16500 27674 16528 27950
rect 16488 27668 16540 27674
rect 16488 27610 16540 27616
rect 16488 26852 16540 26858
rect 16488 26794 16540 26800
rect 16500 26042 16528 26794
rect 16488 26036 16540 26042
rect 16488 25978 16540 25984
rect 16488 25832 16540 25838
rect 16592 25809 16620 31742
rect 16776 31754 16804 32263
rect 16868 32230 16896 33458
rect 17052 32434 17080 40870
rect 17040 32428 17092 32434
rect 17040 32370 17092 32376
rect 16856 32224 16908 32230
rect 16856 32166 16908 32172
rect 16776 31726 16988 31754
rect 16856 30388 16908 30394
rect 16856 30330 16908 30336
rect 16672 30048 16724 30054
rect 16672 29990 16724 29996
rect 16684 29753 16712 29990
rect 16764 29776 16816 29782
rect 16670 29744 16726 29753
rect 16764 29718 16816 29724
rect 16670 29679 16672 29688
rect 16724 29679 16726 29688
rect 16672 29650 16724 29656
rect 16776 29578 16804 29718
rect 16764 29572 16816 29578
rect 16764 29514 16816 29520
rect 16670 29472 16726 29481
rect 16670 29407 16726 29416
rect 16684 29306 16712 29407
rect 16762 29336 16818 29345
rect 16672 29300 16724 29306
rect 16762 29271 16818 29280
rect 16672 29242 16724 29248
rect 16672 29096 16724 29102
rect 16776 29084 16804 29271
rect 16868 29170 16896 30330
rect 16856 29164 16908 29170
rect 16856 29106 16908 29112
rect 16724 29056 16804 29084
rect 16672 29038 16724 29044
rect 16764 28212 16816 28218
rect 16764 28154 16816 28160
rect 16776 27878 16804 28154
rect 16764 27872 16816 27878
rect 16764 27814 16816 27820
rect 16868 26858 16896 29106
rect 16856 26852 16908 26858
rect 16856 26794 16908 26800
rect 16672 26444 16724 26450
rect 16724 26404 16804 26432
rect 16672 26386 16724 26392
rect 16672 26036 16724 26042
rect 16672 25978 16724 25984
rect 16488 25774 16540 25780
rect 16578 25800 16634 25809
rect 16500 25498 16528 25774
rect 16578 25735 16634 25744
rect 16488 25492 16540 25498
rect 16488 25434 16540 25440
rect 16684 23746 16712 25978
rect 16776 25498 16804 26404
rect 16960 26382 16988 31726
rect 17040 28960 17092 28966
rect 17040 28902 17092 28908
rect 16948 26376 17000 26382
rect 16868 26336 16948 26364
rect 16764 25492 16816 25498
rect 16764 25434 16816 25440
rect 16684 23730 16804 23746
rect 16684 23724 16816 23730
rect 16684 23718 16764 23724
rect 16488 22976 16540 22982
rect 16488 22918 16540 22924
rect 16500 21486 16528 22918
rect 16488 21480 16540 21486
rect 16488 21422 16540 21428
rect 16684 19514 16712 23718
rect 16764 23666 16816 23672
rect 16764 23520 16816 23526
rect 16764 23462 16816 23468
rect 16672 19508 16724 19514
rect 16408 19468 16528 19496
rect 16396 19372 16448 19378
rect 16396 19314 16448 19320
rect 16304 18284 16356 18290
rect 16304 18226 16356 18232
rect 16304 17332 16356 17338
rect 16304 17274 16356 17280
rect 16132 16000 16252 16028
rect 16028 13524 16080 13530
rect 16028 13466 16080 13472
rect 16132 13410 16160 16000
rect 16212 15632 16264 15638
rect 16212 15574 16264 15580
rect 16224 14521 16252 15574
rect 16316 15026 16344 17274
rect 16304 15020 16356 15026
rect 16304 14962 16356 14968
rect 16210 14512 16266 14521
rect 16210 14447 16266 14456
rect 16212 14272 16264 14278
rect 16212 14214 16264 14220
rect 16224 13870 16252 14214
rect 16212 13864 16264 13870
rect 16212 13806 16264 13812
rect 16212 13728 16264 13734
rect 16212 13670 16264 13676
rect 16224 13462 16252 13670
rect 16040 13382 16160 13410
rect 16212 13456 16264 13462
rect 16212 13398 16264 13404
rect 15936 12844 15988 12850
rect 15936 12786 15988 12792
rect 15612 12540 15920 12549
rect 15612 12538 15618 12540
rect 15674 12538 15698 12540
rect 15754 12538 15778 12540
rect 15834 12538 15858 12540
rect 15914 12538 15920 12540
rect 15674 12486 15676 12538
rect 15856 12486 15858 12538
rect 15612 12484 15618 12486
rect 15674 12484 15698 12486
rect 15754 12484 15778 12486
rect 15834 12484 15858 12486
rect 15914 12484 15920 12486
rect 15612 12475 15920 12484
rect 15568 12368 15620 12374
rect 15568 12310 15620 12316
rect 15936 12368 15988 12374
rect 15936 12310 15988 12316
rect 15580 12102 15608 12310
rect 15752 12300 15804 12306
rect 15752 12242 15804 12248
rect 15568 12096 15620 12102
rect 15660 12096 15712 12102
rect 15568 12038 15620 12044
rect 15658 12064 15660 12073
rect 15712 12064 15714 12073
rect 15658 11999 15714 12008
rect 15764 11898 15792 12242
rect 15752 11892 15804 11898
rect 15752 11834 15804 11840
rect 15612 11452 15920 11461
rect 15612 11450 15618 11452
rect 15674 11450 15698 11452
rect 15754 11450 15778 11452
rect 15834 11450 15858 11452
rect 15914 11450 15920 11452
rect 15674 11398 15676 11450
rect 15856 11398 15858 11450
rect 15612 11396 15618 11398
rect 15674 11396 15698 11398
rect 15754 11396 15778 11398
rect 15834 11396 15858 11398
rect 15914 11396 15920 11398
rect 15612 11387 15920 11396
rect 15948 11218 15976 12310
rect 15936 11212 15988 11218
rect 15936 11154 15988 11160
rect 15844 11008 15896 11014
rect 15896 10968 15976 10996
rect 15844 10950 15896 10956
rect 15612 10364 15920 10373
rect 15612 10362 15618 10364
rect 15674 10362 15698 10364
rect 15754 10362 15778 10364
rect 15834 10362 15858 10364
rect 15914 10362 15920 10364
rect 15674 10310 15676 10362
rect 15856 10310 15858 10362
rect 15612 10308 15618 10310
rect 15674 10308 15698 10310
rect 15754 10308 15778 10310
rect 15834 10308 15858 10310
rect 15914 10308 15920 10310
rect 15612 10299 15920 10308
rect 15948 10248 15976 10968
rect 15856 10220 15976 10248
rect 15752 10192 15804 10198
rect 15752 10134 15804 10140
rect 15764 10033 15792 10134
rect 15750 10024 15806 10033
rect 15750 9959 15806 9968
rect 15856 9761 15884 10220
rect 15936 9920 15988 9926
rect 15936 9862 15988 9868
rect 15842 9752 15898 9761
rect 15842 9687 15898 9696
rect 15856 9518 15884 9687
rect 15436 9472 15516 9500
rect 15844 9512 15896 9518
rect 15384 9454 15436 9460
rect 15844 9454 15896 9460
rect 15612 9276 15920 9285
rect 15612 9274 15618 9276
rect 15674 9274 15698 9276
rect 15754 9274 15778 9276
rect 15834 9274 15858 9276
rect 15914 9274 15920 9276
rect 15674 9222 15676 9274
rect 15856 9222 15858 9274
rect 15612 9220 15618 9222
rect 15674 9220 15698 9222
rect 15754 9220 15778 9222
rect 15834 9220 15858 9222
rect 15914 9220 15920 9222
rect 15612 9211 15920 9220
rect 15476 8492 15528 8498
rect 15476 8434 15528 8440
rect 15304 7500 15424 7528
rect 15028 7398 15332 7426
rect 15028 7342 15056 7398
rect 15016 7336 15068 7342
rect 15016 7278 15068 7284
rect 15200 7268 15252 7274
rect 15200 7210 15252 7216
rect 15212 7002 15240 7210
rect 15200 6996 15252 7002
rect 15200 6938 15252 6944
rect 15304 5896 15332 7398
rect 15028 5868 15332 5896
rect 15028 5778 15056 5868
rect 15016 5772 15068 5778
rect 15016 5714 15068 5720
rect 15108 5772 15160 5778
rect 15108 5714 15160 5720
rect 15120 5658 15148 5714
rect 15120 5630 15240 5658
rect 14936 5494 15148 5522
rect 15120 5302 15148 5494
rect 15212 5370 15240 5630
rect 15200 5364 15252 5370
rect 15200 5306 15252 5312
rect 15108 5296 15160 5302
rect 15108 5238 15160 5244
rect 14924 5228 14976 5234
rect 14924 5170 14976 5176
rect 14936 5001 14964 5170
rect 14922 4992 14978 5001
rect 14922 4927 14978 4936
rect 15120 4622 15148 5238
rect 15304 4842 15332 5868
rect 15212 4826 15332 4842
rect 15200 4820 15332 4826
rect 15252 4814 15332 4820
rect 15200 4762 15252 4768
rect 15108 4616 15160 4622
rect 15108 4558 15160 4564
rect 14832 4004 14884 4010
rect 14832 3946 14884 3952
rect 14648 3936 14700 3942
rect 14648 3878 14700 3884
rect 14464 2984 14516 2990
rect 14464 2926 14516 2932
rect 14462 2136 14518 2145
rect 14462 2071 14464 2080
rect 14516 2071 14518 2080
rect 14464 2042 14516 2048
rect 14464 1556 14516 1562
rect 14464 1498 14516 1504
rect 14372 604 14424 610
rect 14372 546 14424 552
rect 14476 160 14504 1498
rect 14556 1352 14608 1358
rect 14554 1320 14556 1329
rect 14608 1320 14610 1329
rect 14554 1255 14610 1264
rect 14660 610 14688 3878
rect 15396 2038 15424 7500
rect 15488 6322 15516 8434
rect 15612 8188 15920 8197
rect 15612 8186 15618 8188
rect 15674 8186 15698 8188
rect 15754 8186 15778 8188
rect 15834 8186 15858 8188
rect 15914 8186 15920 8188
rect 15674 8134 15676 8186
rect 15856 8134 15858 8186
rect 15612 8132 15618 8134
rect 15674 8132 15698 8134
rect 15754 8132 15778 8134
rect 15834 8132 15858 8134
rect 15914 8132 15920 8134
rect 15612 8123 15920 8132
rect 15660 7744 15712 7750
rect 15660 7686 15712 7692
rect 15672 7410 15700 7686
rect 15660 7404 15712 7410
rect 15660 7346 15712 7352
rect 15612 7100 15920 7109
rect 15612 7098 15618 7100
rect 15674 7098 15698 7100
rect 15754 7098 15778 7100
rect 15834 7098 15858 7100
rect 15914 7098 15920 7100
rect 15674 7046 15676 7098
rect 15856 7046 15858 7098
rect 15612 7044 15618 7046
rect 15674 7044 15698 7046
rect 15754 7044 15778 7046
rect 15834 7044 15858 7046
rect 15914 7044 15920 7046
rect 15612 7035 15920 7044
rect 15948 6905 15976 9862
rect 16040 9654 16068 13382
rect 16120 12844 16172 12850
rect 16120 12786 16172 12792
rect 16028 9648 16080 9654
rect 16028 9590 16080 9596
rect 16028 9512 16080 9518
rect 16028 9454 16080 9460
rect 16040 7732 16068 9454
rect 16132 7886 16160 12786
rect 16316 12238 16344 14962
rect 16408 13394 16436 19314
rect 16500 19242 16528 19468
rect 16672 19450 16724 19456
rect 16670 19408 16726 19417
rect 16670 19343 16726 19352
rect 16488 19236 16540 19242
rect 16488 19178 16540 19184
rect 16580 18352 16632 18358
rect 16580 18294 16632 18300
rect 16488 17740 16540 17746
rect 16488 17682 16540 17688
rect 16500 17241 16528 17682
rect 16592 17338 16620 18294
rect 16580 17332 16632 17338
rect 16580 17274 16632 17280
rect 16486 17232 16542 17241
rect 16486 17167 16488 17176
rect 16540 17167 16542 17176
rect 16580 17196 16632 17202
rect 16488 17138 16540 17144
rect 16580 17138 16632 17144
rect 16592 17105 16620 17138
rect 16578 17096 16634 17105
rect 16578 17031 16634 17040
rect 16488 16992 16540 16998
rect 16488 16934 16540 16940
rect 16500 16590 16528 16934
rect 16488 16584 16540 16590
rect 16488 16526 16540 16532
rect 16500 16250 16528 16526
rect 16488 16244 16540 16250
rect 16488 16186 16540 16192
rect 16580 15904 16632 15910
rect 16580 15846 16632 15852
rect 16592 15502 16620 15846
rect 16580 15496 16632 15502
rect 16580 15438 16632 15444
rect 16592 15094 16620 15438
rect 16580 15088 16632 15094
rect 16580 15030 16632 15036
rect 16580 14612 16632 14618
rect 16580 14554 16632 14560
rect 16488 13728 16540 13734
rect 16488 13670 16540 13676
rect 16500 13530 16528 13670
rect 16488 13524 16540 13530
rect 16488 13466 16540 13472
rect 16500 13394 16528 13466
rect 16396 13388 16448 13394
rect 16396 13330 16448 13336
rect 16488 13388 16540 13394
rect 16488 13330 16540 13336
rect 16408 13274 16436 13330
rect 16408 13246 16528 13274
rect 16396 13184 16448 13190
rect 16396 13126 16448 13132
rect 16304 12232 16356 12238
rect 16304 12174 16356 12180
rect 16316 11354 16344 12174
rect 16304 11348 16356 11354
rect 16304 11290 16356 11296
rect 16304 11212 16356 11218
rect 16304 11154 16356 11160
rect 16316 10810 16344 11154
rect 16304 10804 16356 10810
rect 16304 10746 16356 10752
rect 16408 9674 16436 13126
rect 16500 9994 16528 13246
rect 16592 11150 16620 14554
rect 16580 11144 16632 11150
rect 16580 11086 16632 11092
rect 16488 9988 16540 9994
rect 16488 9930 16540 9936
rect 16224 9646 16436 9674
rect 16500 9654 16528 9930
rect 16488 9648 16540 9654
rect 16224 9110 16252 9646
rect 16488 9590 16540 9596
rect 16592 9466 16620 11086
rect 16408 9438 16620 9466
rect 16212 9104 16264 9110
rect 16212 9046 16264 9052
rect 16120 7880 16172 7886
rect 16120 7822 16172 7828
rect 16040 7704 16160 7732
rect 16028 7336 16080 7342
rect 16028 7278 16080 7284
rect 15934 6896 15990 6905
rect 15934 6831 15990 6840
rect 15476 6316 15528 6322
rect 15476 6258 15528 6264
rect 16040 6186 16068 7278
rect 15476 6180 15528 6186
rect 15476 6122 15528 6128
rect 16028 6180 16080 6186
rect 16028 6122 16080 6128
rect 15488 5778 15516 6122
rect 15612 6012 15920 6021
rect 15612 6010 15618 6012
rect 15674 6010 15698 6012
rect 15754 6010 15778 6012
rect 15834 6010 15858 6012
rect 15914 6010 15920 6012
rect 15674 5958 15676 6010
rect 15856 5958 15858 6010
rect 15612 5956 15618 5958
rect 15674 5956 15698 5958
rect 15754 5956 15778 5958
rect 15834 5956 15858 5958
rect 15914 5956 15920 5958
rect 15612 5947 15920 5956
rect 15476 5772 15528 5778
rect 15476 5714 15528 5720
rect 16028 5772 16080 5778
rect 16028 5714 16080 5720
rect 15612 4924 15920 4933
rect 15612 4922 15618 4924
rect 15674 4922 15698 4924
rect 15754 4922 15778 4924
rect 15834 4922 15858 4924
rect 15914 4922 15920 4924
rect 15674 4870 15676 4922
rect 15856 4870 15858 4922
rect 15612 4868 15618 4870
rect 15674 4868 15698 4870
rect 15754 4868 15778 4870
rect 15834 4868 15858 4870
rect 15914 4868 15920 4870
rect 15612 4859 15920 4868
rect 16040 4826 16068 5714
rect 16028 4820 16080 4826
rect 16028 4762 16080 4768
rect 15612 3836 15920 3845
rect 15612 3834 15618 3836
rect 15674 3834 15698 3836
rect 15754 3834 15778 3836
rect 15834 3834 15858 3836
rect 15914 3834 15920 3836
rect 15674 3782 15676 3834
rect 15856 3782 15858 3834
rect 15612 3780 15618 3782
rect 15674 3780 15698 3782
rect 15754 3780 15778 3782
rect 15834 3780 15858 3782
rect 15914 3780 15920 3782
rect 15612 3771 15920 3780
rect 16026 3768 16082 3777
rect 16132 3754 16160 7704
rect 16224 7274 16252 9046
rect 16408 9042 16436 9438
rect 16488 9376 16540 9382
rect 16488 9318 16540 9324
rect 16304 9036 16356 9042
rect 16304 8978 16356 8984
rect 16396 9036 16448 9042
rect 16396 8978 16448 8984
rect 16316 8294 16344 8978
rect 16408 8838 16436 8978
rect 16396 8832 16448 8838
rect 16396 8774 16448 8780
rect 16304 8288 16356 8294
rect 16304 8230 16356 8236
rect 16396 7472 16448 7478
rect 16396 7414 16448 7420
rect 16212 7268 16264 7274
rect 16212 7210 16264 7216
rect 16408 7002 16436 7414
rect 16500 7410 16528 9318
rect 16684 7732 16712 19343
rect 16776 18306 16804 23462
rect 16868 22778 16896 26336
rect 16948 26318 17000 26324
rect 16948 25424 17000 25430
rect 16948 25366 17000 25372
rect 16856 22772 16908 22778
rect 16856 22714 16908 22720
rect 16856 21684 16908 21690
rect 16856 21626 16908 21632
rect 16868 19514 16896 21626
rect 16856 19508 16908 19514
rect 16856 19450 16908 19456
rect 16960 18902 16988 25366
rect 17052 23662 17080 28902
rect 17040 23656 17092 23662
rect 17040 23598 17092 23604
rect 17040 22024 17092 22030
rect 17040 21966 17092 21972
rect 17052 21010 17080 21966
rect 17040 21004 17092 21010
rect 17040 20946 17092 20952
rect 17040 19304 17092 19310
rect 17040 19246 17092 19252
rect 16948 18896 17000 18902
rect 16948 18838 17000 18844
rect 16776 18278 16988 18306
rect 16960 17678 16988 18278
rect 16948 17672 17000 17678
rect 16948 17614 17000 17620
rect 16854 14512 16910 14521
rect 16910 14470 16988 14498
rect 16854 14447 16910 14456
rect 16856 11756 16908 11762
rect 16856 11698 16908 11704
rect 16868 11354 16896 11698
rect 16856 11348 16908 11354
rect 16856 11290 16908 11296
rect 16856 11144 16908 11150
rect 16856 11086 16908 11092
rect 16868 10810 16896 11086
rect 16960 11014 16988 14470
rect 17052 13530 17080 19246
rect 17040 13524 17092 13530
rect 17040 13466 17092 13472
rect 17040 12640 17092 12646
rect 17040 12582 17092 12588
rect 16948 11008 17000 11014
rect 16948 10950 17000 10956
rect 16856 10804 16908 10810
rect 16856 10746 16908 10752
rect 16948 10668 17000 10674
rect 16948 10610 17000 10616
rect 16960 10470 16988 10610
rect 16948 10464 17000 10470
rect 16948 10406 17000 10412
rect 17052 10248 17080 12582
rect 16868 10220 17080 10248
rect 16868 9518 16896 10220
rect 17038 10160 17094 10169
rect 16960 10118 17038 10146
rect 16856 9512 16908 9518
rect 16856 9454 16908 9460
rect 16764 9036 16816 9042
rect 16764 8978 16816 8984
rect 16776 8634 16804 8978
rect 16856 8968 16908 8974
rect 16856 8910 16908 8916
rect 16868 8634 16896 8910
rect 16764 8628 16816 8634
rect 16764 8570 16816 8576
rect 16856 8628 16908 8634
rect 16856 8570 16908 8576
rect 16856 7744 16908 7750
rect 16684 7704 16856 7732
rect 16856 7686 16908 7692
rect 16960 7562 16988 10118
rect 17038 10095 17094 10104
rect 17144 7562 17172 42502
rect 17512 42129 17540 42502
rect 17498 42120 17554 42129
rect 17498 42055 17554 42064
rect 17972 41993 18000 42570
rect 18328 42560 18380 42566
rect 18696 42560 18748 42566
rect 18328 42502 18380 42508
rect 18432 42520 18696 42548
rect 18340 41993 18368 42502
rect 17958 41984 18014 41993
rect 17958 41919 18014 41928
rect 18326 41984 18382 41993
rect 18326 41919 18382 41928
rect 18432 41834 18460 42520
rect 18696 42502 18748 42508
rect 18544 42460 18852 42469
rect 18544 42458 18550 42460
rect 18606 42458 18630 42460
rect 18686 42458 18710 42460
rect 18766 42458 18790 42460
rect 18846 42458 18852 42460
rect 18606 42406 18608 42458
rect 18788 42406 18790 42458
rect 18544 42404 18550 42406
rect 18606 42404 18630 42406
rect 18686 42404 18710 42406
rect 18766 42404 18790 42406
rect 18846 42404 18852 42406
rect 18544 42395 18852 42404
rect 19076 42226 19104 43166
rect 19168 43166 19288 43194
rect 19628 43178 19656 43574
rect 19616 43172 19668 43178
rect 19168 42906 19196 43166
rect 19616 43114 19668 43120
rect 19248 43104 19300 43110
rect 19248 43046 19300 43052
rect 19432 43104 19484 43110
rect 19432 43046 19484 43052
rect 19156 42900 19208 42906
rect 19156 42842 19208 42848
rect 19260 42838 19288 43046
rect 19248 42832 19300 42838
rect 19248 42774 19300 42780
rect 19444 42634 19472 43046
rect 19432 42628 19484 42634
rect 19432 42570 19484 42576
rect 19524 42628 19576 42634
rect 19524 42570 19576 42576
rect 19430 42256 19486 42265
rect 18696 42220 18748 42226
rect 18696 42162 18748 42168
rect 19064 42220 19116 42226
rect 19430 42191 19486 42200
rect 19064 42162 19116 42168
rect 18512 42016 18564 42022
rect 18512 41958 18564 41964
rect 18248 41806 18460 41834
rect 18144 36712 18196 36718
rect 18144 36654 18196 36660
rect 17224 35624 17276 35630
rect 17224 35566 17276 35572
rect 17236 35290 17264 35566
rect 17316 35488 17368 35494
rect 17316 35430 17368 35436
rect 17224 35284 17276 35290
rect 17224 35226 17276 35232
rect 17328 35086 17356 35430
rect 17316 35080 17368 35086
rect 17316 35022 17368 35028
rect 17224 34400 17276 34406
rect 17224 34342 17276 34348
rect 17236 33862 17264 34342
rect 17960 33924 18012 33930
rect 17960 33866 18012 33872
rect 18052 33924 18104 33930
rect 18052 33866 18104 33872
rect 17224 33856 17276 33862
rect 17224 33798 17276 33804
rect 17972 33522 18000 33866
rect 17960 33516 18012 33522
rect 17960 33458 18012 33464
rect 17224 33108 17276 33114
rect 17224 33050 17276 33056
rect 17236 33017 17264 33050
rect 17222 33008 17278 33017
rect 17222 32943 17278 32952
rect 17224 32768 17276 32774
rect 17224 32710 17276 32716
rect 17236 27402 17264 32710
rect 17408 32564 17460 32570
rect 17408 32506 17460 32512
rect 17420 32026 17448 32506
rect 17408 32020 17460 32026
rect 17408 31962 17460 31968
rect 17960 32020 18012 32026
rect 17960 31962 18012 31968
rect 17408 31816 17460 31822
rect 17408 31758 17460 31764
rect 17316 31680 17368 31686
rect 17316 31622 17368 31628
rect 17328 30802 17356 31622
rect 17316 30796 17368 30802
rect 17316 30738 17368 30744
rect 17420 30190 17448 31758
rect 17500 31680 17552 31686
rect 17500 31622 17552 31628
rect 17512 31346 17540 31622
rect 17972 31346 18000 31962
rect 17500 31340 17552 31346
rect 17500 31282 17552 31288
rect 17960 31340 18012 31346
rect 17960 31282 18012 31288
rect 17512 30938 17540 31282
rect 17500 30932 17552 30938
rect 17500 30874 17552 30880
rect 17500 30660 17552 30666
rect 17500 30602 17552 30608
rect 17408 30184 17460 30190
rect 17408 30126 17460 30132
rect 17420 29646 17448 30126
rect 17408 29640 17460 29646
rect 17408 29582 17460 29588
rect 17316 29572 17368 29578
rect 17316 29514 17368 29520
rect 17328 29102 17356 29514
rect 17316 29096 17368 29102
rect 17316 29038 17368 29044
rect 17512 27538 17540 30602
rect 17684 29572 17736 29578
rect 17604 29532 17684 29560
rect 17604 29481 17632 29532
rect 17684 29514 17736 29520
rect 17868 29504 17920 29510
rect 17590 29472 17646 29481
rect 17868 29446 17920 29452
rect 17590 29407 17646 29416
rect 17684 29300 17736 29306
rect 17684 29242 17736 29248
rect 17696 29170 17724 29242
rect 17880 29170 17908 29446
rect 17972 29306 18000 31282
rect 17960 29300 18012 29306
rect 17960 29242 18012 29248
rect 17684 29164 17736 29170
rect 17684 29106 17736 29112
rect 17868 29164 17920 29170
rect 17868 29106 17920 29112
rect 17972 28558 18000 29242
rect 18064 28665 18092 33866
rect 18156 31414 18184 36654
rect 18144 31408 18196 31414
rect 18144 31350 18196 31356
rect 18156 30734 18184 31350
rect 18144 30728 18196 30734
rect 18144 30670 18196 30676
rect 18050 28656 18106 28665
rect 18050 28591 18106 28600
rect 17960 28552 18012 28558
rect 17960 28494 18012 28500
rect 17592 28484 17644 28490
rect 17592 28426 17644 28432
rect 17604 28082 17632 28426
rect 17592 28076 17644 28082
rect 17592 28018 17644 28024
rect 17592 27872 17644 27878
rect 17592 27814 17644 27820
rect 17500 27532 17552 27538
rect 17500 27474 17552 27480
rect 17224 27396 17276 27402
rect 17224 27338 17276 27344
rect 17512 26994 17540 27474
rect 17500 26988 17552 26994
rect 17500 26930 17552 26936
rect 17408 26784 17460 26790
rect 17408 26726 17460 26732
rect 17420 26450 17448 26726
rect 17408 26444 17460 26450
rect 17408 26386 17460 26392
rect 17224 26376 17276 26382
rect 17224 26318 17276 26324
rect 17236 26042 17264 26318
rect 17224 26036 17276 26042
rect 17224 25978 17276 25984
rect 17224 25910 17276 25916
rect 17224 25852 17276 25858
rect 17236 21536 17264 25852
rect 17420 25430 17448 26386
rect 17408 25424 17460 25430
rect 17408 25366 17460 25372
rect 17408 24812 17460 24818
rect 17408 24754 17460 24760
rect 17420 24206 17448 24754
rect 17512 24342 17540 26930
rect 17604 25770 17632 27814
rect 17972 27470 18000 28494
rect 17960 27464 18012 27470
rect 17960 27406 18012 27412
rect 17972 26450 18000 27406
rect 17960 26444 18012 26450
rect 17960 26386 18012 26392
rect 17684 26240 17736 26246
rect 17684 26182 17736 26188
rect 17592 25764 17644 25770
rect 17592 25706 17644 25712
rect 17500 24336 17552 24342
rect 17500 24278 17552 24284
rect 17408 24200 17460 24206
rect 17408 24142 17460 24148
rect 17408 23656 17460 23662
rect 17408 23598 17460 23604
rect 17420 22964 17448 23598
rect 17604 23526 17632 25706
rect 17696 23730 17724 26182
rect 17972 25906 18000 26386
rect 17960 25900 18012 25906
rect 17960 25842 18012 25848
rect 17776 25152 17828 25158
rect 17776 25094 17828 25100
rect 17684 23724 17736 23730
rect 17684 23666 17736 23672
rect 17592 23520 17644 23526
rect 17592 23462 17644 23468
rect 17420 22936 17632 22964
rect 17408 22772 17460 22778
rect 17408 22714 17460 22720
rect 17316 22432 17368 22438
rect 17316 22374 17368 22380
rect 17328 22030 17356 22374
rect 17316 22024 17368 22030
rect 17316 21966 17368 21972
rect 17316 21548 17368 21554
rect 17236 21508 17316 21536
rect 17316 21490 17368 21496
rect 17224 20936 17276 20942
rect 17224 20878 17276 20884
rect 17236 18154 17264 20878
rect 17328 20806 17356 21490
rect 17316 20800 17368 20806
rect 17316 20742 17368 20748
rect 17316 19236 17368 19242
rect 17316 19178 17368 19184
rect 17328 18222 17356 19178
rect 17420 18426 17448 22714
rect 17498 19680 17554 19689
rect 17498 19615 17554 19624
rect 17408 18420 17460 18426
rect 17408 18362 17460 18368
rect 17316 18216 17368 18222
rect 17316 18158 17368 18164
rect 17408 18216 17460 18222
rect 17408 18158 17460 18164
rect 17224 18148 17276 18154
rect 17224 18090 17276 18096
rect 17328 17338 17356 18158
rect 17316 17332 17368 17338
rect 17316 17274 17368 17280
rect 17224 15428 17276 15434
rect 17224 15370 17276 15376
rect 17236 9926 17264 15370
rect 17420 14618 17448 18158
rect 17408 14612 17460 14618
rect 17408 14554 17460 14560
rect 17512 14414 17540 19615
rect 17604 18170 17632 22936
rect 17696 21690 17724 23666
rect 17788 23254 17816 25094
rect 17972 24818 18000 25842
rect 17960 24812 18012 24818
rect 17960 24754 18012 24760
rect 17972 24206 18000 24754
rect 17960 24200 18012 24206
rect 17960 24142 18012 24148
rect 17868 23656 17920 23662
rect 17868 23598 17920 23604
rect 17880 23322 17908 23598
rect 17868 23316 17920 23322
rect 17868 23258 17920 23264
rect 17776 23248 17828 23254
rect 17776 23190 17828 23196
rect 17972 22642 18000 24142
rect 17960 22636 18012 22642
rect 17960 22578 18012 22584
rect 17868 22024 17920 22030
rect 17868 21966 17920 21972
rect 17684 21684 17736 21690
rect 17684 21626 17736 21632
rect 17684 21344 17736 21350
rect 17684 21286 17736 21292
rect 17696 21146 17724 21286
rect 17880 21146 17908 21966
rect 17960 21684 18012 21690
rect 17960 21626 18012 21632
rect 17972 21418 18000 21626
rect 18064 21486 18092 28591
rect 18248 27946 18276 41806
rect 18524 41698 18552 41958
rect 18708 41834 18736 42162
rect 19340 42084 19392 42090
rect 19340 42026 19392 42032
rect 18708 41806 18920 41834
rect 19352 41818 19380 42026
rect 18340 41670 18552 41698
rect 18236 27940 18288 27946
rect 18236 27882 18288 27888
rect 18144 26988 18196 26994
rect 18144 26930 18196 26936
rect 18156 23050 18184 26930
rect 18340 26908 18368 41670
rect 18544 41372 18852 41381
rect 18544 41370 18550 41372
rect 18606 41370 18630 41372
rect 18686 41370 18710 41372
rect 18766 41370 18790 41372
rect 18846 41370 18852 41372
rect 18606 41318 18608 41370
rect 18788 41318 18790 41370
rect 18544 41316 18550 41318
rect 18606 41316 18630 41318
rect 18686 41316 18710 41318
rect 18766 41316 18790 41318
rect 18846 41316 18852 41318
rect 18544 41307 18852 41316
rect 18544 40284 18852 40293
rect 18544 40282 18550 40284
rect 18606 40282 18630 40284
rect 18686 40282 18710 40284
rect 18766 40282 18790 40284
rect 18846 40282 18852 40284
rect 18606 40230 18608 40282
rect 18788 40230 18790 40282
rect 18544 40228 18550 40230
rect 18606 40228 18630 40230
rect 18686 40228 18710 40230
rect 18766 40228 18790 40230
rect 18846 40228 18852 40230
rect 18544 40219 18852 40228
rect 18544 39196 18852 39205
rect 18544 39194 18550 39196
rect 18606 39194 18630 39196
rect 18686 39194 18710 39196
rect 18766 39194 18790 39196
rect 18846 39194 18852 39196
rect 18606 39142 18608 39194
rect 18788 39142 18790 39194
rect 18544 39140 18550 39142
rect 18606 39140 18630 39142
rect 18686 39140 18710 39142
rect 18766 39140 18790 39142
rect 18846 39140 18852 39142
rect 18544 39131 18852 39140
rect 18544 38108 18852 38117
rect 18544 38106 18550 38108
rect 18606 38106 18630 38108
rect 18686 38106 18710 38108
rect 18766 38106 18790 38108
rect 18846 38106 18852 38108
rect 18606 38054 18608 38106
rect 18788 38054 18790 38106
rect 18544 38052 18550 38054
rect 18606 38052 18630 38054
rect 18686 38052 18710 38054
rect 18766 38052 18790 38054
rect 18846 38052 18852 38054
rect 18544 38043 18852 38052
rect 18544 37020 18852 37029
rect 18544 37018 18550 37020
rect 18606 37018 18630 37020
rect 18686 37018 18710 37020
rect 18766 37018 18790 37020
rect 18846 37018 18852 37020
rect 18606 36966 18608 37018
rect 18788 36966 18790 37018
rect 18544 36964 18550 36966
rect 18606 36964 18630 36966
rect 18686 36964 18710 36966
rect 18766 36964 18790 36966
rect 18846 36964 18852 36966
rect 18544 36955 18852 36964
rect 18544 35932 18852 35941
rect 18544 35930 18550 35932
rect 18606 35930 18630 35932
rect 18686 35930 18710 35932
rect 18766 35930 18790 35932
rect 18846 35930 18852 35932
rect 18606 35878 18608 35930
rect 18788 35878 18790 35930
rect 18544 35876 18550 35878
rect 18606 35876 18630 35878
rect 18686 35876 18710 35878
rect 18766 35876 18790 35878
rect 18846 35876 18852 35878
rect 18544 35867 18852 35876
rect 18544 34844 18852 34853
rect 18544 34842 18550 34844
rect 18606 34842 18630 34844
rect 18686 34842 18710 34844
rect 18766 34842 18790 34844
rect 18846 34842 18852 34844
rect 18606 34790 18608 34842
rect 18788 34790 18790 34842
rect 18544 34788 18550 34790
rect 18606 34788 18630 34790
rect 18686 34788 18710 34790
rect 18766 34788 18790 34790
rect 18846 34788 18852 34790
rect 18544 34779 18852 34788
rect 18892 34610 18920 41806
rect 19340 41812 19392 41818
rect 19340 41754 19392 41760
rect 19444 41614 19472 42191
rect 19536 41993 19564 42570
rect 19522 41984 19578 41993
rect 19522 41919 19578 41928
rect 19432 41608 19484 41614
rect 19432 41550 19484 41556
rect 19340 41540 19392 41546
rect 19340 41482 19392 41488
rect 19248 41132 19300 41138
rect 19248 41074 19300 41080
rect 19260 40730 19288 41074
rect 19248 40724 19300 40730
rect 19248 40666 19300 40672
rect 19352 40186 19380 41482
rect 19432 41472 19484 41478
rect 19616 41472 19668 41478
rect 19432 41414 19484 41420
rect 19614 41440 19616 41449
rect 19668 41440 19670 41449
rect 19340 40180 19392 40186
rect 19340 40122 19392 40128
rect 19340 36576 19392 36582
rect 19340 36518 19392 36524
rect 19352 36145 19380 36518
rect 19338 36136 19394 36145
rect 19338 36071 19394 36080
rect 19340 35692 19392 35698
rect 19340 35634 19392 35640
rect 19248 35284 19300 35290
rect 19248 35226 19300 35232
rect 19156 35080 19208 35086
rect 19156 35022 19208 35028
rect 19168 34678 19196 35022
rect 19156 34672 19208 34678
rect 19156 34614 19208 34620
rect 18880 34604 18932 34610
rect 18880 34546 18932 34552
rect 18544 33756 18852 33765
rect 18544 33754 18550 33756
rect 18606 33754 18630 33756
rect 18686 33754 18710 33756
rect 18766 33754 18790 33756
rect 18846 33754 18852 33756
rect 18606 33702 18608 33754
rect 18788 33702 18790 33754
rect 18544 33700 18550 33702
rect 18606 33700 18630 33702
rect 18686 33700 18710 33702
rect 18766 33700 18790 33702
rect 18846 33700 18852 33702
rect 18544 33691 18852 33700
rect 18892 33522 18920 34546
rect 18880 33516 18932 33522
rect 18880 33458 18932 33464
rect 18544 32668 18852 32677
rect 18544 32666 18550 32668
rect 18606 32666 18630 32668
rect 18686 32666 18710 32668
rect 18766 32666 18790 32668
rect 18846 32666 18852 32668
rect 18606 32614 18608 32666
rect 18788 32614 18790 32666
rect 18544 32612 18550 32614
rect 18606 32612 18630 32614
rect 18686 32612 18710 32614
rect 18766 32612 18790 32614
rect 18846 32612 18852 32614
rect 18544 32603 18852 32612
rect 18892 32434 18920 33458
rect 19064 33108 19116 33114
rect 19064 33050 19116 33056
rect 18880 32428 18932 32434
rect 18880 32370 18932 32376
rect 18892 32026 18920 32370
rect 18880 32020 18932 32026
rect 18880 31962 18932 31968
rect 18788 31816 18840 31822
rect 18786 31784 18788 31793
rect 18840 31784 18842 31793
rect 18786 31719 18842 31728
rect 18544 31580 18852 31589
rect 18544 31578 18550 31580
rect 18606 31578 18630 31580
rect 18686 31578 18710 31580
rect 18766 31578 18790 31580
rect 18846 31578 18852 31580
rect 18606 31526 18608 31578
rect 18788 31526 18790 31578
rect 18544 31524 18550 31526
rect 18606 31524 18630 31526
rect 18686 31524 18710 31526
rect 18766 31524 18790 31526
rect 18846 31524 18852 31526
rect 18544 31515 18852 31524
rect 18892 31414 18920 31962
rect 18972 31816 19024 31822
rect 18972 31758 19024 31764
rect 18984 31482 19012 31758
rect 18972 31476 19024 31482
rect 18972 31418 19024 31424
rect 18880 31408 18932 31414
rect 18880 31350 18932 31356
rect 19076 31346 19104 33050
rect 19260 32910 19288 35226
rect 19248 32904 19300 32910
rect 19248 32846 19300 32852
rect 19156 32428 19208 32434
rect 19156 32370 19208 32376
rect 19168 31890 19196 32370
rect 19156 31884 19208 31890
rect 19156 31826 19208 31832
rect 19260 31770 19288 32846
rect 19352 32570 19380 35634
rect 19340 32564 19392 32570
rect 19340 32506 19392 32512
rect 19168 31742 19288 31770
rect 19338 31784 19394 31793
rect 19064 31340 19116 31346
rect 19064 31282 19116 31288
rect 18420 31272 18472 31278
rect 18420 31214 18472 31220
rect 18248 26880 18368 26908
rect 18144 23044 18196 23050
rect 18144 22986 18196 22992
rect 18052 21480 18104 21486
rect 18052 21422 18104 21428
rect 17960 21412 18012 21418
rect 17960 21354 18012 21360
rect 17684 21140 17736 21146
rect 17684 21082 17736 21088
rect 17868 21140 17920 21146
rect 17868 21082 17920 21088
rect 17960 20800 18012 20806
rect 17960 20742 18012 20748
rect 17774 19408 17830 19417
rect 17774 19343 17830 19352
rect 17684 19304 17736 19310
rect 17684 19246 17736 19252
rect 17696 18902 17724 19246
rect 17684 18896 17736 18902
rect 17684 18838 17736 18844
rect 17684 18692 17736 18698
rect 17684 18634 17736 18640
rect 17696 18426 17724 18634
rect 17684 18420 17736 18426
rect 17684 18362 17736 18368
rect 17684 18216 17736 18222
rect 17604 18164 17684 18170
rect 17604 18158 17736 18164
rect 17604 18142 17724 18158
rect 17500 14408 17552 14414
rect 17500 14350 17552 14356
rect 17316 13184 17368 13190
rect 17316 13126 17368 13132
rect 17328 12986 17356 13126
rect 17316 12980 17368 12986
rect 17316 12922 17368 12928
rect 17408 12844 17460 12850
rect 17512 12832 17540 14350
rect 17460 12804 17540 12832
rect 17408 12786 17460 12792
rect 17604 12434 17632 18142
rect 17684 15904 17736 15910
rect 17684 15846 17736 15852
rect 17696 14414 17724 15846
rect 17684 14408 17736 14414
rect 17684 14350 17736 14356
rect 17696 14278 17724 14350
rect 17684 14272 17736 14278
rect 17684 14214 17736 14220
rect 17684 13728 17736 13734
rect 17684 13670 17736 13676
rect 17696 13394 17724 13670
rect 17684 13388 17736 13394
rect 17684 13330 17736 13336
rect 17512 12406 17632 12434
rect 17316 11552 17368 11558
rect 17316 11494 17368 11500
rect 17328 11234 17356 11494
rect 17328 11218 17448 11234
rect 17328 11212 17460 11218
rect 17328 11206 17408 11212
rect 17408 11154 17460 11160
rect 17408 11076 17460 11082
rect 17408 11018 17460 11024
rect 17420 10713 17448 11018
rect 17406 10704 17462 10713
rect 17406 10639 17462 10648
rect 17224 9920 17276 9926
rect 17224 9862 17276 9868
rect 17314 9616 17370 9625
rect 17314 9551 17316 9560
rect 17368 9551 17370 9560
rect 17316 9522 17368 9528
rect 17328 8498 17356 9522
rect 17408 9376 17460 9382
rect 17408 9318 17460 9324
rect 17316 8492 17368 8498
rect 17316 8434 17368 8440
rect 17316 7744 17368 7750
rect 17316 7686 17368 7692
rect 16580 7540 16632 7546
rect 16580 7482 16632 7488
rect 16776 7534 16988 7562
rect 17052 7534 17172 7562
rect 16488 7404 16540 7410
rect 16488 7346 16540 7352
rect 16396 6996 16448 7002
rect 16396 6938 16448 6944
rect 16304 6248 16356 6254
rect 16304 6190 16356 6196
rect 16212 6180 16264 6186
rect 16212 6122 16264 6128
rect 16082 3726 16160 3754
rect 16026 3703 16082 3712
rect 15612 2748 15920 2757
rect 15612 2746 15618 2748
rect 15674 2746 15698 2748
rect 15754 2746 15778 2748
rect 15834 2746 15858 2748
rect 15914 2746 15920 2748
rect 15674 2694 15676 2746
rect 15856 2694 15858 2746
rect 15612 2692 15618 2694
rect 15674 2692 15698 2694
rect 15754 2692 15778 2694
rect 15834 2692 15858 2694
rect 15914 2692 15920 2694
rect 15612 2683 15920 2692
rect 16224 2650 16252 6122
rect 16316 5710 16344 6190
rect 16396 6112 16448 6118
rect 16396 6054 16448 6060
rect 16304 5704 16356 5710
rect 16304 5646 16356 5652
rect 16212 2644 16264 2650
rect 16212 2586 16264 2592
rect 16408 2553 16436 6054
rect 16488 3120 16540 3126
rect 16486 3088 16488 3097
rect 16540 3088 16542 3097
rect 16486 3023 16542 3032
rect 16394 2544 16450 2553
rect 16394 2479 16450 2488
rect 16488 2440 16540 2446
rect 15750 2408 15806 2417
rect 16488 2382 16540 2388
rect 15750 2343 15752 2352
rect 15804 2343 15806 2352
rect 15752 2314 15804 2320
rect 16120 2304 16172 2310
rect 16120 2246 16172 2252
rect 15384 2032 15436 2038
rect 15384 1974 15436 1980
rect 16028 1964 16080 1970
rect 16028 1906 16080 1912
rect 15292 1760 15344 1766
rect 15292 1702 15344 1708
rect 15936 1760 15988 1766
rect 15936 1702 15988 1708
rect 14924 1488 14976 1494
rect 14924 1430 14976 1436
rect 14648 604 14700 610
rect 14648 546 14700 552
rect 12806 54 13032 82
rect 12806 -300 12862 54
rect 13082 -300 13138 160
rect 13358 -300 13414 160
rect 13634 -300 13690 160
rect 13910 -300 13966 160
rect 14186 -300 14242 160
rect 14462 -300 14518 160
rect 14738 82 14794 160
rect 14936 82 14964 1430
rect 15200 1352 15252 1358
rect 15198 1320 15200 1329
rect 15252 1320 15254 1329
rect 15198 1255 15254 1264
rect 15108 1216 15160 1222
rect 15108 1158 15160 1164
rect 14738 54 14964 82
rect 15014 82 15070 160
rect 15120 82 15148 1158
rect 15304 160 15332 1702
rect 15612 1660 15920 1669
rect 15612 1658 15618 1660
rect 15674 1658 15698 1660
rect 15754 1658 15778 1660
rect 15834 1658 15858 1660
rect 15914 1658 15920 1660
rect 15674 1606 15676 1658
rect 15856 1606 15858 1658
rect 15612 1604 15618 1606
rect 15674 1604 15698 1606
rect 15754 1604 15778 1606
rect 15834 1604 15858 1606
rect 15914 1604 15920 1606
rect 15612 1595 15920 1604
rect 15948 1544 15976 1702
rect 16040 1562 16068 1906
rect 15764 1516 15976 1544
rect 16028 1556 16080 1562
rect 15014 54 15148 82
rect 14738 -300 14794 54
rect 15014 -300 15070 54
rect 15290 -300 15346 160
rect 15566 82 15622 160
rect 15764 82 15792 1516
rect 16028 1498 16080 1504
rect 15844 1420 15896 1426
rect 15844 1362 15896 1368
rect 15856 160 15884 1362
rect 16132 1358 16160 2246
rect 16304 1964 16356 1970
rect 16304 1906 16356 1912
rect 16120 1352 16172 1358
rect 16120 1294 16172 1300
rect 15566 54 15792 82
rect 15566 -300 15622 54
rect 15842 -300 15898 160
rect 16118 82 16174 160
rect 16316 82 16344 1906
rect 16396 1760 16448 1766
rect 16396 1702 16448 1708
rect 16408 160 16436 1702
rect 16500 1562 16528 2382
rect 16488 1556 16540 1562
rect 16488 1498 16540 1504
rect 16488 1352 16540 1358
rect 16488 1294 16540 1300
rect 16500 542 16528 1294
rect 16592 814 16620 7482
rect 16672 6248 16724 6254
rect 16672 6190 16724 6196
rect 16684 5778 16712 6190
rect 16672 5772 16724 5778
rect 16672 5714 16724 5720
rect 16672 2304 16724 2310
rect 16672 2246 16724 2252
rect 16684 2106 16712 2246
rect 16672 2100 16724 2106
rect 16672 2042 16724 2048
rect 16672 1828 16724 1834
rect 16672 1770 16724 1776
rect 16580 808 16632 814
rect 16580 750 16632 756
rect 16488 536 16540 542
rect 16488 478 16540 484
rect 16684 160 16712 1770
rect 16776 1358 16804 7534
rect 16948 7404 17000 7410
rect 16948 7346 17000 7352
rect 16960 7002 16988 7346
rect 16948 6996 17000 7002
rect 16948 6938 17000 6944
rect 16948 3460 17000 3466
rect 16948 3402 17000 3408
rect 16960 3194 16988 3402
rect 16948 3188 17000 3194
rect 16948 3130 17000 3136
rect 16854 2680 16910 2689
rect 16854 2615 16910 2624
rect 16868 2446 16896 2615
rect 17052 2514 17080 7534
rect 17224 7336 17276 7342
rect 17224 7278 17276 7284
rect 17132 7200 17184 7206
rect 17132 7142 17184 7148
rect 17144 7002 17172 7142
rect 17132 6996 17184 7002
rect 17132 6938 17184 6944
rect 17236 6458 17264 7278
rect 17224 6452 17276 6458
rect 17224 6394 17276 6400
rect 17132 4208 17184 4214
rect 17132 4150 17184 4156
rect 17144 3058 17172 4150
rect 17222 3632 17278 3641
rect 17222 3567 17224 3576
rect 17276 3567 17278 3576
rect 17224 3538 17276 3544
rect 17132 3052 17184 3058
rect 17132 2994 17184 3000
rect 17224 2916 17276 2922
rect 17224 2858 17276 2864
rect 17130 2680 17186 2689
rect 17130 2615 17186 2624
rect 17040 2508 17092 2514
rect 17040 2450 17092 2456
rect 17144 2446 17172 2615
rect 16856 2440 16908 2446
rect 16856 2382 16908 2388
rect 17132 2440 17184 2446
rect 17132 2382 17184 2388
rect 17236 2378 17264 2858
rect 17224 2372 17276 2378
rect 17224 2314 17276 2320
rect 16948 2304 17000 2310
rect 16948 2246 17000 2252
rect 16960 2106 16988 2246
rect 16948 2100 17000 2106
rect 16948 2042 17000 2048
rect 17132 2032 17184 2038
rect 17328 1986 17356 7686
rect 17420 5778 17448 9318
rect 17512 8974 17540 12406
rect 17684 9580 17736 9586
rect 17684 9522 17736 9528
rect 17592 9172 17644 9178
rect 17592 9114 17644 9120
rect 17500 8968 17552 8974
rect 17500 8910 17552 8916
rect 17498 5808 17554 5817
rect 17408 5772 17460 5778
rect 17498 5743 17554 5752
rect 17408 5714 17460 5720
rect 17406 5536 17462 5545
rect 17406 5471 17462 5480
rect 17420 3058 17448 5471
rect 17512 3058 17540 5743
rect 17604 4729 17632 9114
rect 17696 8974 17724 9522
rect 17684 8968 17736 8974
rect 17684 8910 17736 8916
rect 17696 6780 17724 8910
rect 17788 7546 17816 19343
rect 17868 19304 17920 19310
rect 17868 19246 17920 19252
rect 17880 18290 17908 19246
rect 17868 18284 17920 18290
rect 17868 18226 17920 18232
rect 17880 17882 17908 18226
rect 17868 17876 17920 17882
rect 17868 17818 17920 17824
rect 17972 17678 18000 20742
rect 18156 19553 18184 22986
rect 18142 19544 18198 19553
rect 18142 19479 18144 19488
rect 18196 19479 18198 19488
rect 18144 19450 18196 19456
rect 18052 18828 18104 18834
rect 18052 18770 18104 18776
rect 18064 18086 18092 18770
rect 18144 18760 18196 18766
rect 18144 18702 18196 18708
rect 18052 18080 18104 18086
rect 18052 18022 18104 18028
rect 17960 17672 18012 17678
rect 17960 17614 18012 17620
rect 17960 17128 18012 17134
rect 17960 17070 18012 17076
rect 17972 16658 18000 17070
rect 17960 16652 18012 16658
rect 17960 16594 18012 16600
rect 17972 14822 18000 16594
rect 18052 15360 18104 15366
rect 18052 15302 18104 15308
rect 17960 14816 18012 14822
rect 17960 14758 18012 14764
rect 17972 11762 18000 14758
rect 18064 14074 18092 15302
rect 18156 15162 18184 18702
rect 18144 15156 18196 15162
rect 18144 15098 18196 15104
rect 18144 14340 18196 14346
rect 18144 14282 18196 14288
rect 18156 14074 18184 14282
rect 18052 14068 18104 14074
rect 18052 14010 18104 14016
rect 18144 14068 18196 14074
rect 18144 14010 18196 14016
rect 18052 12640 18104 12646
rect 18052 12582 18104 12588
rect 18064 12434 18092 12582
rect 18064 12406 18184 12434
rect 18156 12238 18184 12406
rect 18052 12232 18104 12238
rect 18052 12174 18104 12180
rect 18144 12232 18196 12238
rect 18144 12174 18196 12180
rect 17960 11756 18012 11762
rect 17960 11698 18012 11704
rect 17868 9716 17920 9722
rect 17868 9658 17920 9664
rect 17880 8294 17908 9658
rect 17972 9586 18000 11698
rect 18064 11354 18092 12174
rect 18144 12096 18196 12102
rect 18144 12038 18196 12044
rect 18156 11762 18184 12038
rect 18144 11756 18196 11762
rect 18144 11698 18196 11704
rect 18052 11348 18104 11354
rect 18052 11290 18104 11296
rect 18248 11082 18276 26880
rect 18432 26738 18460 31214
rect 18544 30492 18852 30501
rect 18544 30490 18550 30492
rect 18606 30490 18630 30492
rect 18686 30490 18710 30492
rect 18766 30490 18790 30492
rect 18846 30490 18852 30492
rect 18606 30438 18608 30490
rect 18788 30438 18790 30490
rect 18544 30436 18550 30438
rect 18606 30436 18630 30438
rect 18686 30436 18710 30438
rect 18766 30436 18790 30438
rect 18846 30436 18852 30438
rect 18544 30427 18852 30436
rect 18880 29640 18932 29646
rect 18880 29582 18932 29588
rect 18544 29404 18852 29413
rect 18544 29402 18550 29404
rect 18606 29402 18630 29404
rect 18686 29402 18710 29404
rect 18766 29402 18790 29404
rect 18846 29402 18852 29404
rect 18606 29350 18608 29402
rect 18788 29350 18790 29402
rect 18544 29348 18550 29350
rect 18606 29348 18630 29350
rect 18686 29348 18710 29350
rect 18766 29348 18790 29350
rect 18846 29348 18852 29350
rect 18544 29339 18852 29348
rect 18544 28316 18852 28325
rect 18544 28314 18550 28316
rect 18606 28314 18630 28316
rect 18686 28314 18710 28316
rect 18766 28314 18790 28316
rect 18846 28314 18852 28316
rect 18606 28262 18608 28314
rect 18788 28262 18790 28314
rect 18544 28260 18550 28262
rect 18606 28260 18630 28262
rect 18686 28260 18710 28262
rect 18766 28260 18790 28262
rect 18846 28260 18852 28262
rect 18544 28251 18852 28260
rect 18892 28098 18920 29582
rect 18972 29028 19024 29034
rect 18972 28970 19024 28976
rect 18984 28506 19012 28970
rect 18984 28478 19104 28506
rect 18972 28416 19024 28422
rect 18972 28358 19024 28364
rect 18984 28218 19012 28358
rect 18972 28212 19024 28218
rect 18972 28154 19024 28160
rect 18892 28070 19012 28098
rect 18604 28008 18656 28014
rect 18604 27950 18656 27956
rect 18616 27674 18644 27950
rect 18604 27668 18656 27674
rect 18604 27610 18656 27616
rect 18544 27228 18852 27237
rect 18544 27226 18550 27228
rect 18606 27226 18630 27228
rect 18686 27226 18710 27228
rect 18766 27226 18790 27228
rect 18846 27226 18852 27228
rect 18606 27174 18608 27226
rect 18788 27174 18790 27226
rect 18544 27172 18550 27174
rect 18606 27172 18630 27174
rect 18686 27172 18710 27174
rect 18766 27172 18790 27174
rect 18846 27172 18852 27174
rect 18544 27163 18852 27172
rect 18340 26710 18460 26738
rect 18340 25786 18368 26710
rect 18420 26376 18472 26382
rect 18420 26318 18472 26324
rect 18432 25974 18460 26318
rect 18544 26140 18852 26149
rect 18544 26138 18550 26140
rect 18606 26138 18630 26140
rect 18686 26138 18710 26140
rect 18766 26138 18790 26140
rect 18846 26138 18852 26140
rect 18606 26086 18608 26138
rect 18788 26086 18790 26138
rect 18544 26084 18550 26086
rect 18606 26084 18630 26086
rect 18686 26084 18710 26086
rect 18766 26084 18790 26086
rect 18846 26084 18852 26086
rect 18544 26075 18852 26084
rect 18420 25968 18472 25974
rect 18420 25910 18472 25916
rect 18340 25758 18460 25786
rect 18328 24744 18380 24750
rect 18328 24686 18380 24692
rect 18340 24410 18368 24686
rect 18328 24404 18380 24410
rect 18328 24346 18380 24352
rect 18432 24290 18460 25758
rect 18544 25052 18852 25061
rect 18544 25050 18550 25052
rect 18606 25050 18630 25052
rect 18686 25050 18710 25052
rect 18766 25050 18790 25052
rect 18846 25050 18852 25052
rect 18606 24998 18608 25050
rect 18788 24998 18790 25050
rect 18544 24996 18550 24998
rect 18606 24996 18630 24998
rect 18686 24996 18710 24998
rect 18766 24996 18790 24998
rect 18846 24996 18852 24998
rect 18544 24987 18852 24996
rect 18788 24608 18840 24614
rect 18788 24550 18840 24556
rect 18340 24262 18460 24290
rect 18340 21978 18368 24262
rect 18800 24154 18828 24550
rect 18800 24126 18920 24154
rect 18544 23964 18852 23973
rect 18544 23962 18550 23964
rect 18606 23962 18630 23964
rect 18686 23962 18710 23964
rect 18766 23962 18790 23964
rect 18846 23962 18852 23964
rect 18606 23910 18608 23962
rect 18788 23910 18790 23962
rect 18544 23908 18550 23910
rect 18606 23908 18630 23910
rect 18686 23908 18710 23910
rect 18766 23908 18790 23910
rect 18846 23908 18852 23910
rect 18544 23899 18852 23908
rect 18788 23724 18840 23730
rect 18892 23712 18920 24126
rect 18840 23684 18920 23712
rect 18788 23666 18840 23672
rect 18420 23656 18472 23662
rect 18418 23624 18420 23633
rect 18472 23624 18474 23633
rect 18418 23559 18474 23568
rect 18420 23520 18472 23526
rect 18420 23462 18472 23468
rect 18432 22642 18460 23462
rect 18544 22876 18852 22885
rect 18544 22874 18550 22876
rect 18606 22874 18630 22876
rect 18686 22874 18710 22876
rect 18766 22874 18790 22876
rect 18846 22874 18852 22876
rect 18606 22822 18608 22874
rect 18788 22822 18790 22874
rect 18544 22820 18550 22822
rect 18606 22820 18630 22822
rect 18686 22820 18710 22822
rect 18766 22820 18790 22822
rect 18846 22820 18852 22822
rect 18544 22811 18852 22820
rect 18420 22636 18472 22642
rect 18420 22578 18472 22584
rect 18432 22094 18460 22578
rect 18984 22094 19012 28070
rect 18432 22066 18552 22094
rect 18524 22030 18552 22066
rect 18892 22066 19012 22094
rect 18512 22024 18564 22030
rect 18340 21950 18460 21978
rect 18512 21966 18564 21972
rect 18328 21888 18380 21894
rect 18328 21830 18380 21836
rect 18340 21146 18368 21830
rect 18432 21690 18460 21950
rect 18544 21788 18852 21797
rect 18544 21786 18550 21788
rect 18606 21786 18630 21788
rect 18686 21786 18710 21788
rect 18766 21786 18790 21788
rect 18846 21786 18852 21788
rect 18606 21734 18608 21786
rect 18788 21734 18790 21786
rect 18544 21732 18550 21734
rect 18606 21732 18630 21734
rect 18686 21732 18710 21734
rect 18766 21732 18790 21734
rect 18846 21732 18852 21734
rect 18544 21723 18852 21732
rect 18420 21684 18472 21690
rect 18472 21644 18552 21672
rect 18420 21626 18472 21632
rect 18524 21350 18552 21644
rect 18892 21418 18920 22066
rect 18972 21888 19024 21894
rect 18972 21830 19024 21836
rect 18984 21690 19012 21830
rect 18972 21684 19024 21690
rect 18972 21626 19024 21632
rect 18880 21412 18932 21418
rect 18880 21354 18932 21360
rect 18420 21344 18472 21350
rect 18420 21286 18472 21292
rect 18512 21344 18564 21350
rect 18512 21286 18564 21292
rect 18328 21140 18380 21146
rect 18328 21082 18380 21088
rect 18432 19825 18460 21286
rect 18880 20800 18932 20806
rect 18880 20742 18932 20748
rect 18544 20700 18852 20709
rect 18544 20698 18550 20700
rect 18606 20698 18630 20700
rect 18686 20698 18710 20700
rect 18766 20698 18790 20700
rect 18846 20698 18852 20700
rect 18606 20646 18608 20698
rect 18788 20646 18790 20698
rect 18544 20644 18550 20646
rect 18606 20644 18630 20646
rect 18686 20644 18710 20646
rect 18766 20644 18790 20646
rect 18846 20644 18852 20646
rect 18544 20635 18852 20644
rect 18892 20618 18920 20742
rect 18892 20590 19012 20618
rect 18880 20460 18932 20466
rect 18880 20402 18932 20408
rect 18892 20058 18920 20402
rect 18880 20052 18932 20058
rect 18880 19994 18932 20000
rect 18880 19848 18932 19854
rect 18418 19816 18474 19825
rect 18880 19790 18932 19796
rect 18418 19751 18474 19760
rect 18432 19334 18460 19751
rect 18544 19612 18852 19621
rect 18544 19610 18550 19612
rect 18606 19610 18630 19612
rect 18686 19610 18710 19612
rect 18766 19610 18790 19612
rect 18846 19610 18852 19612
rect 18606 19558 18608 19610
rect 18788 19558 18790 19610
rect 18544 19556 18550 19558
rect 18606 19556 18630 19558
rect 18686 19556 18710 19558
rect 18766 19556 18790 19558
rect 18846 19556 18852 19558
rect 18544 19547 18852 19556
rect 18892 19514 18920 19790
rect 18880 19508 18932 19514
rect 18880 19450 18932 19456
rect 18432 19310 18644 19334
rect 18432 19306 18656 19310
rect 18604 19304 18656 19306
rect 18604 19246 18656 19252
rect 18512 19168 18564 19174
rect 18512 19110 18564 19116
rect 18524 18834 18552 19110
rect 18512 18828 18564 18834
rect 18512 18770 18564 18776
rect 18420 18760 18472 18766
rect 18420 18702 18472 18708
rect 18328 18624 18380 18630
rect 18328 18566 18380 18572
rect 18340 16130 18368 18566
rect 18432 18426 18460 18702
rect 18544 18524 18852 18533
rect 18544 18522 18550 18524
rect 18606 18522 18630 18524
rect 18686 18522 18710 18524
rect 18766 18522 18790 18524
rect 18846 18522 18852 18524
rect 18606 18470 18608 18522
rect 18788 18470 18790 18522
rect 18544 18468 18550 18470
rect 18606 18468 18630 18470
rect 18686 18468 18710 18470
rect 18766 18468 18790 18470
rect 18846 18468 18852 18470
rect 18544 18459 18852 18468
rect 18420 18420 18472 18426
rect 18420 18362 18472 18368
rect 18544 17436 18852 17445
rect 18544 17434 18550 17436
rect 18606 17434 18630 17436
rect 18686 17434 18710 17436
rect 18766 17434 18790 17436
rect 18846 17434 18852 17436
rect 18606 17382 18608 17434
rect 18788 17382 18790 17434
rect 18544 17380 18550 17382
rect 18606 17380 18630 17382
rect 18686 17380 18710 17382
rect 18766 17380 18790 17382
rect 18846 17380 18852 17382
rect 18544 17371 18852 17380
rect 18892 17134 18920 19450
rect 18984 19334 19012 20590
rect 19076 19854 19104 28478
rect 19168 26994 19196 31742
rect 19338 31719 19394 31728
rect 19248 31340 19300 31346
rect 19248 31282 19300 31288
rect 19260 30818 19288 31282
rect 19352 30938 19380 31719
rect 19340 30932 19392 30938
rect 19340 30874 19392 30880
rect 19260 30790 19380 30818
rect 19248 29572 19300 29578
rect 19248 29514 19300 29520
rect 19260 29238 19288 29514
rect 19248 29232 19300 29238
rect 19248 29174 19300 29180
rect 19352 27334 19380 30790
rect 19340 27328 19392 27334
rect 19340 27270 19392 27276
rect 19156 26988 19208 26994
rect 19156 26930 19208 26936
rect 19340 25764 19392 25770
rect 19340 25706 19392 25712
rect 19156 24812 19208 24818
rect 19156 24754 19208 24760
rect 19168 24410 19196 24754
rect 19248 24608 19300 24614
rect 19248 24550 19300 24556
rect 19156 24404 19208 24410
rect 19156 24346 19208 24352
rect 19168 23594 19196 24346
rect 19260 23662 19288 24550
rect 19352 23662 19380 25706
rect 19248 23656 19300 23662
rect 19248 23598 19300 23604
rect 19340 23656 19392 23662
rect 19340 23598 19392 23604
rect 19156 23588 19208 23594
rect 19156 23530 19208 23536
rect 19352 23186 19380 23598
rect 19340 23180 19392 23186
rect 19340 23122 19392 23128
rect 19352 22794 19380 23122
rect 19168 22766 19380 22794
rect 19168 22166 19196 22766
rect 19248 22704 19300 22710
rect 19248 22646 19300 22652
rect 19156 22160 19208 22166
rect 19156 22102 19208 22108
rect 19156 21888 19208 21894
rect 19156 21830 19208 21836
rect 19168 21690 19196 21830
rect 19156 21684 19208 21690
rect 19156 21626 19208 21632
rect 19168 21146 19196 21626
rect 19156 21140 19208 21146
rect 19156 21082 19208 21088
rect 19260 20924 19288 22646
rect 19340 21888 19392 21894
rect 19340 21830 19392 21836
rect 19352 21554 19380 21830
rect 19340 21548 19392 21554
rect 19340 21490 19392 21496
rect 19340 20936 19392 20942
rect 19260 20896 19340 20924
rect 19260 19922 19288 20896
rect 19340 20878 19392 20884
rect 19248 19916 19300 19922
rect 19248 19858 19300 19864
rect 19064 19848 19116 19854
rect 19064 19790 19116 19796
rect 18984 19306 19104 19334
rect 18880 17128 18932 17134
rect 18880 17070 18932 17076
rect 18420 16584 18472 16590
rect 18420 16526 18472 16532
rect 18880 16584 18932 16590
rect 18880 16526 18932 16532
rect 18432 16250 18460 16526
rect 18544 16348 18852 16357
rect 18544 16346 18550 16348
rect 18606 16346 18630 16348
rect 18686 16346 18710 16348
rect 18766 16346 18790 16348
rect 18846 16346 18852 16348
rect 18606 16294 18608 16346
rect 18788 16294 18790 16346
rect 18544 16292 18550 16294
rect 18606 16292 18630 16294
rect 18686 16292 18710 16294
rect 18766 16292 18790 16294
rect 18846 16292 18852 16294
rect 18544 16283 18852 16292
rect 18420 16244 18472 16250
rect 18420 16186 18472 16192
rect 18892 16182 18920 16526
rect 18880 16176 18932 16182
rect 18340 16102 18460 16130
rect 18880 16118 18932 16124
rect 18328 14816 18380 14822
rect 18328 14758 18380 14764
rect 18340 14074 18368 14758
rect 18328 14068 18380 14074
rect 18328 14010 18380 14016
rect 18328 13796 18380 13802
rect 18328 13738 18380 13744
rect 18236 11076 18288 11082
rect 18236 11018 18288 11024
rect 18052 11008 18104 11014
rect 18052 10950 18104 10956
rect 18064 9654 18092 10950
rect 18340 10742 18368 13738
rect 18328 10736 18380 10742
rect 18328 10678 18380 10684
rect 18144 10056 18196 10062
rect 18144 9998 18196 10004
rect 18236 10056 18288 10062
rect 18236 9998 18288 10004
rect 18328 10056 18380 10062
rect 18328 9998 18380 10004
rect 18052 9648 18104 9654
rect 18052 9590 18104 9596
rect 17960 9580 18012 9586
rect 17960 9522 18012 9528
rect 18156 9382 18184 9998
rect 18144 9376 18196 9382
rect 18144 9318 18196 9324
rect 18050 8936 18106 8945
rect 18050 8871 18106 8880
rect 17868 8288 17920 8294
rect 17868 8230 17920 8236
rect 17776 7540 17828 7546
rect 17776 7482 17828 7488
rect 17776 6792 17828 6798
rect 17696 6752 17776 6780
rect 17776 6734 17828 6740
rect 17788 6254 17816 6734
rect 18064 6610 18092 8871
rect 18156 8498 18184 9318
rect 18248 8634 18276 9998
rect 18340 8634 18368 9998
rect 18236 8628 18288 8634
rect 18236 8570 18288 8576
rect 18328 8628 18380 8634
rect 18328 8570 18380 8576
rect 18144 8492 18196 8498
rect 18144 8434 18196 8440
rect 18144 7404 18196 7410
rect 18144 7346 18196 7352
rect 17972 6582 18092 6610
rect 17776 6248 17828 6254
rect 17776 6190 17828 6196
rect 17776 5772 17828 5778
rect 17776 5714 17828 5720
rect 17684 5636 17736 5642
rect 17684 5578 17736 5584
rect 17590 4720 17646 4729
rect 17590 4655 17646 4664
rect 17604 4622 17632 4655
rect 17592 4616 17644 4622
rect 17592 4558 17644 4564
rect 17696 3738 17724 5578
rect 17788 5574 17816 5714
rect 17776 5568 17828 5574
rect 17776 5510 17828 5516
rect 17776 4480 17828 4486
rect 17776 4422 17828 4428
rect 17788 4146 17816 4422
rect 17776 4140 17828 4146
rect 17776 4082 17828 4088
rect 17868 4140 17920 4146
rect 17868 4082 17920 4088
rect 17684 3732 17736 3738
rect 17684 3674 17736 3680
rect 17788 3602 17816 4082
rect 17880 3738 17908 4082
rect 17868 3732 17920 3738
rect 17868 3674 17920 3680
rect 17776 3596 17828 3602
rect 17776 3538 17828 3544
rect 17592 3528 17644 3534
rect 17592 3470 17644 3476
rect 17684 3528 17736 3534
rect 17684 3470 17736 3476
rect 17604 3058 17632 3470
rect 17696 3194 17724 3470
rect 17684 3188 17736 3194
rect 17684 3130 17736 3136
rect 17774 3088 17830 3097
rect 17408 3052 17460 3058
rect 17408 2994 17460 3000
rect 17500 3052 17552 3058
rect 17500 2994 17552 3000
rect 17592 3052 17644 3058
rect 17774 3023 17830 3032
rect 17592 2994 17644 3000
rect 17408 2848 17460 2854
rect 17408 2790 17460 2796
rect 17500 2848 17552 2854
rect 17500 2790 17552 2796
rect 17420 2038 17448 2790
rect 17132 1974 17184 1980
rect 16948 1760 17000 1766
rect 16948 1702 17000 1708
rect 16764 1352 16816 1358
rect 16764 1294 16816 1300
rect 16960 160 16988 1702
rect 17144 882 17172 1974
rect 17236 1958 17356 1986
rect 17408 2032 17460 2038
rect 17408 1974 17460 1980
rect 17132 876 17184 882
rect 17132 818 17184 824
rect 17236 762 17264 1958
rect 17408 1352 17460 1358
rect 17408 1294 17460 1300
rect 17144 746 17264 762
rect 17132 740 17264 746
rect 17184 734 17264 740
rect 17132 682 17184 688
rect 16118 54 16344 82
rect 16118 -300 16174 54
rect 16394 -300 16450 160
rect 16670 -300 16726 160
rect 16946 -300 17002 160
rect 17222 82 17278 160
rect 17420 82 17448 1294
rect 17512 160 17540 2790
rect 17684 2644 17736 2650
rect 17684 2586 17736 2592
rect 17696 1766 17724 2586
rect 17684 1760 17736 1766
rect 17684 1702 17736 1708
rect 17788 160 17816 3023
rect 17972 2650 18000 6582
rect 18156 6458 18184 7346
rect 18236 6928 18288 6934
rect 18432 6882 18460 16102
rect 18512 16108 18564 16114
rect 18512 16050 18564 16056
rect 18524 15502 18552 16050
rect 18512 15496 18564 15502
rect 18512 15438 18564 15444
rect 18544 15260 18852 15269
rect 18544 15258 18550 15260
rect 18606 15258 18630 15260
rect 18686 15258 18710 15260
rect 18766 15258 18790 15260
rect 18846 15258 18852 15260
rect 18606 15206 18608 15258
rect 18788 15206 18790 15258
rect 18544 15204 18550 15206
rect 18606 15204 18630 15206
rect 18686 15204 18710 15206
rect 18766 15204 18790 15206
rect 18846 15204 18852 15206
rect 18544 15195 18852 15204
rect 18972 15156 19024 15162
rect 18972 15098 19024 15104
rect 18696 15020 18748 15026
rect 18696 14962 18748 14968
rect 18880 15020 18932 15026
rect 18880 14962 18932 14968
rect 18708 14618 18736 14962
rect 18788 14816 18840 14822
rect 18788 14758 18840 14764
rect 18800 14618 18828 14758
rect 18696 14612 18748 14618
rect 18696 14554 18748 14560
rect 18788 14612 18840 14618
rect 18788 14554 18840 14560
rect 18544 14172 18852 14181
rect 18544 14170 18550 14172
rect 18606 14170 18630 14172
rect 18686 14170 18710 14172
rect 18766 14170 18790 14172
rect 18846 14170 18852 14172
rect 18606 14118 18608 14170
rect 18788 14118 18790 14170
rect 18544 14116 18550 14118
rect 18606 14116 18630 14118
rect 18686 14116 18710 14118
rect 18766 14116 18790 14118
rect 18846 14116 18852 14118
rect 18544 14107 18852 14116
rect 18892 14074 18920 14962
rect 18880 14068 18932 14074
rect 18880 14010 18932 14016
rect 18984 14006 19012 15098
rect 18972 14000 19024 14006
rect 18972 13942 19024 13948
rect 18544 13084 18852 13093
rect 18544 13082 18550 13084
rect 18606 13082 18630 13084
rect 18686 13082 18710 13084
rect 18766 13082 18790 13084
rect 18846 13082 18852 13084
rect 18606 13030 18608 13082
rect 18788 13030 18790 13082
rect 18544 13028 18550 13030
rect 18606 13028 18630 13030
rect 18686 13028 18710 13030
rect 18766 13028 18790 13030
rect 18846 13028 18852 13030
rect 18544 13019 18852 13028
rect 18984 12986 19012 13942
rect 18972 12980 19024 12986
rect 18972 12922 19024 12928
rect 18880 12232 18932 12238
rect 18880 12174 18932 12180
rect 18544 11996 18852 12005
rect 18544 11994 18550 11996
rect 18606 11994 18630 11996
rect 18686 11994 18710 11996
rect 18766 11994 18790 11996
rect 18846 11994 18852 11996
rect 18606 11942 18608 11994
rect 18788 11942 18790 11994
rect 18544 11940 18550 11942
rect 18606 11940 18630 11942
rect 18686 11940 18710 11942
rect 18766 11940 18790 11942
rect 18846 11940 18852 11942
rect 18544 11931 18852 11940
rect 18788 11756 18840 11762
rect 18788 11698 18840 11704
rect 18800 11626 18828 11698
rect 18788 11620 18840 11626
rect 18788 11562 18840 11568
rect 18892 11354 18920 12174
rect 18880 11348 18932 11354
rect 18880 11290 18932 11296
rect 18880 11076 18932 11082
rect 18880 11018 18932 11024
rect 18544 10908 18852 10917
rect 18544 10906 18550 10908
rect 18606 10906 18630 10908
rect 18686 10906 18710 10908
rect 18766 10906 18790 10908
rect 18846 10906 18852 10908
rect 18606 10854 18608 10906
rect 18788 10854 18790 10906
rect 18544 10852 18550 10854
rect 18606 10852 18630 10854
rect 18686 10852 18710 10854
rect 18766 10852 18790 10854
rect 18846 10852 18852 10854
rect 18544 10843 18852 10852
rect 18544 9820 18852 9829
rect 18544 9818 18550 9820
rect 18606 9818 18630 9820
rect 18686 9818 18710 9820
rect 18766 9818 18790 9820
rect 18846 9818 18852 9820
rect 18606 9766 18608 9818
rect 18788 9766 18790 9818
rect 18544 9764 18550 9766
rect 18606 9764 18630 9766
rect 18686 9764 18710 9766
rect 18766 9764 18790 9766
rect 18846 9764 18852 9766
rect 18544 9755 18852 9764
rect 18604 9512 18656 9518
rect 18510 9480 18566 9489
rect 18604 9454 18656 9460
rect 18510 9415 18566 9424
rect 18524 9382 18552 9415
rect 18512 9376 18564 9382
rect 18512 9318 18564 9324
rect 18616 9110 18644 9454
rect 18604 9104 18656 9110
rect 18604 9046 18656 9052
rect 18544 8732 18852 8741
rect 18544 8730 18550 8732
rect 18606 8730 18630 8732
rect 18686 8730 18710 8732
rect 18766 8730 18790 8732
rect 18846 8730 18852 8732
rect 18606 8678 18608 8730
rect 18788 8678 18790 8730
rect 18544 8676 18550 8678
rect 18606 8676 18630 8678
rect 18686 8676 18710 8678
rect 18766 8676 18790 8678
rect 18846 8676 18852 8678
rect 18544 8667 18852 8676
rect 18544 7644 18852 7653
rect 18544 7642 18550 7644
rect 18606 7642 18630 7644
rect 18686 7642 18710 7644
rect 18766 7642 18790 7644
rect 18846 7642 18852 7644
rect 18606 7590 18608 7642
rect 18788 7590 18790 7642
rect 18544 7588 18550 7590
rect 18606 7588 18630 7590
rect 18686 7588 18710 7590
rect 18766 7588 18790 7590
rect 18846 7588 18852 7590
rect 18544 7579 18852 7588
rect 18236 6870 18288 6876
rect 18248 6458 18276 6870
rect 18340 6854 18460 6882
rect 18144 6452 18196 6458
rect 18144 6394 18196 6400
rect 18236 6452 18288 6458
rect 18236 6394 18288 6400
rect 18052 5568 18104 5574
rect 18052 5510 18104 5516
rect 18064 4010 18092 5510
rect 18236 4616 18288 4622
rect 18236 4558 18288 4564
rect 18248 4282 18276 4558
rect 18236 4276 18288 4282
rect 18236 4218 18288 4224
rect 18236 4140 18288 4146
rect 18236 4082 18288 4088
rect 18052 4004 18104 4010
rect 18052 3946 18104 3952
rect 18248 3738 18276 4082
rect 18236 3732 18288 3738
rect 18236 3674 18288 3680
rect 18064 3454 18276 3482
rect 17960 2644 18012 2650
rect 17960 2586 18012 2592
rect 17960 2304 18012 2310
rect 17960 2246 18012 2252
rect 17972 2038 18000 2246
rect 17960 2032 18012 2038
rect 17960 1974 18012 1980
rect 17960 1216 18012 1222
rect 17960 1158 18012 1164
rect 17972 814 18000 1158
rect 17960 808 18012 814
rect 17960 750 18012 756
rect 18064 160 18092 3454
rect 18248 3398 18276 3454
rect 18144 3392 18196 3398
rect 18144 3334 18196 3340
rect 18236 3392 18288 3398
rect 18236 3334 18288 3340
rect 17222 54 17448 82
rect 17222 -300 17278 54
rect 17498 -300 17554 160
rect 17774 -300 17830 160
rect 18050 -300 18106 160
rect 18156 82 18184 3334
rect 18340 2774 18368 6854
rect 18544 6556 18852 6565
rect 18544 6554 18550 6556
rect 18606 6554 18630 6556
rect 18686 6554 18710 6556
rect 18766 6554 18790 6556
rect 18846 6554 18852 6556
rect 18606 6502 18608 6554
rect 18788 6502 18790 6554
rect 18544 6500 18550 6502
rect 18606 6500 18630 6502
rect 18686 6500 18710 6502
rect 18766 6500 18790 6502
rect 18846 6500 18852 6502
rect 18544 6491 18852 6500
rect 18604 6248 18656 6254
rect 18604 6190 18656 6196
rect 18512 6180 18564 6186
rect 18512 6122 18564 6128
rect 18524 5846 18552 6122
rect 18512 5840 18564 5846
rect 18512 5782 18564 5788
rect 18616 5778 18644 6190
rect 18604 5772 18656 5778
rect 18604 5714 18656 5720
rect 18544 5468 18852 5477
rect 18544 5466 18550 5468
rect 18606 5466 18630 5468
rect 18686 5466 18710 5468
rect 18766 5466 18790 5468
rect 18846 5466 18852 5468
rect 18606 5414 18608 5466
rect 18788 5414 18790 5466
rect 18544 5412 18550 5414
rect 18606 5412 18630 5414
rect 18686 5412 18710 5414
rect 18766 5412 18790 5414
rect 18846 5412 18852 5414
rect 18544 5403 18852 5412
rect 18420 4480 18472 4486
rect 18420 4422 18472 4428
rect 18432 3534 18460 4422
rect 18544 4380 18852 4389
rect 18544 4378 18550 4380
rect 18606 4378 18630 4380
rect 18686 4378 18710 4380
rect 18766 4378 18790 4380
rect 18846 4378 18852 4380
rect 18606 4326 18608 4378
rect 18788 4326 18790 4378
rect 18544 4324 18550 4326
rect 18606 4324 18630 4326
rect 18686 4324 18710 4326
rect 18766 4324 18790 4326
rect 18846 4324 18852 4326
rect 18544 4315 18852 4324
rect 18696 4276 18748 4282
rect 18696 4218 18748 4224
rect 18708 4146 18736 4218
rect 18696 4140 18748 4146
rect 18696 4082 18748 4088
rect 18512 4004 18564 4010
rect 18512 3946 18564 3952
rect 18420 3528 18472 3534
rect 18420 3470 18472 3476
rect 18524 3380 18552 3946
rect 18432 3352 18552 3380
rect 18432 3176 18460 3352
rect 18544 3292 18852 3301
rect 18544 3290 18550 3292
rect 18606 3290 18630 3292
rect 18686 3290 18710 3292
rect 18766 3290 18790 3292
rect 18846 3290 18852 3292
rect 18606 3238 18608 3290
rect 18788 3238 18790 3290
rect 18544 3236 18550 3238
rect 18606 3236 18630 3238
rect 18686 3236 18710 3238
rect 18766 3236 18790 3238
rect 18846 3236 18852 3238
rect 18544 3227 18852 3236
rect 18432 3148 18644 3176
rect 18420 2984 18472 2990
rect 18472 2932 18552 2938
rect 18420 2926 18552 2932
rect 18432 2910 18552 2926
rect 18340 2746 18460 2774
rect 18328 2644 18380 2650
rect 18328 2586 18380 2592
rect 18340 1902 18368 2586
rect 18236 1896 18288 1902
rect 18236 1838 18288 1844
rect 18328 1896 18380 1902
rect 18328 1838 18380 1844
rect 18248 1494 18276 1838
rect 18236 1488 18288 1494
rect 18236 1430 18288 1436
rect 18432 1358 18460 2746
rect 18524 2650 18552 2910
rect 18512 2644 18564 2650
rect 18512 2586 18564 2592
rect 18616 2310 18644 3148
rect 18788 3120 18840 3126
rect 18892 3074 18920 11018
rect 18972 9920 19024 9926
rect 18972 9862 19024 9868
rect 18984 8945 19012 9862
rect 18970 8936 19026 8945
rect 18970 8871 19026 8880
rect 18970 8528 19026 8537
rect 18970 8463 19026 8472
rect 18984 4690 19012 8463
rect 18972 4684 19024 4690
rect 18972 4626 19024 4632
rect 18972 3936 19024 3942
rect 18972 3878 19024 3884
rect 18840 3068 18920 3074
rect 18788 3062 18920 3068
rect 18800 3046 18920 3062
rect 18984 3058 19012 3878
rect 19076 3126 19104 19306
rect 19248 18624 19300 18630
rect 19248 18566 19300 18572
rect 19156 17672 19208 17678
rect 19156 17614 19208 17620
rect 19168 17270 19196 17614
rect 19156 17264 19208 17270
rect 19156 17206 19208 17212
rect 19156 14816 19208 14822
rect 19156 14758 19208 14764
rect 19168 13802 19196 14758
rect 19156 13796 19208 13802
rect 19156 13738 19208 13744
rect 19156 12640 19208 12646
rect 19156 12582 19208 12588
rect 19168 12306 19196 12582
rect 19156 12300 19208 12306
rect 19156 12242 19208 12248
rect 19156 12096 19208 12102
rect 19156 12038 19208 12044
rect 19168 11801 19196 12038
rect 19154 11792 19210 11801
rect 19154 11727 19210 11736
rect 19156 9648 19208 9654
rect 19156 9590 19208 9596
rect 19168 9110 19196 9590
rect 19156 9104 19208 9110
rect 19156 9046 19208 9052
rect 19156 8832 19208 8838
rect 19156 8774 19208 8780
rect 19168 8498 19196 8774
rect 19156 8492 19208 8498
rect 19156 8434 19208 8440
rect 19260 6914 19288 18566
rect 19340 17536 19392 17542
rect 19340 17478 19392 17484
rect 19352 16658 19380 17478
rect 19340 16652 19392 16658
rect 19340 16594 19392 16600
rect 19338 12744 19394 12753
rect 19338 12679 19394 12688
rect 19352 12356 19380 12679
rect 19444 12481 19472 41414
rect 19720 41414 19748 44540
rect 19800 43104 19852 43110
rect 19800 43046 19852 43052
rect 19812 42838 19840 43046
rect 19800 42832 19852 42838
rect 19800 42774 19852 42780
rect 19800 42560 19852 42566
rect 19800 42502 19852 42508
rect 19812 41993 19840 42502
rect 19798 41984 19854 41993
rect 19798 41919 19854 41928
rect 19720 41386 19932 41414
rect 19614 41375 19670 41384
rect 19708 40384 19760 40390
rect 19708 40326 19760 40332
rect 19524 39432 19576 39438
rect 19524 39374 19576 39380
rect 19536 38554 19564 39374
rect 19524 38548 19576 38554
rect 19524 38490 19576 38496
rect 19720 34202 19748 40326
rect 19904 40118 19932 41386
rect 19996 40730 20024 44540
rect 20272 43450 20300 44540
rect 20548 43450 20576 44540
rect 20260 43444 20312 43450
rect 20260 43386 20312 43392
rect 20536 43444 20588 43450
rect 20536 43386 20588 43392
rect 20168 43308 20220 43314
rect 20168 43250 20220 43256
rect 20076 43240 20128 43246
rect 20076 43182 20128 43188
rect 20088 41750 20116 43182
rect 20180 42906 20208 43250
rect 20824 43246 20852 44540
rect 20812 43240 20864 43246
rect 20812 43182 20864 43188
rect 20536 43172 20588 43178
rect 20536 43114 20588 43120
rect 20168 42900 20220 42906
rect 20168 42842 20220 42848
rect 20352 42832 20404 42838
rect 20352 42774 20404 42780
rect 20260 42764 20312 42770
rect 20260 42706 20312 42712
rect 20168 42560 20220 42566
rect 20168 42502 20220 42508
rect 20180 42294 20208 42502
rect 20168 42288 20220 42294
rect 20168 42230 20220 42236
rect 20272 42226 20300 42706
rect 20260 42220 20312 42226
rect 20260 42162 20312 42168
rect 20168 42152 20220 42158
rect 20168 42094 20220 42100
rect 20076 41744 20128 41750
rect 20076 41686 20128 41692
rect 19984 40724 20036 40730
rect 19984 40666 20036 40672
rect 19892 40112 19944 40118
rect 19892 40054 19944 40060
rect 20180 39522 20208 42094
rect 20260 42016 20312 42022
rect 20260 41958 20312 41964
rect 20272 40474 20300 41958
rect 20364 41750 20392 42774
rect 20548 42702 20576 43114
rect 20628 42900 20680 42906
rect 20628 42842 20680 42848
rect 20444 42696 20496 42702
rect 20444 42638 20496 42644
rect 20536 42696 20588 42702
rect 20536 42638 20588 42644
rect 20456 41818 20484 42638
rect 20640 42634 20668 42842
rect 20628 42628 20680 42634
rect 20628 42570 20680 42576
rect 20720 42560 20772 42566
rect 20720 42502 20772 42508
rect 20812 42560 20864 42566
rect 20812 42502 20864 42508
rect 20628 42152 20680 42158
rect 20628 42094 20680 42100
rect 20444 41812 20496 41818
rect 20444 41754 20496 41760
rect 20352 41744 20404 41750
rect 20640 41721 20668 42094
rect 20732 41970 20760 42502
rect 20824 42362 20852 42502
rect 21100 42362 21128 44540
rect 21376 43450 21404 44540
rect 21364 43444 21416 43450
rect 21364 43386 21416 43392
rect 21272 43308 21324 43314
rect 21272 43250 21324 43256
rect 21284 43217 21312 43250
rect 21270 43208 21326 43217
rect 21270 43143 21326 43152
rect 21652 43092 21680 44540
rect 21928 43364 21956 44540
rect 22006 43752 22062 43761
rect 22006 43687 22062 43696
rect 22020 43432 22048 43687
rect 22020 43404 22140 43432
rect 21928 43336 22048 43364
rect 21916 43104 21968 43110
rect 21652 43064 21916 43092
rect 21916 43046 21968 43052
rect 21477 43004 21785 43013
rect 21477 43002 21483 43004
rect 21539 43002 21563 43004
rect 21619 43002 21643 43004
rect 21699 43002 21723 43004
rect 21779 43002 21785 43004
rect 21539 42950 21541 43002
rect 21721 42950 21723 43002
rect 21477 42948 21483 42950
rect 21539 42948 21563 42950
rect 21619 42948 21643 42950
rect 21699 42948 21723 42950
rect 21779 42948 21785 42950
rect 21477 42939 21785 42948
rect 22020 42770 22048 43336
rect 22112 42906 22140 43404
rect 22100 42900 22152 42906
rect 22100 42842 22152 42848
rect 21916 42764 21968 42770
rect 21916 42706 21968 42712
rect 22008 42764 22060 42770
rect 22008 42706 22060 42712
rect 21272 42560 21324 42566
rect 21272 42502 21324 42508
rect 20812 42356 20864 42362
rect 20812 42298 20864 42304
rect 21088 42356 21140 42362
rect 21088 42298 21140 42304
rect 21086 42256 21142 42265
rect 20996 42220 21048 42226
rect 21086 42191 21088 42200
rect 20996 42162 21048 42168
rect 21140 42191 21142 42200
rect 21088 42162 21140 42168
rect 20904 42016 20956 42022
rect 20732 41942 20852 41970
rect 20904 41958 20956 41964
rect 20352 41686 20404 41692
rect 20626 41712 20682 41721
rect 20626 41647 20682 41656
rect 20536 41608 20588 41614
rect 20534 41576 20536 41585
rect 20588 41576 20590 41585
rect 20534 41511 20590 41520
rect 20628 41472 20680 41478
rect 20628 41414 20680 41420
rect 20640 41386 20760 41414
rect 20350 40488 20406 40497
rect 20272 40446 20350 40474
rect 20350 40423 20406 40432
rect 20258 39536 20314 39545
rect 20180 39494 20258 39522
rect 20258 39471 20314 39480
rect 20352 39500 20404 39506
rect 20352 39442 20404 39448
rect 20364 39098 20392 39442
rect 20352 39092 20404 39098
rect 20352 39034 20404 39040
rect 20536 38956 20588 38962
rect 20536 38898 20588 38904
rect 20548 38554 20576 38898
rect 20536 38548 20588 38554
rect 20536 38490 20588 38496
rect 20350 36816 20406 36825
rect 20350 36751 20352 36760
rect 20404 36751 20406 36760
rect 20352 36722 20404 36728
rect 19984 36236 20036 36242
rect 19984 36178 20036 36184
rect 19708 34196 19760 34202
rect 19708 34138 19760 34144
rect 19522 34096 19578 34105
rect 19578 34054 19656 34082
rect 19522 34031 19578 34040
rect 19628 33998 19656 34054
rect 19616 33992 19668 33998
rect 19616 33934 19668 33940
rect 19720 33114 19748 34138
rect 19708 33108 19760 33114
rect 19708 33050 19760 33056
rect 19800 32020 19852 32026
rect 19800 31962 19852 31968
rect 19812 30734 19840 31962
rect 19800 30728 19852 30734
rect 19800 30670 19852 30676
rect 19996 28558 20024 36178
rect 20260 35080 20312 35086
rect 20260 35022 20312 35028
rect 20076 34944 20128 34950
rect 20076 34886 20128 34892
rect 20088 34746 20116 34886
rect 20272 34746 20300 35022
rect 20352 34944 20404 34950
rect 20352 34886 20404 34892
rect 20364 34746 20392 34886
rect 20076 34740 20128 34746
rect 20076 34682 20128 34688
rect 20260 34740 20312 34746
rect 20260 34682 20312 34688
rect 20352 34740 20404 34746
rect 20352 34682 20404 34688
rect 20628 34604 20680 34610
rect 20628 34546 20680 34552
rect 20536 34468 20588 34474
rect 20536 34410 20588 34416
rect 20076 33992 20128 33998
rect 20076 33934 20128 33940
rect 20088 29578 20116 33934
rect 20260 32224 20312 32230
rect 20260 32166 20312 32172
rect 20272 32026 20300 32166
rect 20260 32020 20312 32026
rect 20260 31962 20312 31968
rect 20352 31952 20404 31958
rect 20352 31894 20404 31900
rect 20168 31816 20220 31822
rect 20168 31758 20220 31764
rect 20180 31482 20208 31758
rect 20364 31754 20392 31894
rect 20272 31726 20392 31754
rect 20168 31476 20220 31482
rect 20168 31418 20220 31424
rect 20076 29572 20128 29578
rect 20076 29514 20128 29520
rect 19984 28552 20036 28558
rect 19984 28494 20036 28500
rect 20076 28484 20128 28490
rect 20076 28426 20128 28432
rect 19708 27940 19760 27946
rect 19708 27882 19760 27888
rect 19524 24812 19576 24818
rect 19524 24754 19576 24760
rect 19536 24206 19564 24754
rect 19524 24200 19576 24206
rect 19524 24142 19576 24148
rect 19616 21888 19668 21894
rect 19616 21830 19668 21836
rect 19628 21554 19656 21830
rect 19616 21548 19668 21554
rect 19616 21490 19668 21496
rect 19524 21344 19576 21350
rect 19524 21286 19576 21292
rect 19536 19378 19564 21286
rect 19616 20800 19668 20806
rect 19616 20742 19668 20748
rect 19524 19372 19576 19378
rect 19524 19314 19576 19320
rect 19524 19168 19576 19174
rect 19524 19110 19576 19116
rect 19536 18766 19564 19110
rect 19524 18760 19576 18766
rect 19524 18702 19576 18708
rect 19628 17202 19656 20742
rect 19616 17196 19668 17202
rect 19616 17138 19668 17144
rect 19524 16584 19576 16590
rect 19524 16526 19576 16532
rect 19536 16250 19564 16526
rect 19524 16244 19576 16250
rect 19524 16186 19576 16192
rect 19720 15008 19748 27882
rect 19800 26784 19852 26790
rect 19800 26726 19852 26732
rect 19812 26382 19840 26726
rect 19892 26580 19944 26586
rect 19892 26522 19944 26528
rect 19800 26376 19852 26382
rect 19800 26318 19852 26324
rect 19904 20874 19932 26522
rect 20088 25770 20116 28426
rect 20168 26784 20220 26790
rect 20168 26726 20220 26732
rect 20180 26450 20208 26726
rect 20168 26444 20220 26450
rect 20168 26386 20220 26392
rect 20076 25764 20128 25770
rect 20076 25706 20128 25712
rect 20272 25158 20300 31726
rect 20444 31136 20496 31142
rect 20444 31078 20496 31084
rect 20456 30870 20484 31078
rect 20444 30864 20496 30870
rect 20444 30806 20496 30812
rect 20352 29640 20404 29646
rect 20352 29582 20404 29588
rect 20364 29306 20392 29582
rect 20352 29300 20404 29306
rect 20352 29242 20404 29248
rect 20442 29200 20498 29209
rect 20364 29170 20442 29186
rect 20352 29164 20442 29170
rect 20404 29158 20442 29164
rect 20442 29135 20498 29144
rect 20352 29106 20404 29112
rect 20548 27146 20576 34410
rect 20640 34202 20668 34546
rect 20628 34196 20680 34202
rect 20628 34138 20680 34144
rect 20732 32978 20760 41386
rect 20824 40594 20852 41942
rect 20916 41682 20944 41958
rect 20904 41676 20956 41682
rect 20904 41618 20956 41624
rect 21008 41414 21036 42162
rect 21284 41818 21312 42502
rect 21364 42220 21416 42226
rect 21364 42162 21416 42168
rect 21272 41812 21324 41818
rect 21272 41754 21324 41760
rect 21270 41712 21326 41721
rect 21270 41647 21326 41656
rect 21284 41614 21312 41647
rect 21272 41608 21324 41614
rect 21272 41550 21324 41556
rect 21376 41414 21404 42162
rect 21456 42016 21508 42022
rect 21508 41976 21864 42004
rect 21456 41958 21508 41964
rect 21477 41916 21785 41925
rect 21477 41914 21483 41916
rect 21539 41914 21563 41916
rect 21619 41914 21643 41916
rect 21699 41914 21723 41916
rect 21779 41914 21785 41916
rect 21539 41862 21541 41914
rect 21721 41862 21723 41914
rect 21477 41860 21483 41862
rect 21539 41860 21563 41862
rect 21619 41860 21643 41862
rect 21699 41860 21723 41862
rect 21779 41860 21785 41862
rect 21477 41851 21785 41860
rect 21836 41614 21864 41976
rect 21640 41608 21692 41614
rect 21640 41550 21692 41556
rect 21824 41608 21876 41614
rect 21824 41550 21876 41556
rect 21548 41472 21600 41478
rect 20916 41386 21036 41414
rect 21284 41386 21404 41414
rect 21454 41440 21510 41449
rect 20812 40588 20864 40594
rect 20812 40530 20864 40536
rect 20812 40452 20864 40458
rect 20812 40394 20864 40400
rect 20720 32972 20772 32978
rect 20720 32914 20772 32920
rect 20720 32496 20772 32502
rect 20720 32438 20772 32444
rect 20732 31686 20760 32438
rect 20720 31680 20772 31686
rect 20720 31622 20772 31628
rect 20720 29776 20772 29782
rect 20720 29718 20772 29724
rect 20732 29238 20760 29718
rect 20824 29322 20852 40394
rect 20916 30054 20944 41386
rect 21088 41268 21140 41274
rect 21284 41256 21312 41386
rect 21510 41420 21548 41426
rect 21510 41414 21600 41420
rect 21652 41414 21680 41550
rect 21510 41398 21588 41414
rect 21652 41386 21864 41414
rect 21454 41375 21510 41384
rect 21140 41228 21312 41256
rect 21088 41210 21140 41216
rect 20996 41200 21048 41206
rect 20996 41142 21048 41148
rect 21008 38894 21036 41142
rect 21272 41132 21324 41138
rect 21456 41132 21508 41138
rect 21272 41074 21324 41080
rect 21376 41092 21456 41120
rect 21088 40656 21140 40662
rect 21088 40598 21140 40604
rect 21100 39030 21128 40598
rect 21284 39846 21312 41074
rect 21272 39840 21324 39846
rect 21272 39782 21324 39788
rect 21376 39642 21404 41092
rect 21456 41074 21508 41080
rect 21477 40828 21785 40837
rect 21477 40826 21483 40828
rect 21539 40826 21563 40828
rect 21619 40826 21643 40828
rect 21699 40826 21723 40828
rect 21779 40826 21785 40828
rect 21539 40774 21541 40826
rect 21721 40774 21723 40826
rect 21477 40772 21483 40774
rect 21539 40772 21563 40774
rect 21619 40772 21643 40774
rect 21699 40772 21723 40774
rect 21779 40772 21785 40774
rect 21477 40763 21785 40772
rect 21836 40730 21864 41386
rect 21928 41070 21956 42706
rect 22204 42566 22232 44540
rect 22480 43602 22508 44540
rect 22480 43574 22692 43602
rect 22376 43308 22428 43314
rect 22376 43250 22428 43256
rect 22284 42628 22336 42634
rect 22284 42570 22336 42576
rect 22192 42560 22244 42566
rect 22192 42502 22244 42508
rect 22100 41540 22152 41546
rect 22100 41482 22152 41488
rect 22192 41540 22244 41546
rect 22192 41482 22244 41488
rect 22008 41132 22060 41138
rect 22008 41074 22060 41080
rect 21916 41064 21968 41070
rect 21916 41006 21968 41012
rect 21914 40896 21970 40905
rect 21914 40831 21970 40840
rect 21928 40730 21956 40831
rect 21824 40724 21876 40730
rect 21824 40666 21876 40672
rect 21916 40724 21968 40730
rect 21916 40666 21968 40672
rect 21916 40588 21968 40594
rect 21916 40530 21968 40536
rect 21822 39944 21878 39953
rect 21822 39879 21878 39888
rect 21477 39740 21785 39749
rect 21477 39738 21483 39740
rect 21539 39738 21563 39740
rect 21619 39738 21643 39740
rect 21699 39738 21723 39740
rect 21779 39738 21785 39740
rect 21539 39686 21541 39738
rect 21721 39686 21723 39738
rect 21477 39684 21483 39686
rect 21539 39684 21563 39686
rect 21619 39684 21643 39686
rect 21699 39684 21723 39686
rect 21779 39684 21785 39686
rect 21477 39675 21785 39684
rect 21364 39636 21416 39642
rect 21364 39578 21416 39584
rect 21088 39024 21140 39030
rect 21088 38966 21140 38972
rect 20996 38888 21048 38894
rect 20996 38830 21048 38836
rect 21477 38652 21785 38661
rect 21477 38650 21483 38652
rect 21539 38650 21563 38652
rect 21619 38650 21643 38652
rect 21699 38650 21723 38652
rect 21779 38650 21785 38652
rect 21539 38598 21541 38650
rect 21721 38598 21723 38650
rect 21477 38596 21483 38598
rect 21539 38596 21563 38598
rect 21619 38596 21643 38598
rect 21699 38596 21723 38598
rect 21779 38596 21785 38598
rect 21477 38587 21785 38596
rect 21477 37564 21785 37573
rect 21477 37562 21483 37564
rect 21539 37562 21563 37564
rect 21619 37562 21643 37564
rect 21699 37562 21723 37564
rect 21779 37562 21785 37564
rect 21539 37510 21541 37562
rect 21721 37510 21723 37562
rect 21477 37508 21483 37510
rect 21539 37508 21563 37510
rect 21619 37508 21643 37510
rect 21699 37508 21723 37510
rect 21779 37508 21785 37510
rect 21477 37499 21785 37508
rect 20996 37256 21048 37262
rect 20996 37198 21048 37204
rect 21008 36922 21036 37198
rect 20996 36916 21048 36922
rect 20996 36858 21048 36864
rect 21477 36476 21785 36485
rect 21477 36474 21483 36476
rect 21539 36474 21563 36476
rect 21619 36474 21643 36476
rect 21699 36474 21723 36476
rect 21779 36474 21785 36476
rect 21539 36422 21541 36474
rect 21721 36422 21723 36474
rect 21477 36420 21483 36422
rect 21539 36420 21563 36422
rect 21619 36420 21643 36422
rect 21699 36420 21723 36422
rect 21779 36420 21785 36422
rect 21477 36411 21785 36420
rect 21477 35388 21785 35397
rect 21477 35386 21483 35388
rect 21539 35386 21563 35388
rect 21619 35386 21643 35388
rect 21699 35386 21723 35388
rect 21779 35386 21785 35388
rect 21539 35334 21541 35386
rect 21721 35334 21723 35386
rect 21477 35332 21483 35334
rect 21539 35332 21563 35334
rect 21619 35332 21643 35334
rect 21699 35332 21723 35334
rect 21779 35332 21785 35334
rect 21477 35323 21785 35332
rect 21732 34944 21784 34950
rect 21732 34886 21784 34892
rect 21744 34474 21772 34886
rect 21836 34746 21864 39879
rect 21928 39574 21956 40530
rect 22020 40186 22048 41074
rect 22112 40526 22140 41482
rect 22204 41274 22232 41482
rect 22192 41268 22244 41274
rect 22192 41210 22244 41216
rect 22192 41132 22244 41138
rect 22192 41074 22244 41080
rect 22100 40520 22152 40526
rect 22100 40462 22152 40468
rect 22008 40180 22060 40186
rect 22008 40122 22060 40128
rect 21916 39568 21968 39574
rect 21916 39510 21968 39516
rect 22008 38956 22060 38962
rect 22008 38898 22060 38904
rect 22020 38418 22048 38898
rect 22008 38412 22060 38418
rect 22008 38354 22060 38360
rect 21916 37256 21968 37262
rect 21916 37198 21968 37204
rect 21928 36922 21956 37198
rect 21916 36916 21968 36922
rect 21916 36858 21968 36864
rect 22204 36394 22232 41074
rect 22296 39953 22324 42570
rect 22388 41750 22416 43250
rect 22664 42906 22692 43574
rect 22652 42900 22704 42906
rect 22652 42842 22704 42848
rect 22652 42628 22704 42634
rect 22652 42570 22704 42576
rect 22560 42220 22612 42226
rect 22560 42162 22612 42168
rect 22572 41818 22600 42162
rect 22560 41812 22612 41818
rect 22560 41754 22612 41760
rect 22376 41744 22428 41750
rect 22376 41686 22428 41692
rect 22376 41472 22428 41478
rect 22376 41414 22428 41420
rect 22388 40662 22416 41414
rect 22664 41274 22692 42570
rect 22756 42362 22784 44540
rect 22836 43308 22888 43314
rect 22836 43250 22888 43256
rect 22848 42838 22876 43250
rect 22926 43072 22982 43081
rect 22926 43007 22982 43016
rect 22836 42832 22888 42838
rect 22836 42774 22888 42780
rect 22940 42362 22968 43007
rect 23032 42770 23060 44540
rect 23020 42764 23072 42770
rect 23020 42706 23072 42712
rect 22744 42356 22796 42362
rect 22744 42298 22796 42304
rect 22928 42356 22980 42362
rect 22928 42298 22980 42304
rect 23112 42220 23164 42226
rect 23112 42162 23164 42168
rect 22928 42152 22980 42158
rect 22928 42094 22980 42100
rect 22652 41268 22704 41274
rect 22652 41210 22704 41216
rect 22468 41132 22520 41138
rect 22468 41074 22520 41080
rect 22480 40730 22508 41074
rect 22468 40724 22520 40730
rect 22468 40666 22520 40672
rect 22376 40656 22428 40662
rect 22376 40598 22428 40604
rect 22468 40520 22520 40526
rect 22468 40462 22520 40468
rect 22374 40080 22430 40089
rect 22374 40015 22376 40024
rect 22428 40015 22430 40024
rect 22376 39986 22428 39992
rect 22282 39944 22338 39953
rect 22282 39879 22338 39888
rect 22112 36366 22232 36394
rect 21824 34740 21876 34746
rect 21824 34682 21876 34688
rect 22008 34604 22060 34610
rect 22008 34546 22060 34552
rect 21732 34468 21784 34474
rect 21732 34410 21784 34416
rect 21364 34400 21416 34406
rect 21364 34342 21416 34348
rect 21272 33312 21324 33318
rect 21272 33254 21324 33260
rect 20996 32972 21048 32978
rect 20996 32914 21048 32920
rect 21008 30802 21036 32914
rect 20996 30796 21048 30802
rect 20996 30738 21048 30744
rect 20904 30048 20956 30054
rect 20904 29990 20956 29996
rect 20824 29294 20944 29322
rect 20720 29232 20772 29238
rect 20626 29200 20682 29209
rect 20720 29174 20772 29180
rect 20626 29135 20682 29144
rect 20640 28762 20668 29135
rect 20916 29016 20944 29294
rect 20824 28988 20944 29016
rect 20628 28756 20680 28762
rect 20628 28698 20680 28704
rect 20720 28688 20772 28694
rect 20720 28630 20772 28636
rect 20732 28150 20760 28630
rect 20720 28144 20772 28150
rect 20720 28086 20772 28092
rect 20364 27118 20576 27146
rect 20260 25152 20312 25158
rect 20260 25094 20312 25100
rect 20168 24608 20220 24614
rect 20168 24550 20220 24556
rect 20180 24410 20208 24550
rect 20168 24404 20220 24410
rect 20168 24346 20220 24352
rect 20260 23656 20312 23662
rect 20260 23598 20312 23604
rect 20272 22642 20300 23598
rect 20260 22636 20312 22642
rect 20260 22578 20312 22584
rect 20364 22094 20392 27118
rect 20444 27056 20496 27062
rect 20444 26998 20496 27004
rect 20456 26314 20484 26998
rect 20536 26988 20588 26994
rect 20536 26930 20588 26936
rect 20444 26308 20496 26314
rect 20444 26250 20496 26256
rect 20548 26042 20576 26930
rect 20824 26908 20852 28988
rect 21008 28626 21036 30738
rect 21088 30592 21140 30598
rect 21088 30534 21140 30540
rect 21100 30258 21128 30534
rect 21088 30252 21140 30258
rect 21088 30194 21140 30200
rect 21088 29504 21140 29510
rect 21088 29446 21140 29452
rect 21100 29306 21128 29446
rect 21088 29300 21140 29306
rect 21088 29242 21140 29248
rect 21086 29200 21142 29209
rect 21086 29135 21088 29144
rect 21140 29135 21142 29144
rect 21088 29106 21140 29112
rect 20996 28620 21048 28626
rect 20996 28562 21048 28568
rect 21008 28082 21036 28562
rect 21088 28144 21140 28150
rect 21088 28086 21140 28092
rect 20996 28076 21048 28082
rect 20996 28018 21048 28024
rect 21100 27470 21128 28086
rect 21088 27464 21140 27470
rect 21088 27406 21140 27412
rect 20996 27328 21048 27334
rect 20996 27270 21048 27276
rect 21008 27062 21036 27270
rect 20996 27056 21048 27062
rect 20996 26998 21048 27004
rect 20824 26880 21036 26908
rect 20720 26784 20772 26790
rect 20720 26726 20772 26732
rect 20536 26036 20588 26042
rect 20536 25978 20588 25984
rect 20732 25294 20760 26726
rect 20720 25288 20772 25294
rect 20720 25230 20772 25236
rect 20720 25152 20772 25158
rect 20720 25094 20772 25100
rect 20444 24064 20496 24070
rect 20444 24006 20496 24012
rect 20456 23866 20484 24006
rect 20444 23860 20496 23866
rect 20444 23802 20496 23808
rect 20536 23520 20588 23526
rect 20536 23462 20588 23468
rect 20444 23112 20496 23118
rect 20444 23054 20496 23060
rect 20456 22778 20484 23054
rect 20444 22772 20496 22778
rect 20444 22714 20496 22720
rect 20364 22066 20484 22094
rect 19892 20868 19944 20874
rect 19892 20810 19944 20816
rect 20352 20868 20404 20874
rect 20352 20810 20404 20816
rect 20364 20602 20392 20810
rect 20352 20596 20404 20602
rect 20352 20538 20404 20544
rect 20352 20460 20404 20466
rect 20352 20402 20404 20408
rect 20260 20324 20312 20330
rect 20260 20266 20312 20272
rect 19800 20256 19852 20262
rect 19800 20198 19852 20204
rect 20168 20256 20220 20262
rect 20168 20198 20220 20204
rect 19812 18970 19840 20198
rect 19984 20052 20036 20058
rect 19984 19994 20036 20000
rect 19892 19372 19944 19378
rect 19892 19314 19944 19320
rect 19800 18964 19852 18970
rect 19800 18906 19852 18912
rect 19536 14980 19748 15008
rect 19430 12472 19486 12481
rect 19430 12407 19486 12416
rect 19352 12328 19463 12356
rect 19435 12322 19463 12328
rect 19435 12294 19472 12322
rect 19444 12238 19472 12294
rect 19432 12232 19484 12238
rect 19536 12220 19564 14980
rect 19706 14920 19762 14929
rect 19706 14855 19762 14864
rect 19616 12844 19668 12850
rect 19616 12786 19668 12792
rect 19628 12442 19656 12786
rect 19720 12442 19748 14855
rect 19800 14272 19852 14278
rect 19800 14214 19852 14220
rect 19904 14226 19932 19314
rect 19996 15502 20024 19994
rect 20076 19168 20128 19174
rect 20076 19110 20128 19116
rect 20088 17542 20116 19110
rect 20180 18902 20208 20198
rect 20272 20058 20300 20266
rect 20364 20058 20392 20402
rect 20260 20052 20312 20058
rect 20260 19994 20312 20000
rect 20352 20052 20404 20058
rect 20352 19994 20404 20000
rect 20352 19372 20404 19378
rect 20456 19360 20484 22066
rect 20548 19496 20576 23462
rect 20732 21978 20760 25094
rect 20904 22432 20956 22438
rect 20904 22374 20956 22380
rect 20640 21950 20760 21978
rect 20812 22024 20864 22030
rect 20916 21978 20944 22374
rect 21008 22094 21036 26880
rect 21180 24812 21232 24818
rect 21180 24754 21232 24760
rect 21086 24712 21142 24721
rect 21086 24647 21142 24656
rect 21100 23798 21128 24647
rect 21192 24410 21220 24754
rect 21180 24404 21232 24410
rect 21180 24346 21232 24352
rect 21088 23792 21140 23798
rect 21088 23734 21140 23740
rect 21284 23118 21312 33254
rect 21376 32910 21404 34342
rect 21477 34300 21785 34309
rect 21477 34298 21483 34300
rect 21539 34298 21563 34300
rect 21619 34298 21643 34300
rect 21699 34298 21723 34300
rect 21779 34298 21785 34300
rect 21539 34246 21541 34298
rect 21721 34246 21723 34298
rect 21477 34244 21483 34246
rect 21539 34244 21563 34246
rect 21619 34244 21643 34246
rect 21699 34244 21723 34246
rect 21779 34244 21785 34246
rect 21477 34235 21785 34244
rect 22020 34202 22048 34546
rect 22008 34196 22060 34202
rect 22008 34138 22060 34144
rect 21477 33212 21785 33221
rect 21477 33210 21483 33212
rect 21539 33210 21563 33212
rect 21619 33210 21643 33212
rect 21699 33210 21723 33212
rect 21779 33210 21785 33212
rect 21539 33158 21541 33210
rect 21721 33158 21723 33210
rect 21477 33156 21483 33158
rect 21539 33156 21563 33158
rect 21619 33156 21643 33158
rect 21699 33156 21723 33158
rect 21779 33156 21785 33158
rect 21477 33147 21785 33156
rect 21364 32904 21416 32910
rect 21364 32846 21416 32852
rect 21477 32124 21785 32133
rect 21477 32122 21483 32124
rect 21539 32122 21563 32124
rect 21619 32122 21643 32124
rect 21699 32122 21723 32124
rect 21779 32122 21785 32124
rect 21539 32070 21541 32122
rect 21721 32070 21723 32122
rect 21477 32068 21483 32070
rect 21539 32068 21563 32070
rect 21619 32068 21643 32070
rect 21699 32068 21723 32070
rect 21779 32068 21785 32070
rect 21477 32059 21785 32068
rect 21824 31680 21876 31686
rect 21824 31622 21876 31628
rect 21477 31036 21785 31045
rect 21477 31034 21483 31036
rect 21539 31034 21563 31036
rect 21619 31034 21643 31036
rect 21699 31034 21723 31036
rect 21779 31034 21785 31036
rect 21539 30982 21541 31034
rect 21721 30982 21723 31034
rect 21477 30980 21483 30982
rect 21539 30980 21563 30982
rect 21619 30980 21643 30982
rect 21699 30980 21723 30982
rect 21779 30980 21785 30982
rect 21477 30971 21785 30980
rect 21836 30666 21864 31622
rect 21824 30660 21876 30666
rect 21824 30602 21876 30608
rect 21477 29948 21785 29957
rect 21477 29946 21483 29948
rect 21539 29946 21563 29948
rect 21619 29946 21643 29948
rect 21699 29946 21723 29948
rect 21779 29946 21785 29948
rect 21539 29894 21541 29946
rect 21721 29894 21723 29946
rect 21477 29892 21483 29894
rect 21539 29892 21563 29894
rect 21619 29892 21643 29894
rect 21699 29892 21723 29894
rect 21779 29892 21785 29894
rect 21477 29883 21785 29892
rect 21456 29844 21508 29850
rect 21456 29786 21508 29792
rect 21364 29572 21416 29578
rect 21364 29514 21416 29520
rect 21376 29170 21404 29514
rect 21468 29238 21496 29786
rect 21456 29232 21508 29238
rect 21456 29174 21508 29180
rect 21364 29164 21416 29170
rect 21364 29106 21416 29112
rect 21916 29028 21968 29034
rect 21916 28970 21968 28976
rect 22112 28994 22140 36366
rect 22192 33312 22244 33318
rect 22192 33254 22244 33260
rect 22204 33114 22232 33254
rect 22192 33108 22244 33114
rect 22192 33050 22244 33056
rect 22480 31754 22508 40462
rect 22652 40384 22704 40390
rect 22652 40326 22704 40332
rect 22664 40186 22692 40326
rect 22940 40186 22968 42094
rect 23124 41274 23152 42162
rect 23308 41818 23336 44540
rect 23584 43432 23612 44540
rect 23756 43444 23808 43450
rect 23584 43404 23756 43432
rect 23756 43386 23808 43392
rect 23664 43308 23716 43314
rect 23664 43250 23716 43256
rect 23480 42696 23532 42702
rect 23480 42638 23532 42644
rect 23296 41812 23348 41818
rect 23296 41754 23348 41760
rect 23386 41576 23442 41585
rect 23296 41540 23348 41546
rect 23386 41511 23442 41520
rect 23296 41482 23348 41488
rect 23112 41268 23164 41274
rect 23112 41210 23164 41216
rect 23112 41132 23164 41138
rect 23112 41074 23164 41080
rect 23020 40656 23072 40662
rect 23020 40598 23072 40604
rect 22652 40180 22704 40186
rect 22652 40122 22704 40128
rect 22928 40180 22980 40186
rect 22928 40122 22980 40128
rect 23032 40050 23060 40598
rect 23020 40044 23072 40050
rect 23020 39986 23072 39992
rect 22560 39432 22612 39438
rect 22560 39374 22612 39380
rect 22572 39098 22600 39374
rect 22560 39092 22612 39098
rect 22560 39034 22612 39040
rect 23124 38826 23152 41074
rect 23308 40730 23336 41482
rect 23400 41274 23428 41511
rect 23492 41274 23520 42638
rect 23572 42220 23624 42226
rect 23572 42162 23624 42168
rect 23388 41268 23440 41274
rect 23388 41210 23440 41216
rect 23480 41268 23532 41274
rect 23480 41210 23532 41216
rect 23584 41120 23612 42162
rect 23492 41092 23612 41120
rect 23296 40724 23348 40730
rect 23296 40666 23348 40672
rect 23296 40520 23348 40526
rect 23296 40462 23348 40468
rect 23204 40452 23256 40458
rect 23204 40394 23256 40400
rect 23216 39642 23244 40394
rect 23308 39642 23336 40462
rect 23386 39808 23442 39817
rect 23386 39743 23442 39752
rect 23204 39636 23256 39642
rect 23204 39578 23256 39584
rect 23296 39636 23348 39642
rect 23296 39578 23348 39584
rect 23204 39432 23256 39438
rect 23204 39374 23256 39380
rect 23216 39114 23244 39374
rect 23216 39086 23336 39114
rect 23204 39024 23256 39030
rect 23204 38966 23256 38972
rect 23112 38820 23164 38826
rect 23112 38762 23164 38768
rect 23216 38554 23244 38966
rect 23204 38548 23256 38554
rect 23204 38490 23256 38496
rect 22836 38344 22888 38350
rect 22836 38286 22888 38292
rect 22848 38010 22876 38286
rect 22836 38004 22888 38010
rect 22836 37946 22888 37952
rect 23020 37732 23072 37738
rect 23020 37674 23072 37680
rect 23032 37126 23060 37674
rect 23020 37120 23072 37126
rect 23020 37062 23072 37068
rect 23308 36258 23336 39086
rect 23400 38010 23428 39743
rect 23492 39302 23520 41092
rect 23676 41018 23704 43250
rect 23860 43092 23888 44540
rect 23860 43064 23980 43092
rect 23756 42696 23808 42702
rect 23756 42638 23808 42644
rect 23584 40990 23704 41018
rect 23584 40186 23612 40990
rect 23768 40934 23796 42638
rect 23952 41818 23980 43064
rect 24136 42650 24164 44540
rect 24412 43738 24440 44540
rect 24320 43710 24440 43738
rect 24688 43738 24716 44540
rect 24688 43710 24808 43738
rect 24216 43240 24268 43246
rect 24216 43182 24268 43188
rect 24044 42622 24164 42650
rect 24044 42294 24072 42622
rect 24124 42560 24176 42566
rect 24124 42502 24176 42508
rect 24032 42288 24084 42294
rect 24032 42230 24084 42236
rect 24136 41993 24164 42502
rect 24122 41984 24178 41993
rect 24122 41919 24178 41928
rect 23940 41812 23992 41818
rect 23940 41754 23992 41760
rect 23848 41540 23900 41546
rect 23848 41482 23900 41488
rect 23860 41437 23888 41482
rect 24032 41472 24084 41478
rect 23846 41428 23902 41437
rect 24032 41414 24084 41420
rect 23846 41363 23902 41372
rect 23860 41274 23980 41290
rect 23848 41268 23980 41274
rect 23900 41262 23980 41268
rect 23848 41210 23900 41216
rect 23848 41132 23900 41138
rect 23848 41074 23900 41080
rect 23664 40928 23716 40934
rect 23662 40896 23664 40905
rect 23756 40928 23808 40934
rect 23716 40896 23718 40905
rect 23756 40870 23808 40876
rect 23662 40831 23718 40840
rect 23664 40588 23716 40594
rect 23664 40530 23716 40536
rect 23676 40186 23704 40530
rect 23756 40452 23808 40458
rect 23756 40394 23808 40400
rect 23572 40180 23624 40186
rect 23572 40122 23624 40128
rect 23664 40180 23716 40186
rect 23664 40122 23716 40128
rect 23572 39840 23624 39846
rect 23572 39782 23624 39788
rect 23584 39438 23612 39782
rect 23572 39432 23624 39438
rect 23572 39374 23624 39380
rect 23480 39296 23532 39302
rect 23480 39238 23532 39244
rect 23388 38004 23440 38010
rect 23388 37946 23440 37952
rect 23572 37868 23624 37874
rect 23572 37810 23624 37816
rect 23388 37800 23440 37806
rect 23388 37742 23440 37748
rect 23400 37466 23428 37742
rect 23584 37466 23612 37810
rect 23388 37460 23440 37466
rect 23388 37402 23440 37408
rect 23572 37460 23624 37466
rect 23572 37402 23624 37408
rect 23572 37256 23624 37262
rect 23572 37198 23624 37204
rect 23584 36922 23612 37198
rect 23572 36916 23624 36922
rect 23572 36858 23624 36864
rect 23664 36780 23716 36786
rect 23664 36722 23716 36728
rect 23308 36230 23428 36258
rect 23296 36168 23348 36174
rect 23296 36110 23348 36116
rect 23308 35834 23336 36110
rect 22560 35828 22612 35834
rect 22560 35770 22612 35776
rect 23296 35828 23348 35834
rect 23296 35770 23348 35776
rect 22572 35698 22600 35770
rect 22560 35692 22612 35698
rect 22560 35634 22612 35640
rect 22836 35692 22888 35698
rect 22836 35634 22888 35640
rect 23204 35692 23256 35698
rect 23204 35634 23256 35640
rect 22848 34406 22876 35634
rect 23216 35290 23244 35634
rect 23400 35578 23428 36230
rect 23572 36168 23624 36174
rect 23572 36110 23624 36116
rect 23400 35550 23520 35578
rect 23296 35488 23348 35494
rect 23296 35430 23348 35436
rect 23388 35488 23440 35494
rect 23388 35430 23440 35436
rect 23204 35284 23256 35290
rect 23204 35226 23256 35232
rect 22928 34944 22980 34950
rect 22928 34886 22980 34892
rect 22836 34400 22888 34406
rect 22836 34342 22888 34348
rect 22744 33856 22796 33862
rect 22744 33798 22796 33804
rect 22756 33522 22784 33798
rect 22744 33516 22796 33522
rect 22744 33458 22796 33464
rect 22652 32428 22704 32434
rect 22652 32370 22704 32376
rect 22480 31726 22600 31754
rect 22192 30592 22244 30598
rect 22192 30534 22244 30540
rect 22204 30258 22232 30534
rect 22284 30320 22336 30326
rect 22284 30262 22336 30268
rect 22376 30320 22428 30326
rect 22376 30262 22428 30268
rect 22192 30252 22244 30258
rect 22192 30194 22244 30200
rect 22296 29306 22324 30262
rect 22388 29714 22416 30262
rect 22376 29708 22428 29714
rect 22376 29650 22428 29656
rect 22284 29300 22336 29306
rect 22284 29242 22336 29248
rect 21477 28860 21785 28869
rect 21477 28858 21483 28860
rect 21539 28858 21563 28860
rect 21619 28858 21643 28860
rect 21699 28858 21723 28860
rect 21779 28858 21785 28860
rect 21539 28806 21541 28858
rect 21721 28806 21723 28858
rect 21477 28804 21483 28806
rect 21539 28804 21563 28806
rect 21619 28804 21643 28806
rect 21699 28804 21723 28806
rect 21779 28804 21785 28806
rect 21477 28795 21785 28804
rect 21477 27772 21785 27781
rect 21477 27770 21483 27772
rect 21539 27770 21563 27772
rect 21619 27770 21643 27772
rect 21699 27770 21723 27772
rect 21779 27770 21785 27772
rect 21539 27718 21541 27770
rect 21721 27718 21723 27770
rect 21477 27716 21483 27718
rect 21539 27716 21563 27718
rect 21619 27716 21643 27718
rect 21699 27716 21723 27718
rect 21779 27716 21785 27718
rect 21477 27707 21785 27716
rect 21477 26684 21785 26693
rect 21477 26682 21483 26684
rect 21539 26682 21563 26684
rect 21619 26682 21643 26684
rect 21699 26682 21723 26684
rect 21779 26682 21785 26684
rect 21539 26630 21541 26682
rect 21721 26630 21723 26682
rect 21477 26628 21483 26630
rect 21539 26628 21563 26630
rect 21619 26628 21643 26630
rect 21699 26628 21723 26630
rect 21779 26628 21785 26630
rect 21477 26619 21785 26628
rect 21824 26036 21876 26042
rect 21824 25978 21876 25984
rect 21836 25702 21864 25978
rect 21928 25786 21956 28970
rect 22112 28966 22324 28994
rect 22100 28552 22152 28558
rect 22100 28494 22152 28500
rect 22112 28218 22140 28494
rect 22192 28416 22244 28422
rect 22192 28358 22244 28364
rect 22204 28218 22232 28358
rect 22100 28212 22152 28218
rect 22100 28154 22152 28160
rect 22192 28212 22244 28218
rect 22192 28154 22244 28160
rect 22296 28098 22324 28966
rect 22204 28070 22324 28098
rect 22008 27872 22060 27878
rect 22008 27814 22060 27820
rect 22020 26382 22048 27814
rect 22008 26376 22060 26382
rect 22008 26318 22060 26324
rect 21928 25758 22048 25786
rect 21824 25696 21876 25702
rect 21824 25638 21876 25644
rect 21916 25696 21968 25702
rect 21916 25638 21968 25644
rect 21477 25596 21785 25605
rect 21477 25594 21483 25596
rect 21539 25594 21563 25596
rect 21619 25594 21643 25596
rect 21699 25594 21723 25596
rect 21779 25594 21785 25596
rect 21539 25542 21541 25594
rect 21721 25542 21723 25594
rect 21477 25540 21483 25542
rect 21539 25540 21563 25542
rect 21619 25540 21643 25542
rect 21699 25540 21723 25542
rect 21779 25540 21785 25542
rect 21477 25531 21785 25540
rect 21836 25294 21864 25638
rect 21928 25498 21956 25638
rect 21916 25492 21968 25498
rect 21916 25434 21968 25440
rect 21824 25288 21876 25294
rect 21824 25230 21876 25236
rect 21477 24508 21785 24517
rect 21477 24506 21483 24508
rect 21539 24506 21563 24508
rect 21619 24506 21643 24508
rect 21699 24506 21723 24508
rect 21779 24506 21785 24508
rect 21539 24454 21541 24506
rect 21721 24454 21723 24506
rect 21477 24452 21483 24454
rect 21539 24452 21563 24454
rect 21619 24452 21643 24454
rect 21699 24452 21723 24454
rect 21779 24452 21785 24454
rect 21477 24443 21785 24452
rect 21824 24064 21876 24070
rect 21824 24006 21876 24012
rect 21364 23724 21416 23730
rect 21364 23666 21416 23672
rect 21376 23322 21404 23666
rect 21477 23420 21785 23429
rect 21477 23418 21483 23420
rect 21539 23418 21563 23420
rect 21619 23418 21643 23420
rect 21699 23418 21723 23420
rect 21779 23418 21785 23420
rect 21539 23366 21541 23418
rect 21721 23366 21723 23418
rect 21477 23364 21483 23366
rect 21539 23364 21563 23366
rect 21619 23364 21643 23366
rect 21699 23364 21723 23366
rect 21779 23364 21785 23366
rect 21477 23355 21785 23364
rect 21364 23316 21416 23322
rect 21364 23258 21416 23264
rect 21272 23112 21324 23118
rect 21272 23054 21324 23060
rect 21477 22332 21785 22341
rect 21477 22330 21483 22332
rect 21539 22330 21563 22332
rect 21619 22330 21643 22332
rect 21699 22330 21723 22332
rect 21779 22330 21785 22332
rect 21539 22278 21541 22330
rect 21721 22278 21723 22330
rect 21477 22276 21483 22278
rect 21539 22276 21563 22278
rect 21619 22276 21643 22278
rect 21699 22276 21723 22278
rect 21779 22276 21785 22278
rect 21477 22267 21785 22276
rect 21456 22228 21508 22234
rect 21456 22170 21508 22176
rect 21008 22066 21312 22094
rect 20864 21972 20944 21978
rect 20812 21966 20944 21972
rect 21180 22024 21232 22030
rect 21180 21966 21232 21972
rect 20824 21950 20944 21966
rect 20640 21570 20668 21950
rect 20720 21888 20772 21894
rect 20720 21830 20772 21836
rect 20732 21690 20760 21830
rect 20720 21684 20772 21690
rect 20720 21626 20772 21632
rect 20640 21542 20760 21570
rect 20732 20874 20760 21542
rect 20720 20868 20772 20874
rect 20720 20810 20772 20816
rect 20720 20324 20772 20330
rect 20640 20284 20720 20312
rect 20640 19922 20668 20284
rect 20720 20266 20772 20272
rect 20628 19916 20680 19922
rect 20628 19858 20680 19864
rect 20628 19508 20680 19514
rect 20548 19468 20628 19496
rect 20628 19450 20680 19456
rect 20404 19332 20484 19360
rect 20352 19314 20404 19320
rect 20996 19168 21048 19174
rect 20996 19110 21048 19116
rect 20168 18896 20220 18902
rect 20168 18838 20220 18844
rect 21008 18698 21036 19110
rect 20996 18692 21048 18698
rect 20996 18634 21048 18640
rect 20444 18624 20496 18630
rect 20444 18566 20496 18572
rect 20168 18080 20220 18086
rect 20168 18022 20220 18028
rect 20076 17536 20128 17542
rect 20076 17478 20128 17484
rect 19984 15496 20036 15502
rect 19984 15438 20036 15444
rect 19996 15026 20024 15438
rect 19984 15020 20036 15026
rect 19984 14962 20036 14968
rect 19984 14408 20036 14414
rect 20036 14368 20116 14396
rect 19984 14350 20036 14356
rect 19812 13938 19840 14214
rect 19904 14198 20024 14226
rect 19892 14068 19944 14074
rect 19892 14010 19944 14016
rect 19800 13932 19852 13938
rect 19800 13874 19852 13880
rect 19812 12646 19840 13874
rect 19800 12640 19852 12646
rect 19800 12582 19852 12588
rect 19616 12436 19668 12442
rect 19616 12378 19668 12384
rect 19708 12436 19760 12442
rect 19708 12378 19760 12384
rect 19536 12192 19748 12220
rect 19432 12174 19484 12180
rect 19432 12096 19484 12102
rect 19338 12064 19394 12073
rect 19720 12050 19748 12192
rect 19432 12038 19484 12044
rect 19435 12022 19472 12038
rect 19338 11999 19394 12008
rect 19352 9081 19380 11999
rect 19444 10538 19472 12022
rect 19536 12022 19748 12050
rect 19432 10532 19484 10538
rect 19432 10474 19484 10480
rect 19432 9580 19484 9586
rect 19432 9522 19484 9528
rect 19338 9072 19394 9081
rect 19338 9007 19394 9016
rect 19340 8900 19392 8906
rect 19340 8842 19392 8848
rect 19352 8430 19380 8842
rect 19340 8424 19392 8430
rect 19340 8366 19392 8372
rect 19444 7886 19472 9522
rect 19536 8401 19564 12022
rect 19708 11756 19760 11762
rect 19708 11698 19760 11704
rect 19720 11150 19748 11698
rect 19812 11218 19840 12582
rect 19800 11212 19852 11218
rect 19800 11154 19852 11160
rect 19708 11144 19760 11150
rect 19708 11086 19760 11092
rect 19800 9920 19852 9926
rect 19800 9862 19852 9868
rect 19616 9580 19668 9586
rect 19616 9522 19668 9528
rect 19628 8634 19656 9522
rect 19812 9518 19840 9862
rect 19800 9512 19852 9518
rect 19800 9454 19852 9460
rect 19904 8922 19932 14010
rect 19996 12345 20024 14198
rect 20088 12434 20116 14368
rect 20180 14074 20208 18022
rect 20352 17128 20404 17134
rect 20352 17070 20404 17076
rect 20364 16046 20392 17070
rect 20352 16040 20404 16046
rect 20352 15982 20404 15988
rect 20352 15360 20404 15366
rect 20352 15302 20404 15308
rect 20364 14414 20392 15302
rect 20352 14408 20404 14414
rect 20352 14350 20404 14356
rect 20168 14068 20220 14074
rect 20168 14010 20220 14016
rect 20352 13796 20404 13802
rect 20352 13738 20404 13744
rect 20364 12850 20392 13738
rect 20352 12844 20404 12850
rect 20352 12786 20404 12792
rect 20260 12776 20312 12782
rect 20260 12718 20312 12724
rect 20272 12442 20300 12718
rect 20456 12646 20484 18566
rect 20812 18352 20864 18358
rect 20812 18294 20864 18300
rect 20720 18216 20772 18222
rect 20720 18158 20772 18164
rect 20732 17610 20760 18158
rect 20824 17610 20852 18294
rect 20720 17604 20772 17610
rect 20720 17546 20772 17552
rect 20812 17604 20864 17610
rect 20812 17546 20864 17552
rect 21192 17218 21220 21966
rect 21284 19496 21312 22066
rect 21362 21992 21418 22001
rect 21362 21927 21418 21936
rect 21376 21894 21404 21927
rect 21364 21888 21416 21894
rect 21364 21830 21416 21836
rect 21468 21554 21496 22170
rect 21456 21548 21508 21554
rect 21456 21490 21508 21496
rect 21477 21244 21785 21253
rect 21477 21242 21483 21244
rect 21539 21242 21563 21244
rect 21619 21242 21643 21244
rect 21699 21242 21723 21244
rect 21779 21242 21785 21244
rect 21539 21190 21541 21242
rect 21721 21190 21723 21242
rect 21477 21188 21483 21190
rect 21539 21188 21563 21190
rect 21619 21188 21643 21190
rect 21699 21188 21723 21190
rect 21779 21188 21785 21190
rect 21477 21179 21785 21188
rect 21456 20800 21508 20806
rect 21456 20742 21508 20748
rect 21468 20602 21496 20742
rect 21456 20596 21508 20602
rect 21456 20538 21508 20544
rect 21364 20256 21416 20262
rect 21364 20198 21416 20204
rect 21376 19854 21404 20198
rect 21477 20156 21785 20165
rect 21477 20154 21483 20156
rect 21539 20154 21563 20156
rect 21619 20154 21643 20156
rect 21699 20154 21723 20156
rect 21779 20154 21785 20156
rect 21539 20102 21541 20154
rect 21721 20102 21723 20154
rect 21477 20100 21483 20102
rect 21539 20100 21563 20102
rect 21619 20100 21643 20102
rect 21699 20100 21723 20102
rect 21779 20100 21785 20102
rect 21477 20091 21785 20100
rect 21364 19848 21416 19854
rect 21364 19790 21416 19796
rect 21284 19468 21404 19496
rect 21272 19372 21324 19378
rect 21272 19314 21324 19320
rect 20720 17196 20772 17202
rect 20720 17138 20772 17144
rect 20916 17190 21220 17218
rect 20732 17082 20760 17138
rect 20640 17054 20760 17082
rect 20640 16522 20668 17054
rect 20720 16992 20772 16998
rect 20720 16934 20772 16940
rect 20732 16590 20760 16934
rect 20720 16584 20772 16590
rect 20720 16526 20772 16532
rect 20628 16516 20680 16522
rect 20628 16458 20680 16464
rect 20812 15360 20864 15366
rect 20812 15302 20864 15308
rect 20628 15020 20680 15026
rect 20628 14962 20680 14968
rect 20640 14618 20668 14962
rect 20824 14822 20852 15302
rect 20812 14816 20864 14822
rect 20812 14758 20864 14764
rect 20628 14612 20680 14618
rect 20628 14554 20680 14560
rect 20812 14340 20864 14346
rect 20812 14282 20864 14288
rect 20824 13433 20852 14282
rect 20810 13424 20866 13433
rect 20810 13359 20866 13368
rect 20720 12912 20772 12918
rect 20720 12854 20772 12860
rect 20444 12640 20496 12646
rect 20444 12582 20496 12588
rect 20732 12442 20760 12854
rect 20260 12436 20312 12442
rect 20088 12406 20208 12434
rect 19982 12336 20038 12345
rect 19982 12271 20038 12280
rect 19996 11914 20024 12271
rect 20180 12209 20208 12406
rect 20260 12378 20312 12384
rect 20720 12436 20772 12442
rect 20720 12378 20772 12384
rect 20812 12232 20864 12238
rect 20166 12200 20222 12209
rect 20812 12174 20864 12180
rect 20166 12135 20222 12144
rect 19996 11886 20116 11914
rect 20088 11150 20116 11886
rect 20076 11144 20128 11150
rect 20076 11086 20128 11092
rect 20180 10690 20208 12135
rect 20824 11898 20852 12174
rect 20812 11892 20864 11898
rect 20812 11834 20864 11840
rect 20916 11098 20944 17190
rect 21088 16992 21140 16998
rect 21008 16952 21088 16980
rect 21008 16726 21036 16952
rect 21088 16934 21140 16940
rect 20996 16720 21048 16726
rect 20996 16662 21048 16668
rect 21008 16590 21036 16662
rect 20996 16584 21048 16590
rect 20996 16526 21048 16532
rect 21088 14884 21140 14890
rect 21088 14826 21140 14832
rect 20996 14816 21048 14822
rect 20996 14758 21048 14764
rect 21008 14618 21036 14758
rect 21100 14618 21128 14826
rect 20996 14612 21048 14618
rect 20996 14554 21048 14560
rect 21088 14612 21140 14618
rect 21088 14554 21140 14560
rect 21180 14272 21232 14278
rect 21180 14214 21232 14220
rect 21192 14006 21220 14214
rect 21180 14000 21232 14006
rect 21180 13942 21232 13948
rect 21088 13864 21140 13870
rect 21088 13806 21140 13812
rect 21100 13258 21128 13806
rect 21088 13252 21140 13258
rect 21088 13194 21140 13200
rect 21180 13252 21232 13258
rect 21180 13194 21232 13200
rect 21088 11552 21140 11558
rect 21088 11494 21140 11500
rect 20732 11070 20944 11098
rect 20352 11008 20404 11014
rect 20352 10950 20404 10956
rect 20088 10662 20208 10690
rect 19984 10056 20036 10062
rect 19984 9998 20036 10004
rect 19708 8900 19760 8906
rect 19708 8842 19760 8848
rect 19812 8894 19932 8922
rect 19720 8634 19748 8842
rect 19616 8628 19668 8634
rect 19616 8570 19668 8576
rect 19708 8628 19760 8634
rect 19708 8570 19760 8576
rect 19522 8392 19578 8401
rect 19522 8327 19578 8336
rect 19432 7880 19484 7886
rect 19432 7822 19484 7828
rect 19444 7410 19472 7822
rect 19432 7404 19484 7410
rect 19432 7346 19484 7352
rect 19260 6886 19380 6914
rect 19248 6792 19300 6798
rect 19248 6734 19300 6740
rect 19260 6458 19288 6734
rect 19352 6458 19380 6886
rect 19616 6656 19668 6662
rect 19616 6598 19668 6604
rect 19248 6452 19300 6458
rect 19248 6394 19300 6400
rect 19340 6452 19392 6458
rect 19340 6394 19392 6400
rect 19432 6316 19484 6322
rect 19432 6258 19484 6264
rect 19246 6216 19302 6225
rect 19246 6151 19302 6160
rect 19260 5710 19288 6151
rect 19444 5710 19472 6258
rect 19524 6112 19576 6118
rect 19524 6054 19576 6060
rect 19248 5704 19300 5710
rect 19248 5646 19300 5652
rect 19432 5704 19484 5710
rect 19432 5646 19484 5652
rect 19536 5642 19564 6054
rect 19628 5710 19656 6598
rect 19616 5704 19668 5710
rect 19616 5646 19668 5652
rect 19524 5636 19576 5642
rect 19524 5578 19576 5584
rect 19812 5522 19840 8894
rect 19892 8832 19944 8838
rect 19892 8774 19944 8780
rect 19904 8498 19932 8774
rect 19996 8634 20024 9998
rect 19984 8628 20036 8634
rect 19984 8570 20036 8576
rect 19892 8492 19944 8498
rect 19892 8434 19944 8440
rect 20088 7410 20116 10662
rect 20166 10568 20222 10577
rect 20166 10503 20222 10512
rect 20180 7410 20208 10503
rect 20260 9512 20312 9518
rect 20260 9454 20312 9460
rect 20272 9178 20300 9454
rect 20260 9172 20312 9178
rect 20260 9114 20312 9120
rect 20258 9072 20314 9081
rect 20258 9007 20314 9016
rect 20076 7404 20128 7410
rect 20076 7346 20128 7352
rect 20168 7404 20220 7410
rect 20168 7346 20220 7352
rect 19892 7200 19944 7206
rect 19892 7142 19944 7148
rect 19904 6390 19932 7142
rect 19984 6452 20036 6458
rect 19984 6394 20036 6400
rect 19892 6384 19944 6390
rect 19892 6326 19944 6332
rect 19996 5574 20024 6394
rect 20168 6112 20220 6118
rect 20168 6054 20220 6060
rect 20180 5710 20208 6054
rect 20168 5704 20220 5710
rect 20168 5646 20220 5652
rect 19628 5494 19840 5522
rect 19984 5568 20036 5574
rect 19984 5510 20036 5516
rect 19522 5400 19578 5409
rect 19340 5364 19392 5370
rect 19392 5324 19472 5352
rect 19522 5335 19578 5344
rect 19340 5306 19392 5312
rect 19444 5273 19472 5324
rect 19430 5264 19486 5273
rect 19248 5228 19300 5234
rect 19536 5244 19564 5335
rect 19430 5199 19486 5208
rect 19524 5238 19576 5244
rect 19524 5180 19576 5186
rect 19248 5170 19300 5176
rect 19156 5024 19208 5030
rect 19156 4966 19208 4972
rect 19168 4826 19196 4966
rect 19156 4820 19208 4826
rect 19156 4762 19208 4768
rect 19260 4146 19288 5170
rect 19340 4480 19392 4486
rect 19340 4422 19392 4428
rect 19248 4140 19300 4146
rect 19248 4082 19300 4088
rect 19248 3936 19300 3942
rect 19248 3878 19300 3884
rect 19260 3534 19288 3878
rect 19352 3738 19380 4422
rect 19430 4312 19486 4321
rect 19536 4282 19564 5180
rect 19430 4247 19486 4256
rect 19524 4276 19576 4282
rect 19444 4214 19472 4247
rect 19524 4218 19576 4224
rect 19432 4208 19484 4214
rect 19432 4150 19484 4156
rect 19430 3768 19486 3777
rect 19340 3732 19392 3738
rect 19430 3703 19432 3712
rect 19340 3674 19392 3680
rect 19484 3703 19486 3712
rect 19432 3674 19484 3680
rect 19248 3528 19300 3534
rect 19248 3470 19300 3476
rect 19432 3528 19484 3534
rect 19432 3470 19484 3476
rect 19156 3392 19208 3398
rect 19156 3334 19208 3340
rect 19064 3120 19116 3126
rect 19064 3062 19116 3068
rect 18972 3052 19024 3058
rect 18972 2994 19024 3000
rect 19168 2938 19196 3334
rect 19260 3194 19288 3470
rect 19340 3460 19392 3466
rect 19340 3402 19392 3408
rect 19352 3194 19380 3402
rect 19248 3188 19300 3194
rect 19248 3130 19300 3136
rect 19340 3188 19392 3194
rect 19340 3130 19392 3136
rect 18696 2916 18748 2922
rect 18696 2858 18748 2864
rect 19076 2910 19196 2938
rect 18708 2774 18736 2858
rect 19076 2854 19104 2910
rect 19064 2848 19116 2854
rect 19064 2790 19116 2796
rect 19156 2848 19208 2854
rect 19156 2790 19208 2796
rect 19248 2848 19300 2854
rect 19248 2790 19300 2796
rect 18708 2746 18920 2774
rect 18604 2304 18656 2310
rect 18604 2246 18656 2252
rect 18544 2204 18852 2213
rect 18544 2202 18550 2204
rect 18606 2202 18630 2204
rect 18686 2202 18710 2204
rect 18766 2202 18790 2204
rect 18846 2202 18852 2204
rect 18606 2150 18608 2202
rect 18788 2150 18790 2202
rect 18544 2148 18550 2150
rect 18606 2148 18630 2150
rect 18686 2148 18710 2150
rect 18766 2148 18790 2150
rect 18846 2148 18852 2150
rect 18544 2139 18852 2148
rect 18236 1352 18288 1358
rect 18236 1294 18288 1300
rect 18420 1352 18472 1358
rect 18420 1294 18472 1300
rect 18248 950 18276 1294
rect 18544 1116 18852 1125
rect 18544 1114 18550 1116
rect 18606 1114 18630 1116
rect 18686 1114 18710 1116
rect 18766 1114 18790 1116
rect 18846 1114 18852 1116
rect 18606 1062 18608 1114
rect 18788 1062 18790 1114
rect 18544 1060 18550 1062
rect 18606 1060 18630 1062
rect 18686 1060 18710 1062
rect 18766 1060 18790 1062
rect 18846 1060 18852 1062
rect 18544 1051 18852 1060
rect 18236 944 18288 950
rect 18236 886 18288 892
rect 18892 490 18920 2746
rect 19168 2666 19196 2790
rect 18800 462 18920 490
rect 18984 2638 19196 2666
rect 18326 82 18382 160
rect 18156 54 18382 82
rect 18326 -300 18382 54
rect 18602 82 18658 160
rect 18800 82 18828 462
rect 18984 354 19012 2638
rect 19156 2576 19208 2582
rect 19156 2518 19208 2524
rect 19168 2310 19196 2518
rect 19156 2304 19208 2310
rect 19156 2246 19208 2252
rect 19064 2100 19116 2106
rect 19064 2042 19116 2048
rect 19076 1834 19104 2042
rect 19064 1828 19116 1834
rect 19064 1770 19116 1776
rect 18892 326 19012 354
rect 18892 160 18920 326
rect 18602 54 18828 82
rect 18602 -300 18658 54
rect 18878 -300 18934 160
rect 19154 82 19210 160
rect 19260 82 19288 2790
rect 19340 2372 19392 2378
rect 19340 2314 19392 2320
rect 19352 1970 19380 2314
rect 19340 1964 19392 1970
rect 19340 1906 19392 1912
rect 19444 1358 19472 3470
rect 19524 3392 19576 3398
rect 19524 3334 19576 3340
rect 19432 1352 19484 1358
rect 19432 1294 19484 1300
rect 19340 1216 19392 1222
rect 19340 1158 19392 1164
rect 19352 882 19380 1158
rect 19340 876 19392 882
rect 19340 818 19392 824
rect 19536 796 19564 3334
rect 19628 3126 19656 5494
rect 20272 5386 20300 9007
rect 20364 7478 20392 10950
rect 20732 10010 20760 11070
rect 20812 11008 20864 11014
rect 20812 10950 20864 10956
rect 20996 11008 21048 11014
rect 20996 10950 21048 10956
rect 20824 10130 20852 10950
rect 20812 10124 20864 10130
rect 20812 10066 20864 10072
rect 20640 9982 20760 10010
rect 20640 9722 20668 9982
rect 20720 9920 20772 9926
rect 20720 9862 20772 9868
rect 20628 9716 20680 9722
rect 20628 9658 20680 9664
rect 20640 9466 20668 9658
rect 20732 9586 20760 9862
rect 20824 9722 20852 10066
rect 20904 10056 20956 10062
rect 20904 9998 20956 10004
rect 20916 9722 20944 9998
rect 20812 9716 20864 9722
rect 20812 9658 20864 9664
rect 20904 9716 20956 9722
rect 20904 9658 20956 9664
rect 20720 9580 20772 9586
rect 20720 9522 20772 9528
rect 20640 9438 20852 9466
rect 20536 9172 20588 9178
rect 20536 9114 20588 9120
rect 20352 7472 20404 7478
rect 20352 7414 20404 7420
rect 20364 5409 20392 7414
rect 20548 6202 20576 9114
rect 20628 8832 20680 8838
rect 20628 8774 20680 8780
rect 20718 8800 20774 8809
rect 20640 8634 20668 8774
rect 20718 8735 20774 8744
rect 20628 8628 20680 8634
rect 20628 8570 20680 8576
rect 20732 8430 20760 8735
rect 20720 8424 20772 8430
rect 20720 8366 20772 8372
rect 20718 7576 20774 7585
rect 20628 7540 20680 7546
rect 20718 7511 20774 7520
rect 20628 7482 20680 7488
rect 20640 6798 20668 7482
rect 20732 6866 20760 7511
rect 20824 7342 20852 9438
rect 21008 9058 21036 10950
rect 20916 9030 21036 9058
rect 20812 7336 20864 7342
rect 20812 7278 20864 7284
rect 20812 7200 20864 7206
rect 20812 7142 20864 7148
rect 20824 6866 20852 7142
rect 20720 6860 20772 6866
rect 20720 6802 20772 6808
rect 20812 6860 20864 6866
rect 20812 6802 20864 6808
rect 20628 6792 20680 6798
rect 20628 6734 20680 6740
rect 20628 6656 20680 6662
rect 20628 6598 20680 6604
rect 20810 6624 20866 6633
rect 20640 6458 20668 6598
rect 20810 6559 20866 6568
rect 20628 6452 20680 6458
rect 20628 6394 20680 6400
rect 20548 6174 20668 6202
rect 20536 6112 20588 6118
rect 20536 6054 20588 6060
rect 20548 5710 20576 6054
rect 20444 5704 20496 5710
rect 20444 5646 20496 5652
rect 20536 5704 20588 5710
rect 20536 5646 20588 5652
rect 19720 5358 20300 5386
rect 20350 5400 20406 5409
rect 19720 4162 19748 5358
rect 20350 5335 20406 5344
rect 19798 5264 19854 5273
rect 19798 5199 19800 5208
rect 19852 5199 19854 5208
rect 19800 5170 19852 5176
rect 20168 5160 20220 5166
rect 20168 5102 20220 5108
rect 20180 4826 20208 5102
rect 20260 5092 20312 5098
rect 20260 5034 20312 5040
rect 20168 4820 20220 4826
rect 20168 4762 20220 4768
rect 19996 4678 20208 4706
rect 20272 4690 20300 5034
rect 20352 5024 20404 5030
rect 20352 4966 20404 4972
rect 20364 4690 20392 4966
rect 19800 4616 19852 4622
rect 19996 4604 20024 4678
rect 19852 4576 20024 4604
rect 20076 4616 20128 4622
rect 19800 4558 19852 4564
rect 20076 4558 20128 4564
rect 19800 4480 19852 4486
rect 19982 4448 20038 4457
rect 19852 4428 19982 4434
rect 19800 4422 19982 4428
rect 19812 4406 19982 4422
rect 19982 4383 20038 4392
rect 19720 4134 19932 4162
rect 19706 4040 19762 4049
rect 19762 3998 19840 4026
rect 19706 3975 19762 3984
rect 19708 3936 19760 3942
rect 19708 3878 19760 3884
rect 19616 3120 19668 3126
rect 19616 3062 19668 3068
rect 19614 2680 19670 2689
rect 19614 2615 19670 2624
rect 19628 2446 19656 2615
rect 19616 2440 19668 2446
rect 19616 2382 19668 2388
rect 19616 1284 19668 1290
rect 19616 1226 19668 1232
rect 19628 1018 19656 1226
rect 19616 1012 19668 1018
rect 19616 954 19668 960
rect 19444 768 19564 796
rect 19444 160 19472 768
rect 19720 160 19748 3878
rect 19812 2854 19840 3998
rect 19904 2961 19932 4134
rect 19982 4040 20038 4049
rect 19982 3975 20038 3984
rect 19996 3534 20024 3975
rect 19984 3528 20036 3534
rect 19984 3470 20036 3476
rect 19890 2952 19946 2961
rect 19890 2887 19946 2896
rect 19800 2848 19852 2854
rect 19800 2790 19852 2796
rect 19892 2508 19944 2514
rect 19892 2450 19944 2456
rect 19904 2106 19932 2450
rect 20088 2106 20116 4558
rect 19892 2100 19944 2106
rect 19892 2042 19944 2048
rect 20076 2100 20128 2106
rect 20076 2042 20128 2048
rect 20180 2038 20208 4678
rect 20260 4684 20312 4690
rect 20260 4626 20312 4632
rect 20352 4684 20404 4690
rect 20352 4626 20404 4632
rect 20456 4622 20484 5646
rect 20536 5568 20588 5574
rect 20536 5510 20588 5516
rect 20444 4616 20496 4622
rect 20444 4558 20496 4564
rect 20260 4480 20312 4486
rect 20260 4422 20312 4428
rect 20272 4321 20300 4422
rect 20258 4312 20314 4321
rect 20258 4247 20314 4256
rect 20260 4140 20312 4146
rect 20260 4082 20312 4088
rect 20352 4140 20404 4146
rect 20352 4082 20404 4088
rect 20272 3738 20300 4082
rect 20260 3732 20312 3738
rect 20260 3674 20312 3680
rect 20364 3602 20392 4082
rect 20352 3596 20404 3602
rect 20352 3538 20404 3544
rect 20352 3392 20404 3398
rect 20352 3334 20404 3340
rect 20364 3233 20392 3334
rect 20350 3224 20406 3233
rect 20350 3159 20406 3168
rect 20260 3052 20312 3058
rect 20260 2994 20312 3000
rect 20352 3052 20404 3058
rect 20352 2994 20404 3000
rect 20272 2650 20300 2994
rect 20260 2644 20312 2650
rect 20260 2586 20312 2592
rect 19984 2032 20036 2038
rect 19984 1974 20036 1980
rect 20168 2032 20220 2038
rect 20168 1974 20220 1980
rect 19996 1873 20024 1974
rect 19982 1864 20038 1873
rect 19982 1799 20038 1808
rect 19996 160 20024 1799
rect 20168 1760 20220 1766
rect 20168 1702 20220 1708
rect 20180 1494 20208 1702
rect 20168 1488 20220 1494
rect 20168 1430 20220 1436
rect 19154 54 19288 82
rect 19154 -300 19210 54
rect 19430 -300 19486 160
rect 19706 -300 19762 160
rect 19982 -300 20038 160
rect 20258 82 20314 160
rect 20364 82 20392 2994
rect 20456 2650 20484 4558
rect 20548 4214 20576 5510
rect 20536 4208 20588 4214
rect 20536 4150 20588 4156
rect 20536 3936 20588 3942
rect 20536 3878 20588 3884
rect 20548 3097 20576 3878
rect 20534 3088 20590 3097
rect 20534 3023 20590 3032
rect 20640 2774 20668 6174
rect 20720 6112 20772 6118
rect 20720 6054 20772 6060
rect 20732 3210 20760 6054
rect 20824 3516 20852 6559
rect 20916 5370 20944 9030
rect 20996 8900 21048 8906
rect 20996 8842 21048 8848
rect 21008 8498 21036 8842
rect 20996 8492 21048 8498
rect 20996 8434 21048 8440
rect 20996 6792 21048 6798
rect 20996 6734 21048 6740
rect 21008 6458 21036 6734
rect 21100 6633 21128 11494
rect 21192 11234 21220 13194
rect 21284 12866 21312 19314
rect 21376 15366 21404 19468
rect 21477 19068 21785 19077
rect 21477 19066 21483 19068
rect 21539 19066 21563 19068
rect 21619 19066 21643 19068
rect 21699 19066 21723 19068
rect 21779 19066 21785 19068
rect 21539 19014 21541 19066
rect 21721 19014 21723 19066
rect 21477 19012 21483 19014
rect 21539 19012 21563 19014
rect 21619 19012 21643 19014
rect 21699 19012 21723 19014
rect 21779 19012 21785 19014
rect 21477 19003 21785 19012
rect 21836 18154 21864 24006
rect 21916 23520 21968 23526
rect 21916 23462 21968 23468
rect 21928 22642 21956 23462
rect 22020 23066 22048 25758
rect 22100 25288 22152 25294
rect 22100 25230 22152 25236
rect 22112 23730 22140 25230
rect 22100 23724 22152 23730
rect 22100 23666 22152 23672
rect 22020 23038 22140 23066
rect 22008 22976 22060 22982
rect 22008 22918 22060 22924
rect 22020 22778 22048 22918
rect 22008 22772 22060 22778
rect 22008 22714 22060 22720
rect 22112 22658 22140 23038
rect 21916 22636 21968 22642
rect 21916 22578 21968 22584
rect 22020 22630 22140 22658
rect 22020 22094 22048 22630
rect 21928 22066 22048 22094
rect 21928 21486 21956 22066
rect 22008 21548 22060 21554
rect 22008 21490 22060 21496
rect 21916 21480 21968 21486
rect 21916 21422 21968 21428
rect 22020 20874 22048 21490
rect 22204 21332 22232 28070
rect 22376 26512 22428 26518
rect 22376 26454 22428 26460
rect 22388 25906 22416 26454
rect 22376 25900 22428 25906
rect 22376 25842 22428 25848
rect 22572 24177 22600 31726
rect 22664 28082 22692 32370
rect 22756 28914 22784 33458
rect 22940 31754 22968 34886
rect 23202 34640 23258 34649
rect 23308 34626 23336 35430
rect 23400 35290 23428 35430
rect 23388 35284 23440 35290
rect 23388 35226 23440 35232
rect 23258 34598 23336 34626
rect 23202 34575 23258 34584
rect 23020 33312 23072 33318
rect 23020 33254 23072 33260
rect 23032 32910 23060 33254
rect 23020 32904 23072 32910
rect 23020 32846 23072 32852
rect 23388 31816 23440 31822
rect 23388 31758 23440 31764
rect 22940 31726 23060 31754
rect 22836 30592 22888 30598
rect 22836 30534 22888 30540
rect 22848 30258 22876 30534
rect 22836 30252 22888 30258
rect 22836 30194 22888 30200
rect 22928 30048 22980 30054
rect 22928 29990 22980 29996
rect 22940 29850 22968 29990
rect 22928 29844 22980 29850
rect 22928 29786 22980 29792
rect 22928 29300 22980 29306
rect 22928 29242 22980 29248
rect 22756 28886 22876 28914
rect 22652 28076 22704 28082
rect 22652 28018 22704 28024
rect 22744 27872 22796 27878
rect 22744 27814 22796 27820
rect 22756 27470 22784 27814
rect 22744 27464 22796 27470
rect 22744 27406 22796 27412
rect 22652 25696 22704 25702
rect 22652 25638 22704 25644
rect 22664 25294 22692 25638
rect 22652 25288 22704 25294
rect 22652 25230 22704 25236
rect 22652 24744 22704 24750
rect 22652 24686 22704 24692
rect 22558 24168 22614 24177
rect 22376 24132 22428 24138
rect 22558 24103 22614 24112
rect 22376 24074 22428 24080
rect 22388 23798 22416 24074
rect 22376 23792 22428 23798
rect 22376 23734 22428 23740
rect 22664 23322 22692 24686
rect 22652 23316 22704 23322
rect 22652 23258 22704 23264
rect 22664 22094 22692 23258
rect 22848 23118 22876 28886
rect 22836 23112 22888 23118
rect 22836 23054 22888 23060
rect 22940 22964 22968 29242
rect 22572 22066 22692 22094
rect 22848 22936 22968 22964
rect 22204 21304 22508 21332
rect 22192 20936 22244 20942
rect 22192 20878 22244 20884
rect 21916 20868 21968 20874
rect 21916 20810 21968 20816
rect 22008 20868 22060 20874
rect 22008 20810 22060 20816
rect 21824 18148 21876 18154
rect 21824 18090 21876 18096
rect 21477 17980 21785 17989
rect 21477 17978 21483 17980
rect 21539 17978 21563 17980
rect 21619 17978 21643 17980
rect 21699 17978 21723 17980
rect 21779 17978 21785 17980
rect 21539 17926 21541 17978
rect 21721 17926 21723 17978
rect 21477 17924 21483 17926
rect 21539 17924 21563 17926
rect 21619 17924 21643 17926
rect 21699 17924 21723 17926
rect 21779 17924 21785 17926
rect 21477 17915 21785 17924
rect 21456 17740 21508 17746
rect 21456 17682 21508 17688
rect 21468 17542 21496 17682
rect 21456 17536 21508 17542
rect 21456 17478 21508 17484
rect 21824 17536 21876 17542
rect 21824 17478 21876 17484
rect 21836 17338 21864 17478
rect 21824 17332 21876 17338
rect 21824 17274 21876 17280
rect 21477 16892 21785 16901
rect 21477 16890 21483 16892
rect 21539 16890 21563 16892
rect 21619 16890 21643 16892
rect 21699 16890 21723 16892
rect 21779 16890 21785 16892
rect 21539 16838 21541 16890
rect 21721 16838 21723 16890
rect 21477 16836 21483 16838
rect 21539 16836 21563 16838
rect 21619 16836 21643 16838
rect 21699 16836 21723 16838
rect 21779 16836 21785 16838
rect 21477 16827 21785 16836
rect 21456 16788 21508 16794
rect 21456 16730 21508 16736
rect 21468 16182 21496 16730
rect 21456 16176 21508 16182
rect 21456 16118 21508 16124
rect 21477 15804 21785 15813
rect 21477 15802 21483 15804
rect 21539 15802 21563 15804
rect 21619 15802 21643 15804
rect 21699 15802 21723 15804
rect 21779 15802 21785 15804
rect 21539 15750 21541 15802
rect 21721 15750 21723 15802
rect 21477 15748 21483 15750
rect 21539 15748 21563 15750
rect 21619 15748 21643 15750
rect 21699 15748 21723 15750
rect 21779 15748 21785 15750
rect 21477 15739 21785 15748
rect 21364 15360 21416 15366
rect 21364 15302 21416 15308
rect 21730 15056 21786 15065
rect 21786 15014 21864 15042
rect 21730 14991 21786 15000
rect 21364 14816 21416 14822
rect 21364 14758 21416 14764
rect 21376 14618 21404 14758
rect 21477 14716 21785 14725
rect 21477 14714 21483 14716
rect 21539 14714 21563 14716
rect 21619 14714 21643 14716
rect 21699 14714 21723 14716
rect 21779 14714 21785 14716
rect 21539 14662 21541 14714
rect 21721 14662 21723 14714
rect 21477 14660 21483 14662
rect 21539 14660 21563 14662
rect 21619 14660 21643 14662
rect 21699 14660 21723 14662
rect 21779 14660 21785 14662
rect 21477 14651 21785 14660
rect 21364 14612 21416 14618
rect 21364 14554 21416 14560
rect 21364 13728 21416 13734
rect 21364 13670 21416 13676
rect 21376 12986 21404 13670
rect 21477 13628 21785 13637
rect 21477 13626 21483 13628
rect 21539 13626 21563 13628
rect 21619 13626 21643 13628
rect 21699 13626 21723 13628
rect 21779 13626 21785 13628
rect 21539 13574 21541 13626
rect 21721 13574 21723 13626
rect 21477 13572 21483 13574
rect 21539 13572 21563 13574
rect 21619 13572 21643 13574
rect 21699 13572 21723 13574
rect 21779 13572 21785 13574
rect 21477 13563 21785 13572
rect 21364 12980 21416 12986
rect 21364 12922 21416 12928
rect 21456 12912 21508 12918
rect 21284 12860 21456 12866
rect 21284 12854 21508 12860
rect 21284 12838 21496 12854
rect 21364 12640 21416 12646
rect 21364 12582 21416 12588
rect 21376 12434 21404 12582
rect 21477 12540 21785 12549
rect 21477 12538 21483 12540
rect 21539 12538 21563 12540
rect 21619 12538 21643 12540
rect 21699 12538 21723 12540
rect 21779 12538 21785 12540
rect 21539 12486 21541 12538
rect 21721 12486 21723 12538
rect 21477 12484 21483 12486
rect 21539 12484 21563 12486
rect 21619 12484 21643 12486
rect 21699 12484 21723 12486
rect 21779 12484 21785 12486
rect 21477 12475 21785 12484
rect 21836 12434 21864 15014
rect 21376 12406 21496 12434
rect 21468 12238 21496 12406
rect 21560 12406 21864 12434
rect 21456 12232 21508 12238
rect 21456 12174 21508 12180
rect 21468 11762 21496 12174
rect 21456 11756 21508 11762
rect 21456 11698 21508 11704
rect 21560 11642 21588 12406
rect 21928 12306 21956 20810
rect 22100 20460 22152 20466
rect 22100 20402 22152 20408
rect 22112 20058 22140 20402
rect 22100 20052 22152 20058
rect 22100 19994 22152 20000
rect 22100 19712 22152 19718
rect 22100 19654 22152 19660
rect 22112 19378 22140 19654
rect 22204 19446 22232 20878
rect 22376 20324 22428 20330
rect 22376 20266 22428 20272
rect 22284 20256 22336 20262
rect 22284 20198 22336 20204
rect 22296 20058 22324 20198
rect 22284 20052 22336 20058
rect 22284 19994 22336 20000
rect 22388 19938 22416 20266
rect 22296 19910 22416 19938
rect 22192 19440 22244 19446
rect 22192 19382 22244 19388
rect 22100 19372 22152 19378
rect 22100 19314 22152 19320
rect 22296 18766 22324 19910
rect 22376 19372 22428 19378
rect 22376 19314 22428 19320
rect 22388 18766 22416 19314
rect 22284 18760 22336 18766
rect 22284 18702 22336 18708
rect 22376 18760 22428 18766
rect 22376 18702 22428 18708
rect 22192 18624 22244 18630
rect 22192 18566 22244 18572
rect 22204 18426 22232 18566
rect 22192 18420 22244 18426
rect 22192 18362 22244 18368
rect 22296 18306 22324 18702
rect 22204 18278 22324 18306
rect 22100 18080 22152 18086
rect 22100 18022 22152 18028
rect 22008 17672 22060 17678
rect 22008 17614 22060 17620
rect 22020 15026 22048 17614
rect 22112 16590 22140 18022
rect 22100 16584 22152 16590
rect 22100 16526 22152 16532
rect 22204 16454 22232 18278
rect 22376 17876 22428 17882
rect 22376 17818 22428 17824
rect 22284 16992 22336 16998
rect 22284 16934 22336 16940
rect 22296 16794 22324 16934
rect 22284 16788 22336 16794
rect 22284 16730 22336 16736
rect 22100 16448 22152 16454
rect 22100 16390 22152 16396
rect 22192 16448 22244 16454
rect 22192 16390 22244 16396
rect 22112 16250 22140 16390
rect 22100 16244 22152 16250
rect 22100 16186 22152 16192
rect 22204 15910 22232 16390
rect 22192 15904 22244 15910
rect 22192 15846 22244 15852
rect 22008 15020 22060 15026
rect 22008 14962 22060 14968
rect 22020 13394 22048 14962
rect 22204 14006 22232 15846
rect 22284 14068 22336 14074
rect 22284 14010 22336 14016
rect 22192 14000 22244 14006
rect 22192 13942 22244 13948
rect 22296 13938 22324 14010
rect 22100 13932 22152 13938
rect 22100 13874 22152 13880
rect 22284 13932 22336 13938
rect 22284 13874 22336 13880
rect 22112 13818 22140 13874
rect 22112 13790 22324 13818
rect 22192 13728 22244 13734
rect 22192 13670 22244 13676
rect 22008 13388 22060 13394
rect 22008 13330 22060 13336
rect 22204 12850 22232 13670
rect 22296 13190 22324 13790
rect 22388 13258 22416 17818
rect 22480 17354 22508 21304
rect 22572 20330 22600 22066
rect 22744 21344 22796 21350
rect 22744 21286 22796 21292
rect 22560 20324 22612 20330
rect 22560 20266 22612 20272
rect 22652 19712 22704 19718
rect 22652 19654 22704 19660
rect 22664 19514 22692 19654
rect 22652 19508 22704 19514
rect 22652 19450 22704 19456
rect 22756 18970 22784 21286
rect 22848 19310 22876 22936
rect 22928 22500 22980 22506
rect 22928 22442 22980 22448
rect 22836 19304 22888 19310
rect 22836 19246 22888 19252
rect 22836 19168 22888 19174
rect 22836 19110 22888 19116
rect 22744 18964 22796 18970
rect 22744 18906 22796 18912
rect 22744 18760 22796 18766
rect 22744 18702 22796 18708
rect 22560 18692 22612 18698
rect 22560 18634 22612 18640
rect 22572 18426 22600 18634
rect 22652 18624 22704 18630
rect 22652 18566 22704 18572
rect 22560 18420 22612 18426
rect 22560 18362 22612 18368
rect 22664 18290 22692 18566
rect 22652 18284 22704 18290
rect 22652 18226 22704 18232
rect 22756 17626 22784 18702
rect 22848 18290 22876 19110
rect 22836 18284 22888 18290
rect 22836 18226 22888 18232
rect 22664 17598 22784 17626
rect 22480 17326 22600 17354
rect 22468 16516 22520 16522
rect 22468 16458 22520 16464
rect 22480 16250 22508 16458
rect 22468 16244 22520 16250
rect 22468 16186 22520 16192
rect 22572 15314 22600 17326
rect 22664 15434 22692 17598
rect 22744 17536 22796 17542
rect 22744 17478 22796 17484
rect 22756 17202 22784 17478
rect 22744 17196 22796 17202
rect 22744 17138 22796 17144
rect 22836 16448 22888 16454
rect 22836 16390 22888 16396
rect 22652 15428 22704 15434
rect 22652 15370 22704 15376
rect 22572 15286 22784 15314
rect 22650 15192 22706 15201
rect 22650 15127 22706 15136
rect 22560 13932 22612 13938
rect 22560 13874 22612 13880
rect 22572 13530 22600 13874
rect 22664 13841 22692 15127
rect 22650 13832 22706 13841
rect 22650 13767 22706 13776
rect 22652 13728 22704 13734
rect 22652 13670 22704 13676
rect 22560 13524 22612 13530
rect 22560 13466 22612 13472
rect 22560 13320 22612 13326
rect 22560 13262 22612 13268
rect 22376 13252 22428 13258
rect 22376 13194 22428 13200
rect 22284 13184 22336 13190
rect 22284 13126 22336 13132
rect 22296 12850 22324 13126
rect 22192 12844 22244 12850
rect 22192 12786 22244 12792
rect 22284 12844 22336 12850
rect 22284 12786 22336 12792
rect 22190 12744 22246 12753
rect 22388 12730 22416 13194
rect 22190 12679 22246 12688
rect 22296 12702 22416 12730
rect 22204 12306 22232 12679
rect 21916 12300 21968 12306
rect 21916 12242 21968 12248
rect 22192 12300 22244 12306
rect 22192 12242 22244 12248
rect 21824 12232 21876 12238
rect 21824 12174 21876 12180
rect 22100 12232 22152 12238
rect 22100 12174 22152 12180
rect 21376 11614 21588 11642
rect 21192 11206 21312 11234
rect 21284 11150 21312 11206
rect 21272 11144 21324 11150
rect 21272 11086 21324 11092
rect 21180 9580 21232 9586
rect 21180 9522 21232 9528
rect 21192 8634 21220 9522
rect 21284 8974 21312 11086
rect 21272 8968 21324 8974
rect 21272 8910 21324 8916
rect 21180 8628 21232 8634
rect 21180 8570 21232 8576
rect 21376 7818 21404 11614
rect 21477 11452 21785 11461
rect 21477 11450 21483 11452
rect 21539 11450 21563 11452
rect 21619 11450 21643 11452
rect 21699 11450 21723 11452
rect 21779 11450 21785 11452
rect 21539 11398 21541 11450
rect 21721 11398 21723 11450
rect 21477 11396 21483 11398
rect 21539 11396 21563 11398
rect 21619 11396 21643 11398
rect 21699 11396 21723 11398
rect 21779 11396 21785 11398
rect 21477 11387 21785 11396
rect 21836 10810 21864 12174
rect 22112 11898 22140 12174
rect 22296 11898 22324 12702
rect 22100 11892 22152 11898
rect 22100 11834 22152 11840
rect 22284 11892 22336 11898
rect 22284 11834 22336 11840
rect 22376 11756 22428 11762
rect 22376 11698 22428 11704
rect 22388 11354 22416 11698
rect 22376 11348 22428 11354
rect 22376 11290 22428 11296
rect 22572 11218 22600 13262
rect 22664 12850 22692 13670
rect 22652 12844 22704 12850
rect 22652 12786 22704 12792
rect 22756 12646 22784 15286
rect 22848 15065 22876 16390
rect 22834 15056 22890 15065
rect 22834 14991 22890 15000
rect 22836 14544 22888 14550
rect 22836 14486 22888 14492
rect 22848 13870 22876 14486
rect 22836 13864 22888 13870
rect 22836 13806 22888 13812
rect 22940 13818 22968 22442
rect 23032 15201 23060 31726
rect 23204 31136 23256 31142
rect 23204 31078 23256 31084
rect 23216 30734 23244 31078
rect 23204 30728 23256 30734
rect 23204 30670 23256 30676
rect 23112 29640 23164 29646
rect 23112 29582 23164 29588
rect 23124 29306 23152 29582
rect 23112 29300 23164 29306
rect 23112 29242 23164 29248
rect 23204 29028 23256 29034
rect 23204 28970 23256 28976
rect 23400 28994 23428 31758
rect 23492 29730 23520 35550
rect 23584 35290 23612 36110
rect 23676 35834 23704 36722
rect 23664 35828 23716 35834
rect 23664 35770 23716 35776
rect 23572 35284 23624 35290
rect 23572 35226 23624 35232
rect 23664 32428 23716 32434
rect 23664 32370 23716 32376
rect 23676 32026 23704 32370
rect 23768 32298 23796 40394
rect 23860 36310 23888 41074
rect 23952 39098 23980 41262
rect 23940 39092 23992 39098
rect 23940 39034 23992 39040
rect 23940 38344 23992 38350
rect 23940 38286 23992 38292
rect 23952 38010 23980 38286
rect 23940 38004 23992 38010
rect 23940 37946 23992 37952
rect 23940 36780 23992 36786
rect 23940 36722 23992 36728
rect 23952 36378 23980 36722
rect 24044 36718 24072 41414
rect 24124 39840 24176 39846
rect 24122 39808 24124 39817
rect 24176 39808 24178 39817
rect 24122 39743 24178 39752
rect 24124 38752 24176 38758
rect 24122 38720 24124 38729
rect 24176 38720 24178 38729
rect 24122 38655 24178 38664
rect 24124 37664 24176 37670
rect 24122 37632 24124 37641
rect 24176 37632 24178 37641
rect 24122 37567 24178 37576
rect 24032 36712 24084 36718
rect 24032 36654 24084 36660
rect 24124 36576 24176 36582
rect 24122 36544 24124 36553
rect 24176 36544 24178 36553
rect 24122 36479 24178 36488
rect 23940 36372 23992 36378
rect 23940 36314 23992 36320
rect 23848 36304 23900 36310
rect 23848 36246 23900 36252
rect 24228 35834 24256 43182
rect 24320 41818 24348 43710
rect 24409 43548 24717 43557
rect 24409 43546 24415 43548
rect 24471 43546 24495 43548
rect 24551 43546 24575 43548
rect 24631 43546 24655 43548
rect 24711 43546 24717 43548
rect 24471 43494 24473 43546
rect 24653 43494 24655 43546
rect 24409 43492 24415 43494
rect 24471 43492 24495 43494
rect 24551 43492 24575 43494
rect 24631 43492 24655 43494
rect 24711 43492 24717 43494
rect 24409 43483 24717 43492
rect 24409 42460 24717 42469
rect 24409 42458 24415 42460
rect 24471 42458 24495 42460
rect 24551 42458 24575 42460
rect 24631 42458 24655 42460
rect 24711 42458 24717 42460
rect 24471 42406 24473 42458
rect 24653 42406 24655 42458
rect 24409 42404 24415 42406
rect 24471 42404 24495 42406
rect 24551 42404 24575 42406
rect 24631 42404 24655 42406
rect 24711 42404 24717 42406
rect 24409 42395 24717 42404
rect 24308 41812 24360 41818
rect 24308 41754 24360 41760
rect 24409 41372 24717 41381
rect 24409 41370 24415 41372
rect 24471 41370 24495 41372
rect 24551 41370 24575 41372
rect 24631 41370 24655 41372
rect 24711 41370 24717 41372
rect 24471 41318 24473 41370
rect 24653 41318 24655 41370
rect 24409 41316 24415 41318
rect 24471 41316 24495 41318
rect 24551 41316 24575 41318
rect 24631 41316 24655 41318
rect 24711 41316 24717 41318
rect 24409 41307 24717 41316
rect 24780 41274 24808 43710
rect 24858 42528 24914 42537
rect 24858 42463 24914 42472
rect 24872 42362 24900 42463
rect 24860 42356 24912 42362
rect 24860 42298 24912 42304
rect 24964 41614 24992 44540
rect 25136 41676 25188 41682
rect 25136 41618 25188 41624
rect 24952 41608 25004 41614
rect 24952 41550 25004 41556
rect 24768 41268 24820 41274
rect 24768 41210 24820 41216
rect 24952 40656 25004 40662
rect 24952 40598 25004 40604
rect 24964 40361 24992 40598
rect 25042 40488 25098 40497
rect 25042 40423 25098 40432
rect 24950 40352 25006 40361
rect 24409 40284 24717 40293
rect 24950 40287 25006 40296
rect 24409 40282 24415 40284
rect 24471 40282 24495 40284
rect 24551 40282 24575 40284
rect 24631 40282 24655 40284
rect 24711 40282 24717 40284
rect 24471 40230 24473 40282
rect 24653 40230 24655 40282
rect 24409 40228 24415 40230
rect 24471 40228 24495 40230
rect 24551 40228 24575 40230
rect 24631 40228 24655 40230
rect 24711 40228 24717 40230
rect 24409 40219 24717 40228
rect 24950 39536 25006 39545
rect 24950 39471 25006 39480
rect 24860 39296 24912 39302
rect 24858 39264 24860 39273
rect 24912 39264 24914 39273
rect 24409 39196 24717 39205
rect 24858 39199 24914 39208
rect 24409 39194 24415 39196
rect 24471 39194 24495 39196
rect 24551 39194 24575 39196
rect 24631 39194 24655 39196
rect 24711 39194 24717 39196
rect 24471 39142 24473 39194
rect 24653 39142 24655 39194
rect 24409 39140 24415 39142
rect 24471 39140 24495 39142
rect 24551 39140 24575 39142
rect 24631 39140 24655 39142
rect 24711 39140 24717 39142
rect 24409 39131 24717 39140
rect 24308 38820 24360 38826
rect 24308 38762 24360 38768
rect 24216 35828 24268 35834
rect 24216 35770 24268 35776
rect 24124 35488 24176 35494
rect 24122 35456 24124 35465
rect 24176 35456 24178 35465
rect 24122 35391 24178 35400
rect 24124 34536 24176 34542
rect 24122 34504 24124 34513
rect 24176 34504 24178 34513
rect 24122 34439 24178 34448
rect 23848 33992 23900 33998
rect 23848 33934 23900 33940
rect 23860 33658 23888 33934
rect 23848 33652 23900 33658
rect 23848 33594 23900 33600
rect 24214 33552 24270 33561
rect 24214 33487 24270 33496
rect 24124 33312 24176 33318
rect 24122 33280 24124 33289
rect 24176 33280 24178 33289
rect 24122 33215 24178 33224
rect 23756 32292 23808 32298
rect 23756 32234 23808 32240
rect 24124 32224 24176 32230
rect 24122 32192 24124 32201
rect 24176 32192 24178 32201
rect 24122 32127 24178 32136
rect 23664 32020 23716 32026
rect 23664 31962 23716 31968
rect 23572 31340 23624 31346
rect 23572 31282 23624 31288
rect 23848 31340 23900 31346
rect 23848 31282 23900 31288
rect 23584 30938 23612 31282
rect 23664 31136 23716 31142
rect 23664 31078 23716 31084
rect 23676 30938 23704 31078
rect 23572 30932 23624 30938
rect 23572 30874 23624 30880
rect 23664 30932 23716 30938
rect 23664 30874 23716 30880
rect 23860 30394 23888 31282
rect 24124 31136 24176 31142
rect 24122 31104 24124 31113
rect 24176 31104 24178 31113
rect 24122 31039 24178 31048
rect 24032 30660 24084 30666
rect 24032 30602 24084 30608
rect 23848 30388 23900 30394
rect 23848 30330 23900 30336
rect 23572 30252 23624 30258
rect 23572 30194 23624 30200
rect 23584 29850 23612 30194
rect 23664 30048 23716 30054
rect 23664 29990 23716 29996
rect 23676 29850 23704 29990
rect 23572 29844 23624 29850
rect 23572 29786 23624 29792
rect 23664 29844 23716 29850
rect 23664 29786 23716 29792
rect 23492 29702 23888 29730
rect 23480 29640 23532 29646
rect 23480 29582 23532 29588
rect 23492 29306 23520 29582
rect 23756 29572 23808 29578
rect 23756 29514 23808 29520
rect 23664 29504 23716 29510
rect 23664 29446 23716 29452
rect 23676 29306 23704 29446
rect 23480 29300 23532 29306
rect 23480 29242 23532 29248
rect 23664 29300 23716 29306
rect 23664 29242 23716 29248
rect 23112 28008 23164 28014
rect 23112 27950 23164 27956
rect 23124 27674 23152 27950
rect 23112 27668 23164 27674
rect 23112 27610 23164 27616
rect 23216 27538 23244 28970
rect 23400 28966 23520 28994
rect 23204 27532 23256 27538
rect 23204 27474 23256 27480
rect 23296 27464 23348 27470
rect 23296 27406 23348 27412
rect 23308 27146 23336 27406
rect 23216 27118 23336 27146
rect 23216 27062 23244 27118
rect 23204 27056 23256 27062
rect 23204 26998 23256 27004
rect 23388 25696 23440 25702
rect 23388 25638 23440 25644
rect 23400 25498 23428 25638
rect 23388 25492 23440 25498
rect 23388 25434 23440 25440
rect 23492 25242 23520 28966
rect 23572 27872 23624 27878
rect 23572 27814 23624 27820
rect 23584 25906 23612 27814
rect 23768 25906 23796 29514
rect 23572 25900 23624 25906
rect 23572 25842 23624 25848
rect 23756 25900 23808 25906
rect 23756 25842 23808 25848
rect 23664 25832 23716 25838
rect 23664 25774 23716 25780
rect 23676 25294 23704 25774
rect 23756 25696 23808 25702
rect 23754 25664 23756 25673
rect 23808 25664 23810 25673
rect 23754 25599 23810 25608
rect 23860 25514 23888 29702
rect 23940 28076 23992 28082
rect 23940 28018 23992 28024
rect 23952 27674 23980 28018
rect 23940 27668 23992 27674
rect 23940 27610 23992 27616
rect 24044 26466 24072 30602
rect 24124 30048 24176 30054
rect 24122 30016 24124 30025
rect 24176 30016 24178 30025
rect 24122 29951 24178 29960
rect 24124 29028 24176 29034
rect 24124 28970 24176 28976
rect 24136 28937 24164 28970
rect 24122 28928 24178 28937
rect 24122 28863 24178 28872
rect 24124 27872 24176 27878
rect 24122 27840 24124 27849
rect 24176 27840 24178 27849
rect 24122 27775 24178 27784
rect 24228 26790 24256 33487
rect 24124 26784 24176 26790
rect 24122 26752 24124 26761
rect 24216 26784 24268 26790
rect 24176 26752 24178 26761
rect 24216 26726 24268 26732
rect 24122 26687 24178 26696
rect 24044 26438 24256 26466
rect 24124 26308 24176 26314
rect 24124 26250 24176 26256
rect 24032 25968 24084 25974
rect 24032 25910 24084 25916
rect 23940 25764 23992 25770
rect 23940 25706 23992 25712
rect 23768 25486 23888 25514
rect 23664 25288 23716 25294
rect 23400 25214 23520 25242
rect 23584 25236 23664 25242
rect 23584 25230 23716 25236
rect 23584 25214 23704 25230
rect 23204 24064 23256 24070
rect 23204 24006 23256 24012
rect 23112 23044 23164 23050
rect 23112 22986 23164 22992
rect 23124 22778 23152 22986
rect 23112 22772 23164 22778
rect 23112 22714 23164 22720
rect 23216 22642 23244 24006
rect 23296 23520 23348 23526
rect 23296 23462 23348 23468
rect 23308 22778 23336 23462
rect 23296 22772 23348 22778
rect 23296 22714 23348 22720
rect 23204 22636 23256 22642
rect 23204 22578 23256 22584
rect 23400 22506 23428 25214
rect 23480 25152 23532 25158
rect 23480 25094 23532 25100
rect 23492 24954 23520 25094
rect 23584 24954 23612 25214
rect 23664 25152 23716 25158
rect 23664 25094 23716 25100
rect 23480 24948 23532 24954
rect 23480 24890 23532 24896
rect 23572 24948 23624 24954
rect 23572 24890 23624 24896
rect 23676 24206 23704 25094
rect 23664 24200 23716 24206
rect 23664 24142 23716 24148
rect 23768 24052 23796 25486
rect 23846 24576 23902 24585
rect 23846 24511 23902 24520
rect 23860 24410 23888 24511
rect 23848 24404 23900 24410
rect 23848 24346 23900 24352
rect 23676 24024 23796 24052
rect 23480 22976 23532 22982
rect 23480 22918 23532 22924
rect 23492 22574 23520 22918
rect 23480 22568 23532 22574
rect 23480 22510 23532 22516
rect 23388 22500 23440 22506
rect 23388 22442 23440 22448
rect 23204 21412 23256 21418
rect 23204 21354 23256 21360
rect 23388 21412 23440 21418
rect 23388 21354 23440 21360
rect 23112 19304 23164 19310
rect 23112 19246 23164 19252
rect 23018 15192 23074 15201
rect 23018 15127 23074 15136
rect 23020 15020 23072 15026
rect 23020 14962 23072 14968
rect 23032 14414 23060 14962
rect 23020 14408 23072 14414
rect 23020 14350 23072 14356
rect 23020 14272 23072 14278
rect 23020 14214 23072 14220
rect 23032 14006 23060 14214
rect 23020 14000 23072 14006
rect 23020 13942 23072 13948
rect 22940 13790 23060 13818
rect 22834 13424 22890 13433
rect 22834 13359 22890 13368
rect 22848 13258 22876 13359
rect 22836 13252 22888 13258
rect 22836 13194 22888 13200
rect 22744 12640 22796 12646
rect 22744 12582 22796 12588
rect 22652 11892 22704 11898
rect 22652 11834 22704 11840
rect 22664 11694 22692 11834
rect 22652 11688 22704 11694
rect 22652 11630 22704 11636
rect 22664 11506 22692 11630
rect 22664 11478 22784 11506
rect 22756 11218 22784 11478
rect 22560 11212 22612 11218
rect 22560 11154 22612 11160
rect 22744 11212 22796 11218
rect 22744 11154 22796 11160
rect 22560 11076 22612 11082
rect 22560 11018 22612 11024
rect 22376 11008 22428 11014
rect 22376 10950 22428 10956
rect 21824 10804 21876 10810
rect 21824 10746 21876 10752
rect 21824 10532 21876 10538
rect 21824 10474 21876 10480
rect 21477 10364 21785 10373
rect 21477 10362 21483 10364
rect 21539 10362 21563 10364
rect 21619 10362 21643 10364
rect 21699 10362 21723 10364
rect 21779 10362 21785 10364
rect 21539 10310 21541 10362
rect 21721 10310 21723 10362
rect 21477 10308 21483 10310
rect 21539 10308 21563 10310
rect 21619 10308 21643 10310
rect 21699 10308 21723 10310
rect 21779 10308 21785 10310
rect 21477 10299 21785 10308
rect 21548 9988 21600 9994
rect 21548 9930 21600 9936
rect 21560 9722 21588 9930
rect 21836 9722 21864 10474
rect 22388 10130 22416 10950
rect 22468 10736 22520 10742
rect 22468 10678 22520 10684
rect 22376 10124 22428 10130
rect 22376 10066 22428 10072
rect 21548 9716 21600 9722
rect 21548 9658 21600 9664
rect 21824 9716 21876 9722
rect 21824 9658 21876 9664
rect 22008 9580 22060 9586
rect 22008 9522 22060 9528
rect 21477 9276 21785 9285
rect 21477 9274 21483 9276
rect 21539 9274 21563 9276
rect 21619 9274 21643 9276
rect 21699 9274 21723 9276
rect 21779 9274 21785 9276
rect 21539 9222 21541 9274
rect 21721 9222 21723 9274
rect 21477 9220 21483 9222
rect 21539 9220 21563 9222
rect 21619 9220 21643 9222
rect 21699 9220 21723 9222
rect 21779 9220 21785 9222
rect 21477 9211 21785 9220
rect 22020 9178 22048 9522
rect 22008 9172 22060 9178
rect 22008 9114 22060 9120
rect 22100 9036 22152 9042
rect 22100 8978 22152 8984
rect 22008 8492 22060 8498
rect 22008 8434 22060 8440
rect 21824 8356 21876 8362
rect 21824 8298 21876 8304
rect 21477 8188 21785 8197
rect 21477 8186 21483 8188
rect 21539 8186 21563 8188
rect 21619 8186 21643 8188
rect 21699 8186 21723 8188
rect 21779 8186 21785 8188
rect 21539 8134 21541 8186
rect 21721 8134 21723 8186
rect 21477 8132 21483 8134
rect 21539 8132 21563 8134
rect 21619 8132 21643 8134
rect 21699 8132 21723 8134
rect 21779 8132 21785 8134
rect 21477 8123 21785 8132
rect 21364 7812 21416 7818
rect 21364 7754 21416 7760
rect 21180 7540 21232 7546
rect 21180 7482 21232 7488
rect 21086 6624 21142 6633
rect 21086 6559 21142 6568
rect 20996 6452 21048 6458
rect 20996 6394 21048 6400
rect 21088 6452 21140 6458
rect 21088 6394 21140 6400
rect 20904 5364 20956 5370
rect 20904 5306 20956 5312
rect 20904 5228 20956 5234
rect 20904 5170 20956 5176
rect 20996 5228 21048 5234
rect 20996 5170 21048 5176
rect 20916 4049 20944 5170
rect 20902 4040 20958 4049
rect 20902 3975 20958 3984
rect 20904 3528 20956 3534
rect 20824 3488 20904 3516
rect 20904 3470 20956 3476
rect 20902 3224 20958 3233
rect 20732 3182 20902 3210
rect 20902 3159 20958 3168
rect 20548 2746 20668 2774
rect 20444 2644 20496 2650
rect 20444 2586 20496 2592
rect 20548 882 20576 2746
rect 20628 2576 20680 2582
rect 20626 2544 20628 2553
rect 20680 2544 20682 2553
rect 20626 2479 20682 2488
rect 20812 2440 20864 2446
rect 20812 2382 20864 2388
rect 20628 2372 20680 2378
rect 20628 2314 20680 2320
rect 20720 2372 20772 2378
rect 20720 2314 20772 2320
rect 20536 876 20588 882
rect 20536 818 20588 824
rect 20258 54 20392 82
rect 20534 82 20590 160
rect 20640 82 20668 2314
rect 20732 1902 20760 2314
rect 20720 1896 20772 1902
rect 20720 1838 20772 1844
rect 20720 1352 20772 1358
rect 20720 1294 20772 1300
rect 20732 1193 20760 1294
rect 20718 1184 20774 1193
rect 20718 1119 20774 1128
rect 20824 160 20852 2382
rect 20916 2038 20944 3159
rect 21008 2961 21036 5170
rect 21100 4457 21128 6394
rect 21192 5642 21220 7482
rect 21364 7336 21416 7342
rect 21364 7278 21416 7284
rect 21376 6474 21404 7278
rect 21477 7100 21785 7109
rect 21477 7098 21483 7100
rect 21539 7098 21563 7100
rect 21619 7098 21643 7100
rect 21699 7098 21723 7100
rect 21779 7098 21785 7100
rect 21539 7046 21541 7098
rect 21721 7046 21723 7098
rect 21477 7044 21483 7046
rect 21539 7044 21563 7046
rect 21619 7044 21643 7046
rect 21699 7044 21723 7046
rect 21779 7044 21785 7046
rect 21477 7035 21785 7044
rect 21836 6934 21864 8298
rect 22020 8072 22048 8434
rect 22112 8430 22140 8978
rect 22192 8968 22244 8974
rect 22192 8910 22244 8916
rect 22284 8968 22336 8974
rect 22284 8910 22336 8916
rect 22204 8430 22232 8910
rect 22100 8424 22152 8430
rect 22100 8366 22152 8372
rect 22192 8424 22244 8430
rect 22192 8366 22244 8372
rect 22192 8084 22244 8090
rect 22020 8044 22192 8072
rect 22192 8026 22244 8032
rect 22296 8022 22324 8910
rect 22376 8492 22428 8498
rect 22376 8434 22428 8440
rect 22284 8016 22336 8022
rect 22284 7958 22336 7964
rect 22100 7472 22152 7478
rect 22100 7414 22152 7420
rect 21824 6928 21876 6934
rect 21824 6870 21876 6876
rect 21376 6446 21956 6474
rect 21272 6316 21324 6322
rect 21272 6258 21324 6264
rect 21364 6316 21416 6322
rect 21364 6258 21416 6264
rect 21824 6316 21876 6322
rect 21824 6258 21876 6264
rect 21180 5636 21232 5642
rect 21180 5578 21232 5584
rect 21180 5024 21232 5030
rect 21180 4966 21232 4972
rect 21086 4448 21142 4457
rect 21086 4383 21142 4392
rect 21088 4004 21140 4010
rect 21088 3946 21140 3952
rect 21100 3534 21128 3946
rect 21192 3890 21220 4966
rect 21284 4010 21312 6258
rect 21376 5098 21404 6258
rect 21546 6216 21602 6225
rect 21546 6151 21602 6160
rect 21560 6118 21588 6151
rect 21548 6112 21600 6118
rect 21548 6054 21600 6060
rect 21477 6012 21785 6021
rect 21477 6010 21483 6012
rect 21539 6010 21563 6012
rect 21619 6010 21643 6012
rect 21699 6010 21723 6012
rect 21779 6010 21785 6012
rect 21539 5958 21541 6010
rect 21721 5958 21723 6010
rect 21477 5956 21483 5958
rect 21539 5956 21563 5958
rect 21619 5956 21643 5958
rect 21699 5956 21723 5958
rect 21779 5956 21785 5958
rect 21477 5947 21785 5956
rect 21364 5092 21416 5098
rect 21364 5034 21416 5040
rect 21477 4924 21785 4933
rect 21477 4922 21483 4924
rect 21539 4922 21563 4924
rect 21619 4922 21643 4924
rect 21699 4922 21723 4924
rect 21779 4922 21785 4924
rect 21539 4870 21541 4922
rect 21721 4870 21723 4922
rect 21477 4868 21483 4870
rect 21539 4868 21563 4870
rect 21619 4868 21643 4870
rect 21699 4868 21723 4870
rect 21779 4868 21785 4870
rect 21477 4859 21785 4868
rect 21836 4808 21864 6258
rect 21928 5386 21956 6446
rect 22112 6322 22140 7414
rect 22388 6882 22416 8434
rect 22204 6854 22416 6882
rect 22100 6316 22152 6322
rect 22100 6258 22152 6264
rect 22100 5908 22152 5914
rect 22100 5850 22152 5856
rect 21928 5358 22048 5386
rect 21916 5228 21968 5234
rect 21916 5170 21968 5176
rect 21928 4826 21956 5170
rect 22020 5030 22048 5358
rect 22112 5098 22140 5850
rect 22204 5778 22232 6854
rect 22284 6792 22336 6798
rect 22284 6734 22336 6740
rect 22296 5914 22324 6734
rect 22376 6112 22428 6118
rect 22376 6054 22428 6060
rect 22284 5908 22336 5914
rect 22284 5850 22336 5856
rect 22192 5772 22244 5778
rect 22192 5714 22244 5720
rect 22284 5704 22336 5710
rect 22284 5646 22336 5652
rect 22190 5400 22246 5409
rect 22190 5335 22246 5344
rect 22100 5092 22152 5098
rect 22100 5034 22152 5040
rect 22008 5024 22060 5030
rect 22008 4966 22060 4972
rect 21560 4780 21864 4808
rect 21560 4010 21588 4780
rect 21638 4720 21694 4729
rect 21638 4655 21694 4664
rect 21652 4214 21680 4655
rect 21640 4208 21692 4214
rect 21640 4150 21692 4156
rect 21732 4072 21784 4078
rect 21732 4014 21784 4020
rect 21272 4004 21324 4010
rect 21272 3946 21324 3952
rect 21548 4004 21600 4010
rect 21548 3946 21600 3952
rect 21744 3924 21772 4014
rect 21836 3992 21864 4780
rect 21916 4820 21968 4826
rect 21916 4762 21968 4768
rect 22204 4690 22232 5335
rect 22192 4684 22244 4690
rect 22192 4626 22244 4632
rect 21916 4616 21968 4622
rect 21916 4558 21968 4564
rect 22100 4616 22152 4622
rect 22100 4558 22152 4564
rect 21928 4214 21956 4558
rect 21916 4208 21968 4214
rect 21916 4150 21968 4156
rect 22008 4140 22060 4146
rect 22008 4082 22060 4088
rect 21836 3964 21956 3992
rect 21744 3896 21864 3924
rect 21192 3862 21404 3890
rect 21088 3528 21140 3534
rect 21088 3470 21140 3476
rect 20994 2952 21050 2961
rect 20994 2887 21050 2896
rect 21272 2916 21324 2922
rect 21272 2858 21324 2864
rect 21284 2774 21312 2858
rect 21192 2746 21312 2774
rect 21086 2408 21142 2417
rect 21086 2343 21142 2352
rect 20904 2032 20956 2038
rect 20904 1974 20956 1980
rect 21100 1902 21128 2343
rect 21088 1896 21140 1902
rect 21088 1838 21140 1844
rect 20904 1828 20956 1834
rect 20904 1770 20956 1776
rect 20916 1562 20944 1770
rect 20904 1556 20956 1562
rect 20904 1498 20956 1504
rect 20996 1284 21048 1290
rect 20996 1226 21048 1232
rect 21008 610 21036 1226
rect 20996 604 21048 610
rect 20996 546 21048 552
rect 20534 54 20668 82
rect 20258 -300 20314 54
rect 20534 -300 20590 54
rect 20810 -300 20866 160
rect 21086 82 21142 160
rect 21192 82 21220 2746
rect 21376 2378 21404 3862
rect 21477 3836 21785 3845
rect 21477 3834 21483 3836
rect 21539 3834 21563 3836
rect 21619 3834 21643 3836
rect 21699 3834 21723 3836
rect 21779 3834 21785 3836
rect 21539 3782 21541 3834
rect 21721 3782 21723 3834
rect 21477 3780 21483 3782
rect 21539 3780 21563 3782
rect 21619 3780 21643 3782
rect 21699 3780 21723 3782
rect 21779 3780 21785 3782
rect 21477 3771 21785 3780
rect 21836 3602 21864 3896
rect 21824 3596 21876 3602
rect 21824 3538 21876 3544
rect 21824 3460 21876 3466
rect 21824 3402 21876 3408
rect 21638 3360 21694 3369
rect 21638 3295 21694 3304
rect 21652 3058 21680 3295
rect 21640 3052 21692 3058
rect 21640 2994 21692 3000
rect 21477 2748 21785 2757
rect 21477 2746 21483 2748
rect 21539 2746 21563 2748
rect 21619 2746 21643 2748
rect 21699 2746 21723 2748
rect 21779 2746 21785 2748
rect 21539 2694 21541 2746
rect 21721 2694 21723 2746
rect 21477 2692 21483 2694
rect 21539 2692 21563 2694
rect 21619 2692 21643 2694
rect 21699 2692 21723 2694
rect 21779 2692 21785 2694
rect 21477 2683 21785 2692
rect 21548 2644 21600 2650
rect 21548 2586 21600 2592
rect 21364 2372 21416 2378
rect 21364 2314 21416 2320
rect 21560 1902 21588 2586
rect 21836 2553 21864 3402
rect 21928 3126 21956 3964
rect 21916 3120 21968 3126
rect 21916 3062 21968 3068
rect 21822 2544 21878 2553
rect 21822 2479 21878 2488
rect 21824 2440 21876 2446
rect 21824 2382 21876 2388
rect 21548 1896 21600 1902
rect 21546 1864 21548 1873
rect 21600 1864 21602 1873
rect 21546 1799 21602 1808
rect 21477 1660 21785 1669
rect 21477 1658 21483 1660
rect 21539 1658 21563 1660
rect 21619 1658 21643 1660
rect 21699 1658 21723 1660
rect 21779 1658 21785 1660
rect 21539 1606 21541 1658
rect 21721 1606 21723 1658
rect 21477 1604 21483 1606
rect 21539 1604 21563 1606
rect 21619 1604 21643 1606
rect 21699 1604 21723 1606
rect 21779 1604 21785 1606
rect 21477 1595 21785 1604
rect 21548 1284 21600 1290
rect 21548 1226 21600 1232
rect 21086 54 21220 82
rect 21362 82 21418 160
rect 21560 82 21588 1226
rect 21362 54 21588 82
rect 21638 82 21694 160
rect 21836 82 21864 2382
rect 22020 1737 22048 4082
rect 22112 4078 22140 4558
rect 22296 4196 22324 5646
rect 22388 4298 22416 6054
rect 22480 5930 22508 10678
rect 22572 10674 22600 11018
rect 22756 10742 22784 11154
rect 22928 11144 22980 11150
rect 22928 11086 22980 11092
rect 22744 10736 22796 10742
rect 22744 10678 22796 10684
rect 22560 10668 22612 10674
rect 22560 10610 22612 10616
rect 22572 8022 22600 10610
rect 22652 10464 22704 10470
rect 22652 10406 22704 10412
rect 22664 10062 22692 10406
rect 22652 10056 22704 10062
rect 22652 9998 22704 10004
rect 22756 9518 22784 10678
rect 22836 10668 22888 10674
rect 22836 10610 22888 10616
rect 22744 9512 22796 9518
rect 22744 9454 22796 9460
rect 22756 9110 22784 9454
rect 22744 9104 22796 9110
rect 22744 9046 22796 9052
rect 22560 8016 22612 8022
rect 22560 7958 22612 7964
rect 22560 6792 22612 6798
rect 22560 6734 22612 6740
rect 22572 6118 22600 6734
rect 22848 6322 22876 10610
rect 22836 6316 22888 6322
rect 22836 6258 22888 6264
rect 22560 6112 22612 6118
rect 22560 6054 22612 6060
rect 22480 5902 22600 5930
rect 22468 5840 22520 5846
rect 22466 5808 22468 5817
rect 22520 5808 22522 5817
rect 22466 5743 22522 5752
rect 22388 4270 22508 4298
rect 22296 4168 22416 4196
rect 22100 4072 22152 4078
rect 22100 4014 22152 4020
rect 22284 3664 22336 3670
rect 22190 3632 22246 3641
rect 22284 3606 22336 3612
rect 22190 3567 22246 3576
rect 22204 3534 22232 3567
rect 22192 3528 22244 3534
rect 22296 3505 22324 3606
rect 22192 3470 22244 3476
rect 22282 3496 22338 3505
rect 22282 3431 22338 3440
rect 22100 3052 22152 3058
rect 22100 2994 22152 3000
rect 22284 3052 22336 3058
rect 22284 2994 22336 3000
rect 22112 2938 22140 2994
rect 22112 2922 22232 2938
rect 22112 2916 22244 2922
rect 22112 2910 22192 2916
rect 22192 2858 22244 2864
rect 22190 2680 22246 2689
rect 22296 2650 22324 2994
rect 22190 2615 22246 2624
rect 22284 2644 22336 2650
rect 22100 2576 22152 2582
rect 22100 2518 22152 2524
rect 22006 1728 22062 1737
rect 22006 1663 22062 1672
rect 21916 1352 21968 1358
rect 21916 1294 21968 1300
rect 21928 160 21956 1294
rect 22112 1018 22140 2518
rect 22204 2417 22232 2615
rect 22284 2586 22336 2592
rect 22190 2408 22246 2417
rect 22190 2343 22246 2352
rect 22204 1358 22232 2343
rect 22192 1352 22244 1358
rect 22192 1294 22244 1300
rect 22192 1216 22244 1222
rect 22192 1158 22244 1164
rect 22284 1216 22336 1222
rect 22284 1158 22336 1164
rect 22100 1012 22152 1018
rect 22100 954 22152 960
rect 22204 160 22232 1158
rect 22296 882 22324 1158
rect 22284 876 22336 882
rect 22284 818 22336 824
rect 22388 649 22416 4168
rect 22480 3534 22508 4270
rect 22468 3528 22520 3534
rect 22468 3470 22520 3476
rect 22572 3176 22600 5902
rect 22652 5840 22704 5846
rect 22652 5782 22704 5788
rect 22664 4622 22692 5782
rect 22744 5704 22796 5710
rect 22744 5646 22796 5652
rect 22652 4616 22704 4622
rect 22652 4558 22704 4564
rect 22756 3913 22784 5646
rect 22836 4616 22888 4622
rect 22836 4558 22888 4564
rect 22742 3904 22798 3913
rect 22742 3839 22798 3848
rect 22744 3460 22796 3466
rect 22744 3402 22796 3408
rect 22652 3188 22704 3194
rect 22572 3148 22652 3176
rect 22652 3130 22704 3136
rect 22756 2922 22784 3402
rect 22744 2916 22796 2922
rect 22744 2858 22796 2864
rect 22848 2292 22876 4558
rect 22940 4146 22968 11086
rect 23032 9058 23060 13790
rect 23124 10742 23152 19246
rect 23216 11082 23244 21354
rect 23400 19854 23428 21354
rect 23388 19848 23440 19854
rect 23388 19790 23440 19796
rect 23572 19780 23624 19786
rect 23572 19722 23624 19728
rect 23584 19514 23612 19722
rect 23572 19508 23624 19514
rect 23572 19450 23624 19456
rect 23388 18964 23440 18970
rect 23388 18906 23440 18912
rect 23400 18290 23428 18906
rect 23388 18284 23440 18290
rect 23388 18226 23440 18232
rect 23572 18080 23624 18086
rect 23570 18048 23572 18057
rect 23624 18048 23626 18057
rect 23570 17983 23626 17992
rect 23388 17536 23440 17542
rect 23388 17478 23440 17484
rect 23400 17338 23428 17478
rect 23388 17332 23440 17338
rect 23388 17274 23440 17280
rect 23480 16992 23532 16998
rect 23572 16992 23624 16998
rect 23480 16934 23532 16940
rect 23570 16960 23572 16969
rect 23624 16960 23626 16969
rect 23492 16794 23520 16934
rect 23570 16895 23626 16904
rect 23676 16810 23704 24024
rect 23952 23798 23980 25706
rect 24044 24954 24072 25910
rect 24032 24948 24084 24954
rect 24032 24890 24084 24896
rect 24136 24206 24164 26250
rect 24228 24682 24256 26438
rect 24216 24676 24268 24682
rect 24216 24618 24268 24624
rect 24124 24200 24176 24206
rect 24124 24142 24176 24148
rect 23940 23792 23992 23798
rect 23940 23734 23992 23740
rect 24124 23520 24176 23526
rect 24122 23488 24124 23497
rect 24176 23488 24178 23497
rect 24122 23423 24178 23432
rect 24032 23112 24084 23118
rect 24032 23054 24084 23060
rect 24044 22778 24072 23054
rect 24032 22772 24084 22778
rect 24032 22714 24084 22720
rect 23756 22432 23808 22438
rect 23754 22400 23756 22409
rect 23808 22400 23810 22409
rect 23754 22335 23810 22344
rect 23848 21548 23900 21554
rect 23848 21490 23900 21496
rect 23860 21146 23888 21490
rect 24032 21344 24084 21350
rect 24124 21344 24176 21350
rect 24032 21286 24084 21292
rect 24122 21312 24124 21321
rect 24176 21312 24178 21321
rect 23848 21140 23900 21146
rect 23848 21082 23900 21088
rect 23848 20256 23900 20262
rect 23754 20224 23810 20233
rect 23848 20198 23900 20204
rect 23754 20159 23810 20168
rect 23768 20058 23796 20159
rect 23756 20052 23808 20058
rect 23756 19994 23808 20000
rect 23860 19922 23888 20198
rect 24044 20058 24072 21286
rect 24122 21247 24178 21256
rect 24032 20052 24084 20058
rect 24032 19994 24084 20000
rect 23848 19916 23900 19922
rect 23848 19858 23900 19864
rect 24216 19712 24268 19718
rect 24216 19654 24268 19660
rect 23940 19168 23992 19174
rect 23938 19136 23940 19145
rect 23992 19136 23994 19145
rect 23938 19071 23994 19080
rect 23940 18760 23992 18766
rect 23940 18702 23992 18708
rect 23848 18624 23900 18630
rect 23848 18566 23900 18572
rect 23860 17678 23888 18566
rect 23952 18426 23980 18702
rect 23940 18420 23992 18426
rect 23940 18362 23992 18368
rect 24228 17678 24256 19654
rect 23848 17672 23900 17678
rect 23848 17614 23900 17620
rect 24216 17672 24268 17678
rect 24216 17614 24268 17620
rect 23756 17196 23808 17202
rect 23756 17138 23808 17144
rect 23848 17196 23900 17202
rect 23848 17138 23900 17144
rect 23480 16788 23532 16794
rect 23480 16730 23532 16736
rect 23584 16782 23704 16810
rect 23768 16794 23796 17138
rect 23756 16788 23808 16794
rect 23296 14816 23348 14822
rect 23296 14758 23348 14764
rect 23308 14550 23336 14758
rect 23296 14544 23348 14550
rect 23296 14486 23348 14492
rect 23296 12980 23348 12986
rect 23296 12922 23348 12928
rect 23308 12866 23336 12922
rect 23308 12838 23520 12866
rect 23492 12238 23520 12838
rect 23480 12232 23532 12238
rect 23480 12174 23532 12180
rect 23204 11076 23256 11082
rect 23204 11018 23256 11024
rect 23112 10736 23164 10742
rect 23112 10678 23164 10684
rect 23584 10554 23612 16782
rect 23756 16730 23808 16736
rect 23756 15904 23808 15910
rect 23754 15872 23756 15881
rect 23808 15872 23810 15881
rect 23754 15807 23810 15816
rect 23860 15502 23888 17138
rect 24124 16992 24176 16998
rect 24124 16934 24176 16940
rect 24136 16794 24164 16934
rect 24124 16788 24176 16794
rect 24124 16730 24176 16736
rect 23848 15496 23900 15502
rect 23848 15438 23900 15444
rect 24124 14816 24176 14822
rect 24122 14784 24124 14793
rect 24176 14784 24178 14793
rect 24122 14719 24178 14728
rect 23756 14612 23808 14618
rect 23756 14554 23808 14560
rect 23768 14414 23796 14554
rect 23756 14408 23808 14414
rect 23756 14350 23808 14356
rect 23848 14408 23900 14414
rect 23848 14350 23900 14356
rect 23768 14006 23796 14350
rect 23860 14074 23888 14350
rect 23848 14068 23900 14074
rect 23848 14010 23900 14016
rect 23756 14000 23808 14006
rect 23756 13942 23808 13948
rect 24122 13696 24178 13705
rect 24122 13631 24178 13640
rect 24136 13530 24164 13631
rect 24124 13524 24176 13530
rect 24124 13466 24176 13472
rect 23940 12640 23992 12646
rect 23938 12608 23940 12617
rect 23992 12608 23994 12617
rect 23938 12543 23994 12552
rect 24320 12434 24348 38762
rect 24860 38208 24912 38214
rect 24858 38176 24860 38185
rect 24912 38176 24914 38185
rect 24409 38108 24717 38117
rect 24858 38111 24914 38120
rect 24409 38106 24415 38108
rect 24471 38106 24495 38108
rect 24551 38106 24575 38108
rect 24631 38106 24655 38108
rect 24711 38106 24717 38108
rect 24471 38054 24473 38106
rect 24653 38054 24655 38106
rect 24409 38052 24415 38054
rect 24471 38052 24495 38054
rect 24551 38052 24575 38054
rect 24631 38052 24655 38054
rect 24711 38052 24717 38054
rect 24409 38043 24717 38052
rect 24860 37120 24912 37126
rect 24858 37088 24860 37097
rect 24912 37088 24914 37097
rect 24409 37020 24717 37029
rect 24858 37023 24914 37032
rect 24409 37018 24415 37020
rect 24471 37018 24495 37020
rect 24551 37018 24575 37020
rect 24631 37018 24655 37020
rect 24711 37018 24717 37020
rect 24471 36966 24473 37018
rect 24653 36966 24655 37018
rect 24409 36964 24415 36966
rect 24471 36964 24495 36966
rect 24551 36964 24575 36966
rect 24631 36964 24655 36966
rect 24711 36964 24717 36966
rect 24409 36955 24717 36964
rect 24964 36650 24992 39471
rect 24952 36644 25004 36650
rect 24952 36586 25004 36592
rect 25056 36530 25084 40423
rect 24780 36502 25084 36530
rect 24409 35932 24717 35941
rect 24409 35930 24415 35932
rect 24471 35930 24495 35932
rect 24551 35930 24575 35932
rect 24631 35930 24655 35932
rect 24711 35930 24717 35932
rect 24471 35878 24473 35930
rect 24653 35878 24655 35930
rect 24409 35876 24415 35878
rect 24471 35876 24495 35878
rect 24551 35876 24575 35878
rect 24631 35876 24655 35878
rect 24711 35876 24717 35878
rect 24409 35867 24717 35876
rect 24409 34844 24717 34853
rect 24409 34842 24415 34844
rect 24471 34842 24495 34844
rect 24551 34842 24575 34844
rect 24631 34842 24655 34844
rect 24711 34842 24717 34844
rect 24471 34790 24473 34842
rect 24653 34790 24655 34842
rect 24409 34788 24415 34790
rect 24471 34788 24495 34790
rect 24551 34788 24575 34790
rect 24631 34788 24655 34790
rect 24711 34788 24717 34790
rect 24409 34779 24717 34788
rect 24409 33756 24717 33765
rect 24409 33754 24415 33756
rect 24471 33754 24495 33756
rect 24551 33754 24575 33756
rect 24631 33754 24655 33756
rect 24711 33754 24717 33756
rect 24471 33702 24473 33754
rect 24653 33702 24655 33754
rect 24409 33700 24415 33702
rect 24471 33700 24495 33702
rect 24551 33700 24575 33702
rect 24631 33700 24655 33702
rect 24711 33700 24717 33702
rect 24409 33691 24717 33700
rect 24409 32668 24717 32677
rect 24409 32666 24415 32668
rect 24471 32666 24495 32668
rect 24551 32666 24575 32668
rect 24631 32666 24655 32668
rect 24711 32666 24717 32668
rect 24471 32614 24473 32666
rect 24653 32614 24655 32666
rect 24409 32612 24415 32614
rect 24471 32612 24495 32614
rect 24551 32612 24575 32614
rect 24631 32612 24655 32614
rect 24711 32612 24717 32614
rect 24409 32603 24717 32612
rect 24409 31580 24717 31589
rect 24409 31578 24415 31580
rect 24471 31578 24495 31580
rect 24551 31578 24575 31580
rect 24631 31578 24655 31580
rect 24711 31578 24717 31580
rect 24471 31526 24473 31578
rect 24653 31526 24655 31578
rect 24409 31524 24415 31526
rect 24471 31524 24495 31526
rect 24551 31524 24575 31526
rect 24631 31524 24655 31526
rect 24711 31524 24717 31526
rect 24409 31515 24717 31524
rect 24409 30492 24717 30501
rect 24409 30490 24415 30492
rect 24471 30490 24495 30492
rect 24551 30490 24575 30492
rect 24631 30490 24655 30492
rect 24711 30490 24717 30492
rect 24471 30438 24473 30490
rect 24653 30438 24655 30490
rect 24409 30436 24415 30438
rect 24471 30436 24495 30438
rect 24551 30436 24575 30438
rect 24631 30436 24655 30438
rect 24711 30436 24717 30438
rect 24409 30427 24717 30436
rect 24409 29404 24717 29413
rect 24409 29402 24415 29404
rect 24471 29402 24495 29404
rect 24551 29402 24575 29404
rect 24631 29402 24655 29404
rect 24711 29402 24717 29404
rect 24471 29350 24473 29402
rect 24653 29350 24655 29402
rect 24409 29348 24415 29350
rect 24471 29348 24495 29350
rect 24551 29348 24575 29350
rect 24631 29348 24655 29350
rect 24711 29348 24717 29350
rect 24409 29339 24717 29348
rect 24409 28316 24717 28325
rect 24409 28314 24415 28316
rect 24471 28314 24495 28316
rect 24551 28314 24575 28316
rect 24631 28314 24655 28316
rect 24711 28314 24717 28316
rect 24471 28262 24473 28314
rect 24653 28262 24655 28314
rect 24409 28260 24415 28262
rect 24471 28260 24495 28262
rect 24551 28260 24575 28262
rect 24631 28260 24655 28262
rect 24711 28260 24717 28262
rect 24409 28251 24717 28260
rect 24409 27228 24717 27237
rect 24409 27226 24415 27228
rect 24471 27226 24495 27228
rect 24551 27226 24575 27228
rect 24631 27226 24655 27228
rect 24711 27226 24717 27228
rect 24471 27174 24473 27226
rect 24653 27174 24655 27226
rect 24409 27172 24415 27174
rect 24471 27172 24495 27174
rect 24551 27172 24575 27174
rect 24631 27172 24655 27174
rect 24711 27172 24717 27174
rect 24409 27163 24717 27172
rect 24409 26140 24717 26149
rect 24409 26138 24415 26140
rect 24471 26138 24495 26140
rect 24551 26138 24575 26140
rect 24631 26138 24655 26140
rect 24711 26138 24717 26140
rect 24471 26086 24473 26138
rect 24653 26086 24655 26138
rect 24409 26084 24415 26086
rect 24471 26084 24495 26086
rect 24551 26084 24575 26086
rect 24631 26084 24655 26086
rect 24711 26084 24717 26086
rect 24409 26075 24717 26084
rect 24409 25052 24717 25061
rect 24409 25050 24415 25052
rect 24471 25050 24495 25052
rect 24551 25050 24575 25052
rect 24631 25050 24655 25052
rect 24711 25050 24717 25052
rect 24471 24998 24473 25050
rect 24653 24998 24655 25050
rect 24409 24996 24415 24998
rect 24471 24996 24495 24998
rect 24551 24996 24575 24998
rect 24631 24996 24655 24998
rect 24711 24996 24717 24998
rect 24409 24987 24717 24996
rect 24409 23964 24717 23973
rect 24409 23962 24415 23964
rect 24471 23962 24495 23964
rect 24551 23962 24575 23964
rect 24631 23962 24655 23964
rect 24711 23962 24717 23964
rect 24471 23910 24473 23962
rect 24653 23910 24655 23962
rect 24409 23908 24415 23910
rect 24471 23908 24495 23910
rect 24551 23908 24575 23910
rect 24631 23908 24655 23910
rect 24711 23908 24717 23910
rect 24409 23899 24717 23908
rect 24409 22876 24717 22885
rect 24409 22874 24415 22876
rect 24471 22874 24495 22876
rect 24551 22874 24575 22876
rect 24631 22874 24655 22876
rect 24711 22874 24717 22876
rect 24471 22822 24473 22874
rect 24653 22822 24655 22874
rect 24409 22820 24415 22822
rect 24471 22820 24495 22822
rect 24551 22820 24575 22822
rect 24631 22820 24655 22822
rect 24711 22820 24717 22822
rect 24409 22811 24717 22820
rect 24409 21788 24717 21797
rect 24409 21786 24415 21788
rect 24471 21786 24495 21788
rect 24551 21786 24575 21788
rect 24631 21786 24655 21788
rect 24711 21786 24717 21788
rect 24471 21734 24473 21786
rect 24653 21734 24655 21786
rect 24409 21732 24415 21734
rect 24471 21732 24495 21734
rect 24551 21732 24575 21734
rect 24631 21732 24655 21734
rect 24711 21732 24717 21734
rect 24409 21723 24717 21732
rect 24409 20700 24717 20709
rect 24409 20698 24415 20700
rect 24471 20698 24495 20700
rect 24551 20698 24575 20700
rect 24631 20698 24655 20700
rect 24711 20698 24717 20700
rect 24471 20646 24473 20698
rect 24653 20646 24655 20698
rect 24409 20644 24415 20646
rect 24471 20644 24495 20646
rect 24551 20644 24575 20646
rect 24631 20644 24655 20646
rect 24711 20644 24717 20646
rect 24409 20635 24717 20644
rect 24409 19612 24717 19621
rect 24409 19610 24415 19612
rect 24471 19610 24495 19612
rect 24551 19610 24575 19612
rect 24631 19610 24655 19612
rect 24711 19610 24717 19612
rect 24471 19558 24473 19610
rect 24653 19558 24655 19610
rect 24409 19556 24415 19558
rect 24471 19556 24495 19558
rect 24551 19556 24575 19558
rect 24631 19556 24655 19558
rect 24711 19556 24717 19558
rect 24409 19547 24717 19556
rect 24409 18524 24717 18533
rect 24409 18522 24415 18524
rect 24471 18522 24495 18524
rect 24551 18522 24575 18524
rect 24631 18522 24655 18524
rect 24711 18522 24717 18524
rect 24471 18470 24473 18522
rect 24653 18470 24655 18522
rect 24409 18468 24415 18470
rect 24471 18468 24495 18470
rect 24551 18468 24575 18470
rect 24631 18468 24655 18470
rect 24711 18468 24717 18470
rect 24409 18459 24717 18468
rect 24409 17436 24717 17445
rect 24409 17434 24415 17436
rect 24471 17434 24495 17436
rect 24551 17434 24575 17436
rect 24631 17434 24655 17436
rect 24711 17434 24717 17436
rect 24471 17382 24473 17434
rect 24653 17382 24655 17434
rect 24409 17380 24415 17382
rect 24471 17380 24495 17382
rect 24551 17380 24575 17382
rect 24631 17380 24655 17382
rect 24711 17380 24717 17382
rect 24409 17371 24717 17380
rect 24409 16348 24717 16357
rect 24409 16346 24415 16348
rect 24471 16346 24495 16348
rect 24551 16346 24575 16348
rect 24631 16346 24655 16348
rect 24711 16346 24717 16348
rect 24471 16294 24473 16346
rect 24653 16294 24655 16346
rect 24409 16292 24415 16294
rect 24471 16292 24495 16294
rect 24551 16292 24575 16294
rect 24631 16292 24655 16294
rect 24711 16292 24717 16294
rect 24409 16283 24717 16292
rect 24409 15260 24717 15269
rect 24409 15258 24415 15260
rect 24471 15258 24495 15260
rect 24551 15258 24575 15260
rect 24631 15258 24655 15260
rect 24711 15258 24717 15260
rect 24471 15206 24473 15258
rect 24653 15206 24655 15258
rect 24409 15204 24415 15206
rect 24471 15204 24495 15206
rect 24551 15204 24575 15206
rect 24631 15204 24655 15206
rect 24711 15204 24717 15206
rect 24409 15195 24717 15204
rect 24409 14172 24717 14181
rect 24409 14170 24415 14172
rect 24471 14170 24495 14172
rect 24551 14170 24575 14172
rect 24631 14170 24655 14172
rect 24711 14170 24717 14172
rect 24471 14118 24473 14170
rect 24653 14118 24655 14170
rect 24409 14116 24415 14118
rect 24471 14116 24495 14118
rect 24551 14116 24575 14118
rect 24631 14116 24655 14118
rect 24711 14116 24717 14118
rect 24409 14107 24717 14116
rect 24409 13084 24717 13093
rect 24409 13082 24415 13084
rect 24471 13082 24495 13084
rect 24551 13082 24575 13084
rect 24631 13082 24655 13084
rect 24711 13082 24717 13084
rect 24471 13030 24473 13082
rect 24653 13030 24655 13082
rect 24409 13028 24415 13030
rect 24471 13028 24495 13030
rect 24551 13028 24575 13030
rect 24631 13028 24655 13030
rect 24711 13028 24717 13030
rect 24409 13019 24717 13028
rect 24228 12406 24348 12434
rect 24032 12164 24084 12170
rect 24032 12106 24084 12112
rect 23848 11552 23900 11558
rect 24044 11529 24072 12106
rect 23848 11494 23900 11500
rect 24030 11520 24086 11529
rect 23860 10810 23888 11494
rect 24030 11455 24086 11464
rect 23848 10804 23900 10810
rect 23848 10746 23900 10752
rect 23492 10526 23612 10554
rect 23032 9030 23152 9058
rect 23020 8968 23072 8974
rect 23020 8910 23072 8916
rect 23032 8090 23060 8910
rect 23020 8084 23072 8090
rect 23020 8026 23072 8032
rect 23124 7698 23152 9030
rect 23388 8832 23440 8838
rect 23386 8800 23388 8809
rect 23440 8800 23442 8809
rect 23386 8735 23442 8744
rect 23204 8560 23256 8566
rect 23204 8502 23256 8508
rect 23216 7886 23244 8502
rect 23492 7970 23520 10526
rect 24032 10464 24084 10470
rect 24032 10406 24084 10412
rect 24044 10062 24072 10406
rect 24032 10056 24084 10062
rect 24032 9998 24084 10004
rect 23940 9716 23992 9722
rect 23940 9658 23992 9664
rect 23848 9376 23900 9382
rect 23848 9318 23900 9324
rect 23860 9178 23888 9318
rect 23848 9172 23900 9178
rect 23848 9114 23900 9120
rect 23572 8968 23624 8974
rect 23570 8936 23572 8945
rect 23624 8936 23626 8945
rect 23570 8871 23626 8880
rect 23756 8628 23808 8634
rect 23756 8570 23808 8576
rect 23768 8090 23796 8570
rect 23756 8084 23808 8090
rect 23756 8026 23808 8032
rect 23952 7970 23980 9658
rect 24122 9344 24178 9353
rect 24122 9279 24178 9288
rect 24136 9178 24164 9279
rect 24124 9172 24176 9178
rect 24124 9114 24176 9120
rect 24228 8650 24256 12406
rect 24409 11996 24717 12005
rect 24409 11994 24415 11996
rect 24471 11994 24495 11996
rect 24551 11994 24575 11996
rect 24631 11994 24655 11996
rect 24711 11994 24717 11996
rect 24471 11942 24473 11994
rect 24653 11942 24655 11994
rect 24409 11940 24415 11942
rect 24471 11940 24495 11942
rect 24551 11940 24575 11942
rect 24631 11940 24655 11942
rect 24711 11940 24717 11942
rect 24409 11931 24717 11940
rect 24308 11824 24360 11830
rect 24308 11766 24360 11772
rect 24136 8622 24256 8650
rect 24136 8106 24164 8622
rect 24216 8492 24268 8498
rect 24216 8434 24268 8440
rect 24228 8265 24256 8434
rect 24214 8256 24270 8265
rect 24214 8191 24270 8200
rect 24136 8078 24256 8106
rect 23492 7942 23796 7970
rect 23952 7942 24164 7970
rect 23204 7880 23256 7886
rect 23204 7822 23256 7828
rect 23388 7880 23440 7886
rect 23388 7822 23440 7828
rect 23124 7670 23244 7698
rect 23020 7404 23072 7410
rect 23020 7346 23072 7352
rect 23032 7002 23060 7346
rect 23020 6996 23072 7002
rect 23020 6938 23072 6944
rect 23112 6792 23164 6798
rect 23112 6734 23164 6740
rect 23124 6458 23152 6734
rect 23020 6452 23072 6458
rect 23020 6394 23072 6400
rect 23112 6452 23164 6458
rect 23112 6394 23164 6400
rect 23032 5386 23060 6394
rect 23112 6112 23164 6118
rect 23112 6054 23164 6060
rect 23124 5545 23152 6054
rect 23110 5536 23166 5545
rect 23110 5471 23166 5480
rect 23032 5358 23152 5386
rect 23020 5228 23072 5234
rect 23020 5170 23072 5176
rect 22928 4140 22980 4146
rect 22928 4082 22980 4088
rect 22928 4004 22980 4010
rect 22928 3946 22980 3952
rect 22756 2264 22876 2292
rect 22468 808 22520 814
rect 22468 750 22520 756
rect 22374 640 22430 649
rect 22374 575 22430 584
rect 22480 160 22508 750
rect 22756 160 22784 2264
rect 22940 746 22968 3946
rect 23032 2854 23060 5170
rect 23124 3942 23152 5358
rect 23112 3936 23164 3942
rect 23112 3878 23164 3884
rect 23124 3602 23152 3878
rect 23112 3596 23164 3602
rect 23112 3538 23164 3544
rect 23112 3460 23164 3466
rect 23216 3448 23244 7670
rect 23296 7404 23348 7410
rect 23296 7346 23348 7352
rect 23308 5642 23336 7346
rect 23296 5636 23348 5642
rect 23296 5578 23348 5584
rect 23400 5545 23428 7822
rect 23664 7744 23716 7750
rect 23664 7686 23716 7692
rect 23572 7200 23624 7206
rect 23572 7142 23624 7148
rect 23480 6792 23532 6798
rect 23480 6734 23532 6740
rect 23492 6458 23520 6734
rect 23480 6452 23532 6458
rect 23480 6394 23532 6400
rect 23584 6322 23612 7142
rect 23676 6458 23704 7686
rect 23664 6452 23716 6458
rect 23664 6394 23716 6400
rect 23572 6316 23624 6322
rect 23572 6258 23624 6264
rect 23664 5636 23716 5642
rect 23664 5578 23716 5584
rect 23480 5568 23532 5574
rect 23386 5536 23442 5545
rect 23480 5510 23532 5516
rect 23386 5471 23442 5480
rect 23388 5024 23440 5030
rect 23388 4966 23440 4972
rect 23296 4140 23348 4146
rect 23296 4082 23348 4088
rect 23164 3420 23244 3448
rect 23112 3402 23164 3408
rect 23112 3188 23164 3194
rect 23112 3130 23164 3136
rect 23020 2848 23072 2854
rect 23020 2790 23072 2796
rect 23020 2508 23072 2514
rect 23020 2450 23072 2456
rect 22928 740 22980 746
rect 22928 682 22980 688
rect 23032 160 23060 2450
rect 23124 1562 23152 3130
rect 23112 1556 23164 1562
rect 23112 1498 23164 1504
rect 23308 160 23336 4082
rect 23400 2514 23428 4966
rect 23492 3534 23520 5510
rect 23572 4276 23624 4282
rect 23572 4218 23624 4224
rect 23480 3528 23532 3534
rect 23480 3470 23532 3476
rect 23480 2848 23532 2854
rect 23480 2790 23532 2796
rect 23388 2508 23440 2514
rect 23388 2450 23440 2456
rect 23492 1494 23520 2790
rect 23480 1488 23532 1494
rect 23480 1430 23532 1436
rect 23584 160 23612 4218
rect 23676 4010 23704 5578
rect 23768 4146 23796 7942
rect 23940 7880 23992 7886
rect 24032 7880 24084 7886
rect 23940 7822 23992 7828
rect 24030 7848 24032 7857
rect 24084 7848 24086 7857
rect 23848 7404 23900 7410
rect 23848 7346 23900 7352
rect 23860 6905 23888 7346
rect 23846 6896 23902 6905
rect 23846 6831 23902 6840
rect 23848 6792 23900 6798
rect 23848 6734 23900 6740
rect 23860 6458 23888 6734
rect 23848 6452 23900 6458
rect 23848 6394 23900 6400
rect 23952 5914 23980 7822
rect 24030 7783 24086 7792
rect 24030 7576 24086 7585
rect 24030 7511 24032 7520
rect 24084 7511 24086 7520
rect 24032 7482 24084 7488
rect 24032 7404 24084 7410
rect 24032 7346 24084 7352
rect 24044 7177 24072 7346
rect 24030 7168 24086 7177
rect 24030 7103 24086 7112
rect 24032 6316 24084 6322
rect 24032 6258 24084 6264
rect 23940 5908 23992 5914
rect 23940 5850 23992 5856
rect 23846 5672 23902 5681
rect 23846 5607 23902 5616
rect 23756 4140 23808 4146
rect 23756 4082 23808 4088
rect 23664 4004 23716 4010
rect 23664 3946 23716 3952
rect 23860 3670 23888 5607
rect 24044 5001 24072 6258
rect 24136 5302 24164 7942
rect 24228 5760 24256 8078
rect 24320 6458 24348 11766
rect 24409 10908 24717 10917
rect 24409 10906 24415 10908
rect 24471 10906 24495 10908
rect 24551 10906 24575 10908
rect 24631 10906 24655 10908
rect 24711 10906 24717 10908
rect 24471 10854 24473 10906
rect 24653 10854 24655 10906
rect 24409 10852 24415 10854
rect 24471 10852 24495 10854
rect 24551 10852 24575 10854
rect 24631 10852 24655 10854
rect 24711 10852 24717 10854
rect 24409 10843 24717 10852
rect 24409 9820 24717 9829
rect 24409 9818 24415 9820
rect 24471 9818 24495 9820
rect 24551 9818 24575 9820
rect 24631 9818 24655 9820
rect 24711 9818 24717 9820
rect 24471 9766 24473 9818
rect 24653 9766 24655 9818
rect 24409 9764 24415 9766
rect 24471 9764 24495 9766
rect 24551 9764 24575 9766
rect 24631 9764 24655 9766
rect 24711 9764 24717 9766
rect 24409 9755 24717 9764
rect 24409 8732 24717 8741
rect 24409 8730 24415 8732
rect 24471 8730 24495 8732
rect 24551 8730 24575 8732
rect 24631 8730 24655 8732
rect 24711 8730 24717 8732
rect 24471 8678 24473 8730
rect 24653 8678 24655 8730
rect 24409 8676 24415 8678
rect 24471 8676 24495 8678
rect 24551 8676 24575 8678
rect 24631 8676 24655 8678
rect 24711 8676 24717 8678
rect 24409 8667 24717 8676
rect 24409 7644 24717 7653
rect 24409 7642 24415 7644
rect 24471 7642 24495 7644
rect 24551 7642 24575 7644
rect 24631 7642 24655 7644
rect 24711 7642 24717 7644
rect 24471 7590 24473 7642
rect 24653 7590 24655 7642
rect 24409 7588 24415 7590
rect 24471 7588 24495 7590
rect 24551 7588 24575 7590
rect 24631 7588 24655 7590
rect 24711 7588 24717 7590
rect 24409 7579 24717 7588
rect 24409 6556 24717 6565
rect 24409 6554 24415 6556
rect 24471 6554 24495 6556
rect 24551 6554 24575 6556
rect 24631 6554 24655 6556
rect 24711 6554 24717 6556
rect 24471 6502 24473 6554
rect 24653 6502 24655 6554
rect 24409 6500 24415 6502
rect 24471 6500 24495 6502
rect 24551 6500 24575 6502
rect 24631 6500 24655 6502
rect 24711 6500 24717 6502
rect 24409 6491 24717 6500
rect 24308 6452 24360 6458
rect 24308 6394 24360 6400
rect 24228 5732 24348 5760
rect 24124 5296 24176 5302
rect 24124 5238 24176 5244
rect 24030 4992 24086 5001
rect 24030 4927 24086 4936
rect 24320 4593 24348 5732
rect 24409 5468 24717 5477
rect 24409 5466 24415 5468
rect 24471 5466 24495 5468
rect 24551 5466 24575 5468
rect 24631 5466 24655 5468
rect 24711 5466 24717 5468
rect 24471 5414 24473 5466
rect 24653 5414 24655 5466
rect 24409 5412 24415 5414
rect 24471 5412 24495 5414
rect 24551 5412 24575 5414
rect 24631 5412 24655 5414
rect 24711 5412 24717 5414
rect 24409 5403 24717 5412
rect 24306 4584 24362 4593
rect 24306 4519 24362 4528
rect 24409 4380 24717 4389
rect 24409 4378 24415 4380
rect 24471 4378 24495 4380
rect 24551 4378 24575 4380
rect 24631 4378 24655 4380
rect 24711 4378 24717 4380
rect 24471 4326 24473 4378
rect 24653 4326 24655 4378
rect 24409 4324 24415 4326
rect 24471 4324 24495 4326
rect 24551 4324 24575 4326
rect 24631 4324 24655 4326
rect 24711 4324 24717 4326
rect 24409 4315 24717 4324
rect 24032 4208 24084 4214
rect 24032 4150 24084 4156
rect 23940 3936 23992 3942
rect 23940 3878 23992 3884
rect 23664 3664 23716 3670
rect 23664 3606 23716 3612
rect 23848 3664 23900 3670
rect 23848 3606 23900 3612
rect 23676 2106 23704 3606
rect 23848 3460 23900 3466
rect 23848 3402 23900 3408
rect 23754 3088 23810 3097
rect 23754 3023 23810 3032
rect 23664 2100 23716 2106
rect 23664 2042 23716 2048
rect 23768 1970 23796 3023
rect 23756 1964 23808 1970
rect 23756 1906 23808 1912
rect 23860 678 23888 3402
rect 23952 2990 23980 3878
rect 23940 2984 23992 2990
rect 23940 2926 23992 2932
rect 23848 672 23900 678
rect 23848 614 23900 620
rect 21638 54 21864 82
rect 21086 -300 21142 54
rect 21362 -300 21418 54
rect 21638 -300 21694 54
rect 21914 -300 21970 160
rect 22190 -300 22246 160
rect 22466 -300 22522 160
rect 22742 -300 22798 160
rect 23018 -300 23074 160
rect 23294 -300 23350 160
rect 23570 -300 23626 160
rect 23846 82 23902 160
rect 24044 82 24072 4150
rect 24409 3292 24717 3301
rect 24409 3290 24415 3292
rect 24471 3290 24495 3292
rect 24551 3290 24575 3292
rect 24631 3290 24655 3292
rect 24711 3290 24717 3292
rect 24471 3238 24473 3290
rect 24653 3238 24655 3290
rect 24409 3236 24415 3238
rect 24471 3236 24495 3238
rect 24551 3236 24575 3238
rect 24631 3236 24655 3238
rect 24711 3236 24717 3238
rect 24409 3227 24717 3236
rect 24780 3176 24808 36502
rect 24952 36100 25004 36106
rect 24952 36042 25004 36048
rect 24964 36009 24992 36042
rect 24950 36000 25006 36009
rect 24950 35935 25006 35944
rect 25148 35850 25176 41618
rect 25240 40730 25268 44540
rect 25516 43450 25544 44540
rect 25504 43444 25556 43450
rect 25504 43386 25556 43392
rect 25228 40724 25280 40730
rect 25228 40666 25280 40672
rect 25504 40112 25556 40118
rect 25504 40054 25556 40060
rect 25228 39500 25280 39506
rect 25228 39442 25280 39448
rect 25240 36802 25268 39442
rect 25240 36774 25360 36802
rect 25228 36644 25280 36650
rect 25228 36586 25280 36592
rect 24964 35822 25176 35850
rect 24860 34944 24912 34950
rect 24858 34912 24860 34921
rect 24912 34912 24914 34921
rect 24858 34847 24914 34856
rect 24860 33856 24912 33862
rect 24858 33824 24860 33833
rect 24912 33824 24914 33833
rect 24858 33759 24914 33768
rect 24860 32768 24912 32774
rect 24858 32736 24860 32745
rect 24912 32736 24914 32745
rect 24858 32671 24914 32680
rect 24860 30660 24912 30666
rect 24860 30602 24912 30608
rect 24872 30569 24900 30602
rect 24858 30560 24914 30569
rect 24858 30495 24914 30504
rect 24860 29504 24912 29510
rect 24858 29472 24860 29481
rect 24912 29472 24914 29481
rect 24858 29407 24914 29416
rect 24860 28416 24912 28422
rect 24858 28384 24860 28393
rect 24912 28384 24914 28393
rect 24858 28319 24914 28328
rect 24860 27328 24912 27334
rect 24858 27296 24860 27305
rect 24912 27296 24914 27305
rect 24858 27231 24914 27240
rect 24860 26308 24912 26314
rect 24860 26250 24912 26256
rect 24872 26217 24900 26250
rect 24858 26208 24914 26217
rect 24858 26143 24914 26152
rect 24860 25696 24912 25702
rect 24860 25638 24912 25644
rect 24872 25129 24900 25638
rect 24858 25120 24914 25129
rect 24858 25055 24914 25064
rect 24860 24064 24912 24070
rect 24858 24032 24860 24041
rect 24912 24032 24914 24041
rect 24858 23967 24914 23976
rect 24858 22944 24914 22953
rect 24858 22879 24914 22888
rect 24872 22438 24900 22879
rect 24860 22432 24912 22438
rect 24860 22374 24912 22380
rect 24860 22296 24912 22302
rect 24860 22238 24912 22244
rect 24872 22030 24900 22238
rect 24860 22024 24912 22030
rect 24860 21966 24912 21972
rect 24860 21888 24912 21894
rect 24858 21856 24860 21865
rect 24912 21856 24914 21865
rect 24858 21791 24914 21800
rect 24860 20868 24912 20874
rect 24860 20810 24912 20816
rect 24872 20777 24900 20810
rect 24858 20768 24914 20777
rect 24858 20703 24914 20712
rect 24858 18592 24914 18601
rect 24858 18527 24914 18536
rect 24872 18086 24900 18527
rect 24860 18080 24912 18086
rect 24860 18022 24912 18028
rect 24860 17808 24912 17814
rect 24860 17750 24912 17756
rect 24872 17513 24900 17750
rect 24858 17504 24914 17513
rect 24858 17439 24914 17448
rect 24858 16416 24914 16425
rect 24858 16351 24914 16360
rect 24872 16250 24900 16351
rect 24860 16244 24912 16250
rect 24860 16186 24912 16192
rect 24860 15428 24912 15434
rect 24860 15370 24912 15376
rect 24872 15337 24900 15370
rect 24858 15328 24914 15337
rect 24858 15263 24914 15272
rect 24860 14272 24912 14278
rect 24858 14240 24860 14249
rect 24912 14240 24914 14249
rect 24858 14175 24914 14184
rect 24858 13152 24914 13161
rect 24858 13087 24914 13096
rect 24872 12986 24900 13087
rect 24860 12980 24912 12986
rect 24860 12922 24912 12928
rect 24860 12368 24912 12374
rect 24860 12310 24912 12316
rect 24872 12073 24900 12310
rect 24858 12064 24914 12073
rect 24858 11999 24914 12008
rect 24858 10976 24914 10985
rect 24858 10911 24914 10920
rect 24872 10266 24900 10911
rect 24860 10260 24912 10266
rect 24860 10202 24912 10208
rect 24860 9988 24912 9994
rect 24860 9930 24912 9936
rect 24872 9897 24900 9930
rect 24858 9888 24914 9897
rect 24858 9823 24914 9832
rect 24860 7336 24912 7342
rect 24860 7278 24912 7284
rect 24872 6633 24900 7278
rect 24858 6624 24914 6633
rect 24858 6559 24914 6568
rect 24964 4146 24992 35822
rect 25240 35714 25268 36586
rect 25148 35686 25268 35714
rect 25044 31816 25096 31822
rect 25044 31758 25096 31764
rect 25056 31657 25084 31758
rect 25042 31648 25098 31657
rect 25042 31583 25098 31592
rect 25148 27130 25176 35686
rect 25332 35578 25360 36774
rect 25240 35550 25360 35578
rect 25136 27124 25188 27130
rect 25136 27066 25188 27072
rect 25240 27010 25268 35550
rect 25516 35306 25544 40054
rect 25596 37256 25648 37262
rect 25596 37198 25648 37204
rect 25056 26982 25268 27010
rect 25332 35278 25544 35306
rect 25056 7410 25084 26982
rect 25136 26920 25188 26926
rect 25136 26862 25188 26868
rect 25148 22302 25176 26862
rect 25228 26784 25280 26790
rect 25228 26726 25280 26732
rect 25136 22296 25188 22302
rect 25136 22238 25188 22244
rect 25136 22024 25188 22030
rect 25136 21966 25188 21972
rect 25148 20942 25176 21966
rect 25136 20936 25188 20942
rect 25136 20878 25188 20884
rect 25134 19680 25190 19689
rect 25134 19615 25190 19624
rect 25148 18426 25176 19615
rect 25136 18420 25188 18426
rect 25136 18362 25188 18368
rect 25134 10432 25190 10441
rect 25134 10367 25190 10376
rect 25148 10062 25176 10367
rect 25136 10056 25188 10062
rect 25136 9998 25188 10004
rect 25044 7404 25096 7410
rect 25044 7346 25096 7352
rect 25136 7200 25188 7206
rect 25136 7142 25188 7148
rect 24952 4140 25004 4146
rect 24952 4082 25004 4088
rect 24952 3188 25004 3194
rect 24780 3148 24952 3176
rect 24952 3130 25004 3136
rect 24860 2984 24912 2990
rect 24860 2926 24912 2932
rect 24124 2372 24176 2378
rect 24124 2314 24176 2320
rect 24136 160 24164 2314
rect 24409 2204 24717 2213
rect 24409 2202 24415 2204
rect 24471 2202 24495 2204
rect 24551 2202 24575 2204
rect 24631 2202 24655 2204
rect 24711 2202 24717 2204
rect 24471 2150 24473 2202
rect 24653 2150 24655 2202
rect 24409 2148 24415 2150
rect 24471 2148 24495 2150
rect 24551 2148 24575 2150
rect 24631 2148 24655 2150
rect 24711 2148 24717 2150
rect 24409 2139 24717 2148
rect 24676 1760 24728 1766
rect 24728 1720 24808 1748
rect 24676 1702 24728 1708
rect 24308 1284 24360 1290
rect 24308 1226 24360 1232
rect 24320 626 24348 1226
rect 24409 1116 24717 1125
rect 24409 1114 24415 1116
rect 24471 1114 24495 1116
rect 24551 1114 24575 1116
rect 24631 1114 24655 1116
rect 24711 1114 24717 1116
rect 24471 1062 24473 1114
rect 24653 1062 24655 1114
rect 24409 1060 24415 1062
rect 24471 1060 24495 1062
rect 24551 1060 24575 1062
rect 24631 1060 24655 1062
rect 24711 1060 24717 1062
rect 24409 1051 24717 1060
rect 24320 598 24440 626
rect 24412 160 24440 598
rect 23846 54 24072 82
rect 23846 -300 23902 54
rect 24122 -300 24178 160
rect 24398 -300 24454 160
rect 24674 82 24730 160
rect 24780 82 24808 1720
rect 24674 54 24808 82
rect 24872 82 24900 2926
rect 25148 1562 25176 7142
rect 25240 3466 25268 26726
rect 25228 3460 25280 3466
rect 25228 3402 25280 3408
rect 25228 2984 25280 2990
rect 25228 2926 25280 2932
rect 25136 1556 25188 1562
rect 25136 1498 25188 1504
rect 25240 160 25268 2926
rect 25332 2650 25360 35278
rect 25608 34490 25636 37198
rect 25424 34462 25636 34490
rect 25424 12434 25452 34462
rect 25596 33108 25648 33114
rect 25596 33050 25648 33056
rect 25504 30592 25556 30598
rect 25504 30534 25556 30540
rect 25516 22098 25544 30534
rect 25504 22092 25556 22098
rect 25504 22034 25556 22040
rect 25608 22030 25636 33050
rect 25596 22024 25648 22030
rect 25596 21966 25648 21972
rect 25596 21888 25648 21894
rect 25596 21830 25648 21836
rect 25424 12406 25544 12434
rect 25412 7744 25464 7750
rect 25412 7686 25464 7692
rect 25320 2644 25372 2650
rect 25320 2586 25372 2592
rect 25424 2174 25452 7686
rect 25516 4826 25544 12406
rect 25608 7954 25636 21830
rect 25596 7948 25648 7954
rect 25596 7890 25648 7896
rect 25504 4820 25556 4826
rect 25504 4762 25556 4768
rect 25504 4548 25556 4554
rect 25504 4490 25556 4496
rect 25412 2168 25464 2174
rect 25412 2110 25464 2116
rect 25516 160 25544 4490
rect 25596 3188 25648 3194
rect 25596 3130 25648 3136
rect 25608 542 25636 3130
rect 25596 536 25648 542
rect 25596 478 25648 484
rect 24950 82 25006 160
rect 24872 54 25006 82
rect 24674 -300 24730 54
rect 24950 -300 25006 54
rect 25226 -300 25282 160
rect 25502 -300 25558 160
<< via2 >>
rect 202 40568 258 40624
rect 1398 41384 1454 41440
rect 570 40160 626 40216
rect 386 30368 442 30424
rect 478 28736 534 28792
rect 386 11872 442 11928
rect 202 3440 258 3496
rect 754 38120 810 38176
rect 1766 43152 1822 43208
rect 1674 40468 1676 40488
rect 1676 40468 1728 40488
rect 1728 40468 1730 40488
rect 1674 40432 1730 40468
rect 1398 39344 1454 39400
rect 938 34720 994 34776
rect 754 29688 810 29744
rect 754 28056 810 28112
rect 846 27240 902 27296
rect 846 25336 902 25392
rect 754 24268 810 24304
rect 754 24248 756 24268
rect 756 24248 808 24268
rect 808 24248 810 24268
rect 846 23704 902 23760
rect 754 23432 810 23488
rect 754 22888 810 22944
rect 846 22616 902 22672
rect 938 21800 994 21856
rect 754 21528 810 21584
rect 754 20168 810 20224
rect 754 19080 810 19136
rect 662 13368 718 13424
rect 938 20476 940 20496
rect 940 20476 992 20496
rect 992 20476 994 20496
rect 938 20440 994 20476
rect 846 16940 848 16960
rect 848 16940 900 16960
rect 900 16940 902 16960
rect 846 16904 902 16940
rect 938 15136 994 15192
rect 1582 38528 1638 38584
rect 1214 37440 1270 37496
rect 1122 33496 1178 33552
rect 1398 37168 1454 37224
rect 1398 36760 1454 36816
rect 1582 37304 1638 37360
rect 2042 42220 2098 42256
rect 2042 42200 2044 42220
rect 2044 42200 2096 42220
rect 2096 42200 2098 42220
rect 2042 41384 2098 41440
rect 1950 39888 2006 39944
rect 1766 36896 1822 36952
rect 1398 34040 1454 34096
rect 1306 33768 1362 33824
rect 1306 33224 1362 33280
rect 1674 36624 1730 36680
rect 1674 33496 1730 33552
rect 1398 32544 1454 32600
rect 1398 32308 1400 32328
rect 1400 32308 1452 32328
rect 1452 32308 1454 32328
rect 1398 32272 1454 32308
rect 1306 31864 1362 31920
rect 1306 31728 1362 31784
rect 1582 32816 1638 32872
rect 1674 32136 1730 32192
rect 2686 42628 2742 42664
rect 2686 42608 2688 42628
rect 2688 42608 2740 42628
rect 2740 42608 2742 42628
rect 2502 41556 2504 41576
rect 2504 41556 2556 41576
rect 2556 41556 2558 41576
rect 2502 41520 2558 41556
rect 2318 41012 2320 41032
rect 2320 41012 2372 41032
rect 2372 41012 2374 41032
rect 2318 40976 2374 41012
rect 3330 42336 3386 42392
rect 2962 39480 3018 39536
rect 3238 40296 3294 40352
rect 3888 43002 3944 43004
rect 3968 43002 4024 43004
rect 4048 43002 4104 43004
rect 4128 43002 4184 43004
rect 3888 42950 3934 43002
rect 3934 42950 3944 43002
rect 3968 42950 3998 43002
rect 3998 42950 4010 43002
rect 4010 42950 4024 43002
rect 4048 42950 4062 43002
rect 4062 42950 4074 43002
rect 4074 42950 4104 43002
rect 4128 42950 4138 43002
rect 4138 42950 4184 43002
rect 3888 42948 3944 42950
rect 3968 42948 4024 42950
rect 4048 42948 4104 42950
rect 4128 42948 4184 42950
rect 3974 42744 4030 42800
rect 3882 42336 3938 42392
rect 4158 42336 4214 42392
rect 4434 42472 4490 42528
rect 3888 41914 3944 41916
rect 3968 41914 4024 41916
rect 4048 41914 4104 41916
rect 4128 41914 4184 41916
rect 3888 41862 3934 41914
rect 3934 41862 3944 41914
rect 3968 41862 3998 41914
rect 3998 41862 4010 41914
rect 4010 41862 4024 41914
rect 4048 41862 4062 41914
rect 4062 41862 4074 41914
rect 4074 41862 4104 41914
rect 4128 41862 4138 41914
rect 4138 41862 4184 41914
rect 3888 41860 3944 41862
rect 3968 41860 4024 41862
rect 4048 41860 4104 41862
rect 4128 41860 4184 41862
rect 3888 40826 3944 40828
rect 3968 40826 4024 40828
rect 4048 40826 4104 40828
rect 4128 40826 4184 40828
rect 3888 40774 3934 40826
rect 3934 40774 3944 40826
rect 3968 40774 3998 40826
rect 3998 40774 4010 40826
rect 4010 40774 4024 40826
rect 4048 40774 4062 40826
rect 4062 40774 4074 40826
rect 4074 40774 4104 40826
rect 4128 40774 4138 40826
rect 4138 40774 4184 40826
rect 3888 40772 3944 40774
rect 3968 40772 4024 40774
rect 4048 40772 4104 40774
rect 4128 40772 4184 40774
rect 4342 42064 4398 42120
rect 4434 41656 4490 41712
rect 4434 40840 4490 40896
rect 4802 41928 4858 41984
rect 5722 42744 5778 42800
rect 5630 42336 5686 42392
rect 3606 40024 3662 40080
rect 2778 39072 2834 39128
rect 1950 33088 2006 33144
rect 2134 35536 2190 35592
rect 2410 37984 2466 38040
rect 2778 38392 2834 38448
rect 2318 36352 2374 36408
rect 2226 33632 2282 33688
rect 2410 34992 2466 35048
rect 1306 31340 1362 31376
rect 1306 31320 1308 31340
rect 1308 31320 1360 31340
rect 1360 31320 1362 31340
rect 1490 31048 1546 31104
rect 1306 29996 1308 30016
rect 1308 29996 1360 30016
rect 1360 29996 1362 30016
rect 1306 29960 1362 29996
rect 1306 29416 1362 29472
rect 1306 29180 1308 29200
rect 1308 29180 1360 29200
rect 1360 29180 1362 29200
rect 1306 29144 1362 29180
rect 1858 29416 1914 29472
rect 1858 29280 1914 29336
rect 1398 28464 1454 28520
rect 1306 27820 1308 27840
rect 1308 27820 1360 27840
rect 1360 27820 1362 27840
rect 1306 27784 1362 27820
rect 1306 26968 1362 27024
rect 1214 26696 1270 26752
rect 1306 26424 1362 26480
rect 1306 25608 1362 25664
rect 1306 24792 1362 24848
rect 1214 24520 1270 24576
rect 1306 23976 1362 24032
rect 1306 22344 1362 22400
rect 1122 21256 1178 21312
rect 1766 27784 1822 27840
rect 1674 25200 1730 25256
rect 1674 24792 1730 24848
rect 1582 24676 1638 24712
rect 1582 24656 1584 24676
rect 1584 24656 1636 24676
rect 1636 24656 1638 24676
rect 1674 23432 1730 23488
rect 2042 30776 2098 30832
rect 2410 33088 2466 33144
rect 2962 37168 3018 37224
rect 3146 38256 3202 38312
rect 2870 36216 2926 36272
rect 3054 37032 3110 37088
rect 3054 36916 3110 36952
rect 3054 36896 3056 36916
rect 3056 36896 3108 36916
rect 3108 36896 3110 36916
rect 3146 36216 3202 36272
rect 3054 35128 3110 35184
rect 2778 34856 2834 34912
rect 3238 35672 3294 35728
rect 4802 40704 4858 40760
rect 2594 32136 2650 32192
rect 2502 31728 2558 31784
rect 2870 31220 2872 31240
rect 2872 31220 2924 31240
rect 2924 31220 2926 31240
rect 2870 31184 2926 31220
rect 2410 29552 2466 29608
rect 2410 28872 2466 28928
rect 2318 27920 2374 27976
rect 2042 26460 2044 26480
rect 2044 26460 2096 26480
rect 2096 26460 2098 26480
rect 2042 26424 2098 26460
rect 2594 29008 2650 29064
rect 2778 28600 2834 28656
rect 2686 28192 2742 28248
rect 3146 32680 3202 32736
rect 3054 30232 3110 30288
rect 3606 39208 3662 39264
rect 3888 39738 3944 39740
rect 3968 39738 4024 39740
rect 4048 39738 4104 39740
rect 4128 39738 4184 39740
rect 3888 39686 3934 39738
rect 3934 39686 3944 39738
rect 3968 39686 3998 39738
rect 3998 39686 4010 39738
rect 4010 39686 4024 39738
rect 4048 39686 4062 39738
rect 4062 39686 4074 39738
rect 4074 39686 4104 39738
rect 4128 39686 4138 39738
rect 4138 39686 4184 39738
rect 3888 39684 3944 39686
rect 3968 39684 4024 39686
rect 4048 39684 4104 39686
rect 4128 39684 4184 39686
rect 3698 38700 3700 38720
rect 3700 38700 3752 38720
rect 3752 38700 3754 38720
rect 3698 38664 3754 38700
rect 3698 38528 3754 38584
rect 3882 39072 3938 39128
rect 3974 38956 4030 38992
rect 3974 38936 3976 38956
rect 3976 38936 4028 38956
rect 4028 38936 4030 38956
rect 3888 38650 3944 38652
rect 3968 38650 4024 38652
rect 4048 38650 4104 38652
rect 4128 38650 4184 38652
rect 3888 38598 3934 38650
rect 3934 38598 3944 38650
rect 3968 38598 3998 38650
rect 3998 38598 4010 38650
rect 4010 38598 4024 38650
rect 4048 38598 4062 38650
rect 4062 38598 4074 38650
rect 4074 38598 4104 38650
rect 4128 38598 4138 38650
rect 4138 38598 4184 38650
rect 3888 38596 3944 38598
rect 3968 38596 4024 38598
rect 4048 38596 4104 38598
rect 4128 38596 4184 38598
rect 3882 38120 3938 38176
rect 3888 37562 3944 37564
rect 3968 37562 4024 37564
rect 4048 37562 4104 37564
rect 4128 37562 4184 37564
rect 3888 37510 3934 37562
rect 3934 37510 3944 37562
rect 3968 37510 3998 37562
rect 3998 37510 4010 37562
rect 4010 37510 4024 37562
rect 4048 37510 4062 37562
rect 4062 37510 4074 37562
rect 4074 37510 4104 37562
rect 4128 37510 4138 37562
rect 4138 37510 4184 37562
rect 3888 37508 3944 37510
rect 3968 37508 4024 37510
rect 4048 37508 4104 37510
rect 4128 37508 4184 37510
rect 4342 37712 4398 37768
rect 4250 37304 4306 37360
rect 3882 37168 3938 37224
rect 4158 37032 4214 37088
rect 4526 39380 4528 39400
rect 4528 39380 4580 39400
rect 4580 39380 4582 39400
rect 4526 39344 4582 39380
rect 5722 41520 5778 41576
rect 5906 43152 5962 43208
rect 5446 40432 5502 40488
rect 5354 40024 5410 40080
rect 4986 37848 5042 37904
rect 4894 37304 4950 37360
rect 3888 36474 3944 36476
rect 3968 36474 4024 36476
rect 4048 36474 4104 36476
rect 4128 36474 4184 36476
rect 3888 36422 3934 36474
rect 3934 36422 3944 36474
rect 3968 36422 3998 36474
rect 3998 36422 4010 36474
rect 4010 36422 4024 36474
rect 4048 36422 4062 36474
rect 4062 36422 4074 36474
rect 4074 36422 4104 36474
rect 4128 36422 4138 36474
rect 4138 36422 4184 36474
rect 3888 36420 3944 36422
rect 3968 36420 4024 36422
rect 4048 36420 4104 36422
rect 4128 36420 4184 36422
rect 3790 36080 3846 36136
rect 4710 36488 4766 36544
rect 4986 36488 5042 36544
rect 5262 37440 5318 37496
rect 3606 35400 3662 35456
rect 4434 35808 4490 35864
rect 3888 35386 3944 35388
rect 3968 35386 4024 35388
rect 4048 35386 4104 35388
rect 4128 35386 4184 35388
rect 3888 35334 3934 35386
rect 3934 35334 3944 35386
rect 3968 35334 3998 35386
rect 3998 35334 4010 35386
rect 4010 35334 4024 35386
rect 4048 35334 4062 35386
rect 4062 35334 4074 35386
rect 4074 35334 4104 35386
rect 4128 35334 4138 35386
rect 4138 35334 4184 35386
rect 3888 35332 3944 35334
rect 3968 35332 4024 35334
rect 4048 35332 4104 35334
rect 4128 35332 4184 35334
rect 3882 34584 3938 34640
rect 3790 34448 3846 34504
rect 4342 34992 4398 35048
rect 3888 34298 3944 34300
rect 3968 34298 4024 34300
rect 4048 34298 4104 34300
rect 4128 34298 4184 34300
rect 3888 34246 3934 34298
rect 3934 34246 3944 34298
rect 3968 34246 3998 34298
rect 3998 34246 4010 34298
rect 4010 34246 4024 34298
rect 4048 34246 4062 34298
rect 4062 34246 4074 34298
rect 4074 34246 4104 34298
rect 4128 34246 4138 34298
rect 4138 34246 4184 34298
rect 3888 34244 3944 34246
rect 3968 34244 4024 34246
rect 4048 34244 4104 34246
rect 4128 34244 4184 34246
rect 3698 34060 3754 34096
rect 3698 34040 3700 34060
rect 3700 34040 3752 34060
rect 3752 34040 3754 34060
rect 4158 33904 4214 33960
rect 4158 33804 4160 33824
rect 4160 33804 4212 33824
rect 4212 33804 4214 33824
rect 4158 33768 4214 33804
rect 3606 32952 3662 33008
rect 3974 33360 4030 33416
rect 3888 33210 3944 33212
rect 3968 33210 4024 33212
rect 4048 33210 4104 33212
rect 4128 33210 4184 33212
rect 3888 33158 3934 33210
rect 3934 33158 3944 33210
rect 3968 33158 3998 33210
rect 3998 33158 4010 33210
rect 4010 33158 4024 33210
rect 4048 33158 4062 33210
rect 4062 33158 4074 33210
rect 4074 33158 4104 33210
rect 4128 33158 4138 33210
rect 4138 33158 4184 33210
rect 3888 33156 3944 33158
rect 3968 33156 4024 33158
rect 4048 33156 4104 33158
rect 4128 33156 4184 33158
rect 3888 32122 3944 32124
rect 3968 32122 4024 32124
rect 4048 32122 4104 32124
rect 4128 32122 4184 32124
rect 3888 32070 3934 32122
rect 3934 32070 3944 32122
rect 3968 32070 3998 32122
rect 3998 32070 4010 32122
rect 4010 32070 4024 32122
rect 4048 32070 4062 32122
rect 4062 32070 4074 32122
rect 4074 32070 4104 32122
rect 4128 32070 4138 32122
rect 4138 32070 4184 32122
rect 3888 32068 3944 32070
rect 3968 32068 4024 32070
rect 4048 32068 4104 32070
rect 4128 32068 4184 32070
rect 3514 31456 3570 31512
rect 3422 30504 3478 30560
rect 3606 30776 3662 30832
rect 3514 29552 3570 29608
rect 2502 26832 2558 26888
rect 2410 26016 2466 26072
rect 2042 23024 2098 23080
rect 1306 20984 1362 21040
rect 1490 20848 1546 20904
rect 1490 20712 1546 20768
rect 1582 20440 1638 20496
rect 1950 22072 2006 22128
rect 1674 20032 1730 20088
rect 1122 19352 1178 19408
rect 1398 19896 1454 19952
rect 1306 19624 1362 19680
rect 1306 17448 1362 17504
rect 1766 18672 1822 18728
rect 1582 16088 1638 16144
rect 1122 15816 1178 15872
rect 1306 15544 1362 15600
rect 1214 15272 1270 15328
rect 1122 15000 1178 15056
rect 1490 15952 1546 16008
rect 1306 14728 1362 14784
rect 1306 13776 1362 13832
rect 1214 13096 1270 13152
rect 2134 20748 2136 20768
rect 2136 20748 2188 20768
rect 2188 20748 2190 20768
rect 2134 20712 2190 20748
rect 2042 20596 2098 20632
rect 2870 27412 2872 27432
rect 2872 27412 2924 27432
rect 2924 27412 2926 27432
rect 2870 27376 2926 27412
rect 2870 26152 2926 26208
rect 2778 25880 2834 25936
rect 2870 25200 2926 25256
rect 2502 23740 2504 23760
rect 2504 23740 2556 23760
rect 2556 23740 2558 23760
rect 2502 23704 2558 23740
rect 2778 23568 2834 23624
rect 2502 23432 2558 23488
rect 2686 23296 2742 23352
rect 2410 22072 2466 22128
rect 2042 20576 2044 20596
rect 2044 20576 2096 20596
rect 2096 20576 2098 20596
rect 2042 19760 2098 19816
rect 2870 23024 2926 23080
rect 2594 22092 2650 22128
rect 2594 22072 2596 22092
rect 2596 22072 2648 22092
rect 2648 22072 2650 22092
rect 2134 19624 2190 19680
rect 2226 19488 2282 19544
rect 2134 18400 2190 18456
rect 1766 14320 1822 14376
rect 1582 13912 1638 13968
rect 1306 12008 1362 12064
rect 1490 12180 1492 12200
rect 1492 12180 1544 12200
rect 1544 12180 1546 12200
rect 1490 12144 1546 12180
rect 1582 11464 1638 11520
rect 1490 8372 1492 8392
rect 1492 8372 1544 8392
rect 1544 8372 1546 8392
rect 1490 8336 1546 8372
rect 1766 12552 1822 12608
rect 2226 17312 2282 17368
rect 3514 29008 3570 29064
rect 3888 31034 3944 31036
rect 3968 31034 4024 31036
rect 4048 31034 4104 31036
rect 4128 31034 4184 31036
rect 3888 30982 3934 31034
rect 3934 30982 3944 31034
rect 3968 30982 3998 31034
rect 3998 30982 4010 31034
rect 4010 30982 4024 31034
rect 4048 30982 4062 31034
rect 4062 30982 4074 31034
rect 4074 30982 4104 31034
rect 4128 30982 4138 31034
rect 4138 30982 4184 31034
rect 3888 30980 3944 30982
rect 3968 30980 4024 30982
rect 4048 30980 4104 30982
rect 4128 30980 4184 30982
rect 4158 30368 4214 30424
rect 4342 33224 4398 33280
rect 4434 33088 4490 33144
rect 4802 34448 4858 34504
rect 4434 31048 4490 31104
rect 4342 30912 4398 30968
rect 4066 30096 4122 30152
rect 3888 29946 3944 29948
rect 3968 29946 4024 29948
rect 4048 29946 4104 29948
rect 4128 29946 4184 29948
rect 3888 29894 3934 29946
rect 3934 29894 3944 29946
rect 3968 29894 3998 29946
rect 3998 29894 4010 29946
rect 4010 29894 4024 29946
rect 4048 29894 4062 29946
rect 4062 29894 4074 29946
rect 4074 29894 4104 29946
rect 4128 29894 4138 29946
rect 4138 29894 4184 29946
rect 3888 29892 3944 29894
rect 3968 29892 4024 29894
rect 4048 29892 4104 29894
rect 4128 29892 4184 29894
rect 3888 28858 3944 28860
rect 3968 28858 4024 28860
rect 4048 28858 4104 28860
rect 4128 28858 4184 28860
rect 3888 28806 3934 28858
rect 3934 28806 3944 28858
rect 3968 28806 3998 28858
rect 3998 28806 4010 28858
rect 4010 28806 4024 28858
rect 4048 28806 4062 28858
rect 4062 28806 4074 28858
rect 4074 28806 4104 28858
rect 4128 28806 4138 28858
rect 4138 28806 4184 28858
rect 3888 28804 3944 28806
rect 3968 28804 4024 28806
rect 4048 28804 4104 28806
rect 4128 28804 4184 28806
rect 3698 28328 3754 28384
rect 3698 27512 3754 27568
rect 3888 27770 3944 27772
rect 3968 27770 4024 27772
rect 4048 27770 4104 27772
rect 4128 27770 4184 27772
rect 3888 27718 3934 27770
rect 3934 27718 3944 27770
rect 3968 27718 3998 27770
rect 3998 27718 4010 27770
rect 4010 27718 4024 27770
rect 4048 27718 4062 27770
rect 4062 27718 4074 27770
rect 4074 27718 4104 27770
rect 4128 27718 4138 27770
rect 4138 27718 4184 27770
rect 3888 27716 3944 27718
rect 3968 27716 4024 27718
rect 4048 27716 4104 27718
rect 4128 27716 4184 27718
rect 4066 27512 4122 27568
rect 3882 27376 3938 27432
rect 3888 26682 3944 26684
rect 3968 26682 4024 26684
rect 4048 26682 4104 26684
rect 4128 26682 4184 26684
rect 3888 26630 3934 26682
rect 3934 26630 3944 26682
rect 3968 26630 3998 26682
rect 3998 26630 4010 26682
rect 4010 26630 4024 26682
rect 4048 26630 4062 26682
rect 4062 26630 4074 26682
rect 4074 26630 4104 26682
rect 4128 26630 4138 26682
rect 4138 26630 4184 26682
rect 3888 26628 3944 26630
rect 3968 26628 4024 26630
rect 4048 26628 4104 26630
rect 4128 26628 4184 26630
rect 4158 26288 4214 26344
rect 3422 24656 3478 24712
rect 3422 24248 3478 24304
rect 3698 25608 3754 25664
rect 3888 25594 3944 25596
rect 3968 25594 4024 25596
rect 4048 25594 4104 25596
rect 4128 25594 4184 25596
rect 3888 25542 3934 25594
rect 3934 25542 3944 25594
rect 3968 25542 3998 25594
rect 3998 25542 4010 25594
rect 4010 25542 4024 25594
rect 4048 25542 4062 25594
rect 4062 25542 4074 25594
rect 4074 25542 4104 25594
rect 4128 25542 4138 25594
rect 4138 25542 4184 25594
rect 3888 25540 3944 25542
rect 3968 25540 4024 25542
rect 4048 25540 4104 25542
rect 4128 25540 4184 25542
rect 4894 34176 4950 34232
rect 4894 33768 4950 33824
rect 5354 35944 5410 36000
rect 5262 35692 5318 35728
rect 5262 35672 5264 35692
rect 5264 35672 5316 35692
rect 5316 35672 5318 35692
rect 4618 30640 4674 30696
rect 4802 31048 4858 31104
rect 4802 30776 4858 30832
rect 4802 30368 4858 30424
rect 4526 27784 4582 27840
rect 4342 26560 4398 26616
rect 4250 24928 4306 24984
rect 3888 24506 3944 24508
rect 3968 24506 4024 24508
rect 4048 24506 4104 24508
rect 4128 24506 4184 24508
rect 3888 24454 3934 24506
rect 3934 24454 3944 24506
rect 3968 24454 3998 24506
rect 3998 24454 4010 24506
rect 4010 24454 4024 24506
rect 4048 24454 4062 24506
rect 4062 24454 4074 24506
rect 4074 24454 4104 24506
rect 4128 24454 4138 24506
rect 4138 24454 4184 24506
rect 3888 24452 3944 24454
rect 3968 24452 4024 24454
rect 4048 24452 4104 24454
rect 4128 24452 4184 24454
rect 2594 19216 2650 19272
rect 2594 17448 2650 17504
rect 2318 14320 2374 14376
rect 2778 18808 2834 18864
rect 2778 18264 2834 18320
rect 2962 18264 3018 18320
rect 3054 15272 3110 15328
rect 2962 13912 3018 13968
rect 1858 9968 1914 10024
rect 2318 11600 2374 11656
rect 1950 8472 2006 8528
rect 2134 8608 2190 8664
rect 1858 7928 1914 7984
rect 1490 6724 1546 6760
rect 1490 6704 1492 6724
rect 1492 6704 1544 6724
rect 1544 6704 1546 6724
rect 1674 5480 1730 5536
rect 1766 5344 1822 5400
rect 1306 4936 1362 4992
rect 1674 4664 1730 4720
rect 1582 3984 1638 4040
rect 1674 2896 1730 2952
rect 2594 11056 2650 11112
rect 2962 11192 3018 11248
rect 2870 10784 2926 10840
rect 2778 10512 2834 10568
rect 2870 9832 2926 9888
rect 3238 20848 3294 20904
rect 3422 20440 3478 20496
rect 3514 19896 3570 19952
rect 3422 19624 3478 19680
rect 4158 24112 4214 24168
rect 3888 23418 3944 23420
rect 3968 23418 4024 23420
rect 4048 23418 4104 23420
rect 4128 23418 4184 23420
rect 3888 23366 3934 23418
rect 3934 23366 3944 23418
rect 3968 23366 3998 23418
rect 3998 23366 4010 23418
rect 4010 23366 4024 23418
rect 4048 23366 4062 23418
rect 4062 23366 4074 23418
rect 4074 23366 4104 23418
rect 4128 23366 4138 23418
rect 4138 23366 4184 23418
rect 3888 23364 3944 23366
rect 3968 23364 4024 23366
rect 4048 23364 4104 23366
rect 4128 23364 4184 23366
rect 3888 22330 3944 22332
rect 3968 22330 4024 22332
rect 4048 22330 4104 22332
rect 4128 22330 4184 22332
rect 3888 22278 3934 22330
rect 3934 22278 3944 22330
rect 3968 22278 3998 22330
rect 3998 22278 4010 22330
rect 4010 22278 4024 22330
rect 4048 22278 4062 22330
rect 4062 22278 4074 22330
rect 4074 22278 4104 22330
rect 4128 22278 4138 22330
rect 4138 22278 4184 22330
rect 3888 22276 3944 22278
rect 3968 22276 4024 22278
rect 4048 22276 4104 22278
rect 4128 22276 4184 22278
rect 3238 17720 3294 17776
rect 3422 17176 3478 17232
rect 3330 16360 3386 16416
rect 3238 15680 3294 15736
rect 3606 18028 3608 18048
rect 3608 18028 3660 18048
rect 3660 18028 3662 18048
rect 3606 17992 3662 18028
rect 3974 21528 4030 21584
rect 4158 21392 4214 21448
rect 3888 21242 3944 21244
rect 3968 21242 4024 21244
rect 4048 21242 4104 21244
rect 4128 21242 4184 21244
rect 3888 21190 3934 21242
rect 3934 21190 3944 21242
rect 3968 21190 3998 21242
rect 3998 21190 4010 21242
rect 4010 21190 4024 21242
rect 4048 21190 4062 21242
rect 4062 21190 4074 21242
rect 4074 21190 4104 21242
rect 4128 21190 4138 21242
rect 4138 21190 4184 21242
rect 3888 21188 3944 21190
rect 3968 21188 4024 21190
rect 4048 21188 4104 21190
rect 4128 21188 4184 21190
rect 4434 25744 4490 25800
rect 4434 22072 4490 22128
rect 4434 21956 4490 21992
rect 4434 21936 4436 21956
rect 4436 21936 4488 21956
rect 4488 21936 4490 21956
rect 4342 21528 4398 21584
rect 4250 20984 4306 21040
rect 3888 20154 3944 20156
rect 3968 20154 4024 20156
rect 4048 20154 4104 20156
rect 4128 20154 4184 20156
rect 3888 20102 3934 20154
rect 3934 20102 3944 20154
rect 3968 20102 3998 20154
rect 3998 20102 4010 20154
rect 4010 20102 4024 20154
rect 4048 20102 4062 20154
rect 4062 20102 4074 20154
rect 4074 20102 4104 20154
rect 4128 20102 4138 20154
rect 4138 20102 4184 20154
rect 3888 20100 3944 20102
rect 3968 20100 4024 20102
rect 4048 20100 4104 20102
rect 4128 20100 4184 20102
rect 4066 19760 4122 19816
rect 3790 19352 3846 19408
rect 4342 20576 4398 20632
rect 5630 39908 5686 39944
rect 5630 39888 5632 39908
rect 5632 39888 5684 39908
rect 5684 39888 5686 39908
rect 5814 40160 5870 40216
rect 5538 35808 5594 35864
rect 5722 36896 5778 36952
rect 5354 32408 5410 32464
rect 5354 31748 5410 31784
rect 5354 31728 5356 31748
rect 5356 31728 5408 31748
rect 5408 31728 5410 31748
rect 5354 31592 5410 31648
rect 5262 30776 5318 30832
rect 5538 31456 5594 31512
rect 5170 29280 5226 29336
rect 5170 28328 5226 28384
rect 4986 27104 5042 27160
rect 4986 26968 5042 27024
rect 4802 24656 4858 24712
rect 4710 23432 4766 23488
rect 4618 20848 4674 20904
rect 3888 19066 3944 19068
rect 3968 19066 4024 19068
rect 4048 19066 4104 19068
rect 4128 19066 4184 19068
rect 3888 19014 3934 19066
rect 3934 19014 3944 19066
rect 3968 19014 3998 19066
rect 3998 19014 4010 19066
rect 4010 19014 4024 19066
rect 4048 19014 4062 19066
rect 4062 19014 4074 19066
rect 4074 19014 4104 19066
rect 4128 19014 4138 19066
rect 4138 19014 4184 19066
rect 3888 19012 3944 19014
rect 3968 19012 4024 19014
rect 4048 19012 4104 19014
rect 4128 19012 4184 19014
rect 3790 18536 3846 18592
rect 3698 16632 3754 16688
rect 3888 17978 3944 17980
rect 3968 17978 4024 17980
rect 4048 17978 4104 17980
rect 4128 17978 4184 17980
rect 3888 17926 3934 17978
rect 3934 17926 3944 17978
rect 3968 17926 3998 17978
rect 3998 17926 4010 17978
rect 4010 17926 4024 17978
rect 4048 17926 4062 17978
rect 4062 17926 4074 17978
rect 4074 17926 4104 17978
rect 4128 17926 4138 17978
rect 4138 17926 4184 17978
rect 3888 17924 3944 17926
rect 3968 17924 4024 17926
rect 4048 17924 4104 17926
rect 4128 17924 4184 17926
rect 4066 17196 4122 17232
rect 4066 17176 4068 17196
rect 4068 17176 4120 17196
rect 4120 17176 4122 17196
rect 4526 18944 4582 19000
rect 3888 16890 3944 16892
rect 3968 16890 4024 16892
rect 4048 16890 4104 16892
rect 4128 16890 4184 16892
rect 3888 16838 3934 16890
rect 3934 16838 3944 16890
rect 3968 16838 3998 16890
rect 3998 16838 4010 16890
rect 4010 16838 4024 16890
rect 4048 16838 4062 16890
rect 4062 16838 4074 16890
rect 4074 16838 4104 16890
rect 4128 16838 4138 16890
rect 4138 16838 4184 16890
rect 3888 16836 3944 16838
rect 3968 16836 4024 16838
rect 4048 16836 4104 16838
rect 4128 16836 4184 16838
rect 4250 16496 4306 16552
rect 4158 16224 4214 16280
rect 3888 15802 3944 15804
rect 3968 15802 4024 15804
rect 4048 15802 4104 15804
rect 4128 15802 4184 15804
rect 3888 15750 3934 15802
rect 3934 15750 3944 15802
rect 3968 15750 3998 15802
rect 3998 15750 4010 15802
rect 4010 15750 4024 15802
rect 4048 15750 4062 15802
rect 4062 15750 4074 15802
rect 4074 15750 4104 15802
rect 4128 15750 4138 15802
rect 4138 15750 4184 15802
rect 3888 15748 3944 15750
rect 3968 15748 4024 15750
rect 4048 15748 4104 15750
rect 4128 15748 4184 15750
rect 3882 15544 3938 15600
rect 3606 13640 3662 13696
rect 4158 14884 4214 14920
rect 4158 14864 4160 14884
rect 4160 14864 4212 14884
rect 4212 14864 4214 14884
rect 3888 14714 3944 14716
rect 3968 14714 4024 14716
rect 4048 14714 4104 14716
rect 4128 14714 4184 14716
rect 3888 14662 3934 14714
rect 3934 14662 3944 14714
rect 3968 14662 3998 14714
rect 3998 14662 4010 14714
rect 4010 14662 4024 14714
rect 4048 14662 4062 14714
rect 4062 14662 4074 14714
rect 4074 14662 4104 14714
rect 4128 14662 4138 14714
rect 4138 14662 4184 14714
rect 3888 14660 3944 14662
rect 3968 14660 4024 14662
rect 4048 14660 4104 14662
rect 4128 14660 4184 14662
rect 3974 14456 4030 14512
rect 4158 14320 4214 14376
rect 3888 13626 3944 13628
rect 3968 13626 4024 13628
rect 4048 13626 4104 13628
rect 4128 13626 4184 13628
rect 3888 13574 3934 13626
rect 3934 13574 3944 13626
rect 3968 13574 3998 13626
rect 3998 13574 4010 13626
rect 4010 13574 4024 13626
rect 4048 13574 4062 13626
rect 4062 13574 4074 13626
rect 4074 13574 4104 13626
rect 4128 13574 4138 13626
rect 4138 13574 4184 13626
rect 3888 13572 3944 13574
rect 3968 13572 4024 13574
rect 4048 13572 4104 13574
rect 4128 13572 4184 13574
rect 3606 12824 3662 12880
rect 3422 11736 3478 11792
rect 2410 5072 2466 5128
rect 1950 3884 1952 3904
rect 1952 3884 2004 3904
rect 2004 3884 2006 3904
rect 1950 3848 2006 3884
rect 2134 1164 2136 1184
rect 2136 1164 2188 1184
rect 2188 1164 2190 1184
rect 2134 1128 2190 1164
rect 2594 6432 2650 6488
rect 2870 7792 2926 7848
rect 2870 6568 2926 6624
rect 2594 6296 2650 6352
rect 2778 5752 2834 5808
rect 2686 4256 2742 4312
rect 3054 8200 3110 8256
rect 2962 3848 3018 3904
rect 3698 12280 3754 12336
rect 5170 26152 5226 26208
rect 4618 16668 4620 16688
rect 4620 16668 4672 16688
rect 4672 16668 4674 16688
rect 4618 16632 4674 16668
rect 3888 12538 3944 12540
rect 3968 12538 4024 12540
rect 4048 12538 4104 12540
rect 4128 12538 4184 12540
rect 3888 12486 3934 12538
rect 3934 12486 3944 12538
rect 3968 12486 3998 12538
rect 3998 12486 4010 12538
rect 4010 12486 4024 12538
rect 4048 12486 4062 12538
rect 4062 12486 4074 12538
rect 4074 12486 4104 12538
rect 4128 12486 4138 12538
rect 4138 12486 4184 12538
rect 3888 12484 3944 12486
rect 3968 12484 4024 12486
rect 4048 12484 4104 12486
rect 4128 12484 4184 12486
rect 3698 10648 3754 10704
rect 3606 10376 3662 10432
rect 3888 11450 3944 11452
rect 3968 11450 4024 11452
rect 4048 11450 4104 11452
rect 4128 11450 4184 11452
rect 3888 11398 3934 11450
rect 3934 11398 3944 11450
rect 3968 11398 3998 11450
rect 3998 11398 4010 11450
rect 4010 11398 4024 11450
rect 4048 11398 4062 11450
rect 4062 11398 4074 11450
rect 4074 11398 4104 11450
rect 4128 11398 4138 11450
rect 4138 11398 4184 11450
rect 3888 11396 3944 11398
rect 3968 11396 4024 11398
rect 4048 11396 4104 11398
rect 4128 11396 4184 11398
rect 4434 12552 4490 12608
rect 3974 10956 3976 10976
rect 3976 10956 4028 10976
rect 4028 10956 4030 10976
rect 3974 10920 4030 10956
rect 4158 10920 4214 10976
rect 3888 10362 3944 10364
rect 3968 10362 4024 10364
rect 4048 10362 4104 10364
rect 4128 10362 4184 10364
rect 3888 10310 3934 10362
rect 3934 10310 3944 10362
rect 3968 10310 3998 10362
rect 3998 10310 4010 10362
rect 4010 10310 4024 10362
rect 4048 10310 4062 10362
rect 4062 10310 4074 10362
rect 4074 10310 4104 10362
rect 4128 10310 4138 10362
rect 4138 10310 4184 10362
rect 3888 10308 3944 10310
rect 3968 10308 4024 10310
rect 4048 10308 4104 10310
rect 4128 10308 4184 10310
rect 3698 9832 3754 9888
rect 3422 8880 3478 8936
rect 3238 8508 3240 8528
rect 3240 8508 3292 8528
rect 3292 8508 3294 8528
rect 3238 8472 3294 8508
rect 3146 7248 3202 7304
rect 3238 6180 3294 6216
rect 3514 8744 3570 8800
rect 4066 10104 4122 10160
rect 4066 9560 4122 9616
rect 4342 9560 4398 9616
rect 3888 9274 3944 9276
rect 3968 9274 4024 9276
rect 4048 9274 4104 9276
rect 4128 9274 4184 9276
rect 3888 9222 3934 9274
rect 3934 9222 3944 9274
rect 3968 9222 3998 9274
rect 3998 9222 4010 9274
rect 4010 9222 4024 9274
rect 4048 9222 4062 9274
rect 4062 9222 4074 9274
rect 4074 9222 4104 9274
rect 4128 9222 4138 9274
rect 4138 9222 4184 9274
rect 3888 9220 3944 9222
rect 3968 9220 4024 9222
rect 4048 9220 4104 9222
rect 4128 9220 4184 9222
rect 3606 7948 3662 7984
rect 3606 7928 3608 7948
rect 3608 7928 3660 7948
rect 3660 7928 3662 7948
rect 3514 7112 3570 7168
rect 3238 6160 3240 6180
rect 3240 6160 3292 6180
rect 3292 6160 3294 6180
rect 3422 6160 3478 6216
rect 3238 6024 3294 6080
rect 2778 856 2834 912
rect 3238 4120 3294 4176
rect 3238 4004 3294 4040
rect 3238 3984 3240 4004
rect 3240 3984 3292 4004
rect 3292 3984 3294 4004
rect 3882 8356 3938 8392
rect 3882 8336 3884 8356
rect 3884 8336 3936 8356
rect 3936 8336 3938 8356
rect 3888 8186 3944 8188
rect 3968 8186 4024 8188
rect 4048 8186 4104 8188
rect 4128 8186 4184 8188
rect 3888 8134 3934 8186
rect 3934 8134 3944 8186
rect 3968 8134 3998 8186
rect 3998 8134 4010 8186
rect 4010 8134 4024 8186
rect 4048 8134 4062 8186
rect 4062 8134 4074 8186
rect 4074 8134 4104 8186
rect 4128 8134 4138 8186
rect 4138 8134 4184 8186
rect 3888 8132 3944 8134
rect 3968 8132 4024 8134
rect 4048 8132 4104 8134
rect 4128 8132 4184 8134
rect 4066 7828 4068 7848
rect 4068 7828 4120 7848
rect 4120 7828 4122 7848
rect 4066 7792 4122 7828
rect 4066 7692 4068 7712
rect 4068 7692 4120 7712
rect 4120 7692 4122 7712
rect 4066 7656 4122 7692
rect 4066 7384 4122 7440
rect 5170 20712 5226 20768
rect 4986 14864 5042 14920
rect 6820 43546 6876 43548
rect 6900 43546 6956 43548
rect 6980 43546 7036 43548
rect 7060 43546 7116 43548
rect 6820 43494 6866 43546
rect 6866 43494 6876 43546
rect 6900 43494 6930 43546
rect 6930 43494 6942 43546
rect 6942 43494 6956 43546
rect 6980 43494 6994 43546
rect 6994 43494 7006 43546
rect 7006 43494 7036 43546
rect 7060 43494 7070 43546
rect 7070 43494 7116 43546
rect 6820 43492 6876 43494
rect 6900 43492 6956 43494
rect 6980 43492 7036 43494
rect 7060 43492 7116 43494
rect 6734 42744 6790 42800
rect 7194 42472 7250 42528
rect 6820 42458 6876 42460
rect 6900 42458 6956 42460
rect 6980 42458 7036 42460
rect 7060 42458 7116 42460
rect 6820 42406 6866 42458
rect 6866 42406 6876 42458
rect 6900 42406 6930 42458
rect 6930 42406 6942 42458
rect 6942 42406 6956 42458
rect 6980 42406 6994 42458
rect 6994 42406 7006 42458
rect 7006 42406 7036 42458
rect 7060 42406 7070 42458
rect 7070 42406 7116 42458
rect 6820 42404 6876 42406
rect 6900 42404 6956 42406
rect 6980 42404 7036 42406
rect 7060 42404 7116 42406
rect 6182 40568 6238 40624
rect 6642 41384 6698 41440
rect 6820 41370 6876 41372
rect 6900 41370 6956 41372
rect 6980 41370 7036 41372
rect 7060 41370 7116 41372
rect 6820 41318 6866 41370
rect 6866 41318 6876 41370
rect 6900 41318 6930 41370
rect 6930 41318 6942 41370
rect 6942 41318 6956 41370
rect 6980 41318 6994 41370
rect 6994 41318 7006 41370
rect 7006 41318 7036 41370
rect 7060 41318 7070 41370
rect 7070 41318 7116 41370
rect 6820 41316 6876 41318
rect 6900 41316 6956 41318
rect 6980 41316 7036 41318
rect 7060 41316 7116 41318
rect 7562 41656 7618 41712
rect 7470 40840 7526 40896
rect 6820 40282 6876 40284
rect 6900 40282 6956 40284
rect 6980 40282 7036 40284
rect 7060 40282 7116 40284
rect 6820 40230 6866 40282
rect 6866 40230 6876 40282
rect 6900 40230 6930 40282
rect 6930 40230 6942 40282
rect 6942 40230 6956 40282
rect 6980 40230 6994 40282
rect 6994 40230 7006 40282
rect 7006 40230 7036 40282
rect 7060 40230 7070 40282
rect 7070 40230 7116 40282
rect 6820 40228 6876 40230
rect 6900 40228 6956 40230
rect 6980 40228 7036 40230
rect 7060 40228 7116 40230
rect 6274 38528 6330 38584
rect 6274 37304 6330 37360
rect 6182 37168 6238 37224
rect 6090 34720 6146 34776
rect 6274 34992 6330 35048
rect 5998 33632 6054 33688
rect 5906 32952 5962 33008
rect 5998 31728 6054 31784
rect 5722 31184 5778 31240
rect 5906 31456 5962 31512
rect 5906 30096 5962 30152
rect 5998 29552 6054 29608
rect 6642 37032 6698 37088
rect 6820 39194 6876 39196
rect 6900 39194 6956 39196
rect 6980 39194 7036 39196
rect 7060 39194 7116 39196
rect 6820 39142 6866 39194
rect 6866 39142 6876 39194
rect 6900 39142 6930 39194
rect 6930 39142 6942 39194
rect 6942 39142 6956 39194
rect 6980 39142 6994 39194
rect 6994 39142 7006 39194
rect 7006 39142 7036 39194
rect 7060 39142 7070 39194
rect 7070 39142 7116 39194
rect 6820 39140 6876 39142
rect 6900 39140 6956 39142
rect 6980 39140 7036 39142
rect 7060 39140 7116 39142
rect 6820 38106 6876 38108
rect 6900 38106 6956 38108
rect 6980 38106 7036 38108
rect 7060 38106 7116 38108
rect 6820 38054 6866 38106
rect 6866 38054 6876 38106
rect 6900 38054 6930 38106
rect 6930 38054 6942 38106
rect 6942 38054 6956 38106
rect 6980 38054 6994 38106
rect 6994 38054 7006 38106
rect 7006 38054 7036 38106
rect 7060 38054 7070 38106
rect 7070 38054 7116 38106
rect 6820 38052 6876 38054
rect 6900 38052 6956 38054
rect 6980 38052 7036 38054
rect 7060 38052 7116 38054
rect 6820 37018 6876 37020
rect 6900 37018 6956 37020
rect 6980 37018 7036 37020
rect 7060 37018 7116 37020
rect 6820 36966 6866 37018
rect 6866 36966 6876 37018
rect 6900 36966 6930 37018
rect 6930 36966 6942 37018
rect 6942 36966 6956 37018
rect 6980 36966 6994 37018
rect 6994 36966 7006 37018
rect 7006 36966 7036 37018
rect 7060 36966 7070 37018
rect 7070 36966 7116 37018
rect 6820 36964 6876 36966
rect 6900 36964 6956 36966
rect 6980 36964 7036 36966
rect 7060 36964 7116 36966
rect 6820 35930 6876 35932
rect 6900 35930 6956 35932
rect 6980 35930 7036 35932
rect 7060 35930 7116 35932
rect 6820 35878 6866 35930
rect 6866 35878 6876 35930
rect 6900 35878 6930 35930
rect 6930 35878 6942 35930
rect 6942 35878 6956 35930
rect 6980 35878 6994 35930
rect 6994 35878 7006 35930
rect 7006 35878 7036 35930
rect 7060 35878 7070 35930
rect 7070 35878 7116 35930
rect 6820 35876 6876 35878
rect 6900 35876 6956 35878
rect 6980 35876 7036 35878
rect 7060 35876 7116 35878
rect 6820 34842 6876 34844
rect 6900 34842 6956 34844
rect 6980 34842 7036 34844
rect 7060 34842 7116 34844
rect 6820 34790 6866 34842
rect 6866 34790 6876 34842
rect 6900 34790 6930 34842
rect 6930 34790 6942 34842
rect 6942 34790 6956 34842
rect 6980 34790 6994 34842
rect 6994 34790 7006 34842
rect 7006 34790 7036 34842
rect 7060 34790 7070 34842
rect 7070 34790 7116 34842
rect 6820 34788 6876 34790
rect 6900 34788 6956 34790
rect 6980 34788 7036 34790
rect 7060 34788 7116 34790
rect 6820 33754 6876 33756
rect 6900 33754 6956 33756
rect 6980 33754 7036 33756
rect 7060 33754 7116 33756
rect 6820 33702 6866 33754
rect 6866 33702 6876 33754
rect 6900 33702 6930 33754
rect 6930 33702 6942 33754
rect 6942 33702 6956 33754
rect 6980 33702 6994 33754
rect 6994 33702 7006 33754
rect 7006 33702 7036 33754
rect 7060 33702 7070 33754
rect 7070 33702 7116 33754
rect 6820 33700 6876 33702
rect 6900 33700 6956 33702
rect 6980 33700 7036 33702
rect 7060 33700 7116 33702
rect 7194 33088 7250 33144
rect 6820 32666 6876 32668
rect 6900 32666 6956 32668
rect 6980 32666 7036 32668
rect 7060 32666 7116 32668
rect 6820 32614 6866 32666
rect 6866 32614 6876 32666
rect 6900 32614 6930 32666
rect 6930 32614 6942 32666
rect 6942 32614 6956 32666
rect 6980 32614 6994 32666
rect 6994 32614 7006 32666
rect 7006 32614 7036 32666
rect 7060 32614 7070 32666
rect 7070 32614 7116 32666
rect 6820 32612 6876 32614
rect 6900 32612 6956 32614
rect 6980 32612 7036 32614
rect 7060 32612 7116 32614
rect 5814 26324 5816 26344
rect 5816 26324 5868 26344
rect 5868 26324 5870 26344
rect 5630 24928 5686 24984
rect 5814 26288 5870 26324
rect 6182 29008 6238 29064
rect 6090 27820 6092 27840
rect 6092 27820 6144 27840
rect 6144 27820 6146 27840
rect 6090 27784 6146 27820
rect 5446 21528 5502 21584
rect 6090 24792 6146 24848
rect 6642 29416 6698 29472
rect 6550 28192 6606 28248
rect 6550 25608 6606 25664
rect 6550 25064 6606 25120
rect 6458 24248 6514 24304
rect 6274 22616 6330 22672
rect 6274 22108 6276 22128
rect 6276 22108 6328 22128
rect 6328 22108 6330 22128
rect 6274 22072 6330 22108
rect 5906 21528 5962 21584
rect 6274 21528 6330 21584
rect 5538 19896 5594 19952
rect 5446 19216 5502 19272
rect 5354 18672 5410 18728
rect 5630 17856 5686 17912
rect 5170 17040 5226 17096
rect 5170 14728 5226 14784
rect 4526 10512 4582 10568
rect 3888 7098 3944 7100
rect 3968 7098 4024 7100
rect 4048 7098 4104 7100
rect 4128 7098 4184 7100
rect 3888 7046 3934 7098
rect 3934 7046 3944 7098
rect 3968 7046 3998 7098
rect 3998 7046 4010 7098
rect 4010 7046 4024 7098
rect 4048 7046 4062 7098
rect 4062 7046 4074 7098
rect 4074 7046 4104 7098
rect 4128 7046 4138 7098
rect 4138 7046 4184 7098
rect 3888 7044 3944 7046
rect 3968 7044 4024 7046
rect 4048 7044 4104 7046
rect 4128 7044 4184 7046
rect 3888 6010 3944 6012
rect 3968 6010 4024 6012
rect 4048 6010 4104 6012
rect 4128 6010 4184 6012
rect 3888 5958 3934 6010
rect 3934 5958 3944 6010
rect 3968 5958 3998 6010
rect 3998 5958 4010 6010
rect 4010 5958 4024 6010
rect 4048 5958 4062 6010
rect 4062 5958 4074 6010
rect 4074 5958 4104 6010
rect 4128 5958 4138 6010
rect 4138 5958 4184 6010
rect 3888 5956 3944 5958
rect 3968 5956 4024 5958
rect 4048 5956 4104 5958
rect 4128 5956 4184 5958
rect 4066 5652 4068 5672
rect 4068 5652 4120 5672
rect 4120 5652 4122 5672
rect 4066 5616 4122 5652
rect 3698 5208 3754 5264
rect 4894 10784 4950 10840
rect 4802 9444 4858 9480
rect 4802 9424 4804 9444
rect 4804 9424 4856 9444
rect 4856 9424 4858 9444
rect 5354 15136 5410 15192
rect 5354 13776 5410 13832
rect 4710 6840 4766 6896
rect 3888 4922 3944 4924
rect 3968 4922 4024 4924
rect 4048 4922 4104 4924
rect 4128 4922 4184 4924
rect 3888 4870 3934 4922
rect 3934 4870 3944 4922
rect 3968 4870 3998 4922
rect 3998 4870 4010 4922
rect 4010 4870 4024 4922
rect 4048 4870 4062 4922
rect 4062 4870 4074 4922
rect 4074 4870 4104 4922
rect 4128 4870 4138 4922
rect 4138 4870 4184 4922
rect 3888 4868 3944 4870
rect 3968 4868 4024 4870
rect 4048 4868 4104 4870
rect 4128 4868 4184 4870
rect 3514 4120 3570 4176
rect 3606 3304 3662 3360
rect 3888 3834 3944 3836
rect 3968 3834 4024 3836
rect 4048 3834 4104 3836
rect 4128 3834 4184 3836
rect 3888 3782 3934 3834
rect 3934 3782 3944 3834
rect 3968 3782 3998 3834
rect 3998 3782 4010 3834
rect 4010 3782 4024 3834
rect 4048 3782 4062 3834
rect 4062 3782 4074 3834
rect 4074 3782 4104 3834
rect 4128 3782 4138 3834
rect 4138 3782 4184 3834
rect 3888 3780 3944 3782
rect 3968 3780 4024 3782
rect 4048 3780 4104 3782
rect 4128 3780 4184 3782
rect 3882 3576 3938 3632
rect 4342 3304 4398 3360
rect 5170 8608 5226 8664
rect 5078 5072 5134 5128
rect 4986 4120 5042 4176
rect 4618 3576 4674 3632
rect 4618 3440 4674 3496
rect 3888 2746 3944 2748
rect 3968 2746 4024 2748
rect 4048 2746 4104 2748
rect 4128 2746 4184 2748
rect 3888 2694 3934 2746
rect 3934 2694 3944 2746
rect 3968 2694 3998 2746
rect 3998 2694 4010 2746
rect 4010 2694 4024 2746
rect 4048 2694 4062 2746
rect 4062 2694 4074 2746
rect 4074 2694 4104 2746
rect 4128 2694 4138 2746
rect 4138 2694 4184 2746
rect 3888 2692 3944 2694
rect 3968 2692 4024 2694
rect 4048 2692 4104 2694
rect 4128 2692 4184 2694
rect 3974 2352 4030 2408
rect 3888 1658 3944 1660
rect 3968 1658 4024 1660
rect 4048 1658 4104 1660
rect 4128 1658 4184 1660
rect 3888 1606 3934 1658
rect 3934 1606 3944 1658
rect 3968 1606 3998 1658
rect 3998 1606 4010 1658
rect 4010 1606 4024 1658
rect 4048 1606 4062 1658
rect 4062 1606 4074 1658
rect 4074 1606 4104 1658
rect 4128 1606 4138 1658
rect 4138 1606 4184 1658
rect 3888 1604 3944 1606
rect 3968 1604 4024 1606
rect 4048 1604 4104 1606
rect 4128 1604 4184 1606
rect 3790 1400 3846 1456
rect 4434 1300 4436 1320
rect 4436 1300 4488 1320
rect 4488 1300 4490 1320
rect 4434 1264 4490 1300
rect 4066 720 4122 776
rect 4802 3712 4858 3768
rect 4802 3304 4858 3360
rect 5446 8880 5502 8936
rect 5722 7928 5778 7984
rect 5262 3712 5318 3768
rect 5354 3032 5410 3088
rect 5354 2644 5410 2680
rect 5722 4256 5778 4312
rect 5630 4140 5686 4176
rect 5630 4120 5632 4140
rect 5632 4120 5684 4140
rect 5684 4120 5686 4140
rect 5354 2624 5356 2644
rect 5356 2624 5408 2644
rect 5408 2624 5410 2644
rect 5906 19624 5962 19680
rect 5998 17992 6054 18048
rect 5906 12280 5962 12336
rect 6820 31578 6876 31580
rect 6900 31578 6956 31580
rect 6980 31578 7036 31580
rect 7060 31578 7116 31580
rect 6820 31526 6866 31578
rect 6866 31526 6876 31578
rect 6900 31526 6930 31578
rect 6930 31526 6942 31578
rect 6942 31526 6956 31578
rect 6980 31526 6994 31578
rect 6994 31526 7006 31578
rect 7006 31526 7036 31578
rect 7060 31526 7070 31578
rect 7070 31526 7116 31578
rect 6820 31524 6876 31526
rect 6900 31524 6956 31526
rect 6980 31524 7036 31526
rect 7060 31524 7116 31526
rect 6820 30490 6876 30492
rect 6900 30490 6956 30492
rect 6980 30490 7036 30492
rect 7060 30490 7116 30492
rect 6820 30438 6866 30490
rect 6866 30438 6876 30490
rect 6900 30438 6930 30490
rect 6930 30438 6942 30490
rect 6942 30438 6956 30490
rect 6980 30438 6994 30490
rect 6994 30438 7006 30490
rect 7006 30438 7036 30490
rect 7060 30438 7070 30490
rect 7070 30438 7116 30490
rect 6820 30436 6876 30438
rect 6900 30436 6956 30438
rect 6980 30436 7036 30438
rect 7060 30436 7116 30438
rect 6826 29960 6882 30016
rect 6820 29402 6876 29404
rect 6900 29402 6956 29404
rect 6980 29402 7036 29404
rect 7060 29402 7116 29404
rect 6820 29350 6866 29402
rect 6866 29350 6876 29402
rect 6900 29350 6930 29402
rect 6930 29350 6942 29402
rect 6942 29350 6956 29402
rect 6980 29350 6994 29402
rect 6994 29350 7006 29402
rect 7006 29350 7036 29402
rect 7060 29350 7070 29402
rect 7070 29350 7116 29402
rect 6820 29348 6876 29350
rect 6900 29348 6956 29350
rect 6980 29348 7036 29350
rect 7060 29348 7116 29350
rect 8114 42064 8170 42120
rect 9678 43152 9734 43208
rect 9753 43002 9809 43004
rect 9833 43002 9889 43004
rect 9913 43002 9969 43004
rect 9993 43002 10049 43004
rect 9753 42950 9799 43002
rect 9799 42950 9809 43002
rect 9833 42950 9863 43002
rect 9863 42950 9875 43002
rect 9875 42950 9889 43002
rect 9913 42950 9927 43002
rect 9927 42950 9939 43002
rect 9939 42950 9969 43002
rect 9993 42950 10003 43002
rect 10003 42950 10049 43002
rect 9753 42948 9809 42950
rect 9833 42948 9889 42950
rect 9913 42948 9969 42950
rect 9993 42948 10049 42950
rect 9954 42744 10010 42800
rect 9034 41792 9090 41848
rect 9310 41928 9366 41984
rect 9126 41556 9128 41576
rect 9128 41556 9180 41576
rect 9180 41556 9182 41576
rect 9126 41520 9182 41556
rect 8666 40432 8722 40488
rect 8022 36352 8078 36408
rect 7838 34448 7894 34504
rect 7838 34076 7840 34096
rect 7840 34076 7892 34096
rect 7892 34076 7894 34096
rect 7838 34040 7894 34076
rect 7746 32408 7802 32464
rect 10138 42508 10140 42528
rect 10140 42508 10192 42528
rect 10192 42508 10194 42528
rect 10138 42472 10194 42508
rect 9753 41914 9809 41916
rect 9833 41914 9889 41916
rect 9913 41914 9969 41916
rect 9993 41914 10049 41916
rect 9753 41862 9799 41914
rect 9799 41862 9809 41914
rect 9833 41862 9863 41914
rect 9863 41862 9875 41914
rect 9875 41862 9889 41914
rect 9913 41862 9927 41914
rect 9927 41862 9939 41914
rect 9939 41862 9969 41914
rect 9993 41862 10003 41914
rect 10003 41862 10049 41914
rect 9753 41860 9809 41862
rect 9833 41860 9889 41862
rect 9913 41860 9969 41862
rect 9993 41860 10049 41862
rect 9753 40826 9809 40828
rect 9833 40826 9889 40828
rect 9913 40826 9969 40828
rect 9993 40826 10049 40828
rect 9753 40774 9799 40826
rect 9799 40774 9809 40826
rect 9833 40774 9863 40826
rect 9863 40774 9875 40826
rect 9875 40774 9889 40826
rect 9913 40774 9927 40826
rect 9927 40774 9939 40826
rect 9939 40774 9969 40826
rect 9993 40774 10003 40826
rect 10003 40774 10049 40826
rect 9753 40772 9809 40774
rect 9833 40772 9889 40774
rect 9913 40772 9969 40774
rect 9993 40772 10049 40774
rect 9753 39738 9809 39740
rect 9833 39738 9889 39740
rect 9913 39738 9969 39740
rect 9993 39738 10049 39740
rect 9753 39686 9799 39738
rect 9799 39686 9809 39738
rect 9833 39686 9863 39738
rect 9863 39686 9875 39738
rect 9875 39686 9889 39738
rect 9913 39686 9927 39738
rect 9927 39686 9939 39738
rect 9939 39686 9969 39738
rect 9993 39686 10003 39738
rect 10003 39686 10049 39738
rect 9753 39684 9809 39686
rect 9833 39684 9889 39686
rect 9913 39684 9969 39686
rect 9993 39684 10049 39686
rect 9218 39480 9274 39536
rect 8758 39344 8814 39400
rect 8298 36116 8300 36136
rect 8300 36116 8352 36136
rect 8352 36116 8354 36136
rect 8298 36080 8354 36116
rect 8298 35536 8354 35592
rect 7930 32272 7986 32328
rect 7654 31592 7710 31648
rect 6820 28314 6876 28316
rect 6900 28314 6956 28316
rect 6980 28314 7036 28316
rect 7060 28314 7116 28316
rect 6820 28262 6866 28314
rect 6866 28262 6876 28314
rect 6900 28262 6930 28314
rect 6930 28262 6942 28314
rect 6942 28262 6956 28314
rect 6980 28262 6994 28314
rect 6994 28262 7006 28314
rect 7006 28262 7036 28314
rect 7060 28262 7070 28314
rect 7070 28262 7116 28314
rect 6820 28260 6876 28262
rect 6900 28260 6956 28262
rect 6980 28260 7036 28262
rect 7060 28260 7116 28262
rect 7286 27512 7342 27568
rect 6820 27226 6876 27228
rect 6900 27226 6956 27228
rect 6980 27226 7036 27228
rect 7060 27226 7116 27228
rect 6820 27174 6866 27226
rect 6866 27174 6876 27226
rect 6900 27174 6930 27226
rect 6930 27174 6942 27226
rect 6942 27174 6956 27226
rect 6980 27174 6994 27226
rect 6994 27174 7006 27226
rect 7006 27174 7036 27226
rect 7060 27174 7070 27226
rect 7070 27174 7116 27226
rect 6820 27172 6876 27174
rect 6900 27172 6956 27174
rect 6980 27172 7036 27174
rect 7060 27172 7116 27174
rect 7378 27240 7434 27296
rect 6820 26138 6876 26140
rect 6900 26138 6956 26140
rect 6980 26138 7036 26140
rect 7060 26138 7116 26140
rect 6820 26086 6866 26138
rect 6866 26086 6876 26138
rect 6900 26086 6930 26138
rect 6930 26086 6942 26138
rect 6942 26086 6956 26138
rect 6980 26086 6994 26138
rect 6994 26086 7006 26138
rect 7006 26086 7036 26138
rect 7060 26086 7070 26138
rect 7070 26086 7116 26138
rect 6820 26084 6876 26086
rect 6900 26084 6956 26086
rect 6980 26084 7036 26086
rect 7060 26084 7116 26086
rect 6820 25050 6876 25052
rect 6900 25050 6956 25052
rect 6980 25050 7036 25052
rect 7060 25050 7116 25052
rect 6820 24998 6866 25050
rect 6866 24998 6876 25050
rect 6900 24998 6930 25050
rect 6930 24998 6942 25050
rect 6942 24998 6956 25050
rect 6980 24998 6994 25050
rect 6994 24998 7006 25050
rect 7006 24998 7036 25050
rect 7060 24998 7070 25050
rect 7070 24998 7116 25050
rect 6820 24996 6876 24998
rect 6900 24996 6956 24998
rect 6980 24996 7036 24998
rect 7060 24996 7116 24998
rect 6820 23962 6876 23964
rect 6900 23962 6956 23964
rect 6980 23962 7036 23964
rect 7060 23962 7116 23964
rect 6820 23910 6866 23962
rect 6866 23910 6876 23962
rect 6900 23910 6930 23962
rect 6930 23910 6942 23962
rect 6942 23910 6956 23962
rect 6980 23910 6994 23962
rect 6994 23910 7006 23962
rect 7006 23910 7036 23962
rect 7060 23910 7070 23962
rect 7070 23910 7116 23962
rect 6820 23908 6876 23910
rect 6900 23908 6956 23910
rect 6980 23908 7036 23910
rect 7060 23908 7116 23910
rect 6820 22874 6876 22876
rect 6900 22874 6956 22876
rect 6980 22874 7036 22876
rect 7060 22874 7116 22876
rect 6820 22822 6866 22874
rect 6866 22822 6876 22874
rect 6900 22822 6930 22874
rect 6930 22822 6942 22874
rect 6942 22822 6956 22874
rect 6980 22822 6994 22874
rect 6994 22822 7006 22874
rect 7006 22822 7036 22874
rect 7060 22822 7070 22874
rect 7070 22822 7116 22874
rect 6820 22820 6876 22822
rect 6900 22820 6956 22822
rect 6980 22820 7036 22822
rect 7060 22820 7116 22822
rect 7470 26696 7526 26752
rect 7378 26560 7434 26616
rect 7470 26424 7526 26480
rect 7654 28464 7710 28520
rect 8114 31048 8170 31104
rect 7654 25880 7710 25936
rect 7654 23976 7710 24032
rect 7838 24676 7894 24712
rect 7838 24656 7840 24676
rect 7840 24656 7892 24676
rect 7892 24656 7894 24676
rect 6820 21786 6876 21788
rect 6900 21786 6956 21788
rect 6980 21786 7036 21788
rect 7060 21786 7116 21788
rect 6820 21734 6866 21786
rect 6866 21734 6876 21786
rect 6900 21734 6930 21786
rect 6930 21734 6942 21786
rect 6942 21734 6956 21786
rect 6980 21734 6994 21786
rect 6994 21734 7006 21786
rect 7006 21734 7036 21786
rect 7060 21734 7070 21786
rect 7070 21734 7116 21786
rect 6820 21732 6876 21734
rect 6900 21732 6956 21734
rect 6980 21732 7036 21734
rect 7060 21732 7116 21734
rect 6820 20698 6876 20700
rect 6900 20698 6956 20700
rect 6980 20698 7036 20700
rect 7060 20698 7116 20700
rect 6820 20646 6866 20698
rect 6866 20646 6876 20698
rect 6900 20646 6930 20698
rect 6930 20646 6942 20698
rect 6942 20646 6956 20698
rect 6980 20646 6994 20698
rect 6994 20646 7006 20698
rect 7006 20646 7036 20698
rect 7060 20646 7070 20698
rect 7070 20646 7116 20698
rect 6820 20644 6876 20646
rect 6900 20644 6956 20646
rect 6980 20644 7036 20646
rect 7060 20644 7116 20646
rect 6366 19624 6422 19680
rect 6458 19080 6514 19136
rect 6820 19610 6876 19612
rect 6900 19610 6956 19612
rect 6980 19610 7036 19612
rect 7060 19610 7116 19612
rect 6820 19558 6866 19610
rect 6866 19558 6876 19610
rect 6900 19558 6930 19610
rect 6930 19558 6942 19610
rect 6942 19558 6956 19610
rect 6980 19558 6994 19610
rect 6994 19558 7006 19610
rect 7006 19558 7036 19610
rect 7060 19558 7070 19610
rect 7070 19558 7116 19610
rect 6820 19556 6876 19558
rect 6900 19556 6956 19558
rect 6980 19556 7036 19558
rect 7060 19556 7116 19558
rect 7378 20440 7434 20496
rect 7654 23024 7710 23080
rect 9034 36524 9036 36544
rect 9036 36524 9088 36544
rect 9088 36524 9090 36544
rect 9034 36488 9090 36524
rect 8850 33260 8852 33280
rect 8852 33260 8904 33280
rect 8904 33260 8906 33280
rect 8850 33224 8906 33260
rect 8758 32172 8760 32192
rect 8760 32172 8812 32192
rect 8812 32172 8814 32192
rect 8758 32136 8814 32172
rect 7746 22616 7802 22672
rect 10046 39072 10102 39128
rect 9862 38800 9918 38856
rect 9753 38650 9809 38652
rect 9833 38650 9889 38652
rect 9913 38650 9969 38652
rect 9993 38650 10049 38652
rect 9753 38598 9799 38650
rect 9799 38598 9809 38650
rect 9833 38598 9863 38650
rect 9863 38598 9875 38650
rect 9875 38598 9889 38650
rect 9913 38598 9927 38650
rect 9927 38598 9939 38650
rect 9939 38598 9969 38650
rect 9993 38598 10003 38650
rect 10003 38598 10049 38650
rect 9753 38596 9809 38598
rect 9833 38596 9889 38598
rect 9913 38596 9969 38598
rect 9993 38596 10049 38598
rect 9753 37562 9809 37564
rect 9833 37562 9889 37564
rect 9913 37562 9969 37564
rect 9993 37562 10049 37564
rect 9753 37510 9799 37562
rect 9799 37510 9809 37562
rect 9833 37510 9863 37562
rect 9863 37510 9875 37562
rect 9875 37510 9889 37562
rect 9913 37510 9927 37562
rect 9927 37510 9939 37562
rect 9939 37510 9969 37562
rect 9993 37510 10003 37562
rect 10003 37510 10049 37562
rect 9753 37508 9809 37510
rect 9833 37508 9889 37510
rect 9913 37508 9969 37510
rect 9993 37508 10049 37510
rect 10138 36780 10194 36816
rect 10138 36760 10140 36780
rect 10140 36760 10192 36780
rect 10192 36760 10194 36780
rect 9753 36474 9809 36476
rect 9833 36474 9889 36476
rect 9913 36474 9969 36476
rect 9993 36474 10049 36476
rect 9753 36422 9799 36474
rect 9799 36422 9809 36474
rect 9833 36422 9863 36474
rect 9863 36422 9875 36474
rect 9875 36422 9889 36474
rect 9913 36422 9927 36474
rect 9927 36422 9939 36474
rect 9939 36422 9969 36474
rect 9993 36422 10003 36474
rect 10003 36422 10049 36474
rect 9753 36420 9809 36422
rect 9833 36420 9889 36422
rect 9913 36420 9969 36422
rect 9993 36420 10049 36422
rect 9753 35386 9809 35388
rect 9833 35386 9889 35388
rect 9913 35386 9969 35388
rect 9993 35386 10049 35388
rect 9753 35334 9799 35386
rect 9799 35334 9809 35386
rect 9833 35334 9863 35386
rect 9863 35334 9875 35386
rect 9875 35334 9889 35386
rect 9913 35334 9927 35386
rect 9927 35334 9939 35386
rect 9939 35334 9969 35386
rect 9993 35334 10003 35386
rect 10003 35334 10049 35386
rect 9753 35332 9809 35334
rect 9833 35332 9889 35334
rect 9913 35332 9969 35334
rect 9993 35332 10049 35334
rect 9753 34298 9809 34300
rect 9833 34298 9889 34300
rect 9913 34298 9969 34300
rect 9993 34298 10049 34300
rect 9753 34246 9799 34298
rect 9799 34246 9809 34298
rect 9833 34246 9863 34298
rect 9863 34246 9875 34298
rect 9875 34246 9889 34298
rect 9913 34246 9927 34298
rect 9927 34246 9939 34298
rect 9939 34246 9969 34298
rect 9993 34246 10003 34298
rect 10003 34246 10049 34298
rect 9753 34244 9809 34246
rect 9833 34244 9889 34246
rect 9913 34244 9969 34246
rect 9993 34244 10049 34246
rect 8574 28600 8630 28656
rect 8482 27104 8538 27160
rect 8482 26696 8538 26752
rect 8666 26560 8722 26616
rect 8758 24792 8814 24848
rect 8206 23740 8208 23760
rect 8208 23740 8260 23760
rect 8260 23740 8262 23760
rect 8206 23704 8262 23740
rect 8390 23724 8446 23760
rect 8390 23704 8392 23724
rect 8392 23704 8444 23724
rect 8444 23704 8446 23724
rect 7746 21800 7802 21856
rect 8758 23976 8814 24032
rect 7378 19386 7434 19442
rect 6458 18400 6514 18456
rect 6274 18128 6330 18184
rect 6090 15816 6146 15872
rect 6458 17040 6514 17096
rect 6642 17312 6698 17368
rect 6820 18522 6876 18524
rect 6900 18522 6956 18524
rect 6980 18522 7036 18524
rect 7060 18522 7116 18524
rect 6820 18470 6866 18522
rect 6866 18470 6876 18522
rect 6900 18470 6930 18522
rect 6930 18470 6942 18522
rect 6942 18470 6956 18522
rect 6980 18470 6994 18522
rect 6994 18470 7006 18522
rect 7006 18470 7036 18522
rect 7060 18470 7070 18522
rect 7070 18470 7116 18522
rect 6820 18468 6876 18470
rect 6900 18468 6956 18470
rect 6980 18468 7036 18470
rect 7060 18468 7116 18470
rect 6820 17434 6876 17436
rect 6900 17434 6956 17436
rect 6980 17434 7036 17436
rect 7060 17434 7116 17436
rect 6820 17382 6866 17434
rect 6866 17382 6876 17434
rect 6900 17382 6930 17434
rect 6930 17382 6942 17434
rect 6942 17382 6956 17434
rect 6980 17382 6994 17434
rect 6994 17382 7006 17434
rect 7006 17382 7036 17434
rect 7060 17382 7070 17434
rect 7070 17382 7116 17434
rect 6820 17380 6876 17382
rect 6900 17380 6956 17382
rect 6980 17380 7036 17382
rect 7060 17380 7116 17382
rect 6826 17176 6882 17232
rect 7286 17176 7342 17232
rect 6458 16224 6514 16280
rect 5998 11056 6054 11112
rect 6820 16346 6876 16348
rect 6900 16346 6956 16348
rect 6980 16346 7036 16348
rect 7060 16346 7116 16348
rect 6820 16294 6866 16346
rect 6866 16294 6876 16346
rect 6900 16294 6930 16346
rect 6930 16294 6942 16346
rect 6942 16294 6956 16346
rect 6980 16294 6994 16346
rect 6994 16294 7006 16346
rect 7006 16294 7036 16346
rect 7060 16294 7070 16346
rect 7070 16294 7116 16346
rect 6820 16292 6876 16294
rect 6900 16292 6956 16294
rect 6980 16292 7036 16294
rect 7060 16292 7116 16294
rect 7562 19292 7618 19348
rect 7746 18944 7802 19000
rect 7470 16496 7526 16552
rect 6820 15258 6876 15260
rect 6900 15258 6956 15260
rect 6980 15258 7036 15260
rect 7060 15258 7116 15260
rect 6820 15206 6866 15258
rect 6866 15206 6876 15258
rect 6900 15206 6930 15258
rect 6930 15206 6942 15258
rect 6942 15206 6956 15258
rect 6980 15206 6994 15258
rect 6994 15206 7006 15258
rect 7006 15206 7036 15258
rect 7060 15206 7070 15258
rect 7070 15206 7116 15258
rect 6820 15204 6876 15206
rect 6900 15204 6956 15206
rect 6980 15204 7036 15206
rect 7060 15204 7116 15206
rect 6820 14170 6876 14172
rect 6900 14170 6956 14172
rect 6980 14170 7036 14172
rect 7060 14170 7116 14172
rect 6820 14118 6866 14170
rect 6866 14118 6876 14170
rect 6900 14118 6930 14170
rect 6930 14118 6942 14170
rect 6942 14118 6956 14170
rect 6980 14118 6994 14170
rect 6994 14118 7006 14170
rect 7006 14118 7036 14170
rect 7060 14118 7070 14170
rect 7070 14118 7116 14170
rect 6820 14116 6876 14118
rect 6900 14116 6956 14118
rect 6980 14116 7036 14118
rect 7060 14116 7116 14118
rect 5998 8492 6054 8528
rect 5998 8472 6000 8492
rect 6000 8472 6052 8492
rect 6052 8472 6054 8492
rect 6820 13082 6876 13084
rect 6900 13082 6956 13084
rect 6980 13082 7036 13084
rect 7060 13082 7116 13084
rect 6820 13030 6866 13082
rect 6866 13030 6876 13082
rect 6900 13030 6930 13082
rect 6930 13030 6942 13082
rect 6942 13030 6956 13082
rect 6980 13030 6994 13082
rect 6994 13030 7006 13082
rect 7006 13030 7036 13082
rect 7060 13030 7070 13082
rect 7070 13030 7116 13082
rect 6820 13028 6876 13030
rect 6900 13028 6956 13030
rect 6980 13028 7036 13030
rect 7060 13028 7116 13030
rect 6550 12280 6606 12336
rect 6820 11994 6876 11996
rect 6900 11994 6956 11996
rect 6980 11994 7036 11996
rect 7060 11994 7116 11996
rect 6820 11942 6866 11994
rect 6866 11942 6876 11994
rect 6900 11942 6930 11994
rect 6930 11942 6942 11994
rect 6942 11942 6956 11994
rect 6980 11942 6994 11994
rect 6994 11942 7006 11994
rect 7006 11942 7036 11994
rect 7060 11942 7070 11994
rect 7070 11942 7116 11994
rect 6820 11940 6876 11942
rect 6900 11940 6956 11942
rect 6980 11940 7036 11942
rect 7060 11940 7116 11942
rect 6826 11600 6882 11656
rect 6550 10648 6606 10704
rect 6820 10906 6876 10908
rect 6900 10906 6956 10908
rect 6980 10906 7036 10908
rect 7060 10906 7116 10908
rect 6820 10854 6866 10906
rect 6866 10854 6876 10906
rect 6900 10854 6930 10906
rect 6930 10854 6942 10906
rect 6942 10854 6956 10906
rect 6980 10854 6994 10906
rect 6994 10854 7006 10906
rect 7006 10854 7036 10906
rect 7060 10854 7070 10906
rect 7070 10854 7116 10906
rect 6820 10852 6876 10854
rect 6900 10852 6956 10854
rect 6980 10852 7036 10854
rect 7060 10852 7116 10854
rect 6820 9818 6876 9820
rect 6900 9818 6956 9820
rect 6980 9818 7036 9820
rect 7060 9818 7116 9820
rect 6820 9766 6866 9818
rect 6866 9766 6876 9818
rect 6900 9766 6930 9818
rect 6930 9766 6942 9818
rect 6942 9766 6956 9818
rect 6980 9766 6994 9818
rect 6994 9766 7006 9818
rect 7006 9766 7036 9818
rect 7060 9766 7070 9818
rect 7070 9766 7116 9818
rect 6820 9764 6876 9766
rect 6900 9764 6956 9766
rect 6980 9764 7036 9766
rect 7060 9764 7116 9766
rect 6820 8730 6876 8732
rect 6900 8730 6956 8732
rect 6980 8730 7036 8732
rect 7060 8730 7116 8732
rect 6820 8678 6866 8730
rect 6866 8678 6876 8730
rect 6900 8678 6930 8730
rect 6930 8678 6942 8730
rect 6942 8678 6956 8730
rect 6980 8678 6994 8730
rect 6994 8678 7006 8730
rect 7006 8678 7036 8730
rect 7060 8678 7070 8730
rect 7070 8678 7116 8730
rect 6820 8676 6876 8678
rect 6900 8676 6956 8678
rect 6980 8676 7036 8678
rect 7060 8676 7116 8678
rect 6820 7642 6876 7644
rect 6900 7642 6956 7644
rect 6980 7642 7036 7644
rect 7060 7642 7116 7644
rect 6820 7590 6866 7642
rect 6866 7590 6876 7642
rect 6900 7590 6930 7642
rect 6930 7590 6942 7642
rect 6942 7590 6956 7642
rect 6980 7590 6994 7642
rect 6994 7590 7006 7642
rect 7006 7590 7036 7642
rect 7060 7590 7070 7642
rect 7070 7590 7116 7642
rect 6820 7588 6876 7590
rect 6900 7588 6956 7590
rect 6980 7588 7036 7590
rect 7060 7588 7116 7590
rect 6820 6554 6876 6556
rect 6900 6554 6956 6556
rect 6980 6554 7036 6556
rect 7060 6554 7116 6556
rect 6820 6502 6866 6554
rect 6866 6502 6876 6554
rect 6900 6502 6930 6554
rect 6930 6502 6942 6554
rect 6942 6502 6956 6554
rect 6980 6502 6994 6554
rect 6994 6502 7006 6554
rect 7006 6502 7036 6554
rect 7060 6502 7070 6554
rect 7070 6502 7116 6554
rect 6820 6500 6876 6502
rect 6900 6500 6956 6502
rect 6980 6500 7036 6502
rect 7060 6500 7116 6502
rect 6820 5466 6876 5468
rect 6900 5466 6956 5468
rect 6980 5466 7036 5468
rect 7060 5466 7116 5468
rect 6820 5414 6866 5466
rect 6866 5414 6876 5466
rect 6900 5414 6930 5466
rect 6930 5414 6942 5466
rect 6942 5414 6956 5466
rect 6980 5414 6994 5466
rect 6994 5414 7006 5466
rect 7006 5414 7036 5466
rect 7060 5414 7070 5466
rect 7070 5414 7116 5466
rect 6820 5412 6876 5414
rect 6900 5412 6956 5414
rect 6980 5412 7036 5414
rect 7060 5412 7116 5414
rect 6820 4378 6876 4380
rect 6900 4378 6956 4380
rect 6980 4378 7036 4380
rect 7060 4378 7116 4380
rect 6820 4326 6866 4378
rect 6866 4326 6876 4378
rect 6900 4326 6930 4378
rect 6930 4326 6942 4378
rect 6942 4326 6956 4378
rect 6980 4326 6994 4378
rect 6994 4326 7006 4378
rect 7006 4326 7036 4378
rect 7060 4326 7070 4378
rect 7070 4326 7116 4378
rect 6820 4324 6876 4326
rect 6900 4324 6956 4326
rect 6980 4324 7036 4326
rect 7060 4324 7116 4326
rect 7470 15020 7526 15056
rect 7470 15000 7472 15020
rect 7472 15000 7524 15020
rect 7524 15000 7526 15020
rect 7286 12280 7342 12336
rect 8390 20712 8446 20768
rect 8022 17040 8078 17096
rect 8022 16652 8078 16688
rect 8022 16632 8024 16652
rect 8024 16632 8076 16652
rect 8076 16632 8078 16652
rect 8114 16496 8170 16552
rect 8022 13812 8024 13832
rect 8024 13812 8076 13832
rect 8076 13812 8078 13832
rect 8022 13776 8078 13812
rect 7654 8472 7710 8528
rect 7654 7928 7710 7984
rect 7562 7248 7618 7304
rect 7286 4120 7342 4176
rect 6274 3440 6330 3496
rect 6366 2760 6422 2816
rect 6274 2352 6330 2408
rect 6820 3290 6876 3292
rect 6900 3290 6956 3292
rect 6980 3290 7036 3292
rect 7060 3290 7116 3292
rect 6820 3238 6866 3290
rect 6866 3238 6876 3290
rect 6900 3238 6930 3290
rect 6930 3238 6942 3290
rect 6942 3238 6956 3290
rect 6980 3238 6994 3290
rect 6994 3238 7006 3290
rect 7006 3238 7036 3290
rect 7060 3238 7070 3290
rect 7070 3238 7116 3290
rect 6820 3236 6876 3238
rect 6900 3236 6956 3238
rect 6980 3236 7036 3238
rect 7060 3236 7116 3238
rect 7378 3712 7434 3768
rect 6642 2760 6698 2816
rect 6820 2202 6876 2204
rect 6900 2202 6956 2204
rect 6980 2202 7036 2204
rect 7060 2202 7116 2204
rect 6820 2150 6866 2202
rect 6866 2150 6876 2202
rect 6900 2150 6930 2202
rect 6930 2150 6942 2202
rect 6942 2150 6956 2202
rect 6980 2150 6994 2202
rect 6994 2150 7006 2202
rect 7006 2150 7036 2202
rect 7060 2150 7070 2202
rect 7070 2150 7116 2202
rect 6820 2148 6876 2150
rect 6900 2148 6956 2150
rect 6980 2148 7036 2150
rect 7060 2148 7116 2150
rect 6820 1114 6876 1116
rect 6900 1114 6956 1116
rect 6980 1114 7036 1116
rect 7060 1114 7116 1116
rect 6820 1062 6866 1114
rect 6866 1062 6876 1114
rect 6900 1062 6930 1114
rect 6930 1062 6942 1114
rect 6942 1062 6956 1114
rect 6980 1062 6994 1114
rect 6994 1062 7006 1114
rect 7006 1062 7036 1114
rect 7060 1062 7070 1114
rect 7070 1062 7116 1114
rect 6820 1060 6876 1062
rect 6900 1060 6956 1062
rect 6980 1060 7036 1062
rect 7060 1060 7116 1062
rect 7378 3168 7434 3224
rect 7286 2216 7342 2272
rect 7470 2488 7526 2544
rect 7470 1164 7472 1184
rect 7472 1164 7524 1184
rect 7524 1164 7526 1184
rect 7470 1128 7526 1164
rect 7838 11328 7894 11384
rect 8022 4564 8024 4584
rect 8024 4564 8076 4584
rect 8076 4564 8078 4584
rect 8022 4528 8078 4564
rect 7930 3984 7986 4040
rect 7746 2760 7802 2816
rect 7654 1944 7710 2000
rect 7746 448 7802 504
rect 8298 16108 8354 16144
rect 8298 16088 8300 16108
rect 8300 16088 8352 16108
rect 8352 16088 8354 16108
rect 8298 15408 8354 15464
rect 8206 15136 8262 15192
rect 8298 14900 8300 14920
rect 8300 14900 8352 14920
rect 8352 14900 8354 14920
rect 8298 14864 8354 14900
rect 8574 20984 8630 21040
rect 8574 18536 8630 18592
rect 8574 15544 8630 15600
rect 8758 19080 8814 19136
rect 8758 18808 8814 18864
rect 9126 30912 9182 30968
rect 9034 29824 9090 29880
rect 10230 35556 10286 35592
rect 10230 35536 10232 35556
rect 10232 35536 10284 35556
rect 10284 35536 10286 35556
rect 10414 41520 10470 41576
rect 10322 33924 10378 33960
rect 10322 33904 10324 33924
rect 10324 33904 10376 33924
rect 10376 33904 10378 33924
rect 9753 33210 9809 33212
rect 9833 33210 9889 33212
rect 9913 33210 9969 33212
rect 9993 33210 10049 33212
rect 9753 33158 9799 33210
rect 9799 33158 9809 33210
rect 9833 33158 9863 33210
rect 9863 33158 9875 33210
rect 9875 33158 9889 33210
rect 9913 33158 9927 33210
rect 9927 33158 9939 33210
rect 9939 33158 9969 33210
rect 9993 33158 10003 33210
rect 10003 33158 10049 33210
rect 9753 33156 9809 33158
rect 9833 33156 9889 33158
rect 9913 33156 9969 33158
rect 9993 33156 10049 33158
rect 9753 32122 9809 32124
rect 9833 32122 9889 32124
rect 9913 32122 9969 32124
rect 9993 32122 10049 32124
rect 9753 32070 9799 32122
rect 9799 32070 9809 32122
rect 9833 32070 9863 32122
rect 9863 32070 9875 32122
rect 9875 32070 9889 32122
rect 9913 32070 9927 32122
rect 9927 32070 9939 32122
rect 9939 32070 9969 32122
rect 9993 32070 10003 32122
rect 10003 32070 10049 32122
rect 9753 32068 9809 32070
rect 9833 32068 9889 32070
rect 9913 32068 9969 32070
rect 9993 32068 10049 32070
rect 9586 31320 9642 31376
rect 9862 31864 9918 31920
rect 10230 32816 10286 32872
rect 10690 39344 10746 39400
rect 10690 39208 10746 39264
rect 9753 31034 9809 31036
rect 9833 31034 9889 31036
rect 9913 31034 9969 31036
rect 9993 31034 10049 31036
rect 9753 30982 9799 31034
rect 9799 30982 9809 31034
rect 9833 30982 9863 31034
rect 9863 30982 9875 31034
rect 9875 30982 9889 31034
rect 9913 30982 9927 31034
rect 9927 30982 9939 31034
rect 9939 30982 9969 31034
rect 9993 30982 10003 31034
rect 10003 30982 10049 31034
rect 9753 30980 9809 30982
rect 9833 30980 9889 30982
rect 9913 30980 9969 30982
rect 9993 30980 10049 30982
rect 9310 26424 9366 26480
rect 9753 29946 9809 29948
rect 9833 29946 9889 29948
rect 9913 29946 9969 29948
rect 9993 29946 10049 29948
rect 9753 29894 9799 29946
rect 9799 29894 9809 29946
rect 9833 29894 9863 29946
rect 9863 29894 9875 29946
rect 9875 29894 9889 29946
rect 9913 29894 9927 29946
rect 9927 29894 9939 29946
rect 9939 29894 9969 29946
rect 9993 29894 10003 29946
rect 10003 29894 10049 29946
rect 9753 29892 9809 29894
rect 9833 29892 9889 29894
rect 9913 29892 9969 29894
rect 9993 29892 10049 29894
rect 10138 29144 10194 29200
rect 9753 28858 9809 28860
rect 9833 28858 9889 28860
rect 9913 28858 9969 28860
rect 9993 28858 10049 28860
rect 9753 28806 9799 28858
rect 9799 28806 9809 28858
rect 9833 28806 9863 28858
rect 9863 28806 9875 28858
rect 9875 28806 9889 28858
rect 9913 28806 9927 28858
rect 9927 28806 9939 28858
rect 9939 28806 9969 28858
rect 9993 28806 10003 28858
rect 10003 28806 10049 28858
rect 9753 28804 9809 28806
rect 9833 28804 9889 28806
rect 9913 28804 9969 28806
rect 9993 28804 10049 28806
rect 10138 27820 10140 27840
rect 10140 27820 10192 27840
rect 10192 27820 10194 27840
rect 10138 27784 10194 27820
rect 9753 27770 9809 27772
rect 9833 27770 9889 27772
rect 9913 27770 9969 27772
rect 9993 27770 10049 27772
rect 9753 27718 9799 27770
rect 9799 27718 9809 27770
rect 9833 27718 9863 27770
rect 9863 27718 9875 27770
rect 9875 27718 9889 27770
rect 9913 27718 9927 27770
rect 9927 27718 9939 27770
rect 9939 27718 9969 27770
rect 9993 27718 10003 27770
rect 10003 27718 10049 27770
rect 9753 27716 9809 27718
rect 9833 27716 9889 27718
rect 9913 27716 9969 27718
rect 9993 27716 10049 27718
rect 9753 26682 9809 26684
rect 9833 26682 9889 26684
rect 9913 26682 9969 26684
rect 9993 26682 10049 26684
rect 9753 26630 9799 26682
rect 9799 26630 9809 26682
rect 9833 26630 9863 26682
rect 9863 26630 9875 26682
rect 9875 26630 9889 26682
rect 9913 26630 9927 26682
rect 9927 26630 9939 26682
rect 9939 26630 9969 26682
rect 9993 26630 10003 26682
rect 10003 26630 10049 26682
rect 9753 26628 9809 26630
rect 9833 26628 9889 26630
rect 9913 26628 9969 26630
rect 9993 26628 10049 26630
rect 9862 26152 9918 26208
rect 9126 18944 9182 19000
rect 9753 25594 9809 25596
rect 9833 25594 9889 25596
rect 9913 25594 9969 25596
rect 9993 25594 10049 25596
rect 9753 25542 9799 25594
rect 9799 25542 9809 25594
rect 9833 25542 9863 25594
rect 9863 25542 9875 25594
rect 9875 25542 9889 25594
rect 9913 25542 9927 25594
rect 9927 25542 9939 25594
rect 9939 25542 9969 25594
rect 9993 25542 10003 25594
rect 10003 25542 10049 25594
rect 9753 25540 9809 25542
rect 9833 25540 9889 25542
rect 9913 25540 9969 25542
rect 9993 25540 10049 25542
rect 9753 24506 9809 24508
rect 9833 24506 9889 24508
rect 9913 24506 9969 24508
rect 9993 24506 10049 24508
rect 9753 24454 9799 24506
rect 9799 24454 9809 24506
rect 9833 24454 9863 24506
rect 9863 24454 9875 24506
rect 9875 24454 9889 24506
rect 9913 24454 9927 24506
rect 9927 24454 9939 24506
rect 9939 24454 9969 24506
rect 9993 24454 10003 24506
rect 10003 24454 10049 24506
rect 9753 24452 9809 24454
rect 9833 24452 9889 24454
rect 9913 24452 9969 24454
rect 9993 24452 10049 24454
rect 9678 23840 9734 23896
rect 9586 23568 9642 23624
rect 10046 23604 10048 23624
rect 10048 23604 10100 23624
rect 10100 23604 10102 23624
rect 10046 23568 10102 23604
rect 9753 23418 9809 23420
rect 9833 23418 9889 23420
rect 9913 23418 9969 23420
rect 9993 23418 10049 23420
rect 9753 23366 9799 23418
rect 9799 23366 9809 23418
rect 9833 23366 9863 23418
rect 9863 23366 9875 23418
rect 9875 23366 9889 23418
rect 9913 23366 9927 23418
rect 9927 23366 9939 23418
rect 9939 23366 9969 23418
rect 9993 23366 10003 23418
rect 10003 23366 10049 23418
rect 9753 23364 9809 23366
rect 9833 23364 9889 23366
rect 9913 23364 9969 23366
rect 9993 23364 10049 23366
rect 9753 22330 9809 22332
rect 9833 22330 9889 22332
rect 9913 22330 9969 22332
rect 9993 22330 10049 22332
rect 9753 22278 9799 22330
rect 9799 22278 9809 22330
rect 9833 22278 9863 22330
rect 9863 22278 9875 22330
rect 9875 22278 9889 22330
rect 9913 22278 9927 22330
rect 9927 22278 9939 22330
rect 9939 22278 9969 22330
rect 9993 22278 10003 22330
rect 10003 22278 10049 22330
rect 9753 22276 9809 22278
rect 9833 22276 9889 22278
rect 9913 22276 9969 22278
rect 9993 22276 10049 22278
rect 9753 21242 9809 21244
rect 9833 21242 9889 21244
rect 9913 21242 9969 21244
rect 9993 21242 10049 21244
rect 9753 21190 9799 21242
rect 9799 21190 9809 21242
rect 9833 21190 9863 21242
rect 9863 21190 9875 21242
rect 9875 21190 9889 21242
rect 9913 21190 9927 21242
rect 9927 21190 9939 21242
rect 9939 21190 9969 21242
rect 9993 21190 10003 21242
rect 10003 21190 10049 21242
rect 9753 21188 9809 21190
rect 9833 21188 9889 21190
rect 9913 21188 9969 21190
rect 9993 21188 10049 21190
rect 10322 28872 10378 28928
rect 10598 30368 10654 30424
rect 10782 30504 10838 30560
rect 10230 25336 10286 25392
rect 10230 24520 10286 24576
rect 10690 27648 10746 27704
rect 11794 42880 11850 42936
rect 10966 39480 11022 39536
rect 10966 31184 11022 31240
rect 11058 30640 11114 30696
rect 11518 39072 11574 39128
rect 11242 36624 11298 36680
rect 11058 30368 11114 30424
rect 10966 30268 10968 30288
rect 10968 30268 11020 30288
rect 11020 30268 11022 30288
rect 10966 30232 11022 30268
rect 11058 26968 11114 27024
rect 10966 26560 11022 26616
rect 10782 25880 10838 25936
rect 10598 24792 10654 24848
rect 10414 24384 10470 24440
rect 9494 20576 9550 20632
rect 9862 20984 9918 21040
rect 10138 20304 10194 20360
rect 9753 20154 9809 20156
rect 9833 20154 9889 20156
rect 9913 20154 9969 20156
rect 9993 20154 10049 20156
rect 9753 20102 9799 20154
rect 9799 20102 9809 20154
rect 9833 20102 9863 20154
rect 9863 20102 9875 20154
rect 9875 20102 9889 20154
rect 9913 20102 9927 20154
rect 9927 20102 9939 20154
rect 9939 20102 9969 20154
rect 9993 20102 10003 20154
rect 10003 20102 10049 20154
rect 9753 20100 9809 20102
rect 9833 20100 9889 20102
rect 9913 20100 9969 20102
rect 9993 20100 10049 20102
rect 9753 19066 9809 19068
rect 9833 19066 9889 19068
rect 9913 19066 9969 19068
rect 9993 19066 10049 19068
rect 9753 19014 9799 19066
rect 9799 19014 9809 19066
rect 9833 19014 9863 19066
rect 9863 19014 9875 19066
rect 9875 19014 9889 19066
rect 9913 19014 9927 19066
rect 9927 19014 9939 19066
rect 9939 19014 9969 19066
rect 9993 19014 10003 19066
rect 10003 19014 10049 19066
rect 9753 19012 9809 19014
rect 9833 19012 9889 19014
rect 9913 19012 9969 19014
rect 9993 19012 10049 19014
rect 9954 18808 10010 18864
rect 9402 18400 9458 18456
rect 10230 18536 10286 18592
rect 9310 17196 9366 17232
rect 9310 17176 9312 17196
rect 9312 17176 9364 17196
rect 9364 17176 9366 17196
rect 8758 14456 8814 14512
rect 8758 13096 8814 13152
rect 8390 11056 8446 11112
rect 9494 18128 9550 18184
rect 9753 17978 9809 17980
rect 9833 17978 9889 17980
rect 9913 17978 9969 17980
rect 9993 17978 10049 17980
rect 9753 17926 9799 17978
rect 9799 17926 9809 17978
rect 9833 17926 9863 17978
rect 9863 17926 9875 17978
rect 9875 17926 9889 17978
rect 9913 17926 9927 17978
rect 9927 17926 9939 17978
rect 9939 17926 9969 17978
rect 9993 17926 10003 17978
rect 10003 17926 10049 17978
rect 9753 17924 9809 17926
rect 9833 17924 9889 17926
rect 9913 17924 9969 17926
rect 9993 17924 10049 17926
rect 10598 23840 10654 23896
rect 10506 23568 10562 23624
rect 10782 24248 10838 24304
rect 10414 21528 10470 21584
rect 10598 22616 10654 22672
rect 11426 37712 11482 37768
rect 11242 29144 11298 29200
rect 11242 28600 11298 28656
rect 11702 38700 11704 38720
rect 11704 38700 11756 38720
rect 11756 38700 11758 38720
rect 11702 38664 11758 38700
rect 11702 34584 11758 34640
rect 11702 32272 11758 32328
rect 11610 30776 11666 30832
rect 11518 30096 11574 30152
rect 12685 43546 12741 43548
rect 12765 43546 12821 43548
rect 12845 43546 12901 43548
rect 12925 43546 12981 43548
rect 12685 43494 12731 43546
rect 12731 43494 12741 43546
rect 12765 43494 12795 43546
rect 12795 43494 12807 43546
rect 12807 43494 12821 43546
rect 12845 43494 12859 43546
rect 12859 43494 12871 43546
rect 12871 43494 12901 43546
rect 12925 43494 12935 43546
rect 12935 43494 12981 43546
rect 12685 43492 12741 43494
rect 12765 43492 12821 43494
rect 12845 43492 12901 43494
rect 12925 43492 12981 43494
rect 12162 37340 12164 37360
rect 12164 37340 12216 37360
rect 12216 37340 12218 37360
rect 12162 37304 12218 37340
rect 11978 31184 12034 31240
rect 11886 30368 11942 30424
rect 11518 29552 11574 29608
rect 11518 28872 11574 28928
rect 11702 27920 11758 27976
rect 11702 27376 11758 27432
rect 11334 24792 11390 24848
rect 10506 19896 10562 19952
rect 9753 16890 9809 16892
rect 9833 16890 9889 16892
rect 9913 16890 9969 16892
rect 9993 16890 10049 16892
rect 9753 16838 9799 16890
rect 9799 16838 9809 16890
rect 9833 16838 9863 16890
rect 9863 16838 9875 16890
rect 9875 16838 9889 16890
rect 9913 16838 9927 16890
rect 9927 16838 9939 16890
rect 9939 16838 9969 16890
rect 9993 16838 10003 16890
rect 10003 16838 10049 16890
rect 9753 16836 9809 16838
rect 9833 16836 9889 16838
rect 9913 16836 9969 16838
rect 9993 16836 10049 16838
rect 10046 16632 10102 16688
rect 10322 16768 10378 16824
rect 9753 15802 9809 15804
rect 9833 15802 9889 15804
rect 9913 15802 9969 15804
rect 9993 15802 10049 15804
rect 9753 15750 9799 15802
rect 9799 15750 9809 15802
rect 9833 15750 9863 15802
rect 9863 15750 9875 15802
rect 9875 15750 9889 15802
rect 9913 15750 9927 15802
rect 9927 15750 9939 15802
rect 9939 15750 9969 15802
rect 9993 15750 10003 15802
rect 10003 15750 10049 15802
rect 9753 15748 9809 15750
rect 9833 15748 9889 15750
rect 9913 15748 9969 15750
rect 9993 15748 10049 15750
rect 9753 14714 9809 14716
rect 9833 14714 9889 14716
rect 9913 14714 9969 14716
rect 9993 14714 10049 14716
rect 9753 14662 9799 14714
rect 9799 14662 9809 14714
rect 9833 14662 9863 14714
rect 9863 14662 9875 14714
rect 9875 14662 9889 14714
rect 9913 14662 9927 14714
rect 9927 14662 9939 14714
rect 9939 14662 9969 14714
rect 9993 14662 10003 14714
rect 10003 14662 10049 14714
rect 9753 14660 9809 14662
rect 9833 14660 9889 14662
rect 9913 14660 9969 14662
rect 9993 14660 10049 14662
rect 9753 13626 9809 13628
rect 9833 13626 9889 13628
rect 9913 13626 9969 13628
rect 9993 13626 10049 13628
rect 9753 13574 9799 13626
rect 9799 13574 9809 13626
rect 9833 13574 9863 13626
rect 9863 13574 9875 13626
rect 9875 13574 9889 13626
rect 9913 13574 9927 13626
rect 9927 13574 9939 13626
rect 9939 13574 9969 13626
rect 9993 13574 10003 13626
rect 10003 13574 10049 13626
rect 9753 13572 9809 13574
rect 9833 13572 9889 13574
rect 9913 13572 9969 13574
rect 9993 13572 10049 13574
rect 10322 14320 10378 14376
rect 9494 12860 9496 12880
rect 9496 12860 9548 12880
rect 9548 12860 9550 12880
rect 9494 12824 9550 12860
rect 9753 12538 9809 12540
rect 9833 12538 9889 12540
rect 9913 12538 9969 12540
rect 9993 12538 10049 12540
rect 9753 12486 9799 12538
rect 9799 12486 9809 12538
rect 9833 12486 9863 12538
rect 9863 12486 9875 12538
rect 9875 12486 9889 12538
rect 9913 12486 9927 12538
rect 9927 12486 9939 12538
rect 9939 12486 9969 12538
rect 9993 12486 10003 12538
rect 10003 12486 10049 12538
rect 9753 12484 9809 12486
rect 9833 12484 9889 12486
rect 9913 12484 9969 12486
rect 9993 12484 10049 12486
rect 8206 3440 8262 3496
rect 8942 5208 8998 5264
rect 8850 3052 8906 3088
rect 8850 3032 8852 3052
rect 8852 3032 8904 3052
rect 8904 3032 8906 3052
rect 8114 2216 8170 2272
rect 7930 1300 7932 1320
rect 7932 1300 7984 1320
rect 7984 1300 7986 1320
rect 7930 1264 7986 1300
rect 8390 1828 8446 1864
rect 8390 1808 8392 1828
rect 8392 1808 8444 1828
rect 8444 1808 8446 1828
rect 8850 2216 8906 2272
rect 9753 11450 9809 11452
rect 9833 11450 9889 11452
rect 9913 11450 9969 11452
rect 9993 11450 10049 11452
rect 9753 11398 9799 11450
rect 9799 11398 9809 11450
rect 9833 11398 9863 11450
rect 9863 11398 9875 11450
rect 9875 11398 9889 11450
rect 9913 11398 9927 11450
rect 9927 11398 9939 11450
rect 9939 11398 9969 11450
rect 9993 11398 10003 11450
rect 10003 11398 10049 11450
rect 9753 11396 9809 11398
rect 9833 11396 9889 11398
rect 9913 11396 9969 11398
rect 9993 11396 10049 11398
rect 9753 10362 9809 10364
rect 9833 10362 9889 10364
rect 9913 10362 9969 10364
rect 9993 10362 10049 10364
rect 9753 10310 9799 10362
rect 9799 10310 9809 10362
rect 9833 10310 9863 10362
rect 9863 10310 9875 10362
rect 9875 10310 9889 10362
rect 9913 10310 9927 10362
rect 9927 10310 9939 10362
rect 9939 10310 9969 10362
rect 9993 10310 10003 10362
rect 10003 10310 10049 10362
rect 9753 10308 9809 10310
rect 9833 10308 9889 10310
rect 9913 10308 9969 10310
rect 9993 10308 10049 10310
rect 9753 9274 9809 9276
rect 9833 9274 9889 9276
rect 9913 9274 9969 9276
rect 9993 9274 10049 9276
rect 9753 9222 9799 9274
rect 9799 9222 9809 9274
rect 9833 9222 9863 9274
rect 9863 9222 9875 9274
rect 9875 9222 9889 9274
rect 9913 9222 9927 9274
rect 9927 9222 9939 9274
rect 9939 9222 9969 9274
rect 9993 9222 10003 9274
rect 10003 9222 10049 9274
rect 9753 9220 9809 9222
rect 9833 9220 9889 9222
rect 9913 9220 9969 9222
rect 9993 9220 10049 9222
rect 9753 8186 9809 8188
rect 9833 8186 9889 8188
rect 9913 8186 9969 8188
rect 9993 8186 10049 8188
rect 9753 8134 9799 8186
rect 9799 8134 9809 8186
rect 9833 8134 9863 8186
rect 9863 8134 9875 8186
rect 9875 8134 9889 8186
rect 9913 8134 9927 8186
rect 9927 8134 9939 8186
rect 9939 8134 9969 8186
rect 9993 8134 10003 8186
rect 10003 8134 10049 8186
rect 9753 8132 9809 8134
rect 9833 8132 9889 8134
rect 9913 8132 9969 8134
rect 9993 8132 10049 8134
rect 9770 7928 9826 7984
rect 9126 6316 9182 6352
rect 9126 6296 9128 6316
rect 9128 6296 9180 6316
rect 9180 6296 9182 6316
rect 9126 6160 9182 6216
rect 9753 7098 9809 7100
rect 9833 7098 9889 7100
rect 9913 7098 9969 7100
rect 9993 7098 10049 7100
rect 9753 7046 9799 7098
rect 9799 7046 9809 7098
rect 9833 7046 9863 7098
rect 9863 7046 9875 7098
rect 9875 7046 9889 7098
rect 9913 7046 9927 7098
rect 9927 7046 9939 7098
rect 9939 7046 9969 7098
rect 9993 7046 10003 7098
rect 10003 7046 10049 7098
rect 9753 7044 9809 7046
rect 9833 7044 9889 7046
rect 9913 7044 9969 7046
rect 9993 7044 10049 7046
rect 9678 6704 9734 6760
rect 9753 6010 9809 6012
rect 9833 6010 9889 6012
rect 9913 6010 9969 6012
rect 9993 6010 10049 6012
rect 9753 5958 9799 6010
rect 9799 5958 9809 6010
rect 9833 5958 9863 6010
rect 9863 5958 9875 6010
rect 9875 5958 9889 6010
rect 9913 5958 9927 6010
rect 9927 5958 9939 6010
rect 9939 5958 9969 6010
rect 9993 5958 10003 6010
rect 10003 5958 10049 6010
rect 9753 5956 9809 5958
rect 9833 5956 9889 5958
rect 9913 5956 9969 5958
rect 9993 5956 10049 5958
rect 10230 6568 10286 6624
rect 10506 13368 10562 13424
rect 10966 21392 11022 21448
rect 10874 16768 10930 16824
rect 10690 13776 10746 13832
rect 10782 13096 10838 13152
rect 9753 4922 9809 4924
rect 9833 4922 9889 4924
rect 9913 4922 9969 4924
rect 9993 4922 10049 4924
rect 9753 4870 9799 4922
rect 9799 4870 9809 4922
rect 9833 4870 9863 4922
rect 9863 4870 9875 4922
rect 9875 4870 9889 4922
rect 9913 4870 9927 4922
rect 9927 4870 9939 4922
rect 9939 4870 9969 4922
rect 9993 4870 10003 4922
rect 10003 4870 10049 4922
rect 9753 4868 9809 4870
rect 9833 4868 9889 4870
rect 9913 4868 9969 4870
rect 9993 4868 10049 4870
rect 9753 3834 9809 3836
rect 9833 3834 9889 3836
rect 9913 3834 9969 3836
rect 9993 3834 10049 3836
rect 9753 3782 9799 3834
rect 9799 3782 9809 3834
rect 9833 3782 9863 3834
rect 9863 3782 9875 3834
rect 9875 3782 9889 3834
rect 9913 3782 9927 3834
rect 9927 3782 9939 3834
rect 9939 3782 9969 3834
rect 9993 3782 10003 3834
rect 10003 3782 10049 3834
rect 9753 3780 9809 3782
rect 9833 3780 9889 3782
rect 9913 3780 9969 3782
rect 9993 3780 10049 3782
rect 9218 1128 9274 1184
rect 9494 1944 9550 2000
rect 9753 2746 9809 2748
rect 9833 2746 9889 2748
rect 9913 2746 9969 2748
rect 9993 2746 10049 2748
rect 9753 2694 9799 2746
rect 9799 2694 9809 2746
rect 9833 2694 9863 2746
rect 9863 2694 9875 2746
rect 9875 2694 9889 2746
rect 9913 2694 9927 2746
rect 9927 2694 9939 2746
rect 9939 2694 9969 2746
rect 9993 2694 10003 2746
rect 10003 2694 10049 2746
rect 9753 2692 9809 2694
rect 9833 2692 9889 2694
rect 9913 2692 9969 2694
rect 9993 2692 10049 2694
rect 9678 2216 9734 2272
rect 11242 20984 11298 21040
rect 11150 20848 11206 20904
rect 11150 18672 11206 18728
rect 11242 18264 11298 18320
rect 12070 29280 12126 29336
rect 11978 26832 12034 26888
rect 11978 26424 12034 26480
rect 12070 25372 12072 25392
rect 12072 25372 12124 25392
rect 12124 25372 12126 25392
rect 12070 25336 12126 25372
rect 11886 23724 11942 23760
rect 11886 23704 11888 23724
rect 11888 23704 11940 23724
rect 11940 23704 11942 23724
rect 11518 20340 11520 20360
rect 11520 20340 11572 20360
rect 11572 20340 11574 20360
rect 11518 20304 11574 20340
rect 11702 21936 11758 21992
rect 11794 21664 11850 21720
rect 11058 9424 11114 9480
rect 11610 16652 11666 16688
rect 11610 16632 11612 16652
rect 11612 16632 11664 16652
rect 11664 16632 11666 16652
rect 11518 14864 11574 14920
rect 11610 13368 11666 13424
rect 12530 43052 12532 43072
rect 12532 43052 12584 43072
rect 12584 43052 12586 43072
rect 12530 43016 12586 43052
rect 12685 42458 12741 42460
rect 12765 42458 12821 42460
rect 12845 42458 12901 42460
rect 12925 42458 12981 42460
rect 12685 42406 12731 42458
rect 12731 42406 12741 42458
rect 12765 42406 12795 42458
rect 12795 42406 12807 42458
rect 12807 42406 12821 42458
rect 12845 42406 12859 42458
rect 12859 42406 12871 42458
rect 12871 42406 12901 42458
rect 12925 42406 12935 42458
rect 12935 42406 12981 42458
rect 12685 42404 12741 42406
rect 12765 42404 12821 42406
rect 12845 42404 12901 42406
rect 12925 42404 12981 42406
rect 12438 41384 12494 41440
rect 12685 41370 12741 41372
rect 12765 41370 12821 41372
rect 12845 41370 12901 41372
rect 12925 41370 12981 41372
rect 12685 41318 12731 41370
rect 12731 41318 12741 41370
rect 12765 41318 12795 41370
rect 12795 41318 12807 41370
rect 12807 41318 12821 41370
rect 12845 41318 12859 41370
rect 12859 41318 12871 41370
rect 12871 41318 12901 41370
rect 12925 41318 12935 41370
rect 12935 41318 12981 41370
rect 12685 41316 12741 41318
rect 12765 41316 12821 41318
rect 12845 41316 12901 41318
rect 12925 41316 12981 41318
rect 12685 40282 12741 40284
rect 12765 40282 12821 40284
rect 12845 40282 12901 40284
rect 12925 40282 12981 40284
rect 12685 40230 12731 40282
rect 12731 40230 12741 40282
rect 12765 40230 12795 40282
rect 12795 40230 12807 40282
rect 12807 40230 12821 40282
rect 12845 40230 12859 40282
rect 12859 40230 12871 40282
rect 12871 40230 12901 40282
rect 12925 40230 12935 40282
rect 12935 40230 12981 40282
rect 12685 40228 12741 40230
rect 12765 40228 12821 40230
rect 12845 40228 12901 40230
rect 12925 40228 12981 40230
rect 12685 39194 12741 39196
rect 12765 39194 12821 39196
rect 12845 39194 12901 39196
rect 12925 39194 12981 39196
rect 12685 39142 12731 39194
rect 12731 39142 12741 39194
rect 12765 39142 12795 39194
rect 12795 39142 12807 39194
rect 12807 39142 12821 39194
rect 12845 39142 12859 39194
rect 12859 39142 12871 39194
rect 12871 39142 12901 39194
rect 12925 39142 12935 39194
rect 12935 39142 12981 39194
rect 12685 39140 12741 39142
rect 12765 39140 12821 39142
rect 12845 39140 12901 39142
rect 12925 39140 12981 39142
rect 12685 38106 12741 38108
rect 12765 38106 12821 38108
rect 12845 38106 12901 38108
rect 12925 38106 12981 38108
rect 12685 38054 12731 38106
rect 12731 38054 12741 38106
rect 12765 38054 12795 38106
rect 12795 38054 12807 38106
rect 12807 38054 12821 38106
rect 12845 38054 12859 38106
rect 12859 38054 12871 38106
rect 12871 38054 12901 38106
rect 12925 38054 12935 38106
rect 12935 38054 12981 38106
rect 12685 38052 12741 38054
rect 12765 38052 12821 38054
rect 12845 38052 12901 38054
rect 12925 38052 12981 38054
rect 12685 37018 12741 37020
rect 12765 37018 12821 37020
rect 12845 37018 12901 37020
rect 12925 37018 12981 37020
rect 12685 36966 12731 37018
rect 12731 36966 12741 37018
rect 12765 36966 12795 37018
rect 12795 36966 12807 37018
rect 12807 36966 12821 37018
rect 12845 36966 12859 37018
rect 12859 36966 12871 37018
rect 12871 36966 12901 37018
rect 12925 36966 12935 37018
rect 12935 36966 12981 37018
rect 12685 36964 12741 36966
rect 12765 36964 12821 36966
rect 12845 36964 12901 36966
rect 12925 36964 12981 36966
rect 12685 35930 12741 35932
rect 12765 35930 12821 35932
rect 12845 35930 12901 35932
rect 12925 35930 12981 35932
rect 12685 35878 12731 35930
rect 12731 35878 12741 35930
rect 12765 35878 12795 35930
rect 12795 35878 12807 35930
rect 12807 35878 12821 35930
rect 12845 35878 12859 35930
rect 12859 35878 12871 35930
rect 12871 35878 12901 35930
rect 12925 35878 12935 35930
rect 12935 35878 12981 35930
rect 12685 35876 12741 35878
rect 12765 35876 12821 35878
rect 12845 35876 12901 35878
rect 12925 35876 12981 35878
rect 12685 34842 12741 34844
rect 12765 34842 12821 34844
rect 12845 34842 12901 34844
rect 12925 34842 12981 34844
rect 12685 34790 12731 34842
rect 12731 34790 12741 34842
rect 12765 34790 12795 34842
rect 12795 34790 12807 34842
rect 12807 34790 12821 34842
rect 12845 34790 12859 34842
rect 12859 34790 12871 34842
rect 12871 34790 12901 34842
rect 12925 34790 12935 34842
rect 12935 34790 12981 34842
rect 12685 34788 12741 34790
rect 12765 34788 12821 34790
rect 12845 34788 12901 34790
rect 12925 34788 12981 34790
rect 13082 34584 13138 34640
rect 12254 33360 12310 33416
rect 12685 33754 12741 33756
rect 12765 33754 12821 33756
rect 12845 33754 12901 33756
rect 12925 33754 12981 33756
rect 12685 33702 12731 33754
rect 12731 33702 12741 33754
rect 12765 33702 12795 33754
rect 12795 33702 12807 33754
rect 12807 33702 12821 33754
rect 12845 33702 12859 33754
rect 12859 33702 12871 33754
rect 12871 33702 12901 33754
rect 12925 33702 12935 33754
rect 12935 33702 12981 33754
rect 12685 33700 12741 33702
rect 12765 33700 12821 33702
rect 12845 33700 12901 33702
rect 12925 33700 12981 33702
rect 12438 33516 12494 33552
rect 12438 33496 12440 33516
rect 12440 33496 12492 33516
rect 12492 33496 12494 33516
rect 12806 33224 12862 33280
rect 12254 31184 12310 31240
rect 12685 32666 12741 32668
rect 12765 32666 12821 32668
rect 12845 32666 12901 32668
rect 12925 32666 12981 32668
rect 12685 32614 12731 32666
rect 12731 32614 12741 32666
rect 12765 32614 12795 32666
rect 12795 32614 12807 32666
rect 12807 32614 12821 32666
rect 12845 32614 12859 32666
rect 12859 32614 12871 32666
rect 12871 32614 12901 32666
rect 12925 32614 12935 32666
rect 12935 32614 12981 32666
rect 12685 32612 12741 32614
rect 12765 32612 12821 32614
rect 12845 32612 12901 32614
rect 12925 32612 12981 32614
rect 12685 31578 12741 31580
rect 12765 31578 12821 31580
rect 12845 31578 12901 31580
rect 12925 31578 12981 31580
rect 12685 31526 12731 31578
rect 12731 31526 12741 31578
rect 12765 31526 12795 31578
rect 12795 31526 12807 31578
rect 12807 31526 12821 31578
rect 12845 31526 12859 31578
rect 12859 31526 12871 31578
rect 12871 31526 12901 31578
rect 12925 31526 12935 31578
rect 12935 31526 12981 31578
rect 12685 31524 12741 31526
rect 12765 31524 12821 31526
rect 12845 31524 12901 31526
rect 12925 31524 12981 31526
rect 12806 31220 12808 31240
rect 12808 31220 12860 31240
rect 12860 31220 12862 31240
rect 12806 31184 12862 31220
rect 12530 30540 12532 30560
rect 12532 30540 12584 30560
rect 12584 30540 12586 30560
rect 12530 30504 12586 30540
rect 12685 30490 12741 30492
rect 12765 30490 12821 30492
rect 12845 30490 12901 30492
rect 12925 30490 12981 30492
rect 12685 30438 12731 30490
rect 12731 30438 12741 30490
rect 12765 30438 12795 30490
rect 12795 30438 12807 30490
rect 12807 30438 12821 30490
rect 12845 30438 12859 30490
rect 12859 30438 12871 30490
rect 12871 30438 12901 30490
rect 12925 30438 12935 30490
rect 12935 30438 12981 30490
rect 12685 30436 12741 30438
rect 12765 30436 12821 30438
rect 12845 30436 12901 30438
rect 12925 30436 12981 30438
rect 12438 28076 12494 28112
rect 12438 28056 12440 28076
rect 12440 28056 12492 28076
rect 12492 28056 12494 28076
rect 12254 26324 12256 26344
rect 12256 26324 12308 26344
rect 12308 26324 12310 26344
rect 12254 26288 12310 26324
rect 12685 29402 12741 29404
rect 12765 29402 12821 29404
rect 12845 29402 12901 29404
rect 12925 29402 12981 29404
rect 12685 29350 12731 29402
rect 12731 29350 12741 29402
rect 12765 29350 12795 29402
rect 12795 29350 12807 29402
rect 12807 29350 12821 29402
rect 12845 29350 12859 29402
rect 12859 29350 12871 29402
rect 12871 29350 12901 29402
rect 12925 29350 12935 29402
rect 12935 29350 12981 29402
rect 12685 29348 12741 29350
rect 12765 29348 12821 29350
rect 12845 29348 12901 29350
rect 12925 29348 12981 29350
rect 12685 28314 12741 28316
rect 12765 28314 12821 28316
rect 12845 28314 12901 28316
rect 12925 28314 12981 28316
rect 12685 28262 12731 28314
rect 12731 28262 12741 28314
rect 12765 28262 12795 28314
rect 12795 28262 12807 28314
rect 12807 28262 12821 28314
rect 12845 28262 12859 28314
rect 12859 28262 12871 28314
rect 12871 28262 12901 28314
rect 12925 28262 12935 28314
rect 12935 28262 12981 28314
rect 12685 28260 12741 28262
rect 12765 28260 12821 28262
rect 12845 28260 12901 28262
rect 12925 28260 12981 28262
rect 12990 27940 13046 27976
rect 12990 27920 12992 27940
rect 12992 27920 13044 27940
rect 13044 27920 13046 27940
rect 13082 27648 13138 27704
rect 12685 27226 12741 27228
rect 12765 27226 12821 27228
rect 12845 27226 12901 27228
rect 12925 27226 12981 27228
rect 12685 27174 12731 27226
rect 12731 27174 12741 27226
rect 12765 27174 12795 27226
rect 12795 27174 12807 27226
rect 12807 27174 12821 27226
rect 12845 27174 12859 27226
rect 12859 27174 12871 27226
rect 12871 27174 12901 27226
rect 12925 27174 12935 27226
rect 12935 27174 12981 27226
rect 12685 27172 12741 27174
rect 12765 27172 12821 27174
rect 12845 27172 12901 27174
rect 12925 27172 12981 27174
rect 12685 26138 12741 26140
rect 12765 26138 12821 26140
rect 12845 26138 12901 26140
rect 12925 26138 12981 26140
rect 12685 26086 12731 26138
rect 12731 26086 12741 26138
rect 12765 26086 12795 26138
rect 12795 26086 12807 26138
rect 12807 26086 12821 26138
rect 12845 26086 12859 26138
rect 12859 26086 12871 26138
rect 12871 26086 12901 26138
rect 12925 26086 12935 26138
rect 12935 26086 12981 26138
rect 12685 26084 12741 26086
rect 12765 26084 12821 26086
rect 12845 26084 12901 26086
rect 12925 26084 12981 26086
rect 12530 25356 12586 25392
rect 12530 25336 12532 25356
rect 12532 25336 12584 25356
rect 12584 25336 12586 25356
rect 12685 25050 12741 25052
rect 12765 25050 12821 25052
rect 12845 25050 12901 25052
rect 12925 25050 12981 25052
rect 12685 24998 12731 25050
rect 12731 24998 12741 25050
rect 12765 24998 12795 25050
rect 12795 24998 12807 25050
rect 12807 24998 12821 25050
rect 12845 24998 12859 25050
rect 12859 24998 12871 25050
rect 12871 24998 12901 25050
rect 12925 24998 12935 25050
rect 12935 24998 12981 25050
rect 12685 24996 12741 24998
rect 12765 24996 12821 24998
rect 12845 24996 12901 24998
rect 12925 24996 12981 24998
rect 12685 23962 12741 23964
rect 12765 23962 12821 23964
rect 12845 23962 12901 23964
rect 12925 23962 12981 23964
rect 12685 23910 12731 23962
rect 12731 23910 12741 23962
rect 12765 23910 12795 23962
rect 12795 23910 12807 23962
rect 12807 23910 12821 23962
rect 12845 23910 12859 23962
rect 12859 23910 12871 23962
rect 12871 23910 12901 23962
rect 12925 23910 12935 23962
rect 12935 23910 12981 23962
rect 12685 23908 12741 23910
rect 12765 23908 12821 23910
rect 12845 23908 12901 23910
rect 12925 23908 12981 23910
rect 12162 21800 12218 21856
rect 12685 22874 12741 22876
rect 12765 22874 12821 22876
rect 12845 22874 12901 22876
rect 12925 22874 12981 22876
rect 12685 22822 12731 22874
rect 12731 22822 12741 22874
rect 12765 22822 12795 22874
rect 12795 22822 12807 22874
rect 12807 22822 12821 22874
rect 12845 22822 12859 22874
rect 12859 22822 12871 22874
rect 12871 22822 12901 22874
rect 12925 22822 12935 22874
rect 12935 22822 12981 22874
rect 12685 22820 12741 22822
rect 12765 22820 12821 22822
rect 12845 22820 12901 22822
rect 12925 22820 12981 22822
rect 13266 23432 13322 23488
rect 13266 22108 13268 22128
rect 13268 22108 13320 22128
rect 13320 22108 13322 22128
rect 13266 22072 13322 22108
rect 12685 21786 12741 21788
rect 12765 21786 12821 21788
rect 12845 21786 12901 21788
rect 12925 21786 12981 21788
rect 12685 21734 12731 21786
rect 12731 21734 12741 21786
rect 12765 21734 12795 21786
rect 12795 21734 12807 21786
rect 12807 21734 12821 21786
rect 12845 21734 12859 21786
rect 12859 21734 12871 21786
rect 12871 21734 12901 21786
rect 12925 21734 12935 21786
rect 12935 21734 12981 21786
rect 12685 21732 12741 21734
rect 12765 21732 12821 21734
rect 12845 21732 12901 21734
rect 12925 21732 12981 21734
rect 12070 19372 12126 19408
rect 12070 19352 12072 19372
rect 12072 19352 12124 19372
rect 12124 19352 12126 19372
rect 12346 20460 12402 20496
rect 12346 20440 12348 20460
rect 12348 20440 12400 20460
rect 12400 20440 12402 20460
rect 12685 20698 12741 20700
rect 12765 20698 12821 20700
rect 12845 20698 12901 20700
rect 12925 20698 12981 20700
rect 12685 20646 12731 20698
rect 12731 20646 12741 20698
rect 12765 20646 12795 20698
rect 12795 20646 12807 20698
rect 12807 20646 12821 20698
rect 12845 20646 12859 20698
rect 12859 20646 12871 20698
rect 12871 20646 12901 20698
rect 12925 20646 12935 20698
rect 12935 20646 12981 20698
rect 12685 20644 12741 20646
rect 12765 20644 12821 20646
rect 12845 20644 12901 20646
rect 12925 20644 12981 20646
rect 12685 19610 12741 19612
rect 12765 19610 12821 19612
rect 12845 19610 12901 19612
rect 12925 19610 12981 19612
rect 12685 19558 12731 19610
rect 12731 19558 12741 19610
rect 12765 19558 12795 19610
rect 12795 19558 12807 19610
rect 12807 19558 12821 19610
rect 12845 19558 12859 19610
rect 12859 19558 12871 19610
rect 12871 19558 12901 19610
rect 12925 19558 12935 19610
rect 12935 19558 12981 19610
rect 12685 19556 12741 19558
rect 12765 19556 12821 19558
rect 12845 19556 12901 19558
rect 12925 19556 12981 19558
rect 13634 38256 13690 38312
rect 13818 41112 13874 41168
rect 14094 42200 14150 42256
rect 14002 40976 14058 41032
rect 15014 42880 15070 42936
rect 15618 43002 15674 43004
rect 15698 43002 15754 43004
rect 15778 43002 15834 43004
rect 15858 43002 15914 43004
rect 15618 42950 15664 43002
rect 15664 42950 15674 43002
rect 15698 42950 15728 43002
rect 15728 42950 15740 43002
rect 15740 42950 15754 43002
rect 15778 42950 15792 43002
rect 15792 42950 15804 43002
rect 15804 42950 15834 43002
rect 15858 42950 15868 43002
rect 15868 42950 15914 43002
rect 15618 42948 15674 42950
rect 15698 42948 15754 42950
rect 15778 42948 15834 42950
rect 15858 42948 15914 42950
rect 15474 42880 15530 42936
rect 15618 41914 15674 41916
rect 15698 41914 15754 41916
rect 15778 41914 15834 41916
rect 15858 41914 15914 41916
rect 15618 41862 15664 41914
rect 15664 41862 15674 41914
rect 15698 41862 15728 41914
rect 15728 41862 15740 41914
rect 15740 41862 15754 41914
rect 15778 41862 15792 41914
rect 15792 41862 15804 41914
rect 15804 41862 15834 41914
rect 15858 41862 15868 41914
rect 15868 41862 15914 41914
rect 15618 41860 15674 41862
rect 15698 41860 15754 41862
rect 15778 41860 15834 41862
rect 15858 41860 15914 41862
rect 15618 40826 15674 40828
rect 15698 40826 15754 40828
rect 15778 40826 15834 40828
rect 15858 40826 15914 40828
rect 15618 40774 15664 40826
rect 15664 40774 15674 40826
rect 15698 40774 15728 40826
rect 15728 40774 15740 40826
rect 15740 40774 15754 40826
rect 15778 40774 15792 40826
rect 15792 40774 15804 40826
rect 15804 40774 15834 40826
rect 15858 40774 15868 40826
rect 15868 40774 15914 40826
rect 15618 40772 15674 40774
rect 15698 40772 15754 40774
rect 15778 40772 15834 40774
rect 15858 40772 15914 40774
rect 15618 39738 15674 39740
rect 15698 39738 15754 39740
rect 15778 39738 15834 39740
rect 15858 39738 15914 39740
rect 15618 39686 15664 39738
rect 15664 39686 15674 39738
rect 15698 39686 15728 39738
rect 15728 39686 15740 39738
rect 15740 39686 15754 39738
rect 15778 39686 15792 39738
rect 15792 39686 15804 39738
rect 15804 39686 15834 39738
rect 15858 39686 15868 39738
rect 15868 39686 15914 39738
rect 15618 39684 15674 39686
rect 15698 39684 15754 39686
rect 15778 39684 15834 39686
rect 15858 39684 15914 39686
rect 15198 38936 15254 38992
rect 15618 38650 15674 38652
rect 15698 38650 15754 38652
rect 15778 38650 15834 38652
rect 15858 38650 15914 38652
rect 15618 38598 15664 38650
rect 15664 38598 15674 38650
rect 15698 38598 15728 38650
rect 15728 38598 15740 38650
rect 15740 38598 15754 38650
rect 15778 38598 15792 38650
rect 15792 38598 15804 38650
rect 15804 38598 15834 38650
rect 15858 38598 15868 38650
rect 15868 38598 15914 38650
rect 15618 38596 15674 38598
rect 15698 38596 15754 38598
rect 15778 38596 15834 38598
rect 15858 38596 15914 38598
rect 14370 32816 14426 32872
rect 14278 32272 14334 32328
rect 13450 29008 13506 29064
rect 13450 22636 13506 22672
rect 13450 22616 13452 22636
rect 13452 22616 13504 22636
rect 13504 22616 13506 22636
rect 13542 20712 13598 20768
rect 13174 19624 13230 19680
rect 12685 18522 12741 18524
rect 12765 18522 12821 18524
rect 12845 18522 12901 18524
rect 12925 18522 12981 18524
rect 12685 18470 12731 18522
rect 12731 18470 12741 18522
rect 12765 18470 12795 18522
rect 12795 18470 12807 18522
rect 12807 18470 12821 18522
rect 12845 18470 12859 18522
rect 12859 18470 12871 18522
rect 12871 18470 12901 18522
rect 12925 18470 12935 18522
rect 12935 18470 12981 18522
rect 12685 18468 12741 18470
rect 12765 18468 12821 18470
rect 12845 18468 12901 18470
rect 12925 18468 12981 18470
rect 12685 17434 12741 17436
rect 12765 17434 12821 17436
rect 12845 17434 12901 17436
rect 12925 17434 12981 17436
rect 12685 17382 12731 17434
rect 12731 17382 12741 17434
rect 12765 17382 12795 17434
rect 12795 17382 12807 17434
rect 12807 17382 12821 17434
rect 12845 17382 12859 17434
rect 12859 17382 12871 17434
rect 12871 17382 12901 17434
rect 12925 17382 12935 17434
rect 12935 17382 12981 17434
rect 12685 17380 12741 17382
rect 12765 17380 12821 17382
rect 12845 17380 12901 17382
rect 12925 17380 12981 17382
rect 12685 16346 12741 16348
rect 12765 16346 12821 16348
rect 12845 16346 12901 16348
rect 12925 16346 12981 16348
rect 12685 16294 12731 16346
rect 12731 16294 12741 16346
rect 12765 16294 12795 16346
rect 12795 16294 12807 16346
rect 12807 16294 12821 16346
rect 12845 16294 12859 16346
rect 12859 16294 12871 16346
rect 12871 16294 12901 16346
rect 12925 16294 12935 16346
rect 12935 16294 12981 16346
rect 12685 16292 12741 16294
rect 12765 16292 12821 16294
rect 12845 16292 12901 16294
rect 12925 16292 12981 16294
rect 11242 9016 11298 9072
rect 11150 8880 11206 8936
rect 11978 11872 12034 11928
rect 12530 15408 12586 15464
rect 12346 13912 12402 13968
rect 12438 13776 12494 13832
rect 13174 15952 13230 16008
rect 12685 15258 12741 15260
rect 12765 15258 12821 15260
rect 12845 15258 12901 15260
rect 12925 15258 12981 15260
rect 12685 15206 12731 15258
rect 12731 15206 12741 15258
rect 12765 15206 12795 15258
rect 12795 15206 12807 15258
rect 12807 15206 12821 15258
rect 12845 15206 12859 15258
rect 12859 15206 12871 15258
rect 12871 15206 12901 15258
rect 12925 15206 12935 15258
rect 12935 15206 12981 15258
rect 12685 15204 12741 15206
rect 12765 15204 12821 15206
rect 12845 15204 12901 15206
rect 12925 15204 12981 15206
rect 12685 14170 12741 14172
rect 12765 14170 12821 14172
rect 12845 14170 12901 14172
rect 12925 14170 12981 14172
rect 12685 14118 12731 14170
rect 12731 14118 12741 14170
rect 12765 14118 12795 14170
rect 12795 14118 12807 14170
rect 12807 14118 12821 14170
rect 12845 14118 12859 14170
rect 12859 14118 12871 14170
rect 12871 14118 12901 14170
rect 12925 14118 12935 14170
rect 12935 14118 12981 14170
rect 12685 14116 12741 14118
rect 12765 14116 12821 14118
rect 12845 14116 12901 14118
rect 12925 14116 12981 14118
rect 12685 13082 12741 13084
rect 12765 13082 12821 13084
rect 12845 13082 12901 13084
rect 12925 13082 12981 13084
rect 12685 13030 12731 13082
rect 12731 13030 12741 13082
rect 12765 13030 12795 13082
rect 12795 13030 12807 13082
rect 12807 13030 12821 13082
rect 12845 13030 12859 13082
rect 12859 13030 12871 13082
rect 12871 13030 12901 13082
rect 12925 13030 12935 13082
rect 12935 13030 12981 13082
rect 12685 13028 12741 13030
rect 12765 13028 12821 13030
rect 12845 13028 12901 13030
rect 12925 13028 12981 13030
rect 13358 19352 13414 19408
rect 13358 16632 13414 16688
rect 12438 11736 12494 11792
rect 12685 11994 12741 11996
rect 12765 11994 12821 11996
rect 12845 11994 12901 11996
rect 12925 11994 12981 11996
rect 12685 11942 12731 11994
rect 12731 11942 12741 11994
rect 12765 11942 12795 11994
rect 12795 11942 12807 11994
rect 12807 11942 12821 11994
rect 12845 11942 12859 11994
rect 12859 11942 12871 11994
rect 12871 11942 12901 11994
rect 12925 11942 12935 11994
rect 12935 11942 12981 11994
rect 12685 11940 12741 11942
rect 12765 11940 12821 11942
rect 12845 11940 12901 11942
rect 12925 11940 12981 11942
rect 12346 11192 12402 11248
rect 11794 9832 11850 9888
rect 11610 5480 11666 5536
rect 11426 4936 11482 4992
rect 11150 4528 11206 4584
rect 10230 2488 10286 2544
rect 9954 1828 10010 1864
rect 9954 1808 9956 1828
rect 9956 1808 10008 1828
rect 10008 1808 10010 1828
rect 10230 1672 10286 1728
rect 9753 1658 9809 1660
rect 9833 1658 9889 1660
rect 9913 1658 9969 1660
rect 9993 1658 10049 1660
rect 9753 1606 9799 1658
rect 9799 1606 9809 1658
rect 9833 1606 9863 1658
rect 9863 1606 9875 1658
rect 9875 1606 9889 1658
rect 9913 1606 9927 1658
rect 9927 1606 9939 1658
rect 9939 1606 9969 1658
rect 9993 1606 10003 1658
rect 10003 1606 10049 1658
rect 9753 1604 9809 1606
rect 9833 1604 9889 1606
rect 9913 1604 9969 1606
rect 9993 1604 10049 1606
rect 9632 1264 9688 1320
rect 10046 1264 10102 1320
rect 11334 4528 11390 4584
rect 10874 3984 10930 4040
rect 11242 2352 11298 2408
rect 11150 2216 11206 2272
rect 11610 3984 11666 4040
rect 11794 2896 11850 2952
rect 12162 9560 12218 9616
rect 12162 3304 12218 3360
rect 12685 10906 12741 10908
rect 12765 10906 12821 10908
rect 12845 10906 12901 10908
rect 12925 10906 12981 10908
rect 12685 10854 12731 10906
rect 12731 10854 12741 10906
rect 12765 10854 12795 10906
rect 12795 10854 12807 10906
rect 12807 10854 12821 10906
rect 12845 10854 12859 10906
rect 12859 10854 12871 10906
rect 12871 10854 12901 10906
rect 12925 10854 12935 10906
rect 12935 10854 12981 10906
rect 12685 10852 12741 10854
rect 12765 10852 12821 10854
rect 12845 10852 12901 10854
rect 12925 10852 12981 10854
rect 12685 9818 12741 9820
rect 12765 9818 12821 9820
rect 12845 9818 12901 9820
rect 12925 9818 12981 9820
rect 12685 9766 12731 9818
rect 12731 9766 12741 9818
rect 12765 9766 12795 9818
rect 12795 9766 12807 9818
rect 12807 9766 12821 9818
rect 12845 9766 12859 9818
rect 12859 9766 12871 9818
rect 12871 9766 12901 9818
rect 12925 9766 12935 9818
rect 12935 9766 12981 9818
rect 12685 9764 12741 9766
rect 12765 9764 12821 9766
rect 12845 9764 12901 9766
rect 12925 9764 12981 9766
rect 12685 8730 12741 8732
rect 12765 8730 12821 8732
rect 12845 8730 12901 8732
rect 12925 8730 12981 8732
rect 12685 8678 12731 8730
rect 12731 8678 12741 8730
rect 12765 8678 12795 8730
rect 12795 8678 12807 8730
rect 12807 8678 12821 8730
rect 12845 8678 12859 8730
rect 12859 8678 12871 8730
rect 12871 8678 12901 8730
rect 12925 8678 12935 8730
rect 12935 8678 12981 8730
rect 12685 8676 12741 8678
rect 12765 8676 12821 8678
rect 12845 8676 12901 8678
rect 12925 8676 12981 8678
rect 12438 6568 12494 6624
rect 12685 7642 12741 7644
rect 12765 7642 12821 7644
rect 12845 7642 12901 7644
rect 12925 7642 12981 7644
rect 12685 7590 12731 7642
rect 12731 7590 12741 7642
rect 12765 7590 12795 7642
rect 12795 7590 12807 7642
rect 12807 7590 12821 7642
rect 12845 7590 12859 7642
rect 12859 7590 12871 7642
rect 12871 7590 12901 7642
rect 12925 7590 12935 7642
rect 12935 7590 12981 7642
rect 12685 7588 12741 7590
rect 12765 7588 12821 7590
rect 12845 7588 12901 7590
rect 12925 7588 12981 7590
rect 12806 6740 12808 6760
rect 12808 6740 12860 6760
rect 12860 6740 12862 6760
rect 12806 6704 12862 6740
rect 12685 6554 12741 6556
rect 12765 6554 12821 6556
rect 12845 6554 12901 6556
rect 12925 6554 12981 6556
rect 12685 6502 12731 6554
rect 12731 6502 12741 6554
rect 12765 6502 12795 6554
rect 12795 6502 12807 6554
rect 12807 6502 12821 6554
rect 12845 6502 12859 6554
rect 12859 6502 12871 6554
rect 12871 6502 12901 6554
rect 12925 6502 12935 6554
rect 12935 6502 12981 6554
rect 12685 6500 12741 6502
rect 12765 6500 12821 6502
rect 12845 6500 12901 6502
rect 12925 6500 12981 6502
rect 12685 5466 12741 5468
rect 12765 5466 12821 5468
rect 12845 5466 12901 5468
rect 12925 5466 12981 5468
rect 12685 5414 12731 5466
rect 12731 5414 12741 5466
rect 12765 5414 12795 5466
rect 12795 5414 12807 5466
rect 12807 5414 12821 5466
rect 12845 5414 12859 5466
rect 12859 5414 12871 5466
rect 12871 5414 12901 5466
rect 12925 5414 12935 5466
rect 12935 5414 12981 5466
rect 12685 5412 12741 5414
rect 12765 5412 12821 5414
rect 12845 5412 12901 5414
rect 12925 5412 12981 5414
rect 12685 4378 12741 4380
rect 12765 4378 12821 4380
rect 12845 4378 12901 4380
rect 12925 4378 12981 4380
rect 12685 4326 12731 4378
rect 12731 4326 12741 4378
rect 12765 4326 12795 4378
rect 12795 4326 12807 4378
rect 12807 4326 12821 4378
rect 12845 4326 12859 4378
rect 12859 4326 12871 4378
rect 12871 4326 12901 4378
rect 12925 4326 12935 4378
rect 12935 4326 12981 4378
rect 12685 4324 12741 4326
rect 12765 4324 12821 4326
rect 12845 4324 12901 4326
rect 12925 4324 12981 4326
rect 12990 4120 13046 4176
rect 12685 3290 12741 3292
rect 12765 3290 12821 3292
rect 12845 3290 12901 3292
rect 12925 3290 12981 3292
rect 12685 3238 12731 3290
rect 12731 3238 12741 3290
rect 12765 3238 12795 3290
rect 12795 3238 12807 3290
rect 12807 3238 12821 3290
rect 12845 3238 12859 3290
rect 12859 3238 12871 3290
rect 12871 3238 12901 3290
rect 12925 3238 12935 3290
rect 12935 3238 12981 3290
rect 12685 3236 12741 3238
rect 12765 3236 12821 3238
rect 12845 3236 12901 3238
rect 12925 3236 12981 3238
rect 12530 3168 12586 3224
rect 11794 2624 11850 2680
rect 11886 2352 11942 2408
rect 11518 1672 11574 1728
rect 11978 2216 12034 2272
rect 11058 1400 11114 1456
rect 11058 1300 11060 1320
rect 11060 1300 11112 1320
rect 11112 1300 11114 1320
rect 11058 1264 11114 1300
rect 11518 1164 11520 1184
rect 11520 1164 11572 1184
rect 11572 1164 11574 1184
rect 11518 1128 11574 1164
rect 14094 31220 14096 31240
rect 14096 31220 14148 31240
rect 14148 31220 14150 31240
rect 14094 31184 14150 31220
rect 14646 29688 14702 29744
rect 14646 29008 14702 29064
rect 14094 27412 14096 27432
rect 14096 27412 14148 27432
rect 14148 27412 14150 27432
rect 14094 27376 14150 27412
rect 14002 25200 14058 25256
rect 13818 20304 13874 20360
rect 13910 19760 13966 19816
rect 13818 17176 13874 17232
rect 14186 26560 14242 26616
rect 14186 21528 14242 21584
rect 14186 20576 14242 20632
rect 13910 15136 13966 15192
rect 13542 12144 13598 12200
rect 14554 27376 14610 27432
rect 15014 32952 15070 33008
rect 15618 37562 15674 37564
rect 15698 37562 15754 37564
rect 15778 37562 15834 37564
rect 15858 37562 15914 37564
rect 15618 37510 15664 37562
rect 15664 37510 15674 37562
rect 15698 37510 15728 37562
rect 15728 37510 15740 37562
rect 15740 37510 15754 37562
rect 15778 37510 15792 37562
rect 15792 37510 15804 37562
rect 15804 37510 15834 37562
rect 15858 37510 15868 37562
rect 15868 37510 15914 37562
rect 15618 37508 15674 37510
rect 15698 37508 15754 37510
rect 15778 37508 15834 37510
rect 15858 37508 15914 37510
rect 15618 36474 15674 36476
rect 15698 36474 15754 36476
rect 15778 36474 15834 36476
rect 15858 36474 15914 36476
rect 15618 36422 15664 36474
rect 15664 36422 15674 36474
rect 15698 36422 15728 36474
rect 15728 36422 15740 36474
rect 15740 36422 15754 36474
rect 15778 36422 15792 36474
rect 15792 36422 15804 36474
rect 15804 36422 15834 36474
rect 15858 36422 15868 36474
rect 15868 36422 15914 36474
rect 15618 36420 15674 36422
rect 15698 36420 15754 36422
rect 15778 36420 15834 36422
rect 15858 36420 15914 36422
rect 15618 35386 15674 35388
rect 15698 35386 15754 35388
rect 15778 35386 15834 35388
rect 15858 35386 15914 35388
rect 15618 35334 15664 35386
rect 15664 35334 15674 35386
rect 15698 35334 15728 35386
rect 15728 35334 15740 35386
rect 15740 35334 15754 35386
rect 15778 35334 15792 35386
rect 15792 35334 15804 35386
rect 15804 35334 15834 35386
rect 15858 35334 15868 35386
rect 15868 35334 15914 35386
rect 15618 35332 15674 35334
rect 15698 35332 15754 35334
rect 15778 35332 15834 35334
rect 15858 35332 15914 35334
rect 15618 34298 15674 34300
rect 15698 34298 15754 34300
rect 15778 34298 15834 34300
rect 15858 34298 15914 34300
rect 15618 34246 15664 34298
rect 15664 34246 15674 34298
rect 15698 34246 15728 34298
rect 15728 34246 15740 34298
rect 15740 34246 15754 34298
rect 15778 34246 15792 34298
rect 15792 34246 15804 34298
rect 15804 34246 15834 34298
rect 15858 34246 15868 34298
rect 15868 34246 15914 34298
rect 15618 34244 15674 34246
rect 15698 34244 15754 34246
rect 15778 34244 15834 34246
rect 15858 34244 15914 34246
rect 15290 32852 15292 32872
rect 15292 32852 15344 32872
rect 15344 32852 15346 32872
rect 15290 32816 15346 32852
rect 15106 32408 15162 32464
rect 15014 29008 15070 29064
rect 15618 33210 15674 33212
rect 15698 33210 15754 33212
rect 15778 33210 15834 33212
rect 15858 33210 15914 33212
rect 15618 33158 15664 33210
rect 15664 33158 15674 33210
rect 15698 33158 15728 33210
rect 15728 33158 15740 33210
rect 15740 33158 15754 33210
rect 15778 33158 15792 33210
rect 15792 33158 15804 33210
rect 15804 33158 15834 33210
rect 15858 33158 15868 33210
rect 15868 33158 15914 33210
rect 15618 33156 15674 33158
rect 15698 33156 15754 33158
rect 15778 33156 15834 33158
rect 15858 33156 15914 33158
rect 15842 32972 15898 33008
rect 15842 32952 15844 32972
rect 15844 32952 15896 32972
rect 15896 32952 15898 32972
rect 15618 32122 15674 32124
rect 15698 32122 15754 32124
rect 15778 32122 15834 32124
rect 15858 32122 15914 32124
rect 15618 32070 15664 32122
rect 15664 32070 15674 32122
rect 15698 32070 15728 32122
rect 15728 32070 15740 32122
rect 15740 32070 15754 32122
rect 15778 32070 15792 32122
rect 15792 32070 15804 32122
rect 15804 32070 15834 32122
rect 15858 32070 15868 32122
rect 15868 32070 15914 32122
rect 15618 32068 15674 32070
rect 15698 32068 15754 32070
rect 15778 32068 15834 32070
rect 15858 32068 15914 32070
rect 15618 31034 15674 31036
rect 15698 31034 15754 31036
rect 15778 31034 15834 31036
rect 15858 31034 15914 31036
rect 15618 30982 15664 31034
rect 15664 30982 15674 31034
rect 15698 30982 15728 31034
rect 15728 30982 15740 31034
rect 15740 30982 15754 31034
rect 15778 30982 15792 31034
rect 15792 30982 15804 31034
rect 15804 30982 15834 31034
rect 15858 30982 15868 31034
rect 15868 30982 15914 31034
rect 15618 30980 15674 30982
rect 15698 30980 15754 30982
rect 15778 30980 15834 30982
rect 15858 30980 15914 30982
rect 15618 29946 15674 29948
rect 15698 29946 15754 29948
rect 15778 29946 15834 29948
rect 15858 29946 15914 29948
rect 15618 29894 15664 29946
rect 15664 29894 15674 29946
rect 15698 29894 15728 29946
rect 15728 29894 15740 29946
rect 15740 29894 15754 29946
rect 15778 29894 15792 29946
rect 15792 29894 15804 29946
rect 15804 29894 15834 29946
rect 15858 29894 15868 29946
rect 15868 29894 15914 29946
rect 15618 29892 15674 29894
rect 15698 29892 15754 29894
rect 15778 29892 15834 29894
rect 15858 29892 15914 29894
rect 15658 29688 15714 29744
rect 15934 29280 15990 29336
rect 15618 28858 15674 28860
rect 15698 28858 15754 28860
rect 15778 28858 15834 28860
rect 15858 28858 15914 28860
rect 15618 28806 15664 28858
rect 15664 28806 15674 28858
rect 15698 28806 15728 28858
rect 15728 28806 15740 28858
rect 15740 28806 15754 28858
rect 15778 28806 15792 28858
rect 15792 28806 15804 28858
rect 15804 28806 15834 28858
rect 15858 28806 15868 28858
rect 15868 28806 15914 28858
rect 15618 28804 15674 28806
rect 15698 28804 15754 28806
rect 15778 28804 15834 28806
rect 15858 28804 15914 28806
rect 15198 26968 15254 27024
rect 14554 24520 14610 24576
rect 14462 22616 14518 22672
rect 15618 27770 15674 27772
rect 15698 27770 15754 27772
rect 15778 27770 15834 27772
rect 15858 27770 15914 27772
rect 15618 27718 15664 27770
rect 15664 27718 15674 27770
rect 15698 27718 15728 27770
rect 15728 27718 15740 27770
rect 15740 27718 15754 27770
rect 15778 27718 15792 27770
rect 15792 27718 15804 27770
rect 15804 27718 15834 27770
rect 15858 27718 15868 27770
rect 15868 27718 15914 27770
rect 15618 27716 15674 27718
rect 15698 27716 15754 27718
rect 15778 27716 15834 27718
rect 15858 27716 15914 27718
rect 15618 26682 15674 26684
rect 15698 26682 15754 26684
rect 15778 26682 15834 26684
rect 15858 26682 15914 26684
rect 15618 26630 15664 26682
rect 15664 26630 15674 26682
rect 15698 26630 15728 26682
rect 15728 26630 15740 26682
rect 15740 26630 15754 26682
rect 15778 26630 15792 26682
rect 15792 26630 15804 26682
rect 15804 26630 15834 26682
rect 15858 26630 15868 26682
rect 15868 26630 15914 26682
rect 15618 26628 15674 26630
rect 15698 26628 15754 26630
rect 15778 26628 15834 26630
rect 15858 26628 15914 26630
rect 15618 25594 15674 25596
rect 15698 25594 15754 25596
rect 15778 25594 15834 25596
rect 15858 25594 15914 25596
rect 15618 25542 15664 25594
rect 15664 25542 15674 25594
rect 15698 25542 15728 25594
rect 15728 25542 15740 25594
rect 15740 25542 15754 25594
rect 15778 25542 15792 25594
rect 15792 25542 15804 25594
rect 15804 25542 15834 25594
rect 15858 25542 15868 25594
rect 15868 25542 15914 25594
rect 15618 25540 15674 25542
rect 15698 25540 15754 25542
rect 15778 25540 15834 25542
rect 15858 25540 15914 25542
rect 14554 21392 14610 21448
rect 14278 19352 14334 19408
rect 14738 17720 14794 17776
rect 13726 11056 13782 11112
rect 14002 11192 14058 11248
rect 13358 6316 13414 6352
rect 13358 6296 13360 6316
rect 13360 6296 13412 6316
rect 13412 6296 13414 6316
rect 14278 11736 14334 11792
rect 15198 19488 15254 19544
rect 15618 24506 15674 24508
rect 15698 24506 15754 24508
rect 15778 24506 15834 24508
rect 15858 24506 15914 24508
rect 15618 24454 15664 24506
rect 15664 24454 15674 24506
rect 15698 24454 15728 24506
rect 15728 24454 15740 24506
rect 15740 24454 15754 24506
rect 15778 24454 15792 24506
rect 15792 24454 15804 24506
rect 15804 24454 15834 24506
rect 15858 24454 15868 24506
rect 15868 24454 15914 24506
rect 15618 24452 15674 24454
rect 15698 24452 15754 24454
rect 15778 24452 15834 24454
rect 15858 24452 15914 24454
rect 15618 23418 15674 23420
rect 15698 23418 15754 23420
rect 15778 23418 15834 23420
rect 15858 23418 15914 23420
rect 15618 23366 15664 23418
rect 15664 23366 15674 23418
rect 15698 23366 15728 23418
rect 15728 23366 15740 23418
rect 15740 23366 15754 23418
rect 15778 23366 15792 23418
rect 15792 23366 15804 23418
rect 15804 23366 15834 23418
rect 15858 23366 15868 23418
rect 15868 23366 15914 23418
rect 15618 23364 15674 23366
rect 15698 23364 15754 23366
rect 15778 23364 15834 23366
rect 15858 23364 15914 23366
rect 15618 22330 15674 22332
rect 15698 22330 15754 22332
rect 15778 22330 15834 22332
rect 15858 22330 15914 22332
rect 15618 22278 15664 22330
rect 15664 22278 15674 22330
rect 15698 22278 15728 22330
rect 15728 22278 15740 22330
rect 15740 22278 15754 22330
rect 15778 22278 15792 22330
rect 15792 22278 15804 22330
rect 15804 22278 15834 22330
rect 15858 22278 15868 22330
rect 15868 22278 15914 22330
rect 15618 22276 15674 22278
rect 15698 22276 15754 22278
rect 15778 22276 15834 22278
rect 15858 22276 15914 22278
rect 15618 21242 15674 21244
rect 15698 21242 15754 21244
rect 15778 21242 15834 21244
rect 15858 21242 15914 21244
rect 15618 21190 15664 21242
rect 15664 21190 15674 21242
rect 15698 21190 15728 21242
rect 15728 21190 15740 21242
rect 15740 21190 15754 21242
rect 15778 21190 15792 21242
rect 15792 21190 15804 21242
rect 15804 21190 15834 21242
rect 15858 21190 15868 21242
rect 15868 21190 15914 21242
rect 15618 21188 15674 21190
rect 15698 21188 15754 21190
rect 15778 21188 15834 21190
rect 15858 21188 15914 21190
rect 15618 20154 15674 20156
rect 15698 20154 15754 20156
rect 15778 20154 15834 20156
rect 15858 20154 15914 20156
rect 15618 20102 15664 20154
rect 15664 20102 15674 20154
rect 15698 20102 15728 20154
rect 15728 20102 15740 20154
rect 15740 20102 15754 20154
rect 15778 20102 15792 20154
rect 15792 20102 15804 20154
rect 15804 20102 15834 20154
rect 15858 20102 15868 20154
rect 15868 20102 15914 20154
rect 15618 20100 15674 20102
rect 15698 20100 15754 20102
rect 15778 20100 15834 20102
rect 15858 20100 15914 20102
rect 15618 19066 15674 19068
rect 15698 19066 15754 19068
rect 15778 19066 15834 19068
rect 15858 19066 15914 19068
rect 15618 19014 15664 19066
rect 15664 19014 15674 19066
rect 15698 19014 15728 19066
rect 15728 19014 15740 19066
rect 15740 19014 15754 19066
rect 15778 19014 15792 19066
rect 15792 19014 15804 19066
rect 15804 19014 15834 19066
rect 15858 19014 15868 19066
rect 15868 19014 15914 19066
rect 15618 19012 15674 19014
rect 15698 19012 15754 19014
rect 15778 19012 15834 19014
rect 15858 19012 15914 19014
rect 15618 17978 15674 17980
rect 15698 17978 15754 17980
rect 15778 17978 15834 17980
rect 15858 17978 15914 17980
rect 15618 17926 15664 17978
rect 15664 17926 15674 17978
rect 15698 17926 15728 17978
rect 15728 17926 15740 17978
rect 15740 17926 15754 17978
rect 15778 17926 15792 17978
rect 15792 17926 15804 17978
rect 15804 17926 15834 17978
rect 15858 17926 15868 17978
rect 15868 17926 15914 17978
rect 15618 17924 15674 17926
rect 15698 17924 15754 17926
rect 15778 17924 15834 17926
rect 15858 17924 15914 17926
rect 14738 15428 14794 15464
rect 14738 15408 14740 15428
rect 14740 15408 14792 15428
rect 14792 15408 14794 15428
rect 14738 10104 14794 10160
rect 12254 2080 12310 2136
rect 12685 2202 12741 2204
rect 12765 2202 12821 2204
rect 12845 2202 12901 2204
rect 12925 2202 12981 2204
rect 12685 2150 12731 2202
rect 12731 2150 12741 2202
rect 12765 2150 12795 2202
rect 12795 2150 12807 2202
rect 12807 2150 12821 2202
rect 12845 2150 12859 2202
rect 12859 2150 12871 2202
rect 12871 2150 12901 2202
rect 12925 2150 12935 2202
rect 12935 2150 12981 2202
rect 12685 2148 12741 2150
rect 12765 2148 12821 2150
rect 12845 2148 12901 2150
rect 12925 2148 12981 2150
rect 13634 4936 13690 4992
rect 14370 9968 14426 10024
rect 14646 9968 14702 10024
rect 14554 9696 14610 9752
rect 14370 8336 14426 8392
rect 13910 2508 13966 2544
rect 13910 2488 13912 2508
rect 13912 2488 13964 2508
rect 13964 2488 13966 2508
rect 13082 1808 13138 1864
rect 12714 1300 12716 1320
rect 12716 1300 12768 1320
rect 12768 1300 12770 1320
rect 12714 1264 12770 1300
rect 13450 1300 13452 1320
rect 13452 1300 13504 1320
rect 13504 1300 13506 1320
rect 13450 1264 13506 1300
rect 12685 1114 12741 1116
rect 12765 1114 12821 1116
rect 12845 1114 12901 1116
rect 12925 1114 12981 1116
rect 12685 1062 12731 1114
rect 12731 1062 12741 1114
rect 12765 1062 12795 1114
rect 12795 1062 12807 1114
rect 12807 1062 12821 1114
rect 12845 1062 12859 1114
rect 12859 1062 12871 1114
rect 12871 1062 12901 1114
rect 12925 1062 12935 1114
rect 12935 1062 12981 1114
rect 12685 1060 12741 1062
rect 12765 1060 12821 1062
rect 12845 1060 12901 1062
rect 12925 1060 12981 1062
rect 14094 1300 14096 1320
rect 14096 1300 14148 1320
rect 14148 1300 14150 1320
rect 14094 1264 14150 1300
rect 15290 16108 15346 16144
rect 15290 16088 15292 16108
rect 15292 16088 15344 16108
rect 15344 16088 15346 16108
rect 15198 10104 15254 10160
rect 15618 16890 15674 16892
rect 15698 16890 15754 16892
rect 15778 16890 15834 16892
rect 15858 16890 15914 16892
rect 15618 16838 15664 16890
rect 15664 16838 15674 16890
rect 15698 16838 15728 16890
rect 15728 16838 15740 16890
rect 15740 16838 15754 16890
rect 15778 16838 15792 16890
rect 15792 16838 15804 16890
rect 15804 16838 15834 16890
rect 15858 16838 15868 16890
rect 15868 16838 15914 16890
rect 15618 16836 15674 16838
rect 15698 16836 15754 16838
rect 15778 16836 15834 16838
rect 15858 16836 15914 16838
rect 15618 15802 15674 15804
rect 15698 15802 15754 15804
rect 15778 15802 15834 15804
rect 15858 15802 15914 15804
rect 15618 15750 15664 15802
rect 15664 15750 15674 15802
rect 15698 15750 15728 15802
rect 15728 15750 15740 15802
rect 15740 15750 15754 15802
rect 15778 15750 15792 15802
rect 15792 15750 15804 15802
rect 15804 15750 15834 15802
rect 15858 15750 15868 15802
rect 15868 15750 15914 15802
rect 15618 15748 15674 15750
rect 15698 15748 15754 15750
rect 15778 15748 15834 15750
rect 15858 15748 15914 15750
rect 18550 43546 18606 43548
rect 18630 43546 18686 43548
rect 18710 43546 18766 43548
rect 18790 43546 18846 43548
rect 18550 43494 18596 43546
rect 18596 43494 18606 43546
rect 18630 43494 18660 43546
rect 18660 43494 18672 43546
rect 18672 43494 18686 43546
rect 18710 43494 18724 43546
rect 18724 43494 18736 43546
rect 18736 43494 18766 43546
rect 18790 43494 18800 43546
rect 18800 43494 18846 43546
rect 18550 43492 18606 43494
rect 18630 43492 18686 43494
rect 18710 43492 18766 43494
rect 18790 43492 18846 43494
rect 17590 42880 17646 42936
rect 18326 42644 18328 42664
rect 18328 42644 18380 42664
rect 18380 42644 18382 42664
rect 18326 42608 18382 42644
rect 16762 33904 16818 33960
rect 16762 32272 16818 32328
rect 16578 31864 16634 31920
rect 16486 29008 16542 29064
rect 16486 28056 16542 28112
rect 15618 14714 15674 14716
rect 15698 14714 15754 14716
rect 15778 14714 15834 14716
rect 15858 14714 15914 14716
rect 15618 14662 15664 14714
rect 15664 14662 15674 14714
rect 15698 14662 15728 14714
rect 15728 14662 15740 14714
rect 15740 14662 15754 14714
rect 15778 14662 15792 14714
rect 15792 14662 15804 14714
rect 15804 14662 15834 14714
rect 15858 14662 15868 14714
rect 15868 14662 15914 14714
rect 15618 14660 15674 14662
rect 15698 14660 15754 14662
rect 15778 14660 15834 14662
rect 15858 14660 15914 14662
rect 15106 9052 15108 9072
rect 15108 9052 15160 9072
rect 15160 9052 15162 9072
rect 15106 9016 15162 9052
rect 15618 13626 15674 13628
rect 15698 13626 15754 13628
rect 15778 13626 15834 13628
rect 15858 13626 15914 13628
rect 15618 13574 15664 13626
rect 15664 13574 15674 13626
rect 15698 13574 15728 13626
rect 15728 13574 15740 13626
rect 15740 13574 15754 13626
rect 15778 13574 15792 13626
rect 15792 13574 15804 13626
rect 15804 13574 15834 13626
rect 15858 13574 15868 13626
rect 15868 13574 15914 13626
rect 15618 13572 15674 13574
rect 15698 13572 15754 13574
rect 15778 13572 15834 13574
rect 15858 13572 15914 13574
rect 16670 29708 16726 29744
rect 16670 29688 16672 29708
rect 16672 29688 16724 29708
rect 16724 29688 16726 29708
rect 16670 29416 16726 29472
rect 16762 29280 16818 29336
rect 16578 25744 16634 25800
rect 16210 14456 16266 14512
rect 15618 12538 15674 12540
rect 15698 12538 15754 12540
rect 15778 12538 15834 12540
rect 15858 12538 15914 12540
rect 15618 12486 15664 12538
rect 15664 12486 15674 12538
rect 15698 12486 15728 12538
rect 15728 12486 15740 12538
rect 15740 12486 15754 12538
rect 15778 12486 15792 12538
rect 15792 12486 15804 12538
rect 15804 12486 15834 12538
rect 15858 12486 15868 12538
rect 15868 12486 15914 12538
rect 15618 12484 15674 12486
rect 15698 12484 15754 12486
rect 15778 12484 15834 12486
rect 15858 12484 15914 12486
rect 15658 12044 15660 12064
rect 15660 12044 15712 12064
rect 15712 12044 15714 12064
rect 15658 12008 15714 12044
rect 15618 11450 15674 11452
rect 15698 11450 15754 11452
rect 15778 11450 15834 11452
rect 15858 11450 15914 11452
rect 15618 11398 15664 11450
rect 15664 11398 15674 11450
rect 15698 11398 15728 11450
rect 15728 11398 15740 11450
rect 15740 11398 15754 11450
rect 15778 11398 15792 11450
rect 15792 11398 15804 11450
rect 15804 11398 15834 11450
rect 15858 11398 15868 11450
rect 15868 11398 15914 11450
rect 15618 11396 15674 11398
rect 15698 11396 15754 11398
rect 15778 11396 15834 11398
rect 15858 11396 15914 11398
rect 15618 10362 15674 10364
rect 15698 10362 15754 10364
rect 15778 10362 15834 10364
rect 15858 10362 15914 10364
rect 15618 10310 15664 10362
rect 15664 10310 15674 10362
rect 15698 10310 15728 10362
rect 15728 10310 15740 10362
rect 15740 10310 15754 10362
rect 15778 10310 15792 10362
rect 15792 10310 15804 10362
rect 15804 10310 15834 10362
rect 15858 10310 15868 10362
rect 15868 10310 15914 10362
rect 15618 10308 15674 10310
rect 15698 10308 15754 10310
rect 15778 10308 15834 10310
rect 15858 10308 15914 10310
rect 15750 9968 15806 10024
rect 15842 9696 15898 9752
rect 15618 9274 15674 9276
rect 15698 9274 15754 9276
rect 15778 9274 15834 9276
rect 15858 9274 15914 9276
rect 15618 9222 15664 9274
rect 15664 9222 15674 9274
rect 15698 9222 15728 9274
rect 15728 9222 15740 9274
rect 15740 9222 15754 9274
rect 15778 9222 15792 9274
rect 15792 9222 15804 9274
rect 15804 9222 15834 9274
rect 15858 9222 15868 9274
rect 15868 9222 15914 9274
rect 15618 9220 15674 9222
rect 15698 9220 15754 9222
rect 15778 9220 15834 9222
rect 15858 9220 15914 9222
rect 14922 4936 14978 4992
rect 14462 2100 14518 2136
rect 14462 2080 14464 2100
rect 14464 2080 14516 2100
rect 14516 2080 14518 2100
rect 14554 1300 14556 1320
rect 14556 1300 14608 1320
rect 14608 1300 14610 1320
rect 14554 1264 14610 1300
rect 15618 8186 15674 8188
rect 15698 8186 15754 8188
rect 15778 8186 15834 8188
rect 15858 8186 15914 8188
rect 15618 8134 15664 8186
rect 15664 8134 15674 8186
rect 15698 8134 15728 8186
rect 15728 8134 15740 8186
rect 15740 8134 15754 8186
rect 15778 8134 15792 8186
rect 15792 8134 15804 8186
rect 15804 8134 15834 8186
rect 15858 8134 15868 8186
rect 15868 8134 15914 8186
rect 15618 8132 15674 8134
rect 15698 8132 15754 8134
rect 15778 8132 15834 8134
rect 15858 8132 15914 8134
rect 15618 7098 15674 7100
rect 15698 7098 15754 7100
rect 15778 7098 15834 7100
rect 15858 7098 15914 7100
rect 15618 7046 15664 7098
rect 15664 7046 15674 7098
rect 15698 7046 15728 7098
rect 15728 7046 15740 7098
rect 15740 7046 15754 7098
rect 15778 7046 15792 7098
rect 15792 7046 15804 7098
rect 15804 7046 15834 7098
rect 15858 7046 15868 7098
rect 15868 7046 15914 7098
rect 15618 7044 15674 7046
rect 15698 7044 15754 7046
rect 15778 7044 15834 7046
rect 15858 7044 15914 7046
rect 16670 19352 16726 19408
rect 16486 17196 16542 17232
rect 16486 17176 16488 17196
rect 16488 17176 16540 17196
rect 16540 17176 16542 17196
rect 16578 17040 16634 17096
rect 15934 6840 15990 6896
rect 15618 6010 15674 6012
rect 15698 6010 15754 6012
rect 15778 6010 15834 6012
rect 15858 6010 15914 6012
rect 15618 5958 15664 6010
rect 15664 5958 15674 6010
rect 15698 5958 15728 6010
rect 15728 5958 15740 6010
rect 15740 5958 15754 6010
rect 15778 5958 15792 6010
rect 15792 5958 15804 6010
rect 15804 5958 15834 6010
rect 15858 5958 15868 6010
rect 15868 5958 15914 6010
rect 15618 5956 15674 5958
rect 15698 5956 15754 5958
rect 15778 5956 15834 5958
rect 15858 5956 15914 5958
rect 15618 4922 15674 4924
rect 15698 4922 15754 4924
rect 15778 4922 15834 4924
rect 15858 4922 15914 4924
rect 15618 4870 15664 4922
rect 15664 4870 15674 4922
rect 15698 4870 15728 4922
rect 15728 4870 15740 4922
rect 15740 4870 15754 4922
rect 15778 4870 15792 4922
rect 15792 4870 15804 4922
rect 15804 4870 15834 4922
rect 15858 4870 15868 4922
rect 15868 4870 15914 4922
rect 15618 4868 15674 4870
rect 15698 4868 15754 4870
rect 15778 4868 15834 4870
rect 15858 4868 15914 4870
rect 15618 3834 15674 3836
rect 15698 3834 15754 3836
rect 15778 3834 15834 3836
rect 15858 3834 15914 3836
rect 15618 3782 15664 3834
rect 15664 3782 15674 3834
rect 15698 3782 15728 3834
rect 15728 3782 15740 3834
rect 15740 3782 15754 3834
rect 15778 3782 15792 3834
rect 15792 3782 15804 3834
rect 15804 3782 15834 3834
rect 15858 3782 15868 3834
rect 15868 3782 15914 3834
rect 15618 3780 15674 3782
rect 15698 3780 15754 3782
rect 15778 3780 15834 3782
rect 15858 3780 15914 3782
rect 16026 3712 16082 3768
rect 16854 14456 16910 14512
rect 17038 10104 17094 10160
rect 17498 42064 17554 42120
rect 17958 41928 18014 41984
rect 18326 41928 18382 41984
rect 18550 42458 18606 42460
rect 18630 42458 18686 42460
rect 18710 42458 18766 42460
rect 18790 42458 18846 42460
rect 18550 42406 18596 42458
rect 18596 42406 18606 42458
rect 18630 42406 18660 42458
rect 18660 42406 18672 42458
rect 18672 42406 18686 42458
rect 18710 42406 18724 42458
rect 18724 42406 18736 42458
rect 18736 42406 18766 42458
rect 18790 42406 18800 42458
rect 18800 42406 18846 42458
rect 18550 42404 18606 42406
rect 18630 42404 18686 42406
rect 18710 42404 18766 42406
rect 18790 42404 18846 42406
rect 19430 42200 19486 42256
rect 17222 32952 17278 33008
rect 17590 29416 17646 29472
rect 18050 28600 18106 28656
rect 17498 19624 17554 19680
rect 18550 41370 18606 41372
rect 18630 41370 18686 41372
rect 18710 41370 18766 41372
rect 18790 41370 18846 41372
rect 18550 41318 18596 41370
rect 18596 41318 18606 41370
rect 18630 41318 18660 41370
rect 18660 41318 18672 41370
rect 18672 41318 18686 41370
rect 18710 41318 18724 41370
rect 18724 41318 18736 41370
rect 18736 41318 18766 41370
rect 18790 41318 18800 41370
rect 18800 41318 18846 41370
rect 18550 41316 18606 41318
rect 18630 41316 18686 41318
rect 18710 41316 18766 41318
rect 18790 41316 18846 41318
rect 18550 40282 18606 40284
rect 18630 40282 18686 40284
rect 18710 40282 18766 40284
rect 18790 40282 18846 40284
rect 18550 40230 18596 40282
rect 18596 40230 18606 40282
rect 18630 40230 18660 40282
rect 18660 40230 18672 40282
rect 18672 40230 18686 40282
rect 18710 40230 18724 40282
rect 18724 40230 18736 40282
rect 18736 40230 18766 40282
rect 18790 40230 18800 40282
rect 18800 40230 18846 40282
rect 18550 40228 18606 40230
rect 18630 40228 18686 40230
rect 18710 40228 18766 40230
rect 18790 40228 18846 40230
rect 18550 39194 18606 39196
rect 18630 39194 18686 39196
rect 18710 39194 18766 39196
rect 18790 39194 18846 39196
rect 18550 39142 18596 39194
rect 18596 39142 18606 39194
rect 18630 39142 18660 39194
rect 18660 39142 18672 39194
rect 18672 39142 18686 39194
rect 18710 39142 18724 39194
rect 18724 39142 18736 39194
rect 18736 39142 18766 39194
rect 18790 39142 18800 39194
rect 18800 39142 18846 39194
rect 18550 39140 18606 39142
rect 18630 39140 18686 39142
rect 18710 39140 18766 39142
rect 18790 39140 18846 39142
rect 18550 38106 18606 38108
rect 18630 38106 18686 38108
rect 18710 38106 18766 38108
rect 18790 38106 18846 38108
rect 18550 38054 18596 38106
rect 18596 38054 18606 38106
rect 18630 38054 18660 38106
rect 18660 38054 18672 38106
rect 18672 38054 18686 38106
rect 18710 38054 18724 38106
rect 18724 38054 18736 38106
rect 18736 38054 18766 38106
rect 18790 38054 18800 38106
rect 18800 38054 18846 38106
rect 18550 38052 18606 38054
rect 18630 38052 18686 38054
rect 18710 38052 18766 38054
rect 18790 38052 18846 38054
rect 18550 37018 18606 37020
rect 18630 37018 18686 37020
rect 18710 37018 18766 37020
rect 18790 37018 18846 37020
rect 18550 36966 18596 37018
rect 18596 36966 18606 37018
rect 18630 36966 18660 37018
rect 18660 36966 18672 37018
rect 18672 36966 18686 37018
rect 18710 36966 18724 37018
rect 18724 36966 18736 37018
rect 18736 36966 18766 37018
rect 18790 36966 18800 37018
rect 18800 36966 18846 37018
rect 18550 36964 18606 36966
rect 18630 36964 18686 36966
rect 18710 36964 18766 36966
rect 18790 36964 18846 36966
rect 18550 35930 18606 35932
rect 18630 35930 18686 35932
rect 18710 35930 18766 35932
rect 18790 35930 18846 35932
rect 18550 35878 18596 35930
rect 18596 35878 18606 35930
rect 18630 35878 18660 35930
rect 18660 35878 18672 35930
rect 18672 35878 18686 35930
rect 18710 35878 18724 35930
rect 18724 35878 18736 35930
rect 18736 35878 18766 35930
rect 18790 35878 18800 35930
rect 18800 35878 18846 35930
rect 18550 35876 18606 35878
rect 18630 35876 18686 35878
rect 18710 35876 18766 35878
rect 18790 35876 18846 35878
rect 18550 34842 18606 34844
rect 18630 34842 18686 34844
rect 18710 34842 18766 34844
rect 18790 34842 18846 34844
rect 18550 34790 18596 34842
rect 18596 34790 18606 34842
rect 18630 34790 18660 34842
rect 18660 34790 18672 34842
rect 18672 34790 18686 34842
rect 18710 34790 18724 34842
rect 18724 34790 18736 34842
rect 18736 34790 18766 34842
rect 18790 34790 18800 34842
rect 18800 34790 18846 34842
rect 18550 34788 18606 34790
rect 18630 34788 18686 34790
rect 18710 34788 18766 34790
rect 18790 34788 18846 34790
rect 19522 41928 19578 41984
rect 19614 41420 19616 41440
rect 19616 41420 19668 41440
rect 19668 41420 19670 41440
rect 19338 36080 19394 36136
rect 18550 33754 18606 33756
rect 18630 33754 18686 33756
rect 18710 33754 18766 33756
rect 18790 33754 18846 33756
rect 18550 33702 18596 33754
rect 18596 33702 18606 33754
rect 18630 33702 18660 33754
rect 18660 33702 18672 33754
rect 18672 33702 18686 33754
rect 18710 33702 18724 33754
rect 18724 33702 18736 33754
rect 18736 33702 18766 33754
rect 18790 33702 18800 33754
rect 18800 33702 18846 33754
rect 18550 33700 18606 33702
rect 18630 33700 18686 33702
rect 18710 33700 18766 33702
rect 18790 33700 18846 33702
rect 18550 32666 18606 32668
rect 18630 32666 18686 32668
rect 18710 32666 18766 32668
rect 18790 32666 18846 32668
rect 18550 32614 18596 32666
rect 18596 32614 18606 32666
rect 18630 32614 18660 32666
rect 18660 32614 18672 32666
rect 18672 32614 18686 32666
rect 18710 32614 18724 32666
rect 18724 32614 18736 32666
rect 18736 32614 18766 32666
rect 18790 32614 18800 32666
rect 18800 32614 18846 32666
rect 18550 32612 18606 32614
rect 18630 32612 18686 32614
rect 18710 32612 18766 32614
rect 18790 32612 18846 32614
rect 18786 31764 18788 31784
rect 18788 31764 18840 31784
rect 18840 31764 18842 31784
rect 18786 31728 18842 31764
rect 18550 31578 18606 31580
rect 18630 31578 18686 31580
rect 18710 31578 18766 31580
rect 18790 31578 18846 31580
rect 18550 31526 18596 31578
rect 18596 31526 18606 31578
rect 18630 31526 18660 31578
rect 18660 31526 18672 31578
rect 18672 31526 18686 31578
rect 18710 31526 18724 31578
rect 18724 31526 18736 31578
rect 18736 31526 18766 31578
rect 18790 31526 18800 31578
rect 18800 31526 18846 31578
rect 18550 31524 18606 31526
rect 18630 31524 18686 31526
rect 18710 31524 18766 31526
rect 18790 31524 18846 31526
rect 17774 19352 17830 19408
rect 17406 10648 17462 10704
rect 17314 9580 17370 9616
rect 17314 9560 17316 9580
rect 17316 9560 17368 9580
rect 17368 9560 17370 9580
rect 15618 2746 15674 2748
rect 15698 2746 15754 2748
rect 15778 2746 15834 2748
rect 15858 2746 15914 2748
rect 15618 2694 15664 2746
rect 15664 2694 15674 2746
rect 15698 2694 15728 2746
rect 15728 2694 15740 2746
rect 15740 2694 15754 2746
rect 15778 2694 15792 2746
rect 15792 2694 15804 2746
rect 15804 2694 15834 2746
rect 15858 2694 15868 2746
rect 15868 2694 15914 2746
rect 15618 2692 15674 2694
rect 15698 2692 15754 2694
rect 15778 2692 15834 2694
rect 15858 2692 15914 2694
rect 16486 3068 16488 3088
rect 16488 3068 16540 3088
rect 16540 3068 16542 3088
rect 16486 3032 16542 3068
rect 16394 2488 16450 2544
rect 15750 2372 15806 2408
rect 15750 2352 15752 2372
rect 15752 2352 15804 2372
rect 15804 2352 15806 2372
rect 15198 1300 15200 1320
rect 15200 1300 15252 1320
rect 15252 1300 15254 1320
rect 15198 1264 15254 1300
rect 15618 1658 15674 1660
rect 15698 1658 15754 1660
rect 15778 1658 15834 1660
rect 15858 1658 15914 1660
rect 15618 1606 15664 1658
rect 15664 1606 15674 1658
rect 15698 1606 15728 1658
rect 15728 1606 15740 1658
rect 15740 1606 15754 1658
rect 15778 1606 15792 1658
rect 15792 1606 15804 1658
rect 15804 1606 15834 1658
rect 15858 1606 15868 1658
rect 15868 1606 15914 1658
rect 15618 1604 15674 1606
rect 15698 1604 15754 1606
rect 15778 1604 15834 1606
rect 15858 1604 15914 1606
rect 16854 2624 16910 2680
rect 17222 3596 17278 3632
rect 17222 3576 17224 3596
rect 17224 3576 17276 3596
rect 17276 3576 17278 3596
rect 17130 2624 17186 2680
rect 17498 5752 17554 5808
rect 17406 5480 17462 5536
rect 18142 19508 18198 19544
rect 18142 19488 18144 19508
rect 18144 19488 18196 19508
rect 18196 19488 18198 19508
rect 18550 30490 18606 30492
rect 18630 30490 18686 30492
rect 18710 30490 18766 30492
rect 18790 30490 18846 30492
rect 18550 30438 18596 30490
rect 18596 30438 18606 30490
rect 18630 30438 18660 30490
rect 18660 30438 18672 30490
rect 18672 30438 18686 30490
rect 18710 30438 18724 30490
rect 18724 30438 18736 30490
rect 18736 30438 18766 30490
rect 18790 30438 18800 30490
rect 18800 30438 18846 30490
rect 18550 30436 18606 30438
rect 18630 30436 18686 30438
rect 18710 30436 18766 30438
rect 18790 30436 18846 30438
rect 18550 29402 18606 29404
rect 18630 29402 18686 29404
rect 18710 29402 18766 29404
rect 18790 29402 18846 29404
rect 18550 29350 18596 29402
rect 18596 29350 18606 29402
rect 18630 29350 18660 29402
rect 18660 29350 18672 29402
rect 18672 29350 18686 29402
rect 18710 29350 18724 29402
rect 18724 29350 18736 29402
rect 18736 29350 18766 29402
rect 18790 29350 18800 29402
rect 18800 29350 18846 29402
rect 18550 29348 18606 29350
rect 18630 29348 18686 29350
rect 18710 29348 18766 29350
rect 18790 29348 18846 29350
rect 18550 28314 18606 28316
rect 18630 28314 18686 28316
rect 18710 28314 18766 28316
rect 18790 28314 18846 28316
rect 18550 28262 18596 28314
rect 18596 28262 18606 28314
rect 18630 28262 18660 28314
rect 18660 28262 18672 28314
rect 18672 28262 18686 28314
rect 18710 28262 18724 28314
rect 18724 28262 18736 28314
rect 18736 28262 18766 28314
rect 18790 28262 18800 28314
rect 18800 28262 18846 28314
rect 18550 28260 18606 28262
rect 18630 28260 18686 28262
rect 18710 28260 18766 28262
rect 18790 28260 18846 28262
rect 18550 27226 18606 27228
rect 18630 27226 18686 27228
rect 18710 27226 18766 27228
rect 18790 27226 18846 27228
rect 18550 27174 18596 27226
rect 18596 27174 18606 27226
rect 18630 27174 18660 27226
rect 18660 27174 18672 27226
rect 18672 27174 18686 27226
rect 18710 27174 18724 27226
rect 18724 27174 18736 27226
rect 18736 27174 18766 27226
rect 18790 27174 18800 27226
rect 18800 27174 18846 27226
rect 18550 27172 18606 27174
rect 18630 27172 18686 27174
rect 18710 27172 18766 27174
rect 18790 27172 18846 27174
rect 18550 26138 18606 26140
rect 18630 26138 18686 26140
rect 18710 26138 18766 26140
rect 18790 26138 18846 26140
rect 18550 26086 18596 26138
rect 18596 26086 18606 26138
rect 18630 26086 18660 26138
rect 18660 26086 18672 26138
rect 18672 26086 18686 26138
rect 18710 26086 18724 26138
rect 18724 26086 18736 26138
rect 18736 26086 18766 26138
rect 18790 26086 18800 26138
rect 18800 26086 18846 26138
rect 18550 26084 18606 26086
rect 18630 26084 18686 26086
rect 18710 26084 18766 26086
rect 18790 26084 18846 26086
rect 18550 25050 18606 25052
rect 18630 25050 18686 25052
rect 18710 25050 18766 25052
rect 18790 25050 18846 25052
rect 18550 24998 18596 25050
rect 18596 24998 18606 25050
rect 18630 24998 18660 25050
rect 18660 24998 18672 25050
rect 18672 24998 18686 25050
rect 18710 24998 18724 25050
rect 18724 24998 18736 25050
rect 18736 24998 18766 25050
rect 18790 24998 18800 25050
rect 18800 24998 18846 25050
rect 18550 24996 18606 24998
rect 18630 24996 18686 24998
rect 18710 24996 18766 24998
rect 18790 24996 18846 24998
rect 18550 23962 18606 23964
rect 18630 23962 18686 23964
rect 18710 23962 18766 23964
rect 18790 23962 18846 23964
rect 18550 23910 18596 23962
rect 18596 23910 18606 23962
rect 18630 23910 18660 23962
rect 18660 23910 18672 23962
rect 18672 23910 18686 23962
rect 18710 23910 18724 23962
rect 18724 23910 18736 23962
rect 18736 23910 18766 23962
rect 18790 23910 18800 23962
rect 18800 23910 18846 23962
rect 18550 23908 18606 23910
rect 18630 23908 18686 23910
rect 18710 23908 18766 23910
rect 18790 23908 18846 23910
rect 18418 23604 18420 23624
rect 18420 23604 18472 23624
rect 18472 23604 18474 23624
rect 18418 23568 18474 23604
rect 18550 22874 18606 22876
rect 18630 22874 18686 22876
rect 18710 22874 18766 22876
rect 18790 22874 18846 22876
rect 18550 22822 18596 22874
rect 18596 22822 18606 22874
rect 18630 22822 18660 22874
rect 18660 22822 18672 22874
rect 18672 22822 18686 22874
rect 18710 22822 18724 22874
rect 18724 22822 18736 22874
rect 18736 22822 18766 22874
rect 18790 22822 18800 22874
rect 18800 22822 18846 22874
rect 18550 22820 18606 22822
rect 18630 22820 18686 22822
rect 18710 22820 18766 22822
rect 18790 22820 18846 22822
rect 18550 21786 18606 21788
rect 18630 21786 18686 21788
rect 18710 21786 18766 21788
rect 18790 21786 18846 21788
rect 18550 21734 18596 21786
rect 18596 21734 18606 21786
rect 18630 21734 18660 21786
rect 18660 21734 18672 21786
rect 18672 21734 18686 21786
rect 18710 21734 18724 21786
rect 18724 21734 18736 21786
rect 18736 21734 18766 21786
rect 18790 21734 18800 21786
rect 18800 21734 18846 21786
rect 18550 21732 18606 21734
rect 18630 21732 18686 21734
rect 18710 21732 18766 21734
rect 18790 21732 18846 21734
rect 18550 20698 18606 20700
rect 18630 20698 18686 20700
rect 18710 20698 18766 20700
rect 18790 20698 18846 20700
rect 18550 20646 18596 20698
rect 18596 20646 18606 20698
rect 18630 20646 18660 20698
rect 18660 20646 18672 20698
rect 18672 20646 18686 20698
rect 18710 20646 18724 20698
rect 18724 20646 18736 20698
rect 18736 20646 18766 20698
rect 18790 20646 18800 20698
rect 18800 20646 18846 20698
rect 18550 20644 18606 20646
rect 18630 20644 18686 20646
rect 18710 20644 18766 20646
rect 18790 20644 18846 20646
rect 18418 19760 18474 19816
rect 18550 19610 18606 19612
rect 18630 19610 18686 19612
rect 18710 19610 18766 19612
rect 18790 19610 18846 19612
rect 18550 19558 18596 19610
rect 18596 19558 18606 19610
rect 18630 19558 18660 19610
rect 18660 19558 18672 19610
rect 18672 19558 18686 19610
rect 18710 19558 18724 19610
rect 18724 19558 18736 19610
rect 18736 19558 18766 19610
rect 18790 19558 18800 19610
rect 18800 19558 18846 19610
rect 18550 19556 18606 19558
rect 18630 19556 18686 19558
rect 18710 19556 18766 19558
rect 18790 19556 18846 19558
rect 18550 18522 18606 18524
rect 18630 18522 18686 18524
rect 18710 18522 18766 18524
rect 18790 18522 18846 18524
rect 18550 18470 18596 18522
rect 18596 18470 18606 18522
rect 18630 18470 18660 18522
rect 18660 18470 18672 18522
rect 18672 18470 18686 18522
rect 18710 18470 18724 18522
rect 18724 18470 18736 18522
rect 18736 18470 18766 18522
rect 18790 18470 18800 18522
rect 18800 18470 18846 18522
rect 18550 18468 18606 18470
rect 18630 18468 18686 18470
rect 18710 18468 18766 18470
rect 18790 18468 18846 18470
rect 18550 17434 18606 17436
rect 18630 17434 18686 17436
rect 18710 17434 18766 17436
rect 18790 17434 18846 17436
rect 18550 17382 18596 17434
rect 18596 17382 18606 17434
rect 18630 17382 18660 17434
rect 18660 17382 18672 17434
rect 18672 17382 18686 17434
rect 18710 17382 18724 17434
rect 18724 17382 18736 17434
rect 18736 17382 18766 17434
rect 18790 17382 18800 17434
rect 18800 17382 18846 17434
rect 18550 17380 18606 17382
rect 18630 17380 18686 17382
rect 18710 17380 18766 17382
rect 18790 17380 18846 17382
rect 19338 31728 19394 31784
rect 18550 16346 18606 16348
rect 18630 16346 18686 16348
rect 18710 16346 18766 16348
rect 18790 16346 18846 16348
rect 18550 16294 18596 16346
rect 18596 16294 18606 16346
rect 18630 16294 18660 16346
rect 18660 16294 18672 16346
rect 18672 16294 18686 16346
rect 18710 16294 18724 16346
rect 18724 16294 18736 16346
rect 18736 16294 18766 16346
rect 18790 16294 18800 16346
rect 18800 16294 18846 16346
rect 18550 16292 18606 16294
rect 18630 16292 18686 16294
rect 18710 16292 18766 16294
rect 18790 16292 18846 16294
rect 18050 8880 18106 8936
rect 17590 4664 17646 4720
rect 17774 3032 17830 3088
rect 18550 15258 18606 15260
rect 18630 15258 18686 15260
rect 18710 15258 18766 15260
rect 18790 15258 18846 15260
rect 18550 15206 18596 15258
rect 18596 15206 18606 15258
rect 18630 15206 18660 15258
rect 18660 15206 18672 15258
rect 18672 15206 18686 15258
rect 18710 15206 18724 15258
rect 18724 15206 18736 15258
rect 18736 15206 18766 15258
rect 18790 15206 18800 15258
rect 18800 15206 18846 15258
rect 18550 15204 18606 15206
rect 18630 15204 18686 15206
rect 18710 15204 18766 15206
rect 18790 15204 18846 15206
rect 18550 14170 18606 14172
rect 18630 14170 18686 14172
rect 18710 14170 18766 14172
rect 18790 14170 18846 14172
rect 18550 14118 18596 14170
rect 18596 14118 18606 14170
rect 18630 14118 18660 14170
rect 18660 14118 18672 14170
rect 18672 14118 18686 14170
rect 18710 14118 18724 14170
rect 18724 14118 18736 14170
rect 18736 14118 18766 14170
rect 18790 14118 18800 14170
rect 18800 14118 18846 14170
rect 18550 14116 18606 14118
rect 18630 14116 18686 14118
rect 18710 14116 18766 14118
rect 18790 14116 18846 14118
rect 18550 13082 18606 13084
rect 18630 13082 18686 13084
rect 18710 13082 18766 13084
rect 18790 13082 18846 13084
rect 18550 13030 18596 13082
rect 18596 13030 18606 13082
rect 18630 13030 18660 13082
rect 18660 13030 18672 13082
rect 18672 13030 18686 13082
rect 18710 13030 18724 13082
rect 18724 13030 18736 13082
rect 18736 13030 18766 13082
rect 18790 13030 18800 13082
rect 18800 13030 18846 13082
rect 18550 13028 18606 13030
rect 18630 13028 18686 13030
rect 18710 13028 18766 13030
rect 18790 13028 18846 13030
rect 18550 11994 18606 11996
rect 18630 11994 18686 11996
rect 18710 11994 18766 11996
rect 18790 11994 18846 11996
rect 18550 11942 18596 11994
rect 18596 11942 18606 11994
rect 18630 11942 18660 11994
rect 18660 11942 18672 11994
rect 18672 11942 18686 11994
rect 18710 11942 18724 11994
rect 18724 11942 18736 11994
rect 18736 11942 18766 11994
rect 18790 11942 18800 11994
rect 18800 11942 18846 11994
rect 18550 11940 18606 11942
rect 18630 11940 18686 11942
rect 18710 11940 18766 11942
rect 18790 11940 18846 11942
rect 18550 10906 18606 10908
rect 18630 10906 18686 10908
rect 18710 10906 18766 10908
rect 18790 10906 18846 10908
rect 18550 10854 18596 10906
rect 18596 10854 18606 10906
rect 18630 10854 18660 10906
rect 18660 10854 18672 10906
rect 18672 10854 18686 10906
rect 18710 10854 18724 10906
rect 18724 10854 18736 10906
rect 18736 10854 18766 10906
rect 18790 10854 18800 10906
rect 18800 10854 18846 10906
rect 18550 10852 18606 10854
rect 18630 10852 18686 10854
rect 18710 10852 18766 10854
rect 18790 10852 18846 10854
rect 18550 9818 18606 9820
rect 18630 9818 18686 9820
rect 18710 9818 18766 9820
rect 18790 9818 18846 9820
rect 18550 9766 18596 9818
rect 18596 9766 18606 9818
rect 18630 9766 18660 9818
rect 18660 9766 18672 9818
rect 18672 9766 18686 9818
rect 18710 9766 18724 9818
rect 18724 9766 18736 9818
rect 18736 9766 18766 9818
rect 18790 9766 18800 9818
rect 18800 9766 18846 9818
rect 18550 9764 18606 9766
rect 18630 9764 18686 9766
rect 18710 9764 18766 9766
rect 18790 9764 18846 9766
rect 18510 9424 18566 9480
rect 18550 8730 18606 8732
rect 18630 8730 18686 8732
rect 18710 8730 18766 8732
rect 18790 8730 18846 8732
rect 18550 8678 18596 8730
rect 18596 8678 18606 8730
rect 18630 8678 18660 8730
rect 18660 8678 18672 8730
rect 18672 8678 18686 8730
rect 18710 8678 18724 8730
rect 18724 8678 18736 8730
rect 18736 8678 18766 8730
rect 18790 8678 18800 8730
rect 18800 8678 18846 8730
rect 18550 8676 18606 8678
rect 18630 8676 18686 8678
rect 18710 8676 18766 8678
rect 18790 8676 18846 8678
rect 18550 7642 18606 7644
rect 18630 7642 18686 7644
rect 18710 7642 18766 7644
rect 18790 7642 18846 7644
rect 18550 7590 18596 7642
rect 18596 7590 18606 7642
rect 18630 7590 18660 7642
rect 18660 7590 18672 7642
rect 18672 7590 18686 7642
rect 18710 7590 18724 7642
rect 18724 7590 18736 7642
rect 18736 7590 18766 7642
rect 18790 7590 18800 7642
rect 18800 7590 18846 7642
rect 18550 7588 18606 7590
rect 18630 7588 18686 7590
rect 18710 7588 18766 7590
rect 18790 7588 18846 7590
rect 18550 6554 18606 6556
rect 18630 6554 18686 6556
rect 18710 6554 18766 6556
rect 18790 6554 18846 6556
rect 18550 6502 18596 6554
rect 18596 6502 18606 6554
rect 18630 6502 18660 6554
rect 18660 6502 18672 6554
rect 18672 6502 18686 6554
rect 18710 6502 18724 6554
rect 18724 6502 18736 6554
rect 18736 6502 18766 6554
rect 18790 6502 18800 6554
rect 18800 6502 18846 6554
rect 18550 6500 18606 6502
rect 18630 6500 18686 6502
rect 18710 6500 18766 6502
rect 18790 6500 18846 6502
rect 18550 5466 18606 5468
rect 18630 5466 18686 5468
rect 18710 5466 18766 5468
rect 18790 5466 18846 5468
rect 18550 5414 18596 5466
rect 18596 5414 18606 5466
rect 18630 5414 18660 5466
rect 18660 5414 18672 5466
rect 18672 5414 18686 5466
rect 18710 5414 18724 5466
rect 18724 5414 18736 5466
rect 18736 5414 18766 5466
rect 18790 5414 18800 5466
rect 18800 5414 18846 5466
rect 18550 5412 18606 5414
rect 18630 5412 18686 5414
rect 18710 5412 18766 5414
rect 18790 5412 18846 5414
rect 18550 4378 18606 4380
rect 18630 4378 18686 4380
rect 18710 4378 18766 4380
rect 18790 4378 18846 4380
rect 18550 4326 18596 4378
rect 18596 4326 18606 4378
rect 18630 4326 18660 4378
rect 18660 4326 18672 4378
rect 18672 4326 18686 4378
rect 18710 4326 18724 4378
rect 18724 4326 18736 4378
rect 18736 4326 18766 4378
rect 18790 4326 18800 4378
rect 18800 4326 18846 4378
rect 18550 4324 18606 4326
rect 18630 4324 18686 4326
rect 18710 4324 18766 4326
rect 18790 4324 18846 4326
rect 18550 3290 18606 3292
rect 18630 3290 18686 3292
rect 18710 3290 18766 3292
rect 18790 3290 18846 3292
rect 18550 3238 18596 3290
rect 18596 3238 18606 3290
rect 18630 3238 18660 3290
rect 18660 3238 18672 3290
rect 18672 3238 18686 3290
rect 18710 3238 18724 3290
rect 18724 3238 18736 3290
rect 18736 3238 18766 3290
rect 18790 3238 18800 3290
rect 18800 3238 18846 3290
rect 18550 3236 18606 3238
rect 18630 3236 18686 3238
rect 18710 3236 18766 3238
rect 18790 3236 18846 3238
rect 18970 8880 19026 8936
rect 18970 8472 19026 8528
rect 19154 11736 19210 11792
rect 19338 12688 19394 12744
rect 19614 41384 19670 41420
rect 19798 41928 19854 41984
rect 21270 43152 21326 43208
rect 22006 43696 22062 43752
rect 21483 43002 21539 43004
rect 21563 43002 21619 43004
rect 21643 43002 21699 43004
rect 21723 43002 21779 43004
rect 21483 42950 21529 43002
rect 21529 42950 21539 43002
rect 21563 42950 21593 43002
rect 21593 42950 21605 43002
rect 21605 42950 21619 43002
rect 21643 42950 21657 43002
rect 21657 42950 21669 43002
rect 21669 42950 21699 43002
rect 21723 42950 21733 43002
rect 21733 42950 21779 43002
rect 21483 42948 21539 42950
rect 21563 42948 21619 42950
rect 21643 42948 21699 42950
rect 21723 42948 21779 42950
rect 21086 42220 21142 42256
rect 21086 42200 21088 42220
rect 21088 42200 21140 42220
rect 21140 42200 21142 42220
rect 20626 41656 20682 41712
rect 20534 41556 20536 41576
rect 20536 41556 20588 41576
rect 20588 41556 20590 41576
rect 20534 41520 20590 41556
rect 20350 40432 20406 40488
rect 20258 39480 20314 39536
rect 20350 36780 20406 36816
rect 20350 36760 20352 36780
rect 20352 36760 20404 36780
rect 20404 36760 20406 36780
rect 19522 34040 19578 34096
rect 20442 29144 20498 29200
rect 21270 41656 21326 41712
rect 21483 41914 21539 41916
rect 21563 41914 21619 41916
rect 21643 41914 21699 41916
rect 21723 41914 21779 41916
rect 21483 41862 21529 41914
rect 21529 41862 21539 41914
rect 21563 41862 21593 41914
rect 21593 41862 21605 41914
rect 21605 41862 21619 41914
rect 21643 41862 21657 41914
rect 21657 41862 21669 41914
rect 21669 41862 21699 41914
rect 21723 41862 21733 41914
rect 21733 41862 21779 41914
rect 21483 41860 21539 41862
rect 21563 41860 21619 41862
rect 21643 41860 21699 41862
rect 21723 41860 21779 41862
rect 21454 41384 21510 41440
rect 21483 40826 21539 40828
rect 21563 40826 21619 40828
rect 21643 40826 21699 40828
rect 21723 40826 21779 40828
rect 21483 40774 21529 40826
rect 21529 40774 21539 40826
rect 21563 40774 21593 40826
rect 21593 40774 21605 40826
rect 21605 40774 21619 40826
rect 21643 40774 21657 40826
rect 21657 40774 21669 40826
rect 21669 40774 21699 40826
rect 21723 40774 21733 40826
rect 21733 40774 21779 40826
rect 21483 40772 21539 40774
rect 21563 40772 21619 40774
rect 21643 40772 21699 40774
rect 21723 40772 21779 40774
rect 21914 40840 21970 40896
rect 21822 39888 21878 39944
rect 21483 39738 21539 39740
rect 21563 39738 21619 39740
rect 21643 39738 21699 39740
rect 21723 39738 21779 39740
rect 21483 39686 21529 39738
rect 21529 39686 21539 39738
rect 21563 39686 21593 39738
rect 21593 39686 21605 39738
rect 21605 39686 21619 39738
rect 21643 39686 21657 39738
rect 21657 39686 21669 39738
rect 21669 39686 21699 39738
rect 21723 39686 21733 39738
rect 21733 39686 21779 39738
rect 21483 39684 21539 39686
rect 21563 39684 21619 39686
rect 21643 39684 21699 39686
rect 21723 39684 21779 39686
rect 21483 38650 21539 38652
rect 21563 38650 21619 38652
rect 21643 38650 21699 38652
rect 21723 38650 21779 38652
rect 21483 38598 21529 38650
rect 21529 38598 21539 38650
rect 21563 38598 21593 38650
rect 21593 38598 21605 38650
rect 21605 38598 21619 38650
rect 21643 38598 21657 38650
rect 21657 38598 21669 38650
rect 21669 38598 21699 38650
rect 21723 38598 21733 38650
rect 21733 38598 21779 38650
rect 21483 38596 21539 38598
rect 21563 38596 21619 38598
rect 21643 38596 21699 38598
rect 21723 38596 21779 38598
rect 21483 37562 21539 37564
rect 21563 37562 21619 37564
rect 21643 37562 21699 37564
rect 21723 37562 21779 37564
rect 21483 37510 21529 37562
rect 21529 37510 21539 37562
rect 21563 37510 21593 37562
rect 21593 37510 21605 37562
rect 21605 37510 21619 37562
rect 21643 37510 21657 37562
rect 21657 37510 21669 37562
rect 21669 37510 21699 37562
rect 21723 37510 21733 37562
rect 21733 37510 21779 37562
rect 21483 37508 21539 37510
rect 21563 37508 21619 37510
rect 21643 37508 21699 37510
rect 21723 37508 21779 37510
rect 21483 36474 21539 36476
rect 21563 36474 21619 36476
rect 21643 36474 21699 36476
rect 21723 36474 21779 36476
rect 21483 36422 21529 36474
rect 21529 36422 21539 36474
rect 21563 36422 21593 36474
rect 21593 36422 21605 36474
rect 21605 36422 21619 36474
rect 21643 36422 21657 36474
rect 21657 36422 21669 36474
rect 21669 36422 21699 36474
rect 21723 36422 21733 36474
rect 21733 36422 21779 36474
rect 21483 36420 21539 36422
rect 21563 36420 21619 36422
rect 21643 36420 21699 36422
rect 21723 36420 21779 36422
rect 21483 35386 21539 35388
rect 21563 35386 21619 35388
rect 21643 35386 21699 35388
rect 21723 35386 21779 35388
rect 21483 35334 21529 35386
rect 21529 35334 21539 35386
rect 21563 35334 21593 35386
rect 21593 35334 21605 35386
rect 21605 35334 21619 35386
rect 21643 35334 21657 35386
rect 21657 35334 21669 35386
rect 21669 35334 21699 35386
rect 21723 35334 21733 35386
rect 21733 35334 21779 35386
rect 21483 35332 21539 35334
rect 21563 35332 21619 35334
rect 21643 35332 21699 35334
rect 21723 35332 21779 35334
rect 22926 43016 22982 43072
rect 22374 40044 22430 40080
rect 22374 40024 22376 40044
rect 22376 40024 22428 40044
rect 22428 40024 22430 40044
rect 22282 39888 22338 39944
rect 20626 29144 20682 29200
rect 21086 29164 21142 29200
rect 21086 29144 21088 29164
rect 21088 29144 21140 29164
rect 21140 29144 21142 29164
rect 19430 12416 19486 12472
rect 19706 14864 19762 14920
rect 21086 24656 21142 24712
rect 21483 34298 21539 34300
rect 21563 34298 21619 34300
rect 21643 34298 21699 34300
rect 21723 34298 21779 34300
rect 21483 34246 21529 34298
rect 21529 34246 21539 34298
rect 21563 34246 21593 34298
rect 21593 34246 21605 34298
rect 21605 34246 21619 34298
rect 21643 34246 21657 34298
rect 21657 34246 21669 34298
rect 21669 34246 21699 34298
rect 21723 34246 21733 34298
rect 21733 34246 21779 34298
rect 21483 34244 21539 34246
rect 21563 34244 21619 34246
rect 21643 34244 21699 34246
rect 21723 34244 21779 34246
rect 21483 33210 21539 33212
rect 21563 33210 21619 33212
rect 21643 33210 21699 33212
rect 21723 33210 21779 33212
rect 21483 33158 21529 33210
rect 21529 33158 21539 33210
rect 21563 33158 21593 33210
rect 21593 33158 21605 33210
rect 21605 33158 21619 33210
rect 21643 33158 21657 33210
rect 21657 33158 21669 33210
rect 21669 33158 21699 33210
rect 21723 33158 21733 33210
rect 21733 33158 21779 33210
rect 21483 33156 21539 33158
rect 21563 33156 21619 33158
rect 21643 33156 21699 33158
rect 21723 33156 21779 33158
rect 21483 32122 21539 32124
rect 21563 32122 21619 32124
rect 21643 32122 21699 32124
rect 21723 32122 21779 32124
rect 21483 32070 21529 32122
rect 21529 32070 21539 32122
rect 21563 32070 21593 32122
rect 21593 32070 21605 32122
rect 21605 32070 21619 32122
rect 21643 32070 21657 32122
rect 21657 32070 21669 32122
rect 21669 32070 21699 32122
rect 21723 32070 21733 32122
rect 21733 32070 21779 32122
rect 21483 32068 21539 32070
rect 21563 32068 21619 32070
rect 21643 32068 21699 32070
rect 21723 32068 21779 32070
rect 21483 31034 21539 31036
rect 21563 31034 21619 31036
rect 21643 31034 21699 31036
rect 21723 31034 21779 31036
rect 21483 30982 21529 31034
rect 21529 30982 21539 31034
rect 21563 30982 21593 31034
rect 21593 30982 21605 31034
rect 21605 30982 21619 31034
rect 21643 30982 21657 31034
rect 21657 30982 21669 31034
rect 21669 30982 21699 31034
rect 21723 30982 21733 31034
rect 21733 30982 21779 31034
rect 21483 30980 21539 30982
rect 21563 30980 21619 30982
rect 21643 30980 21699 30982
rect 21723 30980 21779 30982
rect 21483 29946 21539 29948
rect 21563 29946 21619 29948
rect 21643 29946 21699 29948
rect 21723 29946 21779 29948
rect 21483 29894 21529 29946
rect 21529 29894 21539 29946
rect 21563 29894 21593 29946
rect 21593 29894 21605 29946
rect 21605 29894 21619 29946
rect 21643 29894 21657 29946
rect 21657 29894 21669 29946
rect 21669 29894 21699 29946
rect 21723 29894 21733 29946
rect 21733 29894 21779 29946
rect 21483 29892 21539 29894
rect 21563 29892 21619 29894
rect 21643 29892 21699 29894
rect 21723 29892 21779 29894
rect 23386 41520 23442 41576
rect 23386 39752 23442 39808
rect 24122 41928 24178 41984
rect 23846 41372 23902 41428
rect 23662 40876 23664 40896
rect 23664 40876 23716 40896
rect 23716 40876 23718 40896
rect 23662 40840 23718 40876
rect 21483 28858 21539 28860
rect 21563 28858 21619 28860
rect 21643 28858 21699 28860
rect 21723 28858 21779 28860
rect 21483 28806 21529 28858
rect 21529 28806 21539 28858
rect 21563 28806 21593 28858
rect 21593 28806 21605 28858
rect 21605 28806 21619 28858
rect 21643 28806 21657 28858
rect 21657 28806 21669 28858
rect 21669 28806 21699 28858
rect 21723 28806 21733 28858
rect 21733 28806 21779 28858
rect 21483 28804 21539 28806
rect 21563 28804 21619 28806
rect 21643 28804 21699 28806
rect 21723 28804 21779 28806
rect 21483 27770 21539 27772
rect 21563 27770 21619 27772
rect 21643 27770 21699 27772
rect 21723 27770 21779 27772
rect 21483 27718 21529 27770
rect 21529 27718 21539 27770
rect 21563 27718 21593 27770
rect 21593 27718 21605 27770
rect 21605 27718 21619 27770
rect 21643 27718 21657 27770
rect 21657 27718 21669 27770
rect 21669 27718 21699 27770
rect 21723 27718 21733 27770
rect 21733 27718 21779 27770
rect 21483 27716 21539 27718
rect 21563 27716 21619 27718
rect 21643 27716 21699 27718
rect 21723 27716 21779 27718
rect 21483 26682 21539 26684
rect 21563 26682 21619 26684
rect 21643 26682 21699 26684
rect 21723 26682 21779 26684
rect 21483 26630 21529 26682
rect 21529 26630 21539 26682
rect 21563 26630 21593 26682
rect 21593 26630 21605 26682
rect 21605 26630 21619 26682
rect 21643 26630 21657 26682
rect 21657 26630 21669 26682
rect 21669 26630 21699 26682
rect 21723 26630 21733 26682
rect 21733 26630 21779 26682
rect 21483 26628 21539 26630
rect 21563 26628 21619 26630
rect 21643 26628 21699 26630
rect 21723 26628 21779 26630
rect 21483 25594 21539 25596
rect 21563 25594 21619 25596
rect 21643 25594 21699 25596
rect 21723 25594 21779 25596
rect 21483 25542 21529 25594
rect 21529 25542 21539 25594
rect 21563 25542 21593 25594
rect 21593 25542 21605 25594
rect 21605 25542 21619 25594
rect 21643 25542 21657 25594
rect 21657 25542 21669 25594
rect 21669 25542 21699 25594
rect 21723 25542 21733 25594
rect 21733 25542 21779 25594
rect 21483 25540 21539 25542
rect 21563 25540 21619 25542
rect 21643 25540 21699 25542
rect 21723 25540 21779 25542
rect 21483 24506 21539 24508
rect 21563 24506 21619 24508
rect 21643 24506 21699 24508
rect 21723 24506 21779 24508
rect 21483 24454 21529 24506
rect 21529 24454 21539 24506
rect 21563 24454 21593 24506
rect 21593 24454 21605 24506
rect 21605 24454 21619 24506
rect 21643 24454 21657 24506
rect 21657 24454 21669 24506
rect 21669 24454 21699 24506
rect 21723 24454 21733 24506
rect 21733 24454 21779 24506
rect 21483 24452 21539 24454
rect 21563 24452 21619 24454
rect 21643 24452 21699 24454
rect 21723 24452 21779 24454
rect 21483 23418 21539 23420
rect 21563 23418 21619 23420
rect 21643 23418 21699 23420
rect 21723 23418 21779 23420
rect 21483 23366 21529 23418
rect 21529 23366 21539 23418
rect 21563 23366 21593 23418
rect 21593 23366 21605 23418
rect 21605 23366 21619 23418
rect 21643 23366 21657 23418
rect 21657 23366 21669 23418
rect 21669 23366 21699 23418
rect 21723 23366 21733 23418
rect 21733 23366 21779 23418
rect 21483 23364 21539 23366
rect 21563 23364 21619 23366
rect 21643 23364 21699 23366
rect 21723 23364 21779 23366
rect 21483 22330 21539 22332
rect 21563 22330 21619 22332
rect 21643 22330 21699 22332
rect 21723 22330 21779 22332
rect 21483 22278 21529 22330
rect 21529 22278 21539 22330
rect 21563 22278 21593 22330
rect 21593 22278 21605 22330
rect 21605 22278 21619 22330
rect 21643 22278 21657 22330
rect 21657 22278 21669 22330
rect 21669 22278 21699 22330
rect 21723 22278 21733 22330
rect 21733 22278 21779 22330
rect 21483 22276 21539 22278
rect 21563 22276 21619 22278
rect 21643 22276 21699 22278
rect 21723 22276 21779 22278
rect 19338 12008 19394 12064
rect 19338 9016 19394 9072
rect 21362 21936 21418 21992
rect 21483 21242 21539 21244
rect 21563 21242 21619 21244
rect 21643 21242 21699 21244
rect 21723 21242 21779 21244
rect 21483 21190 21529 21242
rect 21529 21190 21539 21242
rect 21563 21190 21593 21242
rect 21593 21190 21605 21242
rect 21605 21190 21619 21242
rect 21643 21190 21657 21242
rect 21657 21190 21669 21242
rect 21669 21190 21699 21242
rect 21723 21190 21733 21242
rect 21733 21190 21779 21242
rect 21483 21188 21539 21190
rect 21563 21188 21619 21190
rect 21643 21188 21699 21190
rect 21723 21188 21779 21190
rect 21483 20154 21539 20156
rect 21563 20154 21619 20156
rect 21643 20154 21699 20156
rect 21723 20154 21779 20156
rect 21483 20102 21529 20154
rect 21529 20102 21539 20154
rect 21563 20102 21593 20154
rect 21593 20102 21605 20154
rect 21605 20102 21619 20154
rect 21643 20102 21657 20154
rect 21657 20102 21669 20154
rect 21669 20102 21699 20154
rect 21723 20102 21733 20154
rect 21733 20102 21779 20154
rect 21483 20100 21539 20102
rect 21563 20100 21619 20102
rect 21643 20100 21699 20102
rect 21723 20100 21779 20102
rect 20810 13368 20866 13424
rect 19982 12280 20038 12336
rect 20166 12144 20222 12200
rect 19522 8336 19578 8392
rect 19246 6160 19302 6216
rect 20166 10512 20222 10568
rect 20258 9016 20314 9072
rect 19522 5344 19578 5400
rect 19430 5208 19486 5264
rect 19430 4256 19486 4312
rect 19430 3732 19486 3768
rect 19430 3712 19432 3732
rect 19432 3712 19484 3732
rect 19484 3712 19486 3732
rect 18550 2202 18606 2204
rect 18630 2202 18686 2204
rect 18710 2202 18766 2204
rect 18790 2202 18846 2204
rect 18550 2150 18596 2202
rect 18596 2150 18606 2202
rect 18630 2150 18660 2202
rect 18660 2150 18672 2202
rect 18672 2150 18686 2202
rect 18710 2150 18724 2202
rect 18724 2150 18736 2202
rect 18736 2150 18766 2202
rect 18790 2150 18800 2202
rect 18800 2150 18846 2202
rect 18550 2148 18606 2150
rect 18630 2148 18686 2150
rect 18710 2148 18766 2150
rect 18790 2148 18846 2150
rect 18550 1114 18606 1116
rect 18630 1114 18686 1116
rect 18710 1114 18766 1116
rect 18790 1114 18846 1116
rect 18550 1062 18596 1114
rect 18596 1062 18606 1114
rect 18630 1062 18660 1114
rect 18660 1062 18672 1114
rect 18672 1062 18686 1114
rect 18710 1062 18724 1114
rect 18724 1062 18736 1114
rect 18736 1062 18766 1114
rect 18790 1062 18800 1114
rect 18800 1062 18846 1114
rect 18550 1060 18606 1062
rect 18630 1060 18686 1062
rect 18710 1060 18766 1062
rect 18790 1060 18846 1062
rect 20718 8744 20774 8800
rect 20718 7520 20774 7576
rect 20810 6568 20866 6624
rect 20350 5344 20406 5400
rect 19798 5228 19854 5264
rect 19798 5208 19800 5228
rect 19800 5208 19852 5228
rect 19852 5208 19854 5228
rect 19982 4392 20038 4448
rect 19706 3984 19762 4040
rect 19614 2624 19670 2680
rect 19982 3984 20038 4040
rect 19890 2896 19946 2952
rect 20258 4256 20314 4312
rect 20350 3168 20406 3224
rect 19982 1808 20038 1864
rect 20534 3032 20590 3088
rect 21483 19066 21539 19068
rect 21563 19066 21619 19068
rect 21643 19066 21699 19068
rect 21723 19066 21779 19068
rect 21483 19014 21529 19066
rect 21529 19014 21539 19066
rect 21563 19014 21593 19066
rect 21593 19014 21605 19066
rect 21605 19014 21619 19066
rect 21643 19014 21657 19066
rect 21657 19014 21669 19066
rect 21669 19014 21699 19066
rect 21723 19014 21733 19066
rect 21733 19014 21779 19066
rect 21483 19012 21539 19014
rect 21563 19012 21619 19014
rect 21643 19012 21699 19014
rect 21723 19012 21779 19014
rect 23202 34584 23258 34640
rect 22558 24112 22614 24168
rect 21483 17978 21539 17980
rect 21563 17978 21619 17980
rect 21643 17978 21699 17980
rect 21723 17978 21779 17980
rect 21483 17926 21529 17978
rect 21529 17926 21539 17978
rect 21563 17926 21593 17978
rect 21593 17926 21605 17978
rect 21605 17926 21619 17978
rect 21643 17926 21657 17978
rect 21657 17926 21669 17978
rect 21669 17926 21699 17978
rect 21723 17926 21733 17978
rect 21733 17926 21779 17978
rect 21483 17924 21539 17926
rect 21563 17924 21619 17926
rect 21643 17924 21699 17926
rect 21723 17924 21779 17926
rect 21483 16890 21539 16892
rect 21563 16890 21619 16892
rect 21643 16890 21699 16892
rect 21723 16890 21779 16892
rect 21483 16838 21529 16890
rect 21529 16838 21539 16890
rect 21563 16838 21593 16890
rect 21593 16838 21605 16890
rect 21605 16838 21619 16890
rect 21643 16838 21657 16890
rect 21657 16838 21669 16890
rect 21669 16838 21699 16890
rect 21723 16838 21733 16890
rect 21733 16838 21779 16890
rect 21483 16836 21539 16838
rect 21563 16836 21619 16838
rect 21643 16836 21699 16838
rect 21723 16836 21779 16838
rect 21483 15802 21539 15804
rect 21563 15802 21619 15804
rect 21643 15802 21699 15804
rect 21723 15802 21779 15804
rect 21483 15750 21529 15802
rect 21529 15750 21539 15802
rect 21563 15750 21593 15802
rect 21593 15750 21605 15802
rect 21605 15750 21619 15802
rect 21643 15750 21657 15802
rect 21657 15750 21669 15802
rect 21669 15750 21699 15802
rect 21723 15750 21733 15802
rect 21733 15750 21779 15802
rect 21483 15748 21539 15750
rect 21563 15748 21619 15750
rect 21643 15748 21699 15750
rect 21723 15748 21779 15750
rect 21730 15000 21786 15056
rect 21483 14714 21539 14716
rect 21563 14714 21619 14716
rect 21643 14714 21699 14716
rect 21723 14714 21779 14716
rect 21483 14662 21529 14714
rect 21529 14662 21539 14714
rect 21563 14662 21593 14714
rect 21593 14662 21605 14714
rect 21605 14662 21619 14714
rect 21643 14662 21657 14714
rect 21657 14662 21669 14714
rect 21669 14662 21699 14714
rect 21723 14662 21733 14714
rect 21733 14662 21779 14714
rect 21483 14660 21539 14662
rect 21563 14660 21619 14662
rect 21643 14660 21699 14662
rect 21723 14660 21779 14662
rect 21483 13626 21539 13628
rect 21563 13626 21619 13628
rect 21643 13626 21699 13628
rect 21723 13626 21779 13628
rect 21483 13574 21529 13626
rect 21529 13574 21539 13626
rect 21563 13574 21593 13626
rect 21593 13574 21605 13626
rect 21605 13574 21619 13626
rect 21643 13574 21657 13626
rect 21657 13574 21669 13626
rect 21669 13574 21699 13626
rect 21723 13574 21733 13626
rect 21733 13574 21779 13626
rect 21483 13572 21539 13574
rect 21563 13572 21619 13574
rect 21643 13572 21699 13574
rect 21723 13572 21779 13574
rect 21483 12538 21539 12540
rect 21563 12538 21619 12540
rect 21643 12538 21699 12540
rect 21723 12538 21779 12540
rect 21483 12486 21529 12538
rect 21529 12486 21539 12538
rect 21563 12486 21593 12538
rect 21593 12486 21605 12538
rect 21605 12486 21619 12538
rect 21643 12486 21657 12538
rect 21657 12486 21669 12538
rect 21669 12486 21699 12538
rect 21723 12486 21733 12538
rect 21733 12486 21779 12538
rect 21483 12484 21539 12486
rect 21563 12484 21619 12486
rect 21643 12484 21699 12486
rect 21723 12484 21779 12486
rect 22650 15136 22706 15192
rect 22650 13776 22706 13832
rect 22190 12688 22246 12744
rect 21483 11450 21539 11452
rect 21563 11450 21619 11452
rect 21643 11450 21699 11452
rect 21723 11450 21779 11452
rect 21483 11398 21529 11450
rect 21529 11398 21539 11450
rect 21563 11398 21593 11450
rect 21593 11398 21605 11450
rect 21605 11398 21619 11450
rect 21643 11398 21657 11450
rect 21657 11398 21669 11450
rect 21669 11398 21699 11450
rect 21723 11398 21733 11450
rect 21733 11398 21779 11450
rect 21483 11396 21539 11398
rect 21563 11396 21619 11398
rect 21643 11396 21699 11398
rect 21723 11396 21779 11398
rect 22834 15000 22890 15056
rect 24122 39788 24124 39808
rect 24124 39788 24176 39808
rect 24176 39788 24178 39808
rect 24122 39752 24178 39788
rect 24122 38700 24124 38720
rect 24124 38700 24176 38720
rect 24176 38700 24178 38720
rect 24122 38664 24178 38700
rect 24122 37612 24124 37632
rect 24124 37612 24176 37632
rect 24176 37612 24178 37632
rect 24122 37576 24178 37612
rect 24122 36524 24124 36544
rect 24124 36524 24176 36544
rect 24176 36524 24178 36544
rect 24122 36488 24178 36524
rect 24415 43546 24471 43548
rect 24495 43546 24551 43548
rect 24575 43546 24631 43548
rect 24655 43546 24711 43548
rect 24415 43494 24461 43546
rect 24461 43494 24471 43546
rect 24495 43494 24525 43546
rect 24525 43494 24537 43546
rect 24537 43494 24551 43546
rect 24575 43494 24589 43546
rect 24589 43494 24601 43546
rect 24601 43494 24631 43546
rect 24655 43494 24665 43546
rect 24665 43494 24711 43546
rect 24415 43492 24471 43494
rect 24495 43492 24551 43494
rect 24575 43492 24631 43494
rect 24655 43492 24711 43494
rect 24415 42458 24471 42460
rect 24495 42458 24551 42460
rect 24575 42458 24631 42460
rect 24655 42458 24711 42460
rect 24415 42406 24461 42458
rect 24461 42406 24471 42458
rect 24495 42406 24525 42458
rect 24525 42406 24537 42458
rect 24537 42406 24551 42458
rect 24575 42406 24589 42458
rect 24589 42406 24601 42458
rect 24601 42406 24631 42458
rect 24655 42406 24665 42458
rect 24665 42406 24711 42458
rect 24415 42404 24471 42406
rect 24495 42404 24551 42406
rect 24575 42404 24631 42406
rect 24655 42404 24711 42406
rect 24415 41370 24471 41372
rect 24495 41370 24551 41372
rect 24575 41370 24631 41372
rect 24655 41370 24711 41372
rect 24415 41318 24461 41370
rect 24461 41318 24471 41370
rect 24495 41318 24525 41370
rect 24525 41318 24537 41370
rect 24537 41318 24551 41370
rect 24575 41318 24589 41370
rect 24589 41318 24601 41370
rect 24601 41318 24631 41370
rect 24655 41318 24665 41370
rect 24665 41318 24711 41370
rect 24415 41316 24471 41318
rect 24495 41316 24551 41318
rect 24575 41316 24631 41318
rect 24655 41316 24711 41318
rect 24858 42472 24914 42528
rect 25042 40432 25098 40488
rect 24950 40296 25006 40352
rect 24415 40282 24471 40284
rect 24495 40282 24551 40284
rect 24575 40282 24631 40284
rect 24655 40282 24711 40284
rect 24415 40230 24461 40282
rect 24461 40230 24471 40282
rect 24495 40230 24525 40282
rect 24525 40230 24537 40282
rect 24537 40230 24551 40282
rect 24575 40230 24589 40282
rect 24589 40230 24601 40282
rect 24601 40230 24631 40282
rect 24655 40230 24665 40282
rect 24665 40230 24711 40282
rect 24415 40228 24471 40230
rect 24495 40228 24551 40230
rect 24575 40228 24631 40230
rect 24655 40228 24711 40230
rect 24950 39480 25006 39536
rect 24858 39244 24860 39264
rect 24860 39244 24912 39264
rect 24912 39244 24914 39264
rect 24858 39208 24914 39244
rect 24415 39194 24471 39196
rect 24495 39194 24551 39196
rect 24575 39194 24631 39196
rect 24655 39194 24711 39196
rect 24415 39142 24461 39194
rect 24461 39142 24471 39194
rect 24495 39142 24525 39194
rect 24525 39142 24537 39194
rect 24537 39142 24551 39194
rect 24575 39142 24589 39194
rect 24589 39142 24601 39194
rect 24601 39142 24631 39194
rect 24655 39142 24665 39194
rect 24665 39142 24711 39194
rect 24415 39140 24471 39142
rect 24495 39140 24551 39142
rect 24575 39140 24631 39142
rect 24655 39140 24711 39142
rect 24122 35436 24124 35456
rect 24124 35436 24176 35456
rect 24176 35436 24178 35456
rect 24122 35400 24178 35436
rect 24122 34484 24124 34504
rect 24124 34484 24176 34504
rect 24176 34484 24178 34504
rect 24122 34448 24178 34484
rect 24214 33496 24270 33552
rect 24122 33260 24124 33280
rect 24124 33260 24176 33280
rect 24176 33260 24178 33280
rect 24122 33224 24178 33260
rect 24122 32172 24124 32192
rect 24124 32172 24176 32192
rect 24176 32172 24178 32192
rect 24122 32136 24178 32172
rect 24122 31084 24124 31104
rect 24124 31084 24176 31104
rect 24176 31084 24178 31104
rect 24122 31048 24178 31084
rect 23754 25644 23756 25664
rect 23756 25644 23808 25664
rect 23808 25644 23810 25664
rect 23754 25608 23810 25644
rect 24122 29996 24124 30016
rect 24124 29996 24176 30016
rect 24176 29996 24178 30016
rect 24122 29960 24178 29996
rect 24122 28872 24178 28928
rect 24122 27820 24124 27840
rect 24124 27820 24176 27840
rect 24176 27820 24178 27840
rect 24122 27784 24178 27820
rect 24122 26732 24124 26752
rect 24124 26732 24176 26752
rect 24176 26732 24178 26752
rect 24122 26696 24178 26732
rect 23846 24520 23902 24576
rect 23018 15136 23074 15192
rect 22834 13368 22890 13424
rect 21483 10362 21539 10364
rect 21563 10362 21619 10364
rect 21643 10362 21699 10364
rect 21723 10362 21779 10364
rect 21483 10310 21529 10362
rect 21529 10310 21539 10362
rect 21563 10310 21593 10362
rect 21593 10310 21605 10362
rect 21605 10310 21619 10362
rect 21643 10310 21657 10362
rect 21657 10310 21669 10362
rect 21669 10310 21699 10362
rect 21723 10310 21733 10362
rect 21733 10310 21779 10362
rect 21483 10308 21539 10310
rect 21563 10308 21619 10310
rect 21643 10308 21699 10310
rect 21723 10308 21779 10310
rect 21483 9274 21539 9276
rect 21563 9274 21619 9276
rect 21643 9274 21699 9276
rect 21723 9274 21779 9276
rect 21483 9222 21529 9274
rect 21529 9222 21539 9274
rect 21563 9222 21593 9274
rect 21593 9222 21605 9274
rect 21605 9222 21619 9274
rect 21643 9222 21657 9274
rect 21657 9222 21669 9274
rect 21669 9222 21699 9274
rect 21723 9222 21733 9274
rect 21733 9222 21779 9274
rect 21483 9220 21539 9222
rect 21563 9220 21619 9222
rect 21643 9220 21699 9222
rect 21723 9220 21779 9222
rect 21483 8186 21539 8188
rect 21563 8186 21619 8188
rect 21643 8186 21699 8188
rect 21723 8186 21779 8188
rect 21483 8134 21529 8186
rect 21529 8134 21539 8186
rect 21563 8134 21593 8186
rect 21593 8134 21605 8186
rect 21605 8134 21619 8186
rect 21643 8134 21657 8186
rect 21657 8134 21669 8186
rect 21669 8134 21699 8186
rect 21723 8134 21733 8186
rect 21733 8134 21779 8186
rect 21483 8132 21539 8134
rect 21563 8132 21619 8134
rect 21643 8132 21699 8134
rect 21723 8132 21779 8134
rect 21086 6568 21142 6624
rect 20902 3984 20958 4040
rect 20902 3168 20958 3224
rect 20626 2524 20628 2544
rect 20628 2524 20680 2544
rect 20680 2524 20682 2544
rect 20626 2488 20682 2524
rect 20718 1128 20774 1184
rect 21483 7098 21539 7100
rect 21563 7098 21619 7100
rect 21643 7098 21699 7100
rect 21723 7098 21779 7100
rect 21483 7046 21529 7098
rect 21529 7046 21539 7098
rect 21563 7046 21593 7098
rect 21593 7046 21605 7098
rect 21605 7046 21619 7098
rect 21643 7046 21657 7098
rect 21657 7046 21669 7098
rect 21669 7046 21699 7098
rect 21723 7046 21733 7098
rect 21733 7046 21779 7098
rect 21483 7044 21539 7046
rect 21563 7044 21619 7046
rect 21643 7044 21699 7046
rect 21723 7044 21779 7046
rect 21086 4392 21142 4448
rect 21546 6160 21602 6216
rect 21483 6010 21539 6012
rect 21563 6010 21619 6012
rect 21643 6010 21699 6012
rect 21723 6010 21779 6012
rect 21483 5958 21529 6010
rect 21529 5958 21539 6010
rect 21563 5958 21593 6010
rect 21593 5958 21605 6010
rect 21605 5958 21619 6010
rect 21643 5958 21657 6010
rect 21657 5958 21669 6010
rect 21669 5958 21699 6010
rect 21723 5958 21733 6010
rect 21733 5958 21779 6010
rect 21483 5956 21539 5958
rect 21563 5956 21619 5958
rect 21643 5956 21699 5958
rect 21723 5956 21779 5958
rect 21483 4922 21539 4924
rect 21563 4922 21619 4924
rect 21643 4922 21699 4924
rect 21723 4922 21779 4924
rect 21483 4870 21529 4922
rect 21529 4870 21539 4922
rect 21563 4870 21593 4922
rect 21593 4870 21605 4922
rect 21605 4870 21619 4922
rect 21643 4870 21657 4922
rect 21657 4870 21669 4922
rect 21669 4870 21699 4922
rect 21723 4870 21733 4922
rect 21733 4870 21779 4922
rect 21483 4868 21539 4870
rect 21563 4868 21619 4870
rect 21643 4868 21699 4870
rect 21723 4868 21779 4870
rect 22190 5344 22246 5400
rect 21638 4664 21694 4720
rect 20994 2896 21050 2952
rect 21086 2352 21142 2408
rect 21483 3834 21539 3836
rect 21563 3834 21619 3836
rect 21643 3834 21699 3836
rect 21723 3834 21779 3836
rect 21483 3782 21529 3834
rect 21529 3782 21539 3834
rect 21563 3782 21593 3834
rect 21593 3782 21605 3834
rect 21605 3782 21619 3834
rect 21643 3782 21657 3834
rect 21657 3782 21669 3834
rect 21669 3782 21699 3834
rect 21723 3782 21733 3834
rect 21733 3782 21779 3834
rect 21483 3780 21539 3782
rect 21563 3780 21619 3782
rect 21643 3780 21699 3782
rect 21723 3780 21779 3782
rect 21638 3304 21694 3360
rect 21483 2746 21539 2748
rect 21563 2746 21619 2748
rect 21643 2746 21699 2748
rect 21723 2746 21779 2748
rect 21483 2694 21529 2746
rect 21529 2694 21539 2746
rect 21563 2694 21593 2746
rect 21593 2694 21605 2746
rect 21605 2694 21619 2746
rect 21643 2694 21657 2746
rect 21657 2694 21669 2746
rect 21669 2694 21699 2746
rect 21723 2694 21733 2746
rect 21733 2694 21779 2746
rect 21483 2692 21539 2694
rect 21563 2692 21619 2694
rect 21643 2692 21699 2694
rect 21723 2692 21779 2694
rect 21822 2488 21878 2544
rect 21546 1844 21548 1864
rect 21548 1844 21600 1864
rect 21600 1844 21602 1864
rect 21546 1808 21602 1844
rect 21483 1658 21539 1660
rect 21563 1658 21619 1660
rect 21643 1658 21699 1660
rect 21723 1658 21779 1660
rect 21483 1606 21529 1658
rect 21529 1606 21539 1658
rect 21563 1606 21593 1658
rect 21593 1606 21605 1658
rect 21605 1606 21619 1658
rect 21643 1606 21657 1658
rect 21657 1606 21669 1658
rect 21669 1606 21699 1658
rect 21723 1606 21733 1658
rect 21733 1606 21779 1658
rect 21483 1604 21539 1606
rect 21563 1604 21619 1606
rect 21643 1604 21699 1606
rect 21723 1604 21779 1606
rect 22466 5788 22468 5808
rect 22468 5788 22520 5808
rect 22520 5788 22522 5808
rect 22466 5752 22522 5788
rect 22190 3576 22246 3632
rect 22282 3440 22338 3496
rect 22190 2624 22246 2680
rect 22006 1672 22062 1728
rect 22190 2352 22246 2408
rect 22742 3848 22798 3904
rect 23570 18028 23572 18048
rect 23572 18028 23624 18048
rect 23624 18028 23626 18048
rect 23570 17992 23626 18028
rect 23570 16940 23572 16960
rect 23572 16940 23624 16960
rect 23624 16940 23626 16960
rect 23570 16904 23626 16940
rect 24122 23468 24124 23488
rect 24124 23468 24176 23488
rect 24176 23468 24178 23488
rect 24122 23432 24178 23468
rect 23754 22380 23756 22400
rect 23756 22380 23808 22400
rect 23808 22380 23810 22400
rect 23754 22344 23810 22380
rect 24122 21292 24124 21312
rect 24124 21292 24176 21312
rect 24176 21292 24178 21312
rect 23754 20168 23810 20224
rect 24122 21256 24178 21292
rect 23938 19116 23940 19136
rect 23940 19116 23992 19136
rect 23992 19116 23994 19136
rect 23938 19080 23994 19116
rect 23754 15852 23756 15872
rect 23756 15852 23808 15872
rect 23808 15852 23810 15872
rect 23754 15816 23810 15852
rect 24122 14764 24124 14784
rect 24124 14764 24176 14784
rect 24176 14764 24178 14784
rect 24122 14728 24178 14764
rect 24122 13640 24178 13696
rect 23938 12588 23940 12608
rect 23940 12588 23992 12608
rect 23992 12588 23994 12608
rect 23938 12552 23994 12588
rect 24858 38156 24860 38176
rect 24860 38156 24912 38176
rect 24912 38156 24914 38176
rect 24858 38120 24914 38156
rect 24415 38106 24471 38108
rect 24495 38106 24551 38108
rect 24575 38106 24631 38108
rect 24655 38106 24711 38108
rect 24415 38054 24461 38106
rect 24461 38054 24471 38106
rect 24495 38054 24525 38106
rect 24525 38054 24537 38106
rect 24537 38054 24551 38106
rect 24575 38054 24589 38106
rect 24589 38054 24601 38106
rect 24601 38054 24631 38106
rect 24655 38054 24665 38106
rect 24665 38054 24711 38106
rect 24415 38052 24471 38054
rect 24495 38052 24551 38054
rect 24575 38052 24631 38054
rect 24655 38052 24711 38054
rect 24858 37068 24860 37088
rect 24860 37068 24912 37088
rect 24912 37068 24914 37088
rect 24858 37032 24914 37068
rect 24415 37018 24471 37020
rect 24495 37018 24551 37020
rect 24575 37018 24631 37020
rect 24655 37018 24711 37020
rect 24415 36966 24461 37018
rect 24461 36966 24471 37018
rect 24495 36966 24525 37018
rect 24525 36966 24537 37018
rect 24537 36966 24551 37018
rect 24575 36966 24589 37018
rect 24589 36966 24601 37018
rect 24601 36966 24631 37018
rect 24655 36966 24665 37018
rect 24665 36966 24711 37018
rect 24415 36964 24471 36966
rect 24495 36964 24551 36966
rect 24575 36964 24631 36966
rect 24655 36964 24711 36966
rect 24415 35930 24471 35932
rect 24495 35930 24551 35932
rect 24575 35930 24631 35932
rect 24655 35930 24711 35932
rect 24415 35878 24461 35930
rect 24461 35878 24471 35930
rect 24495 35878 24525 35930
rect 24525 35878 24537 35930
rect 24537 35878 24551 35930
rect 24575 35878 24589 35930
rect 24589 35878 24601 35930
rect 24601 35878 24631 35930
rect 24655 35878 24665 35930
rect 24665 35878 24711 35930
rect 24415 35876 24471 35878
rect 24495 35876 24551 35878
rect 24575 35876 24631 35878
rect 24655 35876 24711 35878
rect 24415 34842 24471 34844
rect 24495 34842 24551 34844
rect 24575 34842 24631 34844
rect 24655 34842 24711 34844
rect 24415 34790 24461 34842
rect 24461 34790 24471 34842
rect 24495 34790 24525 34842
rect 24525 34790 24537 34842
rect 24537 34790 24551 34842
rect 24575 34790 24589 34842
rect 24589 34790 24601 34842
rect 24601 34790 24631 34842
rect 24655 34790 24665 34842
rect 24665 34790 24711 34842
rect 24415 34788 24471 34790
rect 24495 34788 24551 34790
rect 24575 34788 24631 34790
rect 24655 34788 24711 34790
rect 24415 33754 24471 33756
rect 24495 33754 24551 33756
rect 24575 33754 24631 33756
rect 24655 33754 24711 33756
rect 24415 33702 24461 33754
rect 24461 33702 24471 33754
rect 24495 33702 24525 33754
rect 24525 33702 24537 33754
rect 24537 33702 24551 33754
rect 24575 33702 24589 33754
rect 24589 33702 24601 33754
rect 24601 33702 24631 33754
rect 24655 33702 24665 33754
rect 24665 33702 24711 33754
rect 24415 33700 24471 33702
rect 24495 33700 24551 33702
rect 24575 33700 24631 33702
rect 24655 33700 24711 33702
rect 24415 32666 24471 32668
rect 24495 32666 24551 32668
rect 24575 32666 24631 32668
rect 24655 32666 24711 32668
rect 24415 32614 24461 32666
rect 24461 32614 24471 32666
rect 24495 32614 24525 32666
rect 24525 32614 24537 32666
rect 24537 32614 24551 32666
rect 24575 32614 24589 32666
rect 24589 32614 24601 32666
rect 24601 32614 24631 32666
rect 24655 32614 24665 32666
rect 24665 32614 24711 32666
rect 24415 32612 24471 32614
rect 24495 32612 24551 32614
rect 24575 32612 24631 32614
rect 24655 32612 24711 32614
rect 24415 31578 24471 31580
rect 24495 31578 24551 31580
rect 24575 31578 24631 31580
rect 24655 31578 24711 31580
rect 24415 31526 24461 31578
rect 24461 31526 24471 31578
rect 24495 31526 24525 31578
rect 24525 31526 24537 31578
rect 24537 31526 24551 31578
rect 24575 31526 24589 31578
rect 24589 31526 24601 31578
rect 24601 31526 24631 31578
rect 24655 31526 24665 31578
rect 24665 31526 24711 31578
rect 24415 31524 24471 31526
rect 24495 31524 24551 31526
rect 24575 31524 24631 31526
rect 24655 31524 24711 31526
rect 24415 30490 24471 30492
rect 24495 30490 24551 30492
rect 24575 30490 24631 30492
rect 24655 30490 24711 30492
rect 24415 30438 24461 30490
rect 24461 30438 24471 30490
rect 24495 30438 24525 30490
rect 24525 30438 24537 30490
rect 24537 30438 24551 30490
rect 24575 30438 24589 30490
rect 24589 30438 24601 30490
rect 24601 30438 24631 30490
rect 24655 30438 24665 30490
rect 24665 30438 24711 30490
rect 24415 30436 24471 30438
rect 24495 30436 24551 30438
rect 24575 30436 24631 30438
rect 24655 30436 24711 30438
rect 24415 29402 24471 29404
rect 24495 29402 24551 29404
rect 24575 29402 24631 29404
rect 24655 29402 24711 29404
rect 24415 29350 24461 29402
rect 24461 29350 24471 29402
rect 24495 29350 24525 29402
rect 24525 29350 24537 29402
rect 24537 29350 24551 29402
rect 24575 29350 24589 29402
rect 24589 29350 24601 29402
rect 24601 29350 24631 29402
rect 24655 29350 24665 29402
rect 24665 29350 24711 29402
rect 24415 29348 24471 29350
rect 24495 29348 24551 29350
rect 24575 29348 24631 29350
rect 24655 29348 24711 29350
rect 24415 28314 24471 28316
rect 24495 28314 24551 28316
rect 24575 28314 24631 28316
rect 24655 28314 24711 28316
rect 24415 28262 24461 28314
rect 24461 28262 24471 28314
rect 24495 28262 24525 28314
rect 24525 28262 24537 28314
rect 24537 28262 24551 28314
rect 24575 28262 24589 28314
rect 24589 28262 24601 28314
rect 24601 28262 24631 28314
rect 24655 28262 24665 28314
rect 24665 28262 24711 28314
rect 24415 28260 24471 28262
rect 24495 28260 24551 28262
rect 24575 28260 24631 28262
rect 24655 28260 24711 28262
rect 24415 27226 24471 27228
rect 24495 27226 24551 27228
rect 24575 27226 24631 27228
rect 24655 27226 24711 27228
rect 24415 27174 24461 27226
rect 24461 27174 24471 27226
rect 24495 27174 24525 27226
rect 24525 27174 24537 27226
rect 24537 27174 24551 27226
rect 24575 27174 24589 27226
rect 24589 27174 24601 27226
rect 24601 27174 24631 27226
rect 24655 27174 24665 27226
rect 24665 27174 24711 27226
rect 24415 27172 24471 27174
rect 24495 27172 24551 27174
rect 24575 27172 24631 27174
rect 24655 27172 24711 27174
rect 24415 26138 24471 26140
rect 24495 26138 24551 26140
rect 24575 26138 24631 26140
rect 24655 26138 24711 26140
rect 24415 26086 24461 26138
rect 24461 26086 24471 26138
rect 24495 26086 24525 26138
rect 24525 26086 24537 26138
rect 24537 26086 24551 26138
rect 24575 26086 24589 26138
rect 24589 26086 24601 26138
rect 24601 26086 24631 26138
rect 24655 26086 24665 26138
rect 24665 26086 24711 26138
rect 24415 26084 24471 26086
rect 24495 26084 24551 26086
rect 24575 26084 24631 26086
rect 24655 26084 24711 26086
rect 24415 25050 24471 25052
rect 24495 25050 24551 25052
rect 24575 25050 24631 25052
rect 24655 25050 24711 25052
rect 24415 24998 24461 25050
rect 24461 24998 24471 25050
rect 24495 24998 24525 25050
rect 24525 24998 24537 25050
rect 24537 24998 24551 25050
rect 24575 24998 24589 25050
rect 24589 24998 24601 25050
rect 24601 24998 24631 25050
rect 24655 24998 24665 25050
rect 24665 24998 24711 25050
rect 24415 24996 24471 24998
rect 24495 24996 24551 24998
rect 24575 24996 24631 24998
rect 24655 24996 24711 24998
rect 24415 23962 24471 23964
rect 24495 23962 24551 23964
rect 24575 23962 24631 23964
rect 24655 23962 24711 23964
rect 24415 23910 24461 23962
rect 24461 23910 24471 23962
rect 24495 23910 24525 23962
rect 24525 23910 24537 23962
rect 24537 23910 24551 23962
rect 24575 23910 24589 23962
rect 24589 23910 24601 23962
rect 24601 23910 24631 23962
rect 24655 23910 24665 23962
rect 24665 23910 24711 23962
rect 24415 23908 24471 23910
rect 24495 23908 24551 23910
rect 24575 23908 24631 23910
rect 24655 23908 24711 23910
rect 24415 22874 24471 22876
rect 24495 22874 24551 22876
rect 24575 22874 24631 22876
rect 24655 22874 24711 22876
rect 24415 22822 24461 22874
rect 24461 22822 24471 22874
rect 24495 22822 24525 22874
rect 24525 22822 24537 22874
rect 24537 22822 24551 22874
rect 24575 22822 24589 22874
rect 24589 22822 24601 22874
rect 24601 22822 24631 22874
rect 24655 22822 24665 22874
rect 24665 22822 24711 22874
rect 24415 22820 24471 22822
rect 24495 22820 24551 22822
rect 24575 22820 24631 22822
rect 24655 22820 24711 22822
rect 24415 21786 24471 21788
rect 24495 21786 24551 21788
rect 24575 21786 24631 21788
rect 24655 21786 24711 21788
rect 24415 21734 24461 21786
rect 24461 21734 24471 21786
rect 24495 21734 24525 21786
rect 24525 21734 24537 21786
rect 24537 21734 24551 21786
rect 24575 21734 24589 21786
rect 24589 21734 24601 21786
rect 24601 21734 24631 21786
rect 24655 21734 24665 21786
rect 24665 21734 24711 21786
rect 24415 21732 24471 21734
rect 24495 21732 24551 21734
rect 24575 21732 24631 21734
rect 24655 21732 24711 21734
rect 24415 20698 24471 20700
rect 24495 20698 24551 20700
rect 24575 20698 24631 20700
rect 24655 20698 24711 20700
rect 24415 20646 24461 20698
rect 24461 20646 24471 20698
rect 24495 20646 24525 20698
rect 24525 20646 24537 20698
rect 24537 20646 24551 20698
rect 24575 20646 24589 20698
rect 24589 20646 24601 20698
rect 24601 20646 24631 20698
rect 24655 20646 24665 20698
rect 24665 20646 24711 20698
rect 24415 20644 24471 20646
rect 24495 20644 24551 20646
rect 24575 20644 24631 20646
rect 24655 20644 24711 20646
rect 24415 19610 24471 19612
rect 24495 19610 24551 19612
rect 24575 19610 24631 19612
rect 24655 19610 24711 19612
rect 24415 19558 24461 19610
rect 24461 19558 24471 19610
rect 24495 19558 24525 19610
rect 24525 19558 24537 19610
rect 24537 19558 24551 19610
rect 24575 19558 24589 19610
rect 24589 19558 24601 19610
rect 24601 19558 24631 19610
rect 24655 19558 24665 19610
rect 24665 19558 24711 19610
rect 24415 19556 24471 19558
rect 24495 19556 24551 19558
rect 24575 19556 24631 19558
rect 24655 19556 24711 19558
rect 24415 18522 24471 18524
rect 24495 18522 24551 18524
rect 24575 18522 24631 18524
rect 24655 18522 24711 18524
rect 24415 18470 24461 18522
rect 24461 18470 24471 18522
rect 24495 18470 24525 18522
rect 24525 18470 24537 18522
rect 24537 18470 24551 18522
rect 24575 18470 24589 18522
rect 24589 18470 24601 18522
rect 24601 18470 24631 18522
rect 24655 18470 24665 18522
rect 24665 18470 24711 18522
rect 24415 18468 24471 18470
rect 24495 18468 24551 18470
rect 24575 18468 24631 18470
rect 24655 18468 24711 18470
rect 24415 17434 24471 17436
rect 24495 17434 24551 17436
rect 24575 17434 24631 17436
rect 24655 17434 24711 17436
rect 24415 17382 24461 17434
rect 24461 17382 24471 17434
rect 24495 17382 24525 17434
rect 24525 17382 24537 17434
rect 24537 17382 24551 17434
rect 24575 17382 24589 17434
rect 24589 17382 24601 17434
rect 24601 17382 24631 17434
rect 24655 17382 24665 17434
rect 24665 17382 24711 17434
rect 24415 17380 24471 17382
rect 24495 17380 24551 17382
rect 24575 17380 24631 17382
rect 24655 17380 24711 17382
rect 24415 16346 24471 16348
rect 24495 16346 24551 16348
rect 24575 16346 24631 16348
rect 24655 16346 24711 16348
rect 24415 16294 24461 16346
rect 24461 16294 24471 16346
rect 24495 16294 24525 16346
rect 24525 16294 24537 16346
rect 24537 16294 24551 16346
rect 24575 16294 24589 16346
rect 24589 16294 24601 16346
rect 24601 16294 24631 16346
rect 24655 16294 24665 16346
rect 24665 16294 24711 16346
rect 24415 16292 24471 16294
rect 24495 16292 24551 16294
rect 24575 16292 24631 16294
rect 24655 16292 24711 16294
rect 24415 15258 24471 15260
rect 24495 15258 24551 15260
rect 24575 15258 24631 15260
rect 24655 15258 24711 15260
rect 24415 15206 24461 15258
rect 24461 15206 24471 15258
rect 24495 15206 24525 15258
rect 24525 15206 24537 15258
rect 24537 15206 24551 15258
rect 24575 15206 24589 15258
rect 24589 15206 24601 15258
rect 24601 15206 24631 15258
rect 24655 15206 24665 15258
rect 24665 15206 24711 15258
rect 24415 15204 24471 15206
rect 24495 15204 24551 15206
rect 24575 15204 24631 15206
rect 24655 15204 24711 15206
rect 24415 14170 24471 14172
rect 24495 14170 24551 14172
rect 24575 14170 24631 14172
rect 24655 14170 24711 14172
rect 24415 14118 24461 14170
rect 24461 14118 24471 14170
rect 24495 14118 24525 14170
rect 24525 14118 24537 14170
rect 24537 14118 24551 14170
rect 24575 14118 24589 14170
rect 24589 14118 24601 14170
rect 24601 14118 24631 14170
rect 24655 14118 24665 14170
rect 24665 14118 24711 14170
rect 24415 14116 24471 14118
rect 24495 14116 24551 14118
rect 24575 14116 24631 14118
rect 24655 14116 24711 14118
rect 24415 13082 24471 13084
rect 24495 13082 24551 13084
rect 24575 13082 24631 13084
rect 24655 13082 24711 13084
rect 24415 13030 24461 13082
rect 24461 13030 24471 13082
rect 24495 13030 24525 13082
rect 24525 13030 24537 13082
rect 24537 13030 24551 13082
rect 24575 13030 24589 13082
rect 24589 13030 24601 13082
rect 24601 13030 24631 13082
rect 24655 13030 24665 13082
rect 24665 13030 24711 13082
rect 24415 13028 24471 13030
rect 24495 13028 24551 13030
rect 24575 13028 24631 13030
rect 24655 13028 24711 13030
rect 24030 11464 24086 11520
rect 23386 8780 23388 8800
rect 23388 8780 23440 8800
rect 23440 8780 23442 8800
rect 23386 8744 23442 8780
rect 23570 8916 23572 8936
rect 23572 8916 23624 8936
rect 23624 8916 23626 8936
rect 23570 8880 23626 8916
rect 24122 9288 24178 9344
rect 24415 11994 24471 11996
rect 24495 11994 24551 11996
rect 24575 11994 24631 11996
rect 24655 11994 24711 11996
rect 24415 11942 24461 11994
rect 24461 11942 24471 11994
rect 24495 11942 24525 11994
rect 24525 11942 24537 11994
rect 24537 11942 24551 11994
rect 24575 11942 24589 11994
rect 24589 11942 24601 11994
rect 24601 11942 24631 11994
rect 24655 11942 24665 11994
rect 24665 11942 24711 11994
rect 24415 11940 24471 11942
rect 24495 11940 24551 11942
rect 24575 11940 24631 11942
rect 24655 11940 24711 11942
rect 24214 8200 24270 8256
rect 23110 5480 23166 5536
rect 22374 584 22430 640
rect 23386 5480 23442 5536
rect 24030 7828 24032 7848
rect 24032 7828 24084 7848
rect 24084 7828 24086 7848
rect 23846 6840 23902 6896
rect 24030 7792 24086 7828
rect 24030 7540 24086 7576
rect 24030 7520 24032 7540
rect 24032 7520 24084 7540
rect 24084 7520 24086 7540
rect 24030 7112 24086 7168
rect 23846 5616 23902 5672
rect 24415 10906 24471 10908
rect 24495 10906 24551 10908
rect 24575 10906 24631 10908
rect 24655 10906 24711 10908
rect 24415 10854 24461 10906
rect 24461 10854 24471 10906
rect 24495 10854 24525 10906
rect 24525 10854 24537 10906
rect 24537 10854 24551 10906
rect 24575 10854 24589 10906
rect 24589 10854 24601 10906
rect 24601 10854 24631 10906
rect 24655 10854 24665 10906
rect 24665 10854 24711 10906
rect 24415 10852 24471 10854
rect 24495 10852 24551 10854
rect 24575 10852 24631 10854
rect 24655 10852 24711 10854
rect 24415 9818 24471 9820
rect 24495 9818 24551 9820
rect 24575 9818 24631 9820
rect 24655 9818 24711 9820
rect 24415 9766 24461 9818
rect 24461 9766 24471 9818
rect 24495 9766 24525 9818
rect 24525 9766 24537 9818
rect 24537 9766 24551 9818
rect 24575 9766 24589 9818
rect 24589 9766 24601 9818
rect 24601 9766 24631 9818
rect 24655 9766 24665 9818
rect 24665 9766 24711 9818
rect 24415 9764 24471 9766
rect 24495 9764 24551 9766
rect 24575 9764 24631 9766
rect 24655 9764 24711 9766
rect 24415 8730 24471 8732
rect 24495 8730 24551 8732
rect 24575 8730 24631 8732
rect 24655 8730 24711 8732
rect 24415 8678 24461 8730
rect 24461 8678 24471 8730
rect 24495 8678 24525 8730
rect 24525 8678 24537 8730
rect 24537 8678 24551 8730
rect 24575 8678 24589 8730
rect 24589 8678 24601 8730
rect 24601 8678 24631 8730
rect 24655 8678 24665 8730
rect 24665 8678 24711 8730
rect 24415 8676 24471 8678
rect 24495 8676 24551 8678
rect 24575 8676 24631 8678
rect 24655 8676 24711 8678
rect 24415 7642 24471 7644
rect 24495 7642 24551 7644
rect 24575 7642 24631 7644
rect 24655 7642 24711 7644
rect 24415 7590 24461 7642
rect 24461 7590 24471 7642
rect 24495 7590 24525 7642
rect 24525 7590 24537 7642
rect 24537 7590 24551 7642
rect 24575 7590 24589 7642
rect 24589 7590 24601 7642
rect 24601 7590 24631 7642
rect 24655 7590 24665 7642
rect 24665 7590 24711 7642
rect 24415 7588 24471 7590
rect 24495 7588 24551 7590
rect 24575 7588 24631 7590
rect 24655 7588 24711 7590
rect 24415 6554 24471 6556
rect 24495 6554 24551 6556
rect 24575 6554 24631 6556
rect 24655 6554 24711 6556
rect 24415 6502 24461 6554
rect 24461 6502 24471 6554
rect 24495 6502 24525 6554
rect 24525 6502 24537 6554
rect 24537 6502 24551 6554
rect 24575 6502 24589 6554
rect 24589 6502 24601 6554
rect 24601 6502 24631 6554
rect 24655 6502 24665 6554
rect 24665 6502 24711 6554
rect 24415 6500 24471 6502
rect 24495 6500 24551 6502
rect 24575 6500 24631 6502
rect 24655 6500 24711 6502
rect 24030 4936 24086 4992
rect 24415 5466 24471 5468
rect 24495 5466 24551 5468
rect 24575 5466 24631 5468
rect 24655 5466 24711 5468
rect 24415 5414 24461 5466
rect 24461 5414 24471 5466
rect 24495 5414 24525 5466
rect 24525 5414 24537 5466
rect 24537 5414 24551 5466
rect 24575 5414 24589 5466
rect 24589 5414 24601 5466
rect 24601 5414 24631 5466
rect 24655 5414 24665 5466
rect 24665 5414 24711 5466
rect 24415 5412 24471 5414
rect 24495 5412 24551 5414
rect 24575 5412 24631 5414
rect 24655 5412 24711 5414
rect 24306 4528 24362 4584
rect 24415 4378 24471 4380
rect 24495 4378 24551 4380
rect 24575 4378 24631 4380
rect 24655 4378 24711 4380
rect 24415 4326 24461 4378
rect 24461 4326 24471 4378
rect 24495 4326 24525 4378
rect 24525 4326 24537 4378
rect 24537 4326 24551 4378
rect 24575 4326 24589 4378
rect 24589 4326 24601 4378
rect 24601 4326 24631 4378
rect 24655 4326 24665 4378
rect 24665 4326 24711 4378
rect 24415 4324 24471 4326
rect 24495 4324 24551 4326
rect 24575 4324 24631 4326
rect 24655 4324 24711 4326
rect 23754 3032 23810 3088
rect 24415 3290 24471 3292
rect 24495 3290 24551 3292
rect 24575 3290 24631 3292
rect 24655 3290 24711 3292
rect 24415 3238 24461 3290
rect 24461 3238 24471 3290
rect 24495 3238 24525 3290
rect 24525 3238 24537 3290
rect 24537 3238 24551 3290
rect 24575 3238 24589 3290
rect 24589 3238 24601 3290
rect 24601 3238 24631 3290
rect 24655 3238 24665 3290
rect 24665 3238 24711 3290
rect 24415 3236 24471 3238
rect 24495 3236 24551 3238
rect 24575 3236 24631 3238
rect 24655 3236 24711 3238
rect 24950 35944 25006 36000
rect 24858 34892 24860 34912
rect 24860 34892 24912 34912
rect 24912 34892 24914 34912
rect 24858 34856 24914 34892
rect 24858 33804 24860 33824
rect 24860 33804 24912 33824
rect 24912 33804 24914 33824
rect 24858 33768 24914 33804
rect 24858 32716 24860 32736
rect 24860 32716 24912 32736
rect 24912 32716 24914 32736
rect 24858 32680 24914 32716
rect 24858 30504 24914 30560
rect 24858 29452 24860 29472
rect 24860 29452 24912 29472
rect 24912 29452 24914 29472
rect 24858 29416 24914 29452
rect 24858 28364 24860 28384
rect 24860 28364 24912 28384
rect 24912 28364 24914 28384
rect 24858 28328 24914 28364
rect 24858 27276 24860 27296
rect 24860 27276 24912 27296
rect 24912 27276 24914 27296
rect 24858 27240 24914 27276
rect 24858 26152 24914 26208
rect 24858 25064 24914 25120
rect 24858 24012 24860 24032
rect 24860 24012 24912 24032
rect 24912 24012 24914 24032
rect 24858 23976 24914 24012
rect 24858 22888 24914 22944
rect 24858 21836 24860 21856
rect 24860 21836 24912 21856
rect 24912 21836 24914 21856
rect 24858 21800 24914 21836
rect 24858 20712 24914 20768
rect 24858 18536 24914 18592
rect 24858 17448 24914 17504
rect 24858 16360 24914 16416
rect 24858 15272 24914 15328
rect 24858 14220 24860 14240
rect 24860 14220 24912 14240
rect 24912 14220 24914 14240
rect 24858 14184 24914 14220
rect 24858 13096 24914 13152
rect 24858 12008 24914 12064
rect 24858 10920 24914 10976
rect 24858 9832 24914 9888
rect 24858 6568 24914 6624
rect 25042 31592 25098 31648
rect 25134 19624 25190 19680
rect 25134 10376 25190 10432
rect 24415 2202 24471 2204
rect 24495 2202 24551 2204
rect 24575 2202 24631 2204
rect 24655 2202 24711 2204
rect 24415 2150 24461 2202
rect 24461 2150 24471 2202
rect 24495 2150 24525 2202
rect 24525 2150 24537 2202
rect 24537 2150 24551 2202
rect 24575 2150 24589 2202
rect 24589 2150 24601 2202
rect 24601 2150 24631 2202
rect 24655 2150 24665 2202
rect 24665 2150 24711 2202
rect 24415 2148 24471 2150
rect 24495 2148 24551 2150
rect 24575 2148 24631 2150
rect 24655 2148 24711 2150
rect 24415 1114 24471 1116
rect 24495 1114 24551 1116
rect 24575 1114 24631 1116
rect 24655 1114 24711 1116
rect 24415 1062 24461 1114
rect 24461 1062 24471 1114
rect 24495 1062 24525 1114
rect 24525 1062 24537 1114
rect 24537 1062 24551 1114
rect 24575 1062 24589 1114
rect 24589 1062 24601 1114
rect 24601 1062 24631 1114
rect 24655 1062 24665 1114
rect 24665 1062 24711 1114
rect 24415 1060 24471 1062
rect 24495 1060 24551 1062
rect 24575 1060 24631 1062
rect 24655 1060 24711 1062
<< metal3 >>
rect 22001 43754 22067 43757
rect 22001 43752 24962 43754
rect 22001 43696 22006 43752
rect 22062 43696 24962 43752
rect 22001 43694 24962 43696
rect 22001 43691 22067 43694
rect 24902 43618 24962 43694
rect 25540 43618 26000 43648
rect 24902 43558 26000 43618
rect 6810 43552 7126 43553
rect 6810 43488 6816 43552
rect 6880 43488 6896 43552
rect 6960 43488 6976 43552
rect 7040 43488 7056 43552
rect 7120 43488 7126 43552
rect 6810 43487 7126 43488
rect 12675 43552 12991 43553
rect 12675 43488 12681 43552
rect 12745 43488 12761 43552
rect 12825 43488 12841 43552
rect 12905 43488 12921 43552
rect 12985 43488 12991 43552
rect 12675 43487 12991 43488
rect 18540 43552 18856 43553
rect 18540 43488 18546 43552
rect 18610 43488 18626 43552
rect 18690 43488 18706 43552
rect 18770 43488 18786 43552
rect 18850 43488 18856 43552
rect 18540 43487 18856 43488
rect 24405 43552 24721 43553
rect 24405 43488 24411 43552
rect 24475 43488 24491 43552
rect 24555 43488 24571 43552
rect 24635 43488 24651 43552
rect 24715 43488 24721 43552
rect 25540 43528 26000 43558
rect 24405 43487 24721 43488
rect 1761 43210 1827 43213
rect 5901 43210 5967 43213
rect 1761 43208 5967 43210
rect 1761 43152 1766 43208
rect 1822 43152 5906 43208
rect 5962 43152 5967 43208
rect 1761 43150 5967 43152
rect 1761 43147 1827 43150
rect 5901 43147 5967 43150
rect 9673 43210 9739 43213
rect 21265 43210 21331 43213
rect 21950 43210 21956 43212
rect 9673 43208 10196 43210
rect 9673 43152 9678 43208
rect 9734 43152 10196 43208
rect 9673 43150 10196 43152
rect 9673 43147 9739 43150
rect 3878 43008 4194 43009
rect 3878 42944 3884 43008
rect 3948 42944 3964 43008
rect 4028 42944 4044 43008
rect 4108 42944 4124 43008
rect 4188 42944 4194 43008
rect 3878 42943 4194 42944
rect 9743 43008 10059 43009
rect 9743 42944 9749 43008
rect 9813 42944 9829 43008
rect 9893 42944 9909 43008
rect 9973 42944 9989 43008
rect 10053 42944 10059 43008
rect 9743 42943 10059 42944
rect 974 42740 980 42804
rect 1044 42802 1050 42804
rect 3969 42802 4035 42805
rect 1044 42800 4035 42802
rect 1044 42744 3974 42800
rect 4030 42744 4035 42800
rect 1044 42742 4035 42744
rect 1044 42740 1050 42742
rect 3969 42739 4035 42742
rect 5717 42802 5783 42805
rect 6729 42802 6795 42805
rect 5717 42800 6795 42802
rect 5717 42744 5722 42800
rect 5778 42744 6734 42800
rect 6790 42744 6795 42800
rect 5717 42742 6795 42744
rect 5717 42739 5783 42742
rect 6729 42739 6795 42742
rect 9949 42802 10015 42805
rect 10136 42802 10196 43150
rect 21265 43208 21956 43210
rect 21265 43152 21270 43208
rect 21326 43152 21956 43208
rect 21265 43150 21956 43152
rect 21265 43147 21331 43150
rect 21950 43148 21956 43150
rect 22020 43148 22026 43212
rect 11646 43012 11652 43076
rect 11716 43074 11722 43076
rect 12525 43074 12591 43077
rect 11716 43072 12591 43074
rect 11716 43016 12530 43072
rect 12586 43016 12591 43072
rect 11716 43014 12591 43016
rect 11716 43012 11722 43014
rect 12525 43011 12591 43014
rect 22921 43074 22987 43077
rect 25540 43074 26000 43104
rect 22921 43072 26000 43074
rect 22921 43016 22926 43072
rect 22982 43016 26000 43072
rect 22921 43014 26000 43016
rect 22921 43011 22987 43014
rect 15608 43008 15924 43009
rect 15608 42944 15614 43008
rect 15678 42944 15694 43008
rect 15758 42944 15774 43008
rect 15838 42944 15854 43008
rect 15918 42944 15924 43008
rect 15608 42943 15924 42944
rect 21473 43008 21789 43009
rect 21473 42944 21479 43008
rect 21543 42944 21559 43008
rect 21623 42944 21639 43008
rect 21703 42944 21719 43008
rect 21783 42944 21789 43008
rect 25540 42984 26000 43014
rect 21473 42943 21789 42944
rect 11789 42940 11855 42941
rect 15009 42940 15075 42941
rect 11789 42936 11836 42940
rect 11900 42938 11906 42940
rect 14958 42938 14964 42940
rect 11789 42880 11794 42936
rect 11789 42876 11836 42880
rect 11900 42878 11946 42938
rect 14918 42878 14964 42938
rect 15028 42936 15075 42940
rect 15070 42880 15075 42936
rect 11900 42876 11906 42878
rect 14958 42876 14964 42878
rect 15028 42876 15075 42880
rect 15326 42876 15332 42940
rect 15396 42938 15402 42940
rect 15469 42938 15535 42941
rect 15396 42936 15535 42938
rect 15396 42880 15474 42936
rect 15530 42880 15535 42936
rect 15396 42878 15535 42880
rect 15396 42876 15402 42878
rect 11789 42875 11855 42876
rect 15009 42875 15075 42876
rect 15469 42875 15535 42878
rect 17585 42938 17651 42941
rect 17718 42938 17724 42940
rect 17585 42936 17724 42938
rect 17585 42880 17590 42936
rect 17646 42880 17724 42936
rect 17585 42878 17724 42880
rect 17585 42875 17651 42878
rect 17718 42876 17724 42878
rect 17788 42876 17794 42940
rect 9949 42800 10196 42802
rect 9949 42744 9954 42800
rect 10010 42744 10196 42800
rect 9949 42742 10196 42744
rect 9949 42739 10015 42742
rect 2681 42666 2747 42669
rect 16614 42666 16620 42668
rect 2681 42664 16620 42666
rect 2681 42608 2686 42664
rect 2742 42608 16620 42664
rect 2681 42606 16620 42608
rect 2681 42603 2747 42606
rect 16614 42604 16620 42606
rect 16684 42604 16690 42668
rect 18321 42666 18387 42669
rect 22134 42666 22140 42668
rect 18321 42664 22140 42666
rect 18321 42608 18326 42664
rect 18382 42608 22140 42664
rect 18321 42606 22140 42608
rect 18321 42603 18387 42606
rect 22134 42604 22140 42606
rect 22204 42604 22210 42668
rect 4429 42530 4495 42533
rect 4838 42530 4844 42532
rect 4429 42528 4844 42530
rect 4429 42472 4434 42528
rect 4490 42472 4844 42528
rect 4429 42470 4844 42472
rect 4429 42467 4495 42470
rect 4838 42468 4844 42470
rect 4908 42468 4914 42532
rect 7189 42530 7255 42533
rect 10133 42530 10199 42533
rect 7189 42528 10199 42530
rect 7189 42472 7194 42528
rect 7250 42472 10138 42528
rect 10194 42472 10199 42528
rect 7189 42470 10199 42472
rect 7189 42467 7255 42470
rect 10133 42467 10199 42470
rect 24853 42530 24919 42533
rect 25540 42530 26000 42560
rect 24853 42528 26000 42530
rect 24853 42472 24858 42528
rect 24914 42472 26000 42528
rect 24853 42470 26000 42472
rect 24853 42467 24919 42470
rect 6810 42464 7126 42465
rect 6810 42400 6816 42464
rect 6880 42400 6896 42464
rect 6960 42400 6976 42464
rect 7040 42400 7056 42464
rect 7120 42400 7126 42464
rect 6810 42399 7126 42400
rect 12675 42464 12991 42465
rect 12675 42400 12681 42464
rect 12745 42400 12761 42464
rect 12825 42400 12841 42464
rect 12905 42400 12921 42464
rect 12985 42400 12991 42464
rect 12675 42399 12991 42400
rect 18540 42464 18856 42465
rect 18540 42400 18546 42464
rect 18610 42400 18626 42464
rect 18690 42400 18706 42464
rect 18770 42400 18786 42464
rect 18850 42400 18856 42464
rect 18540 42399 18856 42400
rect 24405 42464 24721 42465
rect 24405 42400 24411 42464
rect 24475 42400 24491 42464
rect 24555 42400 24571 42464
rect 24635 42400 24651 42464
rect 24715 42400 24721 42464
rect 25540 42440 26000 42470
rect 24405 42399 24721 42400
rect 3325 42394 3391 42397
rect 3877 42394 3943 42397
rect 3325 42392 3943 42394
rect 3325 42336 3330 42392
rect 3386 42336 3882 42392
rect 3938 42336 3943 42392
rect 3325 42334 3943 42336
rect 3325 42331 3391 42334
rect 3877 42331 3943 42334
rect 4153 42394 4219 42397
rect 5625 42394 5691 42397
rect 4153 42392 5691 42394
rect 4153 42336 4158 42392
rect 4214 42336 5630 42392
rect 5686 42336 5691 42392
rect 4153 42334 5691 42336
rect 4153 42331 4219 42334
rect 5625 42331 5691 42334
rect 2037 42258 2103 42261
rect 14089 42258 14155 42261
rect 2037 42256 14155 42258
rect 2037 42200 2042 42256
rect 2098 42200 14094 42256
rect 14150 42200 14155 42256
rect 2037 42198 14155 42200
rect 2037 42195 2103 42198
rect 14089 42195 14155 42198
rect 19425 42258 19491 42261
rect 21081 42258 21147 42261
rect 19425 42256 21147 42258
rect 19425 42200 19430 42256
rect 19486 42200 21086 42256
rect 21142 42200 21147 42256
rect 19425 42198 21147 42200
rect 19425 42195 19491 42198
rect 21081 42195 21147 42198
rect 4337 42122 4403 42125
rect 5574 42122 5580 42124
rect 4337 42120 5580 42122
rect 4337 42064 4342 42120
rect 4398 42064 5580 42120
rect 4337 42062 5580 42064
rect 4337 42059 4403 42062
rect 5574 42060 5580 42062
rect 5644 42122 5650 42124
rect 8109 42122 8175 42125
rect 10358 42122 10364 42124
rect 5644 42120 8175 42122
rect 5644 42064 8114 42120
rect 8170 42064 8175 42120
rect 5644 42062 8175 42064
rect 5644 42060 5650 42062
rect 8109 42059 8175 42062
rect 8526 42062 10364 42122
rect 4797 41986 4863 41989
rect 8526 41986 8586 42062
rect 10358 42060 10364 42062
rect 10428 42060 10434 42124
rect 16982 42060 16988 42124
rect 17052 42122 17058 42124
rect 17493 42122 17559 42125
rect 17052 42120 17559 42122
rect 17052 42064 17498 42120
rect 17554 42064 17559 42120
rect 17052 42062 17559 42064
rect 17052 42060 17058 42062
rect 17493 42059 17559 42062
rect 4797 41984 8586 41986
rect 4797 41928 4802 41984
rect 4858 41928 8586 41984
rect 4797 41926 8586 41928
rect 4797 41923 4863 41926
rect 8886 41924 8892 41988
rect 8956 41986 8962 41988
rect 9305 41986 9371 41989
rect 8956 41984 9371 41986
rect 8956 41928 9310 41984
rect 9366 41928 9371 41984
rect 8956 41926 9371 41928
rect 8956 41924 8962 41926
rect 9305 41923 9371 41926
rect 17166 41924 17172 41988
rect 17236 41986 17242 41988
rect 17953 41986 18019 41989
rect 18321 41988 18387 41989
rect 18270 41986 18276 41988
rect 17236 41984 18019 41986
rect 17236 41928 17958 41984
rect 18014 41928 18019 41984
rect 17236 41926 18019 41928
rect 18230 41926 18276 41986
rect 18340 41984 18387 41988
rect 18382 41928 18387 41984
rect 17236 41924 17242 41926
rect 17953 41923 18019 41926
rect 18270 41924 18276 41926
rect 18340 41924 18387 41928
rect 18321 41923 18387 41924
rect 19517 41988 19583 41989
rect 19517 41984 19564 41988
rect 19628 41986 19634 41988
rect 19793 41986 19859 41989
rect 19926 41986 19932 41988
rect 19517 41928 19522 41984
rect 19517 41924 19564 41928
rect 19628 41926 19674 41986
rect 19793 41984 19932 41986
rect 19793 41928 19798 41984
rect 19854 41928 19932 41984
rect 19793 41926 19932 41928
rect 19628 41924 19634 41926
rect 19517 41923 19583 41924
rect 19793 41923 19859 41926
rect 19926 41924 19932 41926
rect 19996 41924 20002 41988
rect 24117 41986 24183 41989
rect 25540 41986 26000 42016
rect 24117 41984 26000 41986
rect 24117 41928 24122 41984
rect 24178 41928 26000 41984
rect 24117 41926 26000 41928
rect 24117 41923 24183 41926
rect 3878 41920 4194 41921
rect 3878 41856 3884 41920
rect 3948 41856 3964 41920
rect 4028 41856 4044 41920
rect 4108 41856 4124 41920
rect 4188 41856 4194 41920
rect 3878 41855 4194 41856
rect 9743 41920 10059 41921
rect 9743 41856 9749 41920
rect 9813 41856 9829 41920
rect 9893 41856 9909 41920
rect 9973 41856 9989 41920
rect 10053 41856 10059 41920
rect 9743 41855 10059 41856
rect 15608 41920 15924 41921
rect 15608 41856 15614 41920
rect 15678 41856 15694 41920
rect 15758 41856 15774 41920
rect 15838 41856 15854 41920
rect 15918 41856 15924 41920
rect 15608 41855 15924 41856
rect 21473 41920 21789 41921
rect 21473 41856 21479 41920
rect 21543 41856 21559 41920
rect 21623 41856 21639 41920
rect 21703 41856 21719 41920
rect 21783 41856 21789 41920
rect 25540 41896 26000 41926
rect 21473 41855 21789 41856
rect 9029 41852 9095 41853
rect 9029 41848 9076 41852
rect 9140 41850 9146 41852
rect 9029 41792 9034 41848
rect 9029 41788 9076 41792
rect 9140 41790 9186 41850
rect 9140 41788 9146 41790
rect 9029 41787 9095 41788
rect 4429 41714 4495 41717
rect 7557 41714 7623 41717
rect 4429 41712 7623 41714
rect 4429 41656 4434 41712
rect 4490 41656 7562 41712
rect 7618 41656 7623 41712
rect 4429 41654 7623 41656
rect 4429 41651 4495 41654
rect 7557 41651 7623 41654
rect 20621 41714 20687 41717
rect 21265 41714 21331 41717
rect 20621 41712 21331 41714
rect 20621 41656 20626 41712
rect 20682 41656 21270 41712
rect 21326 41656 21331 41712
rect 20621 41654 21331 41656
rect 20621 41651 20687 41654
rect 21265 41651 21331 41654
rect 2497 41578 2563 41581
rect 3734 41578 3740 41580
rect 2497 41576 3740 41578
rect 2497 41520 2502 41576
rect 2558 41520 3740 41576
rect 2497 41518 3740 41520
rect 2497 41515 2563 41518
rect 3734 41516 3740 41518
rect 3804 41578 3810 41580
rect 5717 41578 5783 41581
rect 9121 41578 9187 41581
rect 9254 41578 9260 41580
rect 3804 41576 5783 41578
rect 3804 41520 5722 41576
rect 5778 41520 5783 41576
rect 3804 41518 5783 41520
rect 3804 41516 3810 41518
rect 5717 41515 5783 41518
rect 5950 41518 7298 41578
rect 1393 41442 1459 41445
rect 1526 41442 1532 41444
rect 1393 41440 1532 41442
rect 1393 41384 1398 41440
rect 1454 41384 1532 41440
rect 1393 41382 1532 41384
rect 1393 41379 1459 41382
rect 1526 41380 1532 41382
rect 1596 41380 1602 41444
rect 2037 41442 2103 41445
rect 2446 41442 2452 41444
rect 2037 41440 2452 41442
rect 2037 41384 2042 41440
rect 2098 41384 2452 41440
rect 2037 41382 2452 41384
rect 2037 41379 2103 41382
rect 2446 41380 2452 41382
rect 2516 41380 2522 41444
rect 2313 41034 2379 41037
rect 5950 41034 6010 41518
rect 6126 41380 6132 41444
rect 6196 41442 6202 41444
rect 6637 41442 6703 41445
rect 6196 41440 6703 41442
rect 6196 41384 6642 41440
rect 6698 41384 6703 41440
rect 6196 41382 6703 41384
rect 6196 41380 6202 41382
rect 6637 41379 6703 41382
rect 6810 41376 7126 41377
rect 6810 41312 6816 41376
rect 6880 41312 6896 41376
rect 6960 41312 6976 41376
rect 7040 41312 7056 41376
rect 7120 41312 7126 41376
rect 6810 41311 7126 41312
rect 7238 41170 7298 41518
rect 9121 41576 9260 41578
rect 9121 41520 9126 41576
rect 9182 41520 9260 41576
rect 9121 41518 9260 41520
rect 9121 41515 9187 41518
rect 9254 41516 9260 41518
rect 9324 41516 9330 41580
rect 9438 41516 9444 41580
rect 9508 41578 9514 41580
rect 10409 41578 10475 41581
rect 9508 41576 10475 41578
rect 9508 41520 10414 41576
rect 10470 41520 10475 41576
rect 9508 41518 10475 41520
rect 9508 41516 9514 41518
rect 10409 41515 10475 41518
rect 20529 41578 20595 41581
rect 21214 41578 21220 41580
rect 20529 41576 21220 41578
rect 20529 41520 20534 41576
rect 20590 41520 21220 41576
rect 20529 41518 21220 41520
rect 20529 41515 20595 41518
rect 21214 41516 21220 41518
rect 21284 41516 21290 41580
rect 23381 41578 23447 41581
rect 23381 41576 24962 41578
rect 23381 41520 23386 41576
rect 23442 41520 24962 41576
rect 23381 41518 24962 41520
rect 23381 41515 23447 41518
rect 10910 41380 10916 41444
rect 10980 41442 10986 41444
rect 12433 41442 12499 41445
rect 10980 41440 12499 41442
rect 10980 41384 12438 41440
rect 12494 41384 12499 41440
rect 10980 41382 12499 41384
rect 10980 41380 10986 41382
rect 12433 41379 12499 41382
rect 19609 41442 19675 41445
rect 21449 41442 21515 41445
rect 19609 41440 21515 41442
rect 19609 41384 19614 41440
rect 19670 41384 21454 41440
rect 21510 41384 21515 41440
rect 24902 41442 24962 41518
rect 25540 41442 26000 41472
rect 23841 41430 23907 41433
rect 19609 41382 21515 41384
rect 19609 41379 19675 41382
rect 21449 41379 21515 41382
rect 23798 41428 23907 41430
rect 12675 41376 12991 41377
rect 12675 41312 12681 41376
rect 12745 41312 12761 41376
rect 12825 41312 12841 41376
rect 12905 41312 12921 41376
rect 12985 41312 12991 41376
rect 12675 41311 12991 41312
rect 18540 41376 18856 41377
rect 18540 41312 18546 41376
rect 18610 41312 18626 41376
rect 18690 41312 18706 41376
rect 18770 41312 18786 41376
rect 18850 41312 18856 41376
rect 18540 41311 18856 41312
rect 23798 41372 23846 41428
rect 23902 41372 23907 41428
rect 24902 41382 26000 41442
rect 23798 41367 23907 41372
rect 24405 41376 24721 41377
rect 13813 41170 13879 41173
rect 7238 41168 13879 41170
rect 7238 41112 13818 41168
rect 13874 41112 13879 41168
rect 7238 41110 13879 41112
rect 13813 41107 13879 41110
rect 13997 41034 14063 41037
rect 23798 41034 23858 41367
rect 24405 41312 24411 41376
rect 24475 41312 24491 41376
rect 24555 41312 24571 41376
rect 24635 41312 24651 41376
rect 24715 41312 24721 41376
rect 25540 41352 26000 41382
rect 24405 41311 24721 41312
rect 2313 41032 6010 41034
rect 2313 40976 2318 41032
rect 2374 40976 6010 41032
rect 2313 40974 6010 40976
rect 8526 41032 14063 41034
rect 8526 40976 14002 41032
rect 14058 40976 14063 41032
rect 8526 40974 14063 40976
rect 2313 40971 2379 40974
rect 4429 40898 4495 40901
rect 7465 40898 7531 40901
rect 4429 40896 7531 40898
rect 4429 40840 4434 40896
rect 4490 40840 7470 40896
rect 7526 40840 7531 40896
rect 4429 40838 7531 40840
rect 4429 40835 4495 40838
rect 7465 40835 7531 40838
rect 3878 40832 4194 40833
rect 3878 40768 3884 40832
rect 3948 40768 3964 40832
rect 4028 40768 4044 40832
rect 4108 40768 4124 40832
rect 4188 40768 4194 40832
rect 3878 40767 4194 40768
rect 4797 40762 4863 40765
rect 8526 40762 8586 40974
rect 13997 40971 14063 40974
rect 22050 40974 23858 41034
rect 21909 40898 21975 40901
rect 22050 40898 22110 40974
rect 21909 40896 22110 40898
rect 21909 40840 21914 40896
rect 21970 40840 22110 40896
rect 21909 40838 22110 40840
rect 23657 40898 23723 40901
rect 25540 40898 26000 40928
rect 23657 40896 26000 40898
rect 23657 40840 23662 40896
rect 23718 40840 26000 40896
rect 23657 40838 26000 40840
rect 21909 40835 21975 40838
rect 23657 40835 23723 40838
rect 9743 40832 10059 40833
rect 9743 40768 9749 40832
rect 9813 40768 9829 40832
rect 9893 40768 9909 40832
rect 9973 40768 9989 40832
rect 10053 40768 10059 40832
rect 9743 40767 10059 40768
rect 15608 40832 15924 40833
rect 15608 40768 15614 40832
rect 15678 40768 15694 40832
rect 15758 40768 15774 40832
rect 15838 40768 15854 40832
rect 15918 40768 15924 40832
rect 15608 40767 15924 40768
rect 21473 40832 21789 40833
rect 21473 40768 21479 40832
rect 21543 40768 21559 40832
rect 21623 40768 21639 40832
rect 21703 40768 21719 40832
rect 21783 40768 21789 40832
rect 25540 40808 26000 40838
rect 21473 40767 21789 40768
rect 4797 40760 8586 40762
rect 4797 40704 4802 40760
rect 4858 40704 8586 40760
rect 4797 40702 8586 40704
rect 4797 40699 4863 40702
rect 197 40626 263 40629
rect 6177 40626 6243 40629
rect 197 40624 6243 40626
rect 197 40568 202 40624
rect 258 40568 6182 40624
rect 6238 40568 6243 40624
rect 197 40566 6243 40568
rect 197 40563 263 40566
rect 6177 40563 6243 40566
rect 1669 40490 1735 40493
rect 5441 40490 5507 40493
rect 8661 40490 8727 40493
rect 1669 40488 8727 40490
rect 1669 40432 1674 40488
rect 1730 40432 5446 40488
rect 5502 40432 8666 40488
rect 8722 40432 8727 40488
rect 1669 40430 8727 40432
rect 1669 40427 1735 40430
rect 5441 40427 5507 40430
rect 8661 40427 8727 40430
rect 20345 40490 20411 40493
rect 25037 40490 25103 40493
rect 20345 40488 25103 40490
rect 20345 40432 20350 40488
rect 20406 40432 25042 40488
rect 25098 40432 25103 40488
rect 20345 40430 25103 40432
rect 20345 40427 20411 40430
rect 25037 40427 25103 40430
rect 2630 40292 2636 40356
rect 2700 40354 2706 40356
rect 3233 40354 3299 40357
rect 2700 40352 3299 40354
rect 2700 40296 3238 40352
rect 3294 40296 3299 40352
rect 2700 40294 3299 40296
rect 2700 40292 2706 40294
rect 3233 40291 3299 40294
rect 24945 40354 25011 40357
rect 25540 40354 26000 40384
rect 24945 40352 26000 40354
rect 24945 40296 24950 40352
rect 25006 40296 26000 40352
rect 24945 40294 26000 40296
rect 24945 40291 25011 40294
rect 6810 40288 7126 40289
rect 6810 40224 6816 40288
rect 6880 40224 6896 40288
rect 6960 40224 6976 40288
rect 7040 40224 7056 40288
rect 7120 40224 7126 40288
rect 6810 40223 7126 40224
rect 12675 40288 12991 40289
rect 12675 40224 12681 40288
rect 12745 40224 12761 40288
rect 12825 40224 12841 40288
rect 12905 40224 12921 40288
rect 12985 40224 12991 40288
rect 12675 40223 12991 40224
rect 18540 40288 18856 40289
rect 18540 40224 18546 40288
rect 18610 40224 18626 40288
rect 18690 40224 18706 40288
rect 18770 40224 18786 40288
rect 18850 40224 18856 40288
rect 18540 40223 18856 40224
rect 24405 40288 24721 40289
rect 24405 40224 24411 40288
rect 24475 40224 24491 40288
rect 24555 40224 24571 40288
rect 24635 40224 24651 40288
rect 24715 40224 24721 40288
rect 25540 40264 26000 40294
rect 24405 40223 24721 40224
rect 565 40218 631 40221
rect 5809 40218 5875 40221
rect 565 40216 5875 40218
rect 565 40160 570 40216
rect 626 40160 5814 40216
rect 5870 40160 5875 40216
rect 565 40158 5875 40160
rect 565 40155 631 40158
rect 5809 40155 5875 40158
rect 606 40020 612 40084
rect 676 40082 682 40084
rect 3601 40082 3667 40085
rect 676 40080 3667 40082
rect 676 40024 3606 40080
rect 3662 40024 3667 40080
rect 676 40022 3667 40024
rect 676 40020 682 40022
rect 3601 40019 3667 40022
rect 4838 40020 4844 40084
rect 4908 40082 4914 40084
rect 5349 40082 5415 40085
rect 22369 40082 22435 40085
rect 4908 40080 22435 40082
rect 4908 40024 5354 40080
rect 5410 40024 22374 40080
rect 22430 40024 22435 40080
rect 4908 40022 22435 40024
rect 4908 40020 4914 40022
rect 5349 40019 5415 40022
rect 22369 40019 22435 40022
rect 1945 39946 2011 39949
rect 5625 39946 5691 39949
rect 13302 39946 13308 39948
rect 1945 39944 13308 39946
rect 1945 39888 1950 39944
rect 2006 39888 5630 39944
rect 5686 39888 13308 39944
rect 1945 39886 13308 39888
rect 1945 39883 2011 39886
rect 5625 39883 5691 39886
rect 13302 39884 13308 39886
rect 13372 39884 13378 39948
rect 21817 39946 21883 39949
rect 22277 39946 22343 39949
rect 21817 39944 22343 39946
rect 21817 39888 21822 39944
rect 21878 39888 22282 39944
rect 22338 39888 22343 39944
rect 21817 39886 22343 39888
rect 21817 39883 21883 39886
rect 22277 39883 22343 39886
rect 21950 39748 21956 39812
rect 22020 39810 22026 39812
rect 23381 39810 23447 39813
rect 22020 39808 23447 39810
rect 22020 39752 23386 39808
rect 23442 39752 23447 39808
rect 22020 39750 23447 39752
rect 22020 39748 22026 39750
rect 23381 39747 23447 39750
rect 24117 39810 24183 39813
rect 25540 39810 26000 39840
rect 24117 39808 26000 39810
rect 24117 39752 24122 39808
rect 24178 39752 26000 39808
rect 24117 39750 26000 39752
rect 24117 39747 24183 39750
rect 3878 39744 4194 39745
rect 3878 39680 3884 39744
rect 3948 39680 3964 39744
rect 4028 39680 4044 39744
rect 4108 39680 4124 39744
rect 4188 39680 4194 39744
rect 3878 39679 4194 39680
rect 9743 39744 10059 39745
rect 9743 39680 9749 39744
rect 9813 39680 9829 39744
rect 9893 39680 9909 39744
rect 9973 39680 9989 39744
rect 10053 39680 10059 39744
rect 9743 39679 10059 39680
rect 15608 39744 15924 39745
rect 15608 39680 15614 39744
rect 15678 39680 15694 39744
rect 15758 39680 15774 39744
rect 15838 39680 15854 39744
rect 15918 39680 15924 39744
rect 15608 39679 15924 39680
rect 21473 39744 21789 39745
rect 21473 39680 21479 39744
rect 21543 39680 21559 39744
rect 21623 39680 21639 39744
rect 21703 39680 21719 39744
rect 21783 39680 21789 39744
rect 25540 39720 26000 39750
rect 21473 39679 21789 39680
rect 1158 39612 1164 39676
rect 1228 39674 1234 39676
rect 1228 39614 3204 39674
rect 1228 39612 1234 39614
rect -300 39538 160 39568
rect 2957 39538 3023 39541
rect -300 39536 3023 39538
rect -300 39480 2962 39536
rect 3018 39480 3023 39536
rect -300 39478 3023 39480
rect 3144 39538 3204 39614
rect 9213 39538 9279 39541
rect 3144 39536 9279 39538
rect 3144 39480 9218 39536
rect 9274 39480 9279 39536
rect 3144 39478 9279 39480
rect -300 39448 160 39478
rect 2957 39475 3023 39478
rect 9213 39475 9279 39478
rect 10961 39538 11027 39541
rect 19374 39538 19380 39540
rect 10961 39536 19380 39538
rect 10961 39480 10966 39536
rect 11022 39480 19380 39536
rect 10961 39478 19380 39480
rect 10961 39475 11027 39478
rect 19374 39476 19380 39478
rect 19444 39476 19450 39540
rect 20253 39538 20319 39541
rect 24945 39538 25011 39541
rect 20253 39536 25011 39538
rect 20253 39480 20258 39536
rect 20314 39480 24950 39536
rect 25006 39480 25011 39536
rect 20253 39478 25011 39480
rect 20253 39475 20319 39478
rect 24945 39475 25011 39478
rect 1393 39400 1459 39405
rect 1393 39344 1398 39400
rect 1454 39344 1459 39400
rect 1393 39339 1459 39344
rect 4521 39402 4587 39405
rect 8753 39402 8819 39405
rect 10685 39402 10751 39405
rect 21030 39402 21036 39404
rect 4521 39400 10472 39402
rect 4521 39344 4526 39400
rect 4582 39344 8758 39400
rect 8814 39344 10472 39400
rect 4521 39342 10472 39344
rect 4521 39339 4587 39342
rect 8753 39339 8819 39342
rect -300 39266 160 39296
rect 1396 39266 1456 39339
rect -300 39206 1456 39266
rect 3601 39266 3667 39269
rect 3734 39266 3740 39268
rect 3601 39264 3740 39266
rect 3601 39208 3606 39264
rect 3662 39208 3740 39264
rect 3601 39206 3740 39208
rect -300 39176 160 39206
rect 3601 39203 3667 39206
rect 3734 39204 3740 39206
rect 3804 39266 3810 39268
rect 5206 39266 5212 39268
rect 3804 39206 5212 39266
rect 3804 39204 3810 39206
rect 5206 39204 5212 39206
rect 5276 39204 5282 39268
rect 10412 39266 10472 39342
rect 10685 39400 21036 39402
rect 10685 39344 10690 39400
rect 10746 39344 21036 39400
rect 10685 39342 21036 39344
rect 10685 39339 10751 39342
rect 21030 39340 21036 39342
rect 21100 39340 21106 39404
rect 10685 39266 10751 39269
rect 10412 39264 10751 39266
rect 10412 39208 10690 39264
rect 10746 39208 10751 39264
rect 10412 39206 10751 39208
rect 10685 39203 10751 39206
rect 24853 39266 24919 39269
rect 25540 39266 26000 39296
rect 24853 39264 26000 39266
rect 24853 39208 24858 39264
rect 24914 39208 26000 39264
rect 24853 39206 26000 39208
rect 24853 39203 24919 39206
rect 6810 39200 7126 39201
rect 6810 39136 6816 39200
rect 6880 39136 6896 39200
rect 6960 39136 6976 39200
rect 7040 39136 7056 39200
rect 7120 39136 7126 39200
rect 6810 39135 7126 39136
rect 12675 39200 12991 39201
rect 12675 39136 12681 39200
rect 12745 39136 12761 39200
rect 12825 39136 12841 39200
rect 12905 39136 12921 39200
rect 12985 39136 12991 39200
rect 12675 39135 12991 39136
rect 18540 39200 18856 39201
rect 18540 39136 18546 39200
rect 18610 39136 18626 39200
rect 18690 39136 18706 39200
rect 18770 39136 18786 39200
rect 18850 39136 18856 39200
rect 18540 39135 18856 39136
rect 24405 39200 24721 39201
rect 24405 39136 24411 39200
rect 24475 39136 24491 39200
rect 24555 39136 24571 39200
rect 24635 39136 24651 39200
rect 24715 39136 24721 39200
rect 25540 39176 26000 39206
rect 24405 39135 24721 39136
rect 2773 39130 2839 39133
rect 2730 39128 2839 39130
rect 2730 39072 2778 39128
rect 2834 39072 2839 39128
rect 2730 39067 2839 39072
rect 3877 39130 3943 39133
rect 6310 39130 6316 39132
rect 3877 39128 6316 39130
rect 3877 39072 3882 39128
rect 3938 39072 6316 39128
rect 3877 39070 6316 39072
rect 3877 39067 3943 39070
rect 6310 39068 6316 39070
rect 6380 39130 6386 39132
rect 10041 39130 10107 39133
rect 11513 39130 11579 39133
rect 6380 39070 6746 39130
rect 6380 39068 6386 39070
rect -300 38994 160 39024
rect 2730 38994 2790 39067
rect -300 38934 2790 38994
rect -300 38904 160 38934
rect 3734 38932 3740 38996
rect 3804 38994 3810 38996
rect 3969 38994 4035 38997
rect 3804 38992 4035 38994
rect 3804 38936 3974 38992
rect 4030 38936 4035 38992
rect 3804 38934 4035 38936
rect 6686 38994 6746 39070
rect 10041 39128 11579 39130
rect 10041 39072 10046 39128
rect 10102 39072 11518 39128
rect 11574 39072 11579 39128
rect 10041 39070 11579 39072
rect 10041 39067 10107 39070
rect 11513 39067 11579 39070
rect 15193 38994 15259 38997
rect 6686 38992 15259 38994
rect 6686 38936 15198 38992
rect 15254 38936 15259 38992
rect 6686 38934 15259 38936
rect 3804 38932 3810 38934
rect 3969 38931 4035 38934
rect 15193 38931 15259 38934
rect 790 38796 796 38860
rect 860 38858 866 38860
rect 9857 38858 9923 38861
rect 860 38856 9923 38858
rect 860 38800 9862 38856
rect 9918 38800 9923 38856
rect 860 38798 9923 38800
rect 860 38796 866 38798
rect 9857 38795 9923 38798
rect -300 38722 160 38752
rect 3693 38722 3759 38725
rect -300 38720 3759 38722
rect -300 38664 3698 38720
rect 3754 38664 3759 38720
rect -300 38662 3759 38664
rect -300 38632 160 38662
rect 3693 38659 3759 38662
rect 11462 38660 11468 38724
rect 11532 38722 11538 38724
rect 11697 38722 11763 38725
rect 11532 38720 11763 38722
rect 11532 38664 11702 38720
rect 11758 38664 11763 38720
rect 11532 38662 11763 38664
rect 11532 38660 11538 38662
rect 11697 38659 11763 38662
rect 24117 38722 24183 38725
rect 25540 38722 26000 38752
rect 24117 38720 26000 38722
rect 24117 38664 24122 38720
rect 24178 38664 26000 38720
rect 24117 38662 26000 38664
rect 24117 38659 24183 38662
rect 3878 38656 4194 38657
rect 3878 38592 3884 38656
rect 3948 38592 3964 38656
rect 4028 38592 4044 38656
rect 4108 38592 4124 38656
rect 4188 38592 4194 38656
rect 3878 38591 4194 38592
rect 9743 38656 10059 38657
rect 9743 38592 9749 38656
rect 9813 38592 9829 38656
rect 9893 38592 9909 38656
rect 9973 38592 9989 38656
rect 10053 38592 10059 38656
rect 9743 38591 10059 38592
rect 15608 38656 15924 38657
rect 15608 38592 15614 38656
rect 15678 38592 15694 38656
rect 15758 38592 15774 38656
rect 15838 38592 15854 38656
rect 15918 38592 15924 38656
rect 15608 38591 15924 38592
rect 21473 38656 21789 38657
rect 21473 38592 21479 38656
rect 21543 38592 21559 38656
rect 21623 38592 21639 38656
rect 21703 38592 21719 38656
rect 21783 38592 21789 38656
rect 25540 38632 26000 38662
rect 21473 38591 21789 38592
rect 1577 38586 1643 38589
rect 3693 38586 3759 38589
rect 6269 38586 6335 38589
rect 1577 38584 3759 38586
rect 1577 38528 1582 38584
rect 1638 38528 3698 38584
rect 3754 38528 3759 38584
rect 1577 38526 3759 38528
rect 1577 38523 1643 38526
rect 3693 38523 3759 38526
rect 4294 38584 6335 38586
rect 4294 38528 6274 38584
rect 6330 38528 6335 38584
rect 4294 38526 6335 38528
rect -300 38450 160 38480
rect 2773 38450 2839 38453
rect -300 38448 2839 38450
rect -300 38392 2778 38448
rect 2834 38392 2839 38448
rect -300 38390 2839 38392
rect -300 38360 160 38390
rect 2773 38387 2839 38390
rect 3550 38388 3556 38452
rect 3620 38450 3626 38452
rect 4294 38450 4354 38526
rect 6269 38523 6335 38526
rect 3620 38390 4354 38450
rect 3620 38388 3626 38390
rect 2446 38252 2452 38316
rect 2516 38314 2522 38316
rect 3141 38314 3207 38317
rect 13629 38314 13695 38317
rect 2516 38312 13695 38314
rect 2516 38256 3146 38312
rect 3202 38256 13634 38312
rect 13690 38256 13695 38312
rect 2516 38254 13695 38256
rect 2516 38252 2522 38254
rect 3141 38251 3207 38254
rect -300 38178 160 38208
rect 749 38178 815 38181
rect -300 38176 815 38178
rect -300 38120 754 38176
rect 810 38120 815 38176
rect -300 38118 815 38120
rect -300 38088 160 38118
rect 749 38115 815 38118
rect 3366 38116 3372 38180
rect 3436 38178 3442 38180
rect 3877 38178 3943 38181
rect 4294 38180 4354 38254
rect 13629 38251 13695 38254
rect 3436 38176 3943 38178
rect 3436 38120 3882 38176
rect 3938 38120 3943 38176
rect 3436 38118 3943 38120
rect 3436 38116 3442 38118
rect 3877 38115 3943 38118
rect 4286 38116 4292 38180
rect 4356 38116 4362 38180
rect 24853 38178 24919 38181
rect 25540 38178 26000 38208
rect 24853 38176 26000 38178
rect 24853 38120 24858 38176
rect 24914 38120 26000 38176
rect 24853 38118 26000 38120
rect 24853 38115 24919 38118
rect 6810 38112 7126 38113
rect 6810 38048 6816 38112
rect 6880 38048 6896 38112
rect 6960 38048 6976 38112
rect 7040 38048 7056 38112
rect 7120 38048 7126 38112
rect 6810 38047 7126 38048
rect 12675 38112 12991 38113
rect 12675 38048 12681 38112
rect 12745 38048 12761 38112
rect 12825 38048 12841 38112
rect 12905 38048 12921 38112
rect 12985 38048 12991 38112
rect 12675 38047 12991 38048
rect 18540 38112 18856 38113
rect 18540 38048 18546 38112
rect 18610 38048 18626 38112
rect 18690 38048 18706 38112
rect 18770 38048 18786 38112
rect 18850 38048 18856 38112
rect 18540 38047 18856 38048
rect 24405 38112 24721 38113
rect 24405 38048 24411 38112
rect 24475 38048 24491 38112
rect 24555 38048 24571 38112
rect 24635 38048 24651 38112
rect 24715 38048 24721 38112
rect 25540 38088 26000 38118
rect 24405 38047 24721 38048
rect 2405 38042 2471 38045
rect 2405 38040 6746 38042
rect 2405 37984 2410 38040
rect 2466 37984 6746 38040
rect 2405 37982 6746 37984
rect 2405 37979 2471 37982
rect -300 37906 160 37936
rect 4981 37906 5047 37909
rect -300 37904 5047 37906
rect -300 37848 4986 37904
rect 5042 37848 5047 37904
rect -300 37846 5047 37848
rect -300 37816 160 37846
rect 4981 37843 5047 37846
rect 4337 37770 4403 37773
rect 2730 37768 4403 37770
rect 2730 37712 4342 37768
rect 4398 37712 4403 37768
rect 2730 37710 4403 37712
rect 6686 37770 6746 37982
rect 11421 37770 11487 37773
rect 6686 37768 11487 37770
rect 6686 37712 11426 37768
rect 11482 37712 11487 37768
rect 6686 37710 11487 37712
rect -300 37634 160 37664
rect 2730 37634 2790 37710
rect 4337 37707 4403 37710
rect 11421 37707 11487 37710
rect -300 37574 2790 37634
rect 24117 37634 24183 37637
rect 25540 37634 26000 37664
rect 24117 37632 26000 37634
rect 24117 37576 24122 37632
rect 24178 37576 26000 37632
rect 24117 37574 26000 37576
rect -300 37544 160 37574
rect 24117 37571 24183 37574
rect 3878 37568 4194 37569
rect 3878 37504 3884 37568
rect 3948 37504 3964 37568
rect 4028 37504 4044 37568
rect 4108 37504 4124 37568
rect 4188 37504 4194 37568
rect 3878 37503 4194 37504
rect 9743 37568 10059 37569
rect 9743 37504 9749 37568
rect 9813 37504 9829 37568
rect 9893 37504 9909 37568
rect 9973 37504 9989 37568
rect 10053 37504 10059 37568
rect 9743 37503 10059 37504
rect 15608 37568 15924 37569
rect 15608 37504 15614 37568
rect 15678 37504 15694 37568
rect 15758 37504 15774 37568
rect 15838 37504 15854 37568
rect 15918 37504 15924 37568
rect 15608 37503 15924 37504
rect 21473 37568 21789 37569
rect 21473 37504 21479 37568
rect 21543 37504 21559 37568
rect 21623 37504 21639 37568
rect 21703 37504 21719 37568
rect 21783 37504 21789 37568
rect 25540 37544 26000 37574
rect 21473 37503 21789 37504
rect 1209 37498 1275 37501
rect 5257 37498 5323 37501
rect 5390 37498 5396 37500
rect 1209 37496 1778 37498
rect 1209 37440 1214 37496
rect 1270 37440 1778 37496
rect 1209 37438 1778 37440
rect 1209 37435 1275 37438
rect -300 37362 160 37392
rect 1577 37362 1643 37365
rect -300 37360 1643 37362
rect -300 37304 1582 37360
rect 1638 37304 1643 37360
rect -300 37302 1643 37304
rect 1718 37362 1778 37438
rect 5257 37496 5396 37498
rect 5257 37440 5262 37496
rect 5318 37440 5396 37496
rect 5257 37438 5396 37440
rect 5257 37435 5323 37438
rect 5390 37436 5396 37438
rect 5460 37436 5466 37500
rect 4245 37362 4311 37365
rect 1718 37360 4311 37362
rect 1718 37304 4250 37360
rect 4306 37304 4311 37360
rect 1718 37302 4311 37304
rect -300 37272 160 37302
rect 1577 37299 1643 37302
rect 4245 37299 4311 37302
rect 4889 37362 4955 37365
rect 6269 37362 6335 37365
rect 4889 37360 6335 37362
rect 4889 37304 4894 37360
rect 4950 37304 6274 37360
rect 6330 37304 6335 37360
rect 4889 37302 6335 37304
rect 4889 37299 4955 37302
rect 6269 37299 6335 37302
rect 12157 37362 12223 37365
rect 13670 37362 13676 37364
rect 12157 37360 13676 37362
rect 12157 37304 12162 37360
rect 12218 37304 13676 37360
rect 12157 37302 13676 37304
rect 12157 37299 12223 37302
rect 13670 37300 13676 37302
rect 13740 37300 13746 37364
rect 1393 37226 1459 37229
rect 2957 37226 3023 37229
rect 1393 37224 3023 37226
rect 1393 37168 1398 37224
rect 1454 37168 2962 37224
rect 3018 37168 3023 37224
rect 1393 37166 3023 37168
rect 1393 37163 1459 37166
rect 2957 37163 3023 37166
rect 3877 37226 3943 37229
rect 6177 37226 6243 37229
rect 3877 37224 6243 37226
rect 3877 37168 3882 37224
rect 3938 37168 6182 37224
rect 6238 37168 6243 37224
rect 3877 37166 6243 37168
rect 3877 37163 3943 37166
rect 6177 37163 6243 37166
rect -300 37090 160 37120
rect 3049 37090 3115 37093
rect -300 37088 3115 37090
rect -300 37032 3054 37088
rect 3110 37032 3115 37088
rect -300 37030 3115 37032
rect -300 37000 160 37030
rect 3049 37027 3115 37030
rect 4153 37090 4219 37093
rect 4654 37090 4660 37092
rect 4153 37088 4660 37090
rect 4153 37032 4158 37088
rect 4214 37032 4660 37088
rect 4153 37030 4660 37032
rect 4153 37027 4219 37030
rect 4654 37028 4660 37030
rect 4724 37090 4730 37092
rect 6637 37090 6703 37093
rect 4724 37088 6703 37090
rect 4724 37032 6642 37088
rect 6698 37032 6703 37088
rect 4724 37030 6703 37032
rect 4724 37028 4730 37030
rect 6637 37027 6703 37030
rect 24853 37090 24919 37093
rect 25540 37090 26000 37120
rect 24853 37088 26000 37090
rect 24853 37032 24858 37088
rect 24914 37032 26000 37088
rect 24853 37030 26000 37032
rect 24853 37027 24919 37030
rect 6810 37024 7126 37025
rect 6810 36960 6816 37024
rect 6880 36960 6896 37024
rect 6960 36960 6976 37024
rect 7040 36960 7056 37024
rect 7120 36960 7126 37024
rect 6810 36959 7126 36960
rect 12675 37024 12991 37025
rect 12675 36960 12681 37024
rect 12745 36960 12761 37024
rect 12825 36960 12841 37024
rect 12905 36960 12921 37024
rect 12985 36960 12991 37024
rect 12675 36959 12991 36960
rect 18540 37024 18856 37025
rect 18540 36960 18546 37024
rect 18610 36960 18626 37024
rect 18690 36960 18706 37024
rect 18770 36960 18786 37024
rect 18850 36960 18856 37024
rect 18540 36959 18856 36960
rect 24405 37024 24721 37025
rect 24405 36960 24411 37024
rect 24475 36960 24491 37024
rect 24555 36960 24571 37024
rect 24635 36960 24651 37024
rect 24715 36960 24721 37024
rect 25540 37000 26000 37030
rect 24405 36959 24721 36960
rect 1761 36954 1827 36957
rect 1534 36952 1827 36954
rect 1534 36896 1766 36952
rect 1822 36896 1827 36952
rect 1534 36894 1827 36896
rect -300 36818 160 36848
rect 1393 36818 1459 36821
rect -300 36816 1459 36818
rect -300 36760 1398 36816
rect 1454 36760 1459 36816
rect -300 36758 1459 36760
rect -300 36728 160 36758
rect 1393 36755 1459 36758
rect -300 36546 160 36576
rect 1534 36546 1594 36894
rect 1761 36891 1827 36894
rect 3049 36954 3115 36957
rect 5717 36954 5783 36957
rect 3049 36952 5783 36954
rect 3049 36896 3054 36952
rect 3110 36896 5722 36952
rect 5778 36896 5783 36952
rect 3049 36894 5783 36896
rect 3049 36891 3115 36894
rect 5717 36891 5783 36894
rect 3734 36756 3740 36820
rect 3804 36818 3810 36820
rect 10133 36818 10199 36821
rect 20345 36818 20411 36821
rect 3804 36816 10199 36818
rect 3804 36760 10138 36816
rect 10194 36760 10199 36816
rect 3804 36758 10199 36760
rect 3804 36756 3810 36758
rect 10133 36755 10199 36758
rect 12390 36816 20411 36818
rect 12390 36760 20350 36816
rect 20406 36760 20411 36816
rect 12390 36758 20411 36760
rect 1669 36682 1735 36685
rect 11237 36682 11303 36685
rect 12390 36682 12450 36758
rect 20345 36755 20411 36758
rect 1669 36680 12450 36682
rect 1669 36624 1674 36680
rect 1730 36624 11242 36680
rect 11298 36624 12450 36680
rect 1669 36622 12450 36624
rect 1669 36619 1735 36622
rect 11237 36619 11303 36622
rect -300 36486 1594 36546
rect -300 36456 160 36486
rect 4470 36484 4476 36548
rect 4540 36546 4546 36548
rect 4705 36546 4771 36549
rect 4981 36546 5047 36549
rect 9029 36546 9095 36549
rect 4540 36544 9095 36546
rect 4540 36488 4710 36544
rect 4766 36488 4986 36544
rect 5042 36488 9034 36544
rect 9090 36488 9095 36544
rect 4540 36486 9095 36488
rect 4540 36484 4546 36486
rect 4705 36483 4771 36486
rect 4981 36483 5047 36486
rect 9029 36483 9095 36486
rect 24117 36546 24183 36549
rect 25540 36546 26000 36576
rect 24117 36544 26000 36546
rect 24117 36488 24122 36544
rect 24178 36488 26000 36544
rect 24117 36486 26000 36488
rect 24117 36483 24183 36486
rect 3878 36480 4194 36481
rect 3878 36416 3884 36480
rect 3948 36416 3964 36480
rect 4028 36416 4044 36480
rect 4108 36416 4124 36480
rect 4188 36416 4194 36480
rect 3878 36415 4194 36416
rect 9743 36480 10059 36481
rect 9743 36416 9749 36480
rect 9813 36416 9829 36480
rect 9893 36416 9909 36480
rect 9973 36416 9989 36480
rect 10053 36416 10059 36480
rect 9743 36415 10059 36416
rect 15608 36480 15924 36481
rect 15608 36416 15614 36480
rect 15678 36416 15694 36480
rect 15758 36416 15774 36480
rect 15838 36416 15854 36480
rect 15918 36416 15924 36480
rect 15608 36415 15924 36416
rect 21473 36480 21789 36481
rect 21473 36416 21479 36480
rect 21543 36416 21559 36480
rect 21623 36416 21639 36480
rect 21703 36416 21719 36480
rect 21783 36416 21789 36480
rect 25540 36456 26000 36486
rect 21473 36415 21789 36416
rect 2313 36410 2379 36413
rect 8017 36410 8083 36413
rect 2313 36408 3802 36410
rect 2313 36352 2318 36408
rect 2374 36352 3802 36408
rect 2313 36350 3802 36352
rect 2313 36347 2379 36350
rect -300 36274 160 36304
rect 2865 36274 2931 36277
rect -300 36272 2931 36274
rect -300 36216 2870 36272
rect 2926 36216 2931 36272
rect -300 36214 2931 36216
rect -300 36184 160 36214
rect 2865 36211 2931 36214
rect 3141 36274 3207 36277
rect 3550 36274 3556 36276
rect 3141 36272 3556 36274
rect 3141 36216 3146 36272
rect 3202 36216 3556 36272
rect 3141 36214 3556 36216
rect 3141 36211 3207 36214
rect 3550 36212 3556 36214
rect 3620 36212 3626 36276
rect 3742 36274 3802 36350
rect 4294 36408 8083 36410
rect 4294 36352 8022 36408
rect 8078 36352 8083 36408
rect 4294 36350 8083 36352
rect 4294 36274 4354 36350
rect 8017 36347 8083 36350
rect 3742 36214 4354 36274
rect 3550 36076 3556 36140
rect 3620 36138 3626 36140
rect 3785 36138 3851 36141
rect 8293 36138 8359 36141
rect 3620 36136 8359 36138
rect 3620 36080 3790 36136
rect 3846 36080 8298 36136
rect 8354 36080 8359 36136
rect 3620 36078 8359 36080
rect 3620 36076 3626 36078
rect 3785 36075 3851 36078
rect 8293 36075 8359 36078
rect 10174 36076 10180 36140
rect 10244 36138 10250 36140
rect 19333 36138 19399 36141
rect 10244 36136 19399 36138
rect 10244 36080 19338 36136
rect 19394 36080 19399 36136
rect 10244 36078 19399 36080
rect 10244 36076 10250 36078
rect 19333 36075 19399 36078
rect -300 36002 160 36032
rect 5349 36002 5415 36005
rect -300 36000 5415 36002
rect -300 35944 5354 36000
rect 5410 35944 5415 36000
rect -300 35942 5415 35944
rect -300 35912 160 35942
rect 5349 35939 5415 35942
rect 24945 36002 25011 36005
rect 25540 36002 26000 36032
rect 24945 36000 26000 36002
rect 24945 35944 24950 36000
rect 25006 35944 26000 36000
rect 24945 35942 26000 35944
rect 24945 35939 25011 35942
rect 6810 35936 7126 35937
rect 6810 35872 6816 35936
rect 6880 35872 6896 35936
rect 6960 35872 6976 35936
rect 7040 35872 7056 35936
rect 7120 35872 7126 35936
rect 6810 35871 7126 35872
rect 12675 35936 12991 35937
rect 12675 35872 12681 35936
rect 12745 35872 12761 35936
rect 12825 35872 12841 35936
rect 12905 35872 12921 35936
rect 12985 35872 12991 35936
rect 12675 35871 12991 35872
rect 18540 35936 18856 35937
rect 18540 35872 18546 35936
rect 18610 35872 18626 35936
rect 18690 35872 18706 35936
rect 18770 35872 18786 35936
rect 18850 35872 18856 35936
rect 18540 35871 18856 35872
rect 24405 35936 24721 35937
rect 24405 35872 24411 35936
rect 24475 35872 24491 35936
rect 24555 35872 24571 35936
rect 24635 35872 24651 35936
rect 24715 35872 24721 35936
rect 25540 35912 26000 35942
rect 24405 35871 24721 35872
rect 4429 35866 4495 35869
rect 5533 35866 5599 35869
rect 4429 35864 5599 35866
rect 4429 35808 4434 35864
rect 4490 35808 5538 35864
rect 5594 35808 5599 35864
rect 4429 35806 5599 35808
rect 4429 35803 4495 35806
rect 5533 35803 5599 35806
rect -300 35730 160 35760
rect 3233 35730 3299 35733
rect 5257 35732 5323 35733
rect -300 35728 3299 35730
rect -300 35672 3238 35728
rect 3294 35672 3299 35728
rect -300 35670 3299 35672
rect -300 35640 160 35670
rect 3233 35667 3299 35670
rect 5206 35668 5212 35732
rect 5276 35730 5323 35732
rect 5942 35730 5948 35732
rect 5276 35728 5948 35730
rect 5318 35672 5948 35728
rect 5276 35670 5948 35672
rect 5276 35668 5323 35670
rect 5942 35668 5948 35670
rect 6012 35668 6018 35732
rect 5257 35667 5323 35668
rect 2129 35594 2195 35597
rect 8293 35594 8359 35597
rect 2129 35592 8359 35594
rect 2129 35536 2134 35592
rect 2190 35536 8298 35592
rect 8354 35536 8359 35592
rect 2129 35534 8359 35536
rect 2129 35531 2195 35534
rect 8293 35531 8359 35534
rect 10225 35594 10291 35597
rect 22502 35594 22508 35596
rect 10225 35592 22508 35594
rect 10225 35536 10230 35592
rect 10286 35536 22508 35592
rect 10225 35534 22508 35536
rect 10225 35531 10291 35534
rect 22502 35532 22508 35534
rect 22572 35532 22578 35596
rect -300 35458 160 35488
rect 3601 35458 3667 35461
rect -300 35456 3667 35458
rect -300 35400 3606 35456
rect 3662 35400 3667 35456
rect -300 35398 3667 35400
rect -300 35368 160 35398
rect 3601 35395 3667 35398
rect 24117 35458 24183 35461
rect 25540 35458 26000 35488
rect 24117 35456 26000 35458
rect 24117 35400 24122 35456
rect 24178 35400 26000 35456
rect 24117 35398 26000 35400
rect 24117 35395 24183 35398
rect 3878 35392 4194 35393
rect 3878 35328 3884 35392
rect 3948 35328 3964 35392
rect 4028 35328 4044 35392
rect 4108 35328 4124 35392
rect 4188 35328 4194 35392
rect 3878 35327 4194 35328
rect 9743 35392 10059 35393
rect 9743 35328 9749 35392
rect 9813 35328 9829 35392
rect 9893 35328 9909 35392
rect 9973 35328 9989 35392
rect 10053 35328 10059 35392
rect 9743 35327 10059 35328
rect 15608 35392 15924 35393
rect 15608 35328 15614 35392
rect 15678 35328 15694 35392
rect 15758 35328 15774 35392
rect 15838 35328 15854 35392
rect 15918 35328 15924 35392
rect 15608 35327 15924 35328
rect 21473 35392 21789 35393
rect 21473 35328 21479 35392
rect 21543 35328 21559 35392
rect 21623 35328 21639 35392
rect 21703 35328 21719 35392
rect 21783 35328 21789 35392
rect 25540 35368 26000 35398
rect 21473 35327 21789 35328
rect -300 35186 160 35216
rect 3049 35186 3115 35189
rect -300 35184 3115 35186
rect -300 35128 3054 35184
rect 3110 35128 3115 35184
rect -300 35126 3115 35128
rect -300 35096 160 35126
rect 3049 35123 3115 35126
rect 2405 35050 2471 35053
rect 4337 35050 4403 35053
rect 2405 35048 4403 35050
rect 2405 34992 2410 35048
rect 2466 34992 4342 35048
rect 4398 34992 4403 35048
rect 2405 34990 4403 34992
rect 2405 34987 2471 34990
rect 4337 34987 4403 34990
rect 6269 35050 6335 35053
rect 17902 35050 17908 35052
rect 6269 35048 17908 35050
rect 6269 34992 6274 35048
rect 6330 34992 17908 35048
rect 6269 34990 17908 34992
rect 6269 34987 6335 34990
rect 17902 34988 17908 34990
rect 17972 34988 17978 35052
rect -300 34914 160 34944
rect 2773 34914 2839 34917
rect -300 34912 2839 34914
rect -300 34856 2778 34912
rect 2834 34856 2839 34912
rect -300 34854 2839 34856
rect -300 34824 160 34854
rect 2773 34851 2839 34854
rect 24853 34914 24919 34917
rect 25540 34914 26000 34944
rect 24853 34912 26000 34914
rect 24853 34856 24858 34912
rect 24914 34856 26000 34912
rect 24853 34854 26000 34856
rect 24853 34851 24919 34854
rect 6810 34848 7126 34849
rect 6810 34784 6816 34848
rect 6880 34784 6896 34848
rect 6960 34784 6976 34848
rect 7040 34784 7056 34848
rect 7120 34784 7126 34848
rect 6810 34783 7126 34784
rect 12675 34848 12991 34849
rect 12675 34784 12681 34848
rect 12745 34784 12761 34848
rect 12825 34784 12841 34848
rect 12905 34784 12921 34848
rect 12985 34784 12991 34848
rect 12675 34783 12991 34784
rect 18540 34848 18856 34849
rect 18540 34784 18546 34848
rect 18610 34784 18626 34848
rect 18690 34784 18706 34848
rect 18770 34784 18786 34848
rect 18850 34784 18856 34848
rect 18540 34783 18856 34784
rect 24405 34848 24721 34849
rect 24405 34784 24411 34848
rect 24475 34784 24491 34848
rect 24555 34784 24571 34848
rect 24635 34784 24651 34848
rect 24715 34784 24721 34848
rect 25540 34824 26000 34854
rect 24405 34783 24721 34784
rect 933 34778 999 34781
rect 6085 34778 6151 34781
rect 933 34776 6151 34778
rect 933 34720 938 34776
rect 994 34720 6090 34776
rect 6146 34720 6151 34776
rect 933 34718 6151 34720
rect 933 34715 999 34718
rect 6085 34715 6151 34718
rect -300 34642 160 34672
rect 3877 34642 3943 34645
rect -300 34640 3943 34642
rect -300 34584 3882 34640
rect 3938 34584 3943 34640
rect -300 34582 3943 34584
rect -300 34552 160 34582
rect 3877 34579 3943 34582
rect 11697 34642 11763 34645
rect 13077 34642 13143 34645
rect 11697 34640 13143 34642
rect 11697 34584 11702 34640
rect 11758 34584 13082 34640
rect 13138 34584 13143 34640
rect 11697 34582 13143 34584
rect 11697 34579 11763 34582
rect 13077 34579 13143 34582
rect 22318 34580 22324 34644
rect 22388 34642 22394 34644
rect 23197 34642 23263 34645
rect 22388 34640 23263 34642
rect 22388 34584 23202 34640
rect 23258 34584 23263 34640
rect 22388 34582 23263 34584
rect 22388 34580 22394 34582
rect 23197 34579 23263 34582
rect 3785 34506 3851 34509
rect 2730 34504 3851 34506
rect 2730 34448 3790 34504
rect 3846 34448 3851 34504
rect 2730 34446 3851 34448
rect -300 34370 160 34400
rect 2730 34370 2790 34446
rect 3785 34443 3851 34446
rect 4797 34506 4863 34509
rect 6126 34506 6132 34508
rect 4797 34504 6132 34506
rect 4797 34448 4802 34504
rect 4858 34448 6132 34504
rect 4797 34446 6132 34448
rect 4797 34443 4863 34446
rect 6126 34444 6132 34446
rect 6196 34444 6202 34508
rect 7833 34506 7899 34509
rect 7966 34506 7972 34508
rect 7833 34504 7972 34506
rect 7833 34448 7838 34504
rect 7894 34448 7972 34504
rect 7833 34446 7972 34448
rect 7833 34443 7899 34446
rect 7966 34444 7972 34446
rect 8036 34506 8042 34508
rect 24117 34506 24183 34509
rect 8036 34446 12450 34506
rect 8036 34444 8042 34446
rect -300 34310 2790 34370
rect -300 34280 160 34310
rect 3878 34304 4194 34305
rect 3878 34240 3884 34304
rect 3948 34240 3964 34304
rect 4028 34240 4044 34304
rect 4108 34240 4124 34304
rect 4188 34240 4194 34304
rect 3878 34239 4194 34240
rect 9743 34304 10059 34305
rect 9743 34240 9749 34304
rect 9813 34240 9829 34304
rect 9893 34240 9909 34304
rect 9973 34240 9989 34304
rect 10053 34240 10059 34304
rect 9743 34239 10059 34240
rect 4889 34234 4955 34237
rect 5206 34234 5212 34236
rect 4889 34232 5212 34234
rect 4889 34176 4894 34232
rect 4950 34176 5212 34232
rect 4889 34174 5212 34176
rect 4889 34171 4955 34174
rect 5206 34172 5212 34174
rect 5276 34172 5282 34236
rect -300 34098 160 34128
rect 1393 34098 1459 34101
rect -300 34096 1459 34098
rect -300 34040 1398 34096
rect 1454 34040 1459 34096
rect -300 34038 1459 34040
rect -300 34008 160 34038
rect 1393 34035 1459 34038
rect 3693 34098 3759 34101
rect 7598 34098 7604 34100
rect 3693 34096 7604 34098
rect 3693 34040 3698 34096
rect 3754 34040 7604 34096
rect 3693 34038 7604 34040
rect 3693 34035 3759 34038
rect 7598 34036 7604 34038
rect 7668 34098 7674 34100
rect 7833 34098 7899 34101
rect 7668 34096 7899 34098
rect 7668 34040 7838 34096
rect 7894 34040 7899 34096
rect 7668 34038 7899 34040
rect 12390 34098 12450 34446
rect 24117 34504 24778 34506
rect 24117 34448 24122 34504
rect 24178 34448 24778 34504
rect 24117 34446 24778 34448
rect 24117 34443 24183 34446
rect 24718 34370 24778 34446
rect 25540 34370 26000 34400
rect 24718 34310 26000 34370
rect 15608 34304 15924 34305
rect 15608 34240 15614 34304
rect 15678 34240 15694 34304
rect 15758 34240 15774 34304
rect 15838 34240 15854 34304
rect 15918 34240 15924 34304
rect 15608 34239 15924 34240
rect 21473 34304 21789 34305
rect 21473 34240 21479 34304
rect 21543 34240 21559 34304
rect 21623 34240 21639 34304
rect 21703 34240 21719 34304
rect 21783 34240 21789 34304
rect 25540 34280 26000 34310
rect 21473 34239 21789 34240
rect 19517 34098 19583 34101
rect 12390 34096 19583 34098
rect 12390 34040 19522 34096
rect 19578 34040 19583 34096
rect 12390 34038 19583 34040
rect 7668 34036 7674 34038
rect 7833 34035 7899 34038
rect 19517 34035 19583 34038
rect 4153 33962 4219 33965
rect 4470 33962 4476 33964
rect 4153 33960 4476 33962
rect 4153 33904 4158 33960
rect 4214 33904 4476 33960
rect 4153 33902 4476 33904
rect 4153 33899 4219 33902
rect 4470 33900 4476 33902
rect 4540 33900 4546 33964
rect 10317 33962 10383 33965
rect 16757 33962 16823 33965
rect 10317 33960 16823 33962
rect 10317 33904 10322 33960
rect 10378 33904 16762 33960
rect 16818 33904 16823 33960
rect 10317 33902 16823 33904
rect 10317 33899 10383 33902
rect 16757 33899 16823 33902
rect -300 33826 160 33856
rect 1301 33826 1367 33829
rect -300 33824 1367 33826
rect -300 33768 1306 33824
rect 1362 33768 1367 33824
rect -300 33766 1367 33768
rect -300 33736 160 33766
rect 1301 33763 1367 33766
rect 4153 33826 4219 33829
rect 4889 33826 4955 33829
rect 4153 33824 4955 33826
rect 4153 33768 4158 33824
rect 4214 33768 4894 33824
rect 4950 33768 4955 33824
rect 4153 33766 4955 33768
rect 4153 33763 4219 33766
rect 4889 33763 4955 33766
rect 24853 33826 24919 33829
rect 25540 33826 26000 33856
rect 24853 33824 26000 33826
rect 24853 33768 24858 33824
rect 24914 33768 26000 33824
rect 24853 33766 26000 33768
rect 24853 33763 24919 33766
rect 6810 33760 7126 33761
rect 6810 33696 6816 33760
rect 6880 33696 6896 33760
rect 6960 33696 6976 33760
rect 7040 33696 7056 33760
rect 7120 33696 7126 33760
rect 6810 33695 7126 33696
rect 12675 33760 12991 33761
rect 12675 33696 12681 33760
rect 12745 33696 12761 33760
rect 12825 33696 12841 33760
rect 12905 33696 12921 33760
rect 12985 33696 12991 33760
rect 12675 33695 12991 33696
rect 18540 33760 18856 33761
rect 18540 33696 18546 33760
rect 18610 33696 18626 33760
rect 18690 33696 18706 33760
rect 18770 33696 18786 33760
rect 18850 33696 18856 33760
rect 18540 33695 18856 33696
rect 24405 33760 24721 33761
rect 24405 33696 24411 33760
rect 24475 33696 24491 33760
rect 24555 33696 24571 33760
rect 24635 33696 24651 33760
rect 24715 33696 24721 33760
rect 25540 33736 26000 33766
rect 24405 33695 24721 33696
rect 2221 33690 2287 33693
rect 5993 33690 6059 33693
rect 2221 33688 6059 33690
rect 2221 33632 2226 33688
rect 2282 33632 5998 33688
rect 6054 33632 6059 33688
rect 2221 33630 6059 33632
rect 2221 33627 2287 33630
rect 5993 33627 6059 33630
rect -300 33554 160 33584
rect 1117 33554 1183 33557
rect -300 33552 1183 33554
rect -300 33496 1122 33552
rect 1178 33496 1183 33552
rect -300 33494 1183 33496
rect -300 33464 160 33494
rect 1117 33491 1183 33494
rect 1669 33554 1735 33557
rect 3366 33554 3372 33556
rect 1669 33552 3372 33554
rect 1669 33496 1674 33552
rect 1730 33496 3372 33552
rect 1669 33494 3372 33496
rect 1669 33491 1735 33494
rect 3366 33492 3372 33494
rect 3436 33554 3442 33556
rect 6494 33554 6500 33556
rect 3436 33494 6500 33554
rect 3436 33492 3442 33494
rect 6494 33492 6500 33494
rect 6564 33492 6570 33556
rect 12433 33554 12499 33557
rect 24209 33554 24275 33557
rect 12433 33552 24275 33554
rect 12433 33496 12438 33552
rect 12494 33496 24214 33552
rect 24270 33496 24275 33552
rect 12433 33494 24275 33496
rect 12433 33491 12499 33494
rect 24209 33491 24275 33494
rect 3969 33418 4035 33421
rect 12249 33418 12315 33421
rect 3969 33416 12450 33418
rect 3969 33360 3974 33416
rect 4030 33360 12254 33416
rect 12310 33360 12450 33416
rect 3969 33358 12450 33360
rect 3969 33355 4035 33358
rect 12249 33355 12315 33358
rect -300 33282 160 33312
rect 1301 33282 1367 33285
rect -300 33280 1367 33282
rect -300 33224 1306 33280
rect 1362 33224 1367 33280
rect -300 33222 1367 33224
rect -300 33192 160 33222
rect 1301 33219 1367 33222
rect 4337 33282 4403 33285
rect 8845 33282 8911 33285
rect 4337 33280 8911 33282
rect 4337 33224 4342 33280
rect 4398 33224 8850 33280
rect 8906 33224 8911 33280
rect 4337 33222 8911 33224
rect 12390 33282 12450 33358
rect 12801 33282 12867 33285
rect 12390 33280 12867 33282
rect 12390 33224 12806 33280
rect 12862 33224 12867 33280
rect 12390 33222 12867 33224
rect 4337 33219 4403 33222
rect 8845 33219 8911 33222
rect 12801 33219 12867 33222
rect 24117 33282 24183 33285
rect 25540 33282 26000 33312
rect 24117 33280 26000 33282
rect 24117 33224 24122 33280
rect 24178 33224 26000 33280
rect 24117 33222 26000 33224
rect 24117 33219 24183 33222
rect 3878 33216 4194 33217
rect 3878 33152 3884 33216
rect 3948 33152 3964 33216
rect 4028 33152 4044 33216
rect 4108 33152 4124 33216
rect 4188 33152 4194 33216
rect 3878 33151 4194 33152
rect 9743 33216 10059 33217
rect 9743 33152 9749 33216
rect 9813 33152 9829 33216
rect 9893 33152 9909 33216
rect 9973 33152 9989 33216
rect 10053 33152 10059 33216
rect 9743 33151 10059 33152
rect 15608 33216 15924 33217
rect 15608 33152 15614 33216
rect 15678 33152 15694 33216
rect 15758 33152 15774 33216
rect 15838 33152 15854 33216
rect 15918 33152 15924 33216
rect 15608 33151 15924 33152
rect 21473 33216 21789 33217
rect 21473 33152 21479 33216
rect 21543 33152 21559 33216
rect 21623 33152 21639 33216
rect 21703 33152 21719 33216
rect 21783 33152 21789 33216
rect 25540 33192 26000 33222
rect 21473 33151 21789 33152
rect 1945 33146 2011 33149
rect 982 33144 2011 33146
rect 982 33088 1950 33144
rect 2006 33088 2011 33144
rect 982 33086 2011 33088
rect -300 33010 160 33040
rect 982 33010 1042 33086
rect 1945 33083 2011 33086
rect 2405 33146 2471 33149
rect 3734 33146 3740 33148
rect 2405 33144 3740 33146
rect 2405 33088 2410 33144
rect 2466 33088 3740 33144
rect 2405 33086 3740 33088
rect 2405 33083 2471 33086
rect 3734 33084 3740 33086
rect 3804 33084 3810 33148
rect 4286 33084 4292 33148
rect 4356 33146 4362 33148
rect 4429 33146 4495 33149
rect 4356 33144 4495 33146
rect 4356 33088 4434 33144
rect 4490 33088 4495 33144
rect 4356 33086 4495 33088
rect 4356 33084 4362 33086
rect 4429 33083 4495 33086
rect 6126 33084 6132 33148
rect 6196 33146 6202 33148
rect 7189 33146 7255 33149
rect 6196 33144 7255 33146
rect 6196 33088 7194 33144
rect 7250 33088 7255 33144
rect 6196 33086 7255 33088
rect 6196 33084 6202 33086
rect 7189 33083 7255 33086
rect -300 32950 1042 33010
rect 3601 33010 3667 33013
rect 5901 33010 5967 33013
rect 3601 33008 5967 33010
rect 3601 32952 3606 33008
rect 3662 32952 5906 33008
rect 5962 32952 5967 33008
rect 3601 32950 5967 32952
rect -300 32920 160 32950
rect 3601 32947 3667 32950
rect 5901 32947 5967 32950
rect 15009 33010 15075 33013
rect 15837 33010 15903 33013
rect 17217 33010 17283 33013
rect 15009 33008 17283 33010
rect 15009 32952 15014 33008
rect 15070 32952 15842 33008
rect 15898 32952 17222 33008
rect 17278 32952 17283 33008
rect 15009 32950 17283 32952
rect 15009 32947 15075 32950
rect 15837 32947 15903 32950
rect 17217 32947 17283 32950
rect 1577 32874 1643 32877
rect 2078 32874 2084 32876
rect 1577 32872 2084 32874
rect 1577 32816 1582 32872
rect 1638 32816 2084 32872
rect 1577 32814 2084 32816
rect 1577 32811 1643 32814
rect 2078 32812 2084 32814
rect 2148 32874 2154 32876
rect 10225 32874 10291 32877
rect 2148 32872 10291 32874
rect 2148 32816 10230 32872
rect 10286 32816 10291 32872
rect 2148 32814 10291 32816
rect 2148 32812 2154 32814
rect 10225 32811 10291 32814
rect 14365 32874 14431 32877
rect 15285 32874 15351 32877
rect 14365 32872 15351 32874
rect 14365 32816 14370 32872
rect 14426 32816 15290 32872
rect 15346 32816 15351 32872
rect 14365 32814 15351 32816
rect 14365 32811 14431 32814
rect 15285 32811 15351 32814
rect -300 32738 160 32768
rect 3141 32738 3207 32741
rect -300 32736 3207 32738
rect -300 32680 3146 32736
rect 3202 32680 3207 32736
rect -300 32678 3207 32680
rect -300 32648 160 32678
rect 3141 32675 3207 32678
rect 24853 32738 24919 32741
rect 25540 32738 26000 32768
rect 24853 32736 26000 32738
rect 24853 32680 24858 32736
rect 24914 32680 26000 32736
rect 24853 32678 26000 32680
rect 24853 32675 24919 32678
rect 6810 32672 7126 32673
rect 6810 32608 6816 32672
rect 6880 32608 6896 32672
rect 6960 32608 6976 32672
rect 7040 32608 7056 32672
rect 7120 32608 7126 32672
rect 6810 32607 7126 32608
rect 12675 32672 12991 32673
rect 12675 32608 12681 32672
rect 12745 32608 12761 32672
rect 12825 32608 12841 32672
rect 12905 32608 12921 32672
rect 12985 32608 12991 32672
rect 12675 32607 12991 32608
rect 18540 32672 18856 32673
rect 18540 32608 18546 32672
rect 18610 32608 18626 32672
rect 18690 32608 18706 32672
rect 18770 32608 18786 32672
rect 18850 32608 18856 32672
rect 18540 32607 18856 32608
rect 24405 32672 24721 32673
rect 24405 32608 24411 32672
rect 24475 32608 24491 32672
rect 24555 32608 24571 32672
rect 24635 32608 24651 32672
rect 24715 32608 24721 32672
rect 25540 32648 26000 32678
rect 24405 32607 24721 32608
rect 1393 32600 1459 32605
rect 10174 32602 10180 32604
rect 1393 32544 1398 32600
rect 1454 32544 1459 32600
rect 1393 32539 1459 32544
rect 7192 32542 10180 32602
rect -300 32466 160 32496
rect 1396 32466 1456 32539
rect -300 32406 1456 32466
rect 5349 32466 5415 32469
rect 7192 32466 7252 32542
rect 10174 32540 10180 32542
rect 10244 32540 10250 32604
rect 7741 32468 7807 32469
rect 7741 32466 7788 32468
rect 5349 32464 7252 32466
rect 5349 32408 5354 32464
rect 5410 32408 7252 32464
rect 5349 32406 7252 32408
rect 7700 32464 7788 32466
rect 7852 32466 7858 32468
rect 15101 32466 15167 32469
rect 7852 32464 15167 32466
rect 7700 32408 7746 32464
rect 7852 32408 15106 32464
rect 15162 32408 15167 32464
rect 7700 32406 7788 32408
rect -300 32376 160 32406
rect 5349 32403 5415 32406
rect 7741 32404 7788 32406
rect 7852 32406 15167 32408
rect 7852 32404 7858 32406
rect 7741 32403 7807 32404
rect 15101 32403 15167 32406
rect 1393 32330 1459 32333
rect 2446 32330 2452 32332
rect 1393 32328 2452 32330
rect 1393 32272 1398 32328
rect 1454 32272 2452 32328
rect 1393 32270 2452 32272
rect 1393 32267 1459 32270
rect 2446 32268 2452 32270
rect 2516 32330 2522 32332
rect 7925 32330 7991 32333
rect 8150 32330 8156 32332
rect 2516 32270 2790 32330
rect 2516 32268 2522 32270
rect -300 32194 160 32224
rect 1669 32194 1735 32197
rect 2589 32194 2655 32197
rect -300 32134 1594 32194
rect -300 32104 160 32134
rect -300 31922 160 31952
rect 1301 31922 1367 31925
rect -300 31920 1367 31922
rect -300 31864 1306 31920
rect 1362 31864 1367 31920
rect -300 31862 1367 31864
rect -300 31832 160 31862
rect 1301 31859 1367 31862
rect 1301 31786 1367 31789
rect 1534 31786 1594 32134
rect 1669 32192 2655 32194
rect 1669 32136 1674 32192
rect 1730 32136 2594 32192
rect 2650 32136 2655 32192
rect 1669 32134 2655 32136
rect 1669 32131 1735 32134
rect 2589 32131 2655 32134
rect 2730 31922 2790 32270
rect 7925 32328 8156 32330
rect 7925 32272 7930 32328
rect 7986 32272 8156 32328
rect 7925 32270 8156 32272
rect 7925 32267 7991 32270
rect 8150 32268 8156 32270
rect 8220 32330 8226 32332
rect 8220 32270 10242 32330
rect 8220 32268 8226 32270
rect 5942 32132 5948 32196
rect 6012 32194 6018 32196
rect 8753 32194 8819 32197
rect 6012 32192 8819 32194
rect 6012 32136 8758 32192
rect 8814 32136 8819 32192
rect 6012 32134 8819 32136
rect 6012 32132 6018 32134
rect 8753 32131 8819 32134
rect 3878 32128 4194 32129
rect 3878 32064 3884 32128
rect 3948 32064 3964 32128
rect 4028 32064 4044 32128
rect 4108 32064 4124 32128
rect 4188 32064 4194 32128
rect 3878 32063 4194 32064
rect 9743 32128 10059 32129
rect 9743 32064 9749 32128
rect 9813 32064 9829 32128
rect 9893 32064 9909 32128
rect 9973 32064 9989 32128
rect 10053 32064 10059 32128
rect 9743 32063 10059 32064
rect 10182 32058 10242 32270
rect 11094 32268 11100 32332
rect 11164 32330 11170 32332
rect 11697 32330 11763 32333
rect 11164 32328 11763 32330
rect 11164 32272 11702 32328
rect 11758 32272 11763 32328
rect 11164 32270 11763 32272
rect 11164 32268 11170 32270
rect 11697 32267 11763 32270
rect 14273 32330 14339 32333
rect 16757 32330 16823 32333
rect 14273 32328 16823 32330
rect 14273 32272 14278 32328
rect 14334 32272 16762 32328
rect 16818 32272 16823 32328
rect 14273 32270 16823 32272
rect 14273 32267 14339 32270
rect 16757 32267 16823 32270
rect 24117 32194 24183 32197
rect 25540 32194 26000 32224
rect 24117 32192 26000 32194
rect 24117 32136 24122 32192
rect 24178 32136 26000 32192
rect 24117 32134 26000 32136
rect 24117 32131 24183 32134
rect 15608 32128 15924 32129
rect 15608 32064 15614 32128
rect 15678 32064 15694 32128
rect 15758 32064 15774 32128
rect 15838 32064 15854 32128
rect 15918 32064 15924 32128
rect 15608 32063 15924 32064
rect 21473 32128 21789 32129
rect 21473 32064 21479 32128
rect 21543 32064 21559 32128
rect 21623 32064 21639 32128
rect 21703 32064 21719 32128
rect 21783 32064 21789 32128
rect 25540 32104 26000 32134
rect 21473 32063 21789 32064
rect 10182 31998 15394 32058
rect 9857 31922 9923 31925
rect 15142 31922 15148 31924
rect 2730 31920 9923 31922
rect 2730 31864 9862 31920
rect 9918 31864 9923 31920
rect 2730 31862 9923 31864
rect 9857 31859 9923 31862
rect 12390 31862 15148 31922
rect 1301 31784 1594 31786
rect 1301 31728 1306 31784
rect 1362 31728 1594 31784
rect 1301 31726 1594 31728
rect 2497 31786 2563 31789
rect 2814 31786 2820 31788
rect 2497 31784 2820 31786
rect 2497 31728 2502 31784
rect 2558 31728 2820 31784
rect 2497 31726 2820 31728
rect 1301 31723 1367 31726
rect 2497 31723 2563 31726
rect 2814 31724 2820 31726
rect 2884 31724 2890 31788
rect 5349 31786 5415 31789
rect 5574 31786 5580 31788
rect 5349 31784 5580 31786
rect 5349 31728 5354 31784
rect 5410 31728 5580 31784
rect 5349 31726 5580 31728
rect 5349 31723 5415 31726
rect 5574 31724 5580 31726
rect 5644 31724 5650 31788
rect 5993 31786 6059 31789
rect 12390 31786 12450 31862
rect 15142 31860 15148 31862
rect 15212 31860 15218 31924
rect 15334 31922 15394 31998
rect 16573 31922 16639 31925
rect 15334 31920 16639 31922
rect 15334 31864 16578 31920
rect 16634 31864 16639 31920
rect 15334 31862 16639 31864
rect 16573 31859 16639 31862
rect 5993 31784 8034 31786
rect 5993 31728 5998 31784
rect 6054 31770 8034 31784
rect 8526 31770 12450 31786
rect 6054 31728 12450 31770
rect 5993 31726 12450 31728
rect 18781 31786 18847 31789
rect 19333 31786 19399 31789
rect 18781 31784 19399 31786
rect 18781 31728 18786 31784
rect 18842 31728 19338 31784
rect 19394 31728 19399 31784
rect 18781 31726 19399 31728
rect 5993 31723 6059 31726
rect 7974 31710 8586 31726
rect 18781 31723 18847 31726
rect 19333 31723 19399 31726
rect -300 31650 160 31680
rect 5349 31650 5415 31653
rect 7649 31652 7715 31653
rect -300 31648 5415 31650
rect -300 31592 5354 31648
rect 5410 31592 5415 31648
rect -300 31590 5415 31592
rect -300 31560 160 31590
rect 5349 31587 5415 31590
rect 7598 31588 7604 31652
rect 7668 31650 7715 31652
rect 25037 31650 25103 31653
rect 25540 31650 26000 31680
rect 7668 31648 7760 31650
rect 7710 31592 7760 31648
rect 7668 31590 7760 31592
rect 25037 31648 26000 31650
rect 25037 31592 25042 31648
rect 25098 31592 26000 31648
rect 25037 31590 26000 31592
rect 7668 31588 7715 31590
rect 7649 31587 7715 31588
rect 25037 31587 25103 31590
rect 6810 31584 7126 31585
rect 6810 31520 6816 31584
rect 6880 31520 6896 31584
rect 6960 31520 6976 31584
rect 7040 31520 7056 31584
rect 7120 31520 7126 31584
rect 6810 31519 7126 31520
rect 12675 31584 12991 31585
rect 12675 31520 12681 31584
rect 12745 31520 12761 31584
rect 12825 31520 12841 31584
rect 12905 31520 12921 31584
rect 12985 31520 12991 31584
rect 12675 31519 12991 31520
rect 18540 31584 18856 31585
rect 18540 31520 18546 31584
rect 18610 31520 18626 31584
rect 18690 31520 18706 31584
rect 18770 31520 18786 31584
rect 18850 31520 18856 31584
rect 18540 31519 18856 31520
rect 24405 31584 24721 31585
rect 24405 31520 24411 31584
rect 24475 31520 24491 31584
rect 24555 31520 24571 31584
rect 24635 31520 24651 31584
rect 24715 31520 24721 31584
rect 25540 31560 26000 31590
rect 24405 31519 24721 31520
rect 2630 31452 2636 31516
rect 2700 31514 2706 31516
rect 3509 31514 3575 31517
rect 5533 31516 5599 31517
rect 5533 31514 5580 31516
rect 2700 31512 3575 31514
rect 2700 31456 3514 31512
rect 3570 31456 3575 31512
rect 2700 31454 3575 31456
rect 5452 31512 5580 31514
rect 5644 31514 5650 31516
rect 5901 31514 5967 31517
rect 5644 31512 5967 31514
rect 5452 31456 5538 31512
rect 5644 31456 5906 31512
rect 5962 31456 5967 31512
rect 5452 31454 5580 31456
rect 2700 31452 2706 31454
rect 3509 31451 3575 31454
rect 5533 31452 5580 31454
rect 5644 31454 5967 31456
rect 5644 31452 5650 31454
rect 5533 31451 5599 31452
rect 5901 31451 5967 31454
rect -300 31378 160 31408
rect 1301 31378 1367 31381
rect -300 31376 1367 31378
rect -300 31320 1306 31376
rect 1362 31320 1367 31376
rect -300 31318 1367 31320
rect -300 31288 160 31318
rect 1301 31315 1367 31318
rect 2630 31316 2636 31380
rect 2700 31378 2706 31380
rect 9581 31378 9647 31381
rect 2700 31376 9647 31378
rect 2700 31320 9586 31376
rect 9642 31320 9647 31376
rect 2700 31318 9647 31320
rect 2700 31316 2706 31318
rect 9581 31315 9647 31318
rect 2865 31242 2931 31245
rect 5717 31242 5783 31245
rect 2865 31240 5783 31242
rect 2865 31184 2870 31240
rect 2926 31184 5722 31240
rect 5778 31184 5783 31240
rect 2865 31182 5783 31184
rect 2865 31179 2931 31182
rect 5717 31179 5783 31182
rect 10174 31180 10180 31244
rect 10244 31242 10250 31244
rect 10961 31242 11027 31245
rect 10244 31240 11027 31242
rect 10244 31184 10966 31240
rect 11022 31184 11027 31240
rect 10244 31182 11027 31184
rect 10244 31180 10250 31182
rect 10961 31179 11027 31182
rect 11973 31242 12039 31245
rect 12249 31242 12315 31245
rect 11973 31240 12315 31242
rect 11973 31184 11978 31240
rect 12034 31184 12254 31240
rect 12310 31184 12315 31240
rect 11973 31182 12315 31184
rect 11973 31179 12039 31182
rect 12249 31179 12315 31182
rect 12801 31242 12867 31245
rect 14089 31242 14155 31245
rect 12801 31240 14155 31242
rect 12801 31184 12806 31240
rect 12862 31184 14094 31240
rect 14150 31184 14155 31240
rect 12801 31182 14155 31184
rect 12801 31179 12867 31182
rect 14089 31179 14155 31182
rect -300 31106 160 31136
rect 1485 31106 1551 31109
rect -300 31104 1551 31106
rect -300 31048 1490 31104
rect 1546 31048 1551 31104
rect -300 31046 1551 31048
rect -300 31016 160 31046
rect 1485 31043 1551 31046
rect 4429 31106 4495 31109
rect 4797 31106 4863 31109
rect 8109 31106 8175 31109
rect 4429 31104 8175 31106
rect 4429 31048 4434 31104
rect 4490 31048 4802 31104
rect 4858 31048 8114 31104
rect 8170 31048 8175 31104
rect 4429 31046 8175 31048
rect 4429 31043 4495 31046
rect 4797 31043 4863 31046
rect 8109 31043 8175 31046
rect 24117 31106 24183 31109
rect 25540 31106 26000 31136
rect 24117 31104 26000 31106
rect 24117 31048 24122 31104
rect 24178 31048 26000 31104
rect 24117 31046 26000 31048
rect 24117 31043 24183 31046
rect 3878 31040 4194 31041
rect 3878 30976 3884 31040
rect 3948 30976 3964 31040
rect 4028 30976 4044 31040
rect 4108 30976 4124 31040
rect 4188 30976 4194 31040
rect 3878 30975 4194 30976
rect 9743 31040 10059 31041
rect 9743 30976 9749 31040
rect 9813 30976 9829 31040
rect 9893 30976 9909 31040
rect 9973 30976 9989 31040
rect 10053 30976 10059 31040
rect 9743 30975 10059 30976
rect 15608 31040 15924 31041
rect 15608 30976 15614 31040
rect 15678 30976 15694 31040
rect 15758 30976 15774 31040
rect 15838 30976 15854 31040
rect 15918 30976 15924 31040
rect 15608 30975 15924 30976
rect 21473 31040 21789 31041
rect 21473 30976 21479 31040
rect 21543 30976 21559 31040
rect 21623 30976 21639 31040
rect 21703 30976 21719 31040
rect 21783 30976 21789 31040
rect 25540 31016 26000 31046
rect 21473 30975 21789 30976
rect 4337 30970 4403 30973
rect 9121 30970 9187 30973
rect 4337 30968 9187 30970
rect 4337 30912 4342 30968
rect 4398 30912 9126 30968
rect 9182 30912 9187 30968
rect 4337 30910 9187 30912
rect 4337 30907 4403 30910
rect 9121 30907 9187 30910
rect -300 30834 160 30864
rect 2037 30834 2103 30837
rect -300 30832 2103 30834
rect -300 30776 2042 30832
rect 2098 30776 2103 30832
rect -300 30774 2103 30776
rect -300 30744 160 30774
rect 2037 30771 2103 30774
rect 3601 30834 3667 30837
rect 4797 30834 4863 30837
rect 3601 30832 4863 30834
rect 3601 30776 3606 30832
rect 3662 30776 4802 30832
rect 4858 30776 4863 30832
rect 3601 30774 4863 30776
rect 3601 30771 3667 30774
rect 4797 30771 4863 30774
rect 5257 30834 5323 30837
rect 11605 30834 11671 30837
rect 5257 30832 11671 30834
rect 5257 30776 5262 30832
rect 5318 30776 11610 30832
rect 11666 30776 11671 30832
rect 5257 30774 11671 30776
rect 5257 30771 5323 30774
rect 11605 30771 11671 30774
rect 4613 30698 4679 30701
rect 11053 30698 11119 30701
rect 4613 30696 11119 30698
rect 4613 30640 4618 30696
rect 4674 30640 11058 30696
rect 11114 30640 11119 30696
rect 4613 30638 11119 30640
rect 4613 30635 4679 30638
rect 11053 30635 11119 30638
rect -300 30562 160 30592
rect 3417 30562 3483 30565
rect -300 30560 3483 30562
rect -300 30504 3422 30560
rect 3478 30504 3483 30560
rect -300 30502 3483 30504
rect -300 30472 160 30502
rect 3417 30499 3483 30502
rect 10777 30562 10843 30565
rect 12525 30562 12591 30565
rect 10777 30560 12591 30562
rect 10777 30504 10782 30560
rect 10838 30504 12530 30560
rect 12586 30504 12591 30560
rect 10777 30502 12591 30504
rect 10777 30499 10843 30502
rect 12525 30499 12591 30502
rect 24853 30562 24919 30565
rect 25540 30562 26000 30592
rect 24853 30560 26000 30562
rect 24853 30504 24858 30560
rect 24914 30504 26000 30560
rect 24853 30502 26000 30504
rect 24853 30499 24919 30502
rect 6810 30496 7126 30497
rect 6810 30432 6816 30496
rect 6880 30432 6896 30496
rect 6960 30432 6976 30496
rect 7040 30432 7056 30496
rect 7120 30432 7126 30496
rect 6810 30431 7126 30432
rect 12675 30496 12991 30497
rect 12675 30432 12681 30496
rect 12745 30432 12761 30496
rect 12825 30432 12841 30496
rect 12905 30432 12921 30496
rect 12985 30432 12991 30496
rect 12675 30431 12991 30432
rect 18540 30496 18856 30497
rect 18540 30432 18546 30496
rect 18610 30432 18626 30496
rect 18690 30432 18706 30496
rect 18770 30432 18786 30496
rect 18850 30432 18856 30496
rect 18540 30431 18856 30432
rect 24405 30496 24721 30497
rect 24405 30432 24411 30496
rect 24475 30432 24491 30496
rect 24555 30432 24571 30496
rect 24635 30432 24651 30496
rect 24715 30432 24721 30496
rect 25540 30472 26000 30502
rect 24405 30431 24721 30432
rect 381 30426 447 30429
rect 4153 30426 4219 30429
rect 4797 30426 4863 30429
rect 381 30424 4863 30426
rect 381 30368 386 30424
rect 442 30368 4158 30424
rect 4214 30368 4802 30424
rect 4858 30368 4863 30424
rect 381 30366 4863 30368
rect 381 30363 447 30366
rect 4153 30363 4219 30366
rect 4797 30363 4863 30366
rect 10174 30364 10180 30428
rect 10244 30426 10250 30428
rect 10593 30426 10659 30429
rect 10244 30424 10659 30426
rect 10244 30368 10598 30424
rect 10654 30368 10659 30424
rect 10244 30366 10659 30368
rect 10244 30364 10250 30366
rect 10593 30363 10659 30366
rect 11053 30426 11119 30429
rect 11462 30426 11468 30428
rect 11053 30424 11468 30426
rect 11053 30368 11058 30424
rect 11114 30368 11468 30424
rect 11053 30366 11468 30368
rect 11053 30363 11119 30366
rect 11462 30364 11468 30366
rect 11532 30364 11538 30428
rect 11881 30426 11947 30429
rect 12014 30426 12020 30428
rect 11881 30424 12020 30426
rect 11881 30368 11886 30424
rect 11942 30368 12020 30424
rect 11881 30366 12020 30368
rect 11881 30363 11947 30366
rect 12014 30364 12020 30366
rect 12084 30364 12090 30428
rect -300 30290 160 30320
rect 3049 30290 3115 30293
rect -300 30288 3115 30290
rect -300 30232 3054 30288
rect 3110 30232 3115 30288
rect -300 30230 3115 30232
rect -300 30200 160 30230
rect 3049 30227 3115 30230
rect 5206 30228 5212 30292
rect 5276 30290 5282 30292
rect 10961 30290 11027 30293
rect 5276 30288 11027 30290
rect 5276 30232 10966 30288
rect 11022 30232 11027 30288
rect 5276 30230 11027 30232
rect 5276 30228 5282 30230
rect 10961 30227 11027 30230
rect 1526 30092 1532 30156
rect 1596 30154 1602 30156
rect 4061 30154 4127 30157
rect 1596 30152 4127 30154
rect 1596 30096 4066 30152
rect 4122 30096 4127 30152
rect 1596 30094 4127 30096
rect 1596 30092 1602 30094
rect 4061 30091 4127 30094
rect 5901 30154 5967 30157
rect 11513 30154 11579 30157
rect 5901 30152 11579 30154
rect 5901 30096 5906 30152
rect 5962 30096 11518 30152
rect 11574 30096 11579 30152
rect 5901 30094 11579 30096
rect 5901 30091 5967 30094
rect 11513 30091 11579 30094
rect -300 30018 160 30048
rect 1301 30018 1367 30021
rect -300 30016 1367 30018
rect -300 29960 1306 30016
rect 1362 29960 1367 30016
rect -300 29958 1367 29960
rect -300 29928 160 29958
rect 1301 29955 1367 29958
rect 6821 30018 6887 30021
rect 7966 30018 7972 30020
rect 6821 30016 7972 30018
rect 6821 29960 6826 30016
rect 6882 29960 7972 30016
rect 6821 29958 7972 29960
rect 6821 29955 6887 29958
rect 7966 29956 7972 29958
rect 8036 29956 8042 30020
rect 24117 30018 24183 30021
rect 25540 30018 26000 30048
rect 24117 30016 26000 30018
rect 24117 29960 24122 30016
rect 24178 29960 26000 30016
rect 24117 29958 26000 29960
rect 24117 29955 24183 29958
rect 3878 29952 4194 29953
rect 3878 29888 3884 29952
rect 3948 29888 3964 29952
rect 4028 29888 4044 29952
rect 4108 29888 4124 29952
rect 4188 29888 4194 29952
rect 3878 29887 4194 29888
rect 9743 29952 10059 29953
rect 9743 29888 9749 29952
rect 9813 29888 9829 29952
rect 9893 29888 9909 29952
rect 9973 29888 9989 29952
rect 10053 29888 10059 29952
rect 9743 29887 10059 29888
rect 15608 29952 15924 29953
rect 15608 29888 15614 29952
rect 15678 29888 15694 29952
rect 15758 29888 15774 29952
rect 15838 29888 15854 29952
rect 15918 29888 15924 29952
rect 15608 29887 15924 29888
rect 21473 29952 21789 29953
rect 21473 29888 21479 29952
rect 21543 29888 21559 29952
rect 21623 29888 21639 29952
rect 21703 29888 21719 29952
rect 21783 29888 21789 29952
rect 25540 29928 26000 29958
rect 21473 29887 21789 29888
rect 5022 29820 5028 29884
rect 5092 29882 5098 29884
rect 8702 29882 8708 29884
rect 5092 29822 8708 29882
rect 5092 29820 5098 29822
rect 8702 29820 8708 29822
rect 8772 29882 8778 29884
rect 9029 29882 9095 29885
rect 8772 29880 9095 29882
rect 8772 29824 9034 29880
rect 9090 29824 9095 29880
rect 8772 29822 9095 29824
rect 8772 29820 8778 29822
rect 9029 29819 9095 29822
rect -300 29746 160 29776
rect 749 29746 815 29749
rect 14641 29746 14707 29749
rect -300 29744 815 29746
rect -300 29688 754 29744
rect 810 29688 815 29744
rect -300 29686 815 29688
rect -300 29656 160 29686
rect 749 29683 815 29686
rect 2730 29744 14707 29746
rect 2730 29688 14646 29744
rect 14702 29688 14707 29744
rect 2730 29686 14707 29688
rect 2405 29610 2471 29613
rect 2730 29610 2790 29686
rect 14641 29683 14707 29686
rect 15653 29746 15719 29749
rect 16665 29746 16731 29749
rect 15653 29744 16731 29746
rect 15653 29688 15658 29744
rect 15714 29688 16670 29744
rect 16726 29688 16731 29744
rect 15653 29686 16731 29688
rect 15653 29683 15719 29686
rect 16665 29683 16731 29686
rect 2405 29608 2790 29610
rect 2405 29552 2410 29608
rect 2466 29552 2790 29608
rect 2405 29550 2790 29552
rect 3509 29610 3575 29613
rect 5993 29610 6059 29613
rect 3509 29608 6059 29610
rect 3509 29552 3514 29608
rect 3570 29552 5998 29608
rect 6054 29552 6059 29608
rect 3509 29550 6059 29552
rect 2405 29547 2471 29550
rect 3509 29547 3575 29550
rect 5993 29547 6059 29550
rect 11513 29610 11579 29613
rect 16430 29610 16436 29612
rect 11513 29608 16436 29610
rect 11513 29552 11518 29608
rect 11574 29552 16436 29608
rect 11513 29550 16436 29552
rect 11513 29547 11579 29550
rect 16430 29548 16436 29550
rect 16500 29548 16506 29612
rect -300 29474 160 29504
rect 1301 29474 1367 29477
rect -300 29472 1367 29474
rect -300 29416 1306 29472
rect 1362 29416 1367 29472
rect -300 29414 1367 29416
rect -300 29384 160 29414
rect 1301 29411 1367 29414
rect 1710 29412 1716 29476
rect 1780 29474 1786 29476
rect 1853 29474 1919 29477
rect 6637 29474 6703 29477
rect 1780 29472 6703 29474
rect 1780 29416 1858 29472
rect 1914 29416 6642 29472
rect 6698 29416 6703 29472
rect 1780 29414 6703 29416
rect 1780 29412 1786 29414
rect 1853 29411 1919 29414
rect 6637 29411 6703 29414
rect 16665 29474 16731 29477
rect 17585 29474 17651 29477
rect 16665 29472 17651 29474
rect 16665 29416 16670 29472
rect 16726 29416 17590 29472
rect 17646 29416 17651 29472
rect 16665 29414 17651 29416
rect 16665 29411 16731 29414
rect 17585 29411 17651 29414
rect 24853 29474 24919 29477
rect 25540 29474 26000 29504
rect 24853 29472 26000 29474
rect 24853 29416 24858 29472
rect 24914 29416 26000 29472
rect 24853 29414 26000 29416
rect 24853 29411 24919 29414
rect 6810 29408 7126 29409
rect 6810 29344 6816 29408
rect 6880 29344 6896 29408
rect 6960 29344 6976 29408
rect 7040 29344 7056 29408
rect 7120 29344 7126 29408
rect 6810 29343 7126 29344
rect 12675 29408 12991 29409
rect 12675 29344 12681 29408
rect 12745 29344 12761 29408
rect 12825 29344 12841 29408
rect 12905 29344 12921 29408
rect 12985 29344 12991 29408
rect 12675 29343 12991 29344
rect 18540 29408 18856 29409
rect 18540 29344 18546 29408
rect 18610 29344 18626 29408
rect 18690 29344 18706 29408
rect 18770 29344 18786 29408
rect 18850 29344 18856 29408
rect 18540 29343 18856 29344
rect 24405 29408 24721 29409
rect 24405 29344 24411 29408
rect 24475 29344 24491 29408
rect 24555 29344 24571 29408
rect 24635 29344 24651 29408
rect 24715 29344 24721 29408
rect 25540 29384 26000 29414
rect 24405 29343 24721 29344
rect 1853 29338 1919 29341
rect 5165 29338 5231 29341
rect 12065 29338 12131 29341
rect 1853 29336 5231 29338
rect 1853 29280 1858 29336
rect 1914 29280 5170 29336
rect 5226 29280 5231 29336
rect 1853 29278 5231 29280
rect 1853 29275 1919 29278
rect 5165 29275 5231 29278
rect 9630 29336 12131 29338
rect 9630 29280 12070 29336
rect 12126 29280 12131 29336
rect 9630 29278 12131 29280
rect -300 29202 160 29232
rect 1301 29202 1367 29205
rect 9630 29202 9690 29278
rect 12065 29275 12131 29278
rect 15929 29338 15995 29341
rect 16757 29338 16823 29341
rect 15929 29336 16823 29338
rect 15929 29280 15934 29336
rect 15990 29280 16762 29336
rect 16818 29280 16823 29336
rect 15929 29278 16823 29280
rect 15929 29275 15995 29278
rect 16757 29275 16823 29278
rect -300 29200 1367 29202
rect -300 29144 1306 29200
rect 1362 29144 1367 29200
rect -300 29142 1367 29144
rect -300 29112 160 29142
rect 1301 29139 1367 29142
rect 2730 29142 9690 29202
rect 10133 29200 10199 29205
rect 10133 29144 10138 29200
rect 10194 29144 10199 29200
rect 2589 29066 2655 29069
rect 2730 29066 2790 29142
rect 10133 29139 10199 29144
rect 11237 29202 11303 29205
rect 18086 29202 18092 29204
rect 11237 29200 18092 29202
rect 11237 29144 11242 29200
rect 11298 29144 18092 29200
rect 11237 29142 18092 29144
rect 11237 29139 11303 29142
rect 18086 29140 18092 29142
rect 18156 29140 18162 29204
rect 20437 29202 20503 29205
rect 20621 29202 20687 29205
rect 21081 29202 21147 29205
rect 20437 29200 21147 29202
rect 20437 29144 20442 29200
rect 20498 29144 20626 29200
rect 20682 29144 21086 29200
rect 21142 29144 21147 29200
rect 20437 29142 21147 29144
rect 20437 29139 20503 29142
rect 20621 29139 20687 29142
rect 21081 29139 21147 29142
rect 2589 29064 2790 29066
rect 2589 29008 2594 29064
rect 2650 29008 2790 29064
rect 2589 29006 2790 29008
rect 3509 29066 3575 29069
rect 5574 29066 5580 29068
rect 3509 29064 5580 29066
rect 3509 29008 3514 29064
rect 3570 29008 5580 29064
rect 3509 29006 5580 29008
rect 2589 29003 2655 29006
rect 3509 29003 3575 29006
rect 5574 29004 5580 29006
rect 5644 29004 5650 29068
rect 6177 29066 6243 29069
rect 6494 29066 6500 29068
rect 6177 29064 6500 29066
rect 6177 29008 6182 29064
rect 6238 29008 6500 29064
rect 6177 29006 6500 29008
rect 6177 29003 6243 29006
rect 6494 29004 6500 29006
rect 6564 29004 6570 29068
rect 10136 29066 10196 29139
rect 10136 29006 10242 29066
rect -300 28930 160 28960
rect 2405 28930 2471 28933
rect -300 28928 2471 28930
rect -300 28872 2410 28928
rect 2466 28872 2471 28928
rect -300 28870 2471 28872
rect 10182 28930 10242 29006
rect 13118 29004 13124 29068
rect 13188 29066 13194 29068
rect 13445 29066 13511 29069
rect 13188 29064 13511 29066
rect 13188 29008 13450 29064
rect 13506 29008 13511 29064
rect 13188 29006 13511 29008
rect 13188 29004 13194 29006
rect 13445 29003 13511 29006
rect 14641 29066 14707 29069
rect 15009 29066 15075 29069
rect 14641 29064 15075 29066
rect 14641 29008 14646 29064
rect 14702 29008 15014 29064
rect 15070 29008 15075 29064
rect 14641 29006 15075 29008
rect 14641 29003 14707 29006
rect 15009 29003 15075 29006
rect 16481 29066 16547 29069
rect 20846 29066 20852 29068
rect 16481 29064 20852 29066
rect 16481 29008 16486 29064
rect 16542 29008 20852 29064
rect 16481 29006 20852 29008
rect 16481 29003 16547 29006
rect 20846 29004 20852 29006
rect 20916 29004 20922 29068
rect 10317 28930 10383 28933
rect 11513 28930 11579 28933
rect 10182 28928 11579 28930
rect 10182 28872 10322 28928
rect 10378 28872 11518 28928
rect 11574 28872 11579 28928
rect 10182 28870 11579 28872
rect -300 28840 160 28870
rect 2405 28867 2471 28870
rect 10317 28867 10383 28870
rect 11513 28867 11579 28870
rect 24117 28930 24183 28933
rect 25540 28930 26000 28960
rect 24117 28928 26000 28930
rect 24117 28872 24122 28928
rect 24178 28872 26000 28928
rect 24117 28870 26000 28872
rect 24117 28867 24183 28870
rect 3878 28864 4194 28865
rect 3878 28800 3884 28864
rect 3948 28800 3964 28864
rect 4028 28800 4044 28864
rect 4108 28800 4124 28864
rect 4188 28800 4194 28864
rect 3878 28799 4194 28800
rect 9743 28864 10059 28865
rect 9743 28800 9749 28864
rect 9813 28800 9829 28864
rect 9893 28800 9909 28864
rect 9973 28800 9989 28864
rect 10053 28800 10059 28864
rect 9743 28799 10059 28800
rect 15608 28864 15924 28865
rect 15608 28800 15614 28864
rect 15678 28800 15694 28864
rect 15758 28800 15774 28864
rect 15838 28800 15854 28864
rect 15918 28800 15924 28864
rect 15608 28799 15924 28800
rect 21473 28864 21789 28865
rect 21473 28800 21479 28864
rect 21543 28800 21559 28864
rect 21623 28800 21639 28864
rect 21703 28800 21719 28864
rect 21783 28800 21789 28864
rect 25540 28840 26000 28870
rect 21473 28799 21789 28800
rect 473 28794 539 28797
rect 473 28792 3618 28794
rect 473 28736 478 28792
rect 534 28736 3618 28792
rect 473 28734 3618 28736
rect 473 28731 539 28734
rect -300 28658 160 28688
rect 2773 28658 2839 28661
rect -300 28656 2839 28658
rect -300 28600 2778 28656
rect 2834 28600 2839 28656
rect -300 28598 2839 28600
rect 3558 28658 3618 28734
rect 8569 28658 8635 28661
rect 3558 28656 8635 28658
rect 3558 28600 8574 28656
rect 8630 28600 8635 28656
rect 3558 28598 8635 28600
rect -300 28568 160 28598
rect 2773 28595 2839 28598
rect 8569 28595 8635 28598
rect 11237 28658 11303 28661
rect 18045 28658 18111 28661
rect 11237 28656 18111 28658
rect 11237 28600 11242 28656
rect 11298 28600 18050 28656
rect 18106 28600 18111 28656
rect 11237 28598 18111 28600
rect 11237 28595 11303 28598
rect 18045 28595 18111 28598
rect 1393 28522 1459 28525
rect 798 28520 1459 28522
rect 798 28464 1398 28520
rect 1454 28464 1459 28520
rect 798 28462 1459 28464
rect -300 28386 160 28416
rect 798 28386 858 28462
rect 1393 28459 1459 28462
rect 6310 28460 6316 28524
rect 6380 28522 6386 28524
rect 7649 28522 7715 28525
rect 6380 28520 7715 28522
rect 6380 28464 7654 28520
rect 7710 28464 7715 28520
rect 6380 28462 7715 28464
rect 6380 28460 6386 28462
rect 7649 28459 7715 28462
rect 8702 28460 8708 28524
rect 8772 28522 8778 28524
rect 14038 28522 14044 28524
rect 8772 28462 14044 28522
rect 8772 28460 8778 28462
rect 14038 28460 14044 28462
rect 14108 28460 14114 28524
rect -300 28326 858 28386
rect 3693 28386 3759 28389
rect 5165 28386 5231 28389
rect 3693 28384 5231 28386
rect 3693 28328 3698 28384
rect 3754 28328 5170 28384
rect 5226 28328 5231 28384
rect 3693 28326 5231 28328
rect -300 28296 160 28326
rect 3693 28323 3759 28326
rect 5165 28323 5231 28326
rect 24853 28386 24919 28389
rect 25540 28386 26000 28416
rect 24853 28384 26000 28386
rect 24853 28328 24858 28384
rect 24914 28328 26000 28384
rect 24853 28326 26000 28328
rect 24853 28323 24919 28326
rect 6810 28320 7126 28321
rect 6810 28256 6816 28320
rect 6880 28256 6896 28320
rect 6960 28256 6976 28320
rect 7040 28256 7056 28320
rect 7120 28256 7126 28320
rect 6810 28255 7126 28256
rect 12675 28320 12991 28321
rect 12675 28256 12681 28320
rect 12745 28256 12761 28320
rect 12825 28256 12841 28320
rect 12905 28256 12921 28320
rect 12985 28256 12991 28320
rect 12675 28255 12991 28256
rect 18540 28320 18856 28321
rect 18540 28256 18546 28320
rect 18610 28256 18626 28320
rect 18690 28256 18706 28320
rect 18770 28256 18786 28320
rect 18850 28256 18856 28320
rect 18540 28255 18856 28256
rect 24405 28320 24721 28321
rect 24405 28256 24411 28320
rect 24475 28256 24491 28320
rect 24555 28256 24571 28320
rect 24635 28256 24651 28320
rect 24715 28256 24721 28320
rect 25540 28296 26000 28326
rect 24405 28255 24721 28256
rect 2681 28250 2747 28253
rect 6545 28250 6611 28253
rect 2681 28248 6611 28250
rect 2681 28192 2686 28248
rect 2742 28192 6550 28248
rect 6606 28192 6611 28248
rect 2681 28190 6611 28192
rect 2681 28187 2747 28190
rect 6545 28187 6611 28190
rect -300 28114 160 28144
rect 749 28114 815 28117
rect 12433 28114 12499 28117
rect -300 28112 815 28114
rect -300 28056 754 28112
rect 810 28056 815 28112
rect -300 28054 815 28056
rect -300 28024 160 28054
rect 749 28051 815 28054
rect 2454 28112 12499 28114
rect 2454 28056 12438 28112
rect 12494 28056 12499 28112
rect 2454 28054 12499 28056
rect 2313 27978 2379 27981
rect 2454 27978 2514 28054
rect 12433 28051 12499 28054
rect 15142 28052 15148 28116
rect 15212 28114 15218 28116
rect 16246 28114 16252 28116
rect 15212 28054 16252 28114
rect 15212 28052 15218 28054
rect 16246 28052 16252 28054
rect 16316 28114 16322 28116
rect 16481 28114 16547 28117
rect 16316 28112 16547 28114
rect 16316 28056 16486 28112
rect 16542 28056 16547 28112
rect 16316 28054 16547 28056
rect 16316 28052 16322 28054
rect 16481 28051 16547 28054
rect 11697 27978 11763 27981
rect 2313 27976 2514 27978
rect 2313 27920 2318 27976
rect 2374 27920 2514 27976
rect 2313 27918 2514 27920
rect 2592 27976 11763 27978
rect 2592 27920 11702 27976
rect 11758 27920 11763 27976
rect 2592 27918 11763 27920
rect 2313 27915 2379 27918
rect -300 27842 160 27872
rect 1301 27842 1367 27845
rect -300 27840 1367 27842
rect -300 27784 1306 27840
rect 1362 27784 1367 27840
rect -300 27782 1367 27784
rect -300 27752 160 27782
rect 1301 27779 1367 27782
rect 1761 27842 1827 27845
rect 2592 27842 2652 27918
rect 11697 27915 11763 27918
rect 12985 27978 13051 27981
rect 22686 27978 22692 27980
rect 12985 27976 22692 27978
rect 12985 27920 12990 27976
rect 13046 27920 22692 27976
rect 12985 27918 22692 27920
rect 12985 27915 13051 27918
rect 22686 27916 22692 27918
rect 22756 27916 22762 27980
rect 1761 27840 2652 27842
rect 1761 27784 1766 27840
rect 1822 27784 2652 27840
rect 1761 27782 2652 27784
rect 4521 27842 4587 27845
rect 6085 27842 6151 27845
rect 4521 27840 6151 27842
rect 4521 27784 4526 27840
rect 4582 27784 6090 27840
rect 6146 27784 6151 27840
rect 4521 27782 6151 27784
rect 1761 27779 1827 27782
rect 4521 27779 4587 27782
rect 6085 27779 6151 27782
rect 10133 27842 10199 27845
rect 24117 27842 24183 27845
rect 25540 27842 26000 27872
rect 10133 27840 10610 27842
rect 10133 27784 10138 27840
rect 10194 27784 10610 27840
rect 10133 27782 10610 27784
rect 10133 27779 10199 27782
rect 3878 27776 4194 27777
rect 3878 27712 3884 27776
rect 3948 27712 3964 27776
rect 4028 27712 4044 27776
rect 4108 27712 4124 27776
rect 4188 27712 4194 27776
rect 3878 27711 4194 27712
rect 9743 27776 10059 27777
rect 9743 27712 9749 27776
rect 9813 27712 9829 27776
rect 9893 27712 9909 27776
rect 9973 27712 9989 27776
rect 10053 27712 10059 27776
rect 9743 27711 10059 27712
rect 5758 27644 5764 27708
rect 5828 27706 5834 27708
rect 6126 27706 6132 27708
rect 5828 27646 6132 27706
rect 5828 27644 5834 27646
rect 6126 27644 6132 27646
rect 6196 27644 6202 27708
rect -300 27570 160 27600
rect 3693 27570 3759 27573
rect -300 27568 3759 27570
rect -300 27512 3698 27568
rect 3754 27512 3759 27568
rect -300 27510 3759 27512
rect -300 27480 160 27510
rect 3693 27507 3759 27510
rect 4061 27570 4127 27573
rect 4286 27570 4292 27572
rect 4061 27568 4292 27570
rect 4061 27512 4066 27568
rect 4122 27512 4292 27568
rect 4061 27510 4292 27512
rect 4061 27507 4127 27510
rect 4286 27508 4292 27510
rect 4356 27570 4362 27572
rect 7281 27570 7347 27573
rect 10550 27572 10610 27782
rect 24117 27840 26000 27842
rect 24117 27784 24122 27840
rect 24178 27784 26000 27840
rect 24117 27782 26000 27784
rect 24117 27779 24183 27782
rect 15608 27776 15924 27777
rect 15608 27712 15614 27776
rect 15678 27712 15694 27776
rect 15758 27712 15774 27776
rect 15838 27712 15854 27776
rect 15918 27712 15924 27776
rect 15608 27711 15924 27712
rect 21473 27776 21789 27777
rect 21473 27712 21479 27776
rect 21543 27712 21559 27776
rect 21623 27712 21639 27776
rect 21703 27712 21719 27776
rect 21783 27712 21789 27776
rect 25540 27752 26000 27782
rect 21473 27711 21789 27712
rect 10685 27706 10751 27709
rect 13077 27706 13143 27709
rect 10685 27704 13143 27706
rect 10685 27648 10690 27704
rect 10746 27648 13082 27704
rect 13138 27648 13143 27704
rect 10685 27646 13143 27648
rect 10685 27643 10751 27646
rect 13077 27643 13143 27646
rect 4356 27568 7347 27570
rect 4356 27512 7286 27568
rect 7342 27512 7347 27568
rect 4356 27510 7347 27512
rect 4356 27508 4362 27510
rect 7281 27507 7347 27510
rect 10542 27508 10548 27572
rect 10612 27508 10618 27572
rect 2865 27434 2931 27437
rect 3877 27434 3943 27437
rect 11697 27434 11763 27437
rect 2865 27432 3943 27434
rect 2865 27376 2870 27432
rect 2926 27376 3882 27432
rect 3938 27376 3943 27432
rect 2865 27374 3943 27376
rect 2865 27371 2931 27374
rect 3877 27371 3943 27374
rect 4662 27432 11763 27434
rect 4662 27376 11702 27432
rect 11758 27376 11763 27432
rect 4662 27374 11763 27376
rect -300 27298 160 27328
rect 841 27298 907 27301
rect 4662 27300 4722 27374
rect 11697 27371 11763 27374
rect 14089 27434 14155 27437
rect 14549 27434 14615 27437
rect 14089 27432 14615 27434
rect 14089 27376 14094 27432
rect 14150 27376 14554 27432
rect 14610 27376 14615 27432
rect 14089 27374 14615 27376
rect 14089 27371 14155 27374
rect 14549 27371 14615 27374
rect -300 27296 907 27298
rect -300 27240 846 27296
rect 902 27240 907 27296
rect -300 27238 907 27240
rect -300 27208 160 27238
rect 841 27235 907 27238
rect 4654 27236 4660 27300
rect 4724 27236 4730 27300
rect 7373 27298 7439 27301
rect 7598 27298 7604 27300
rect 7373 27296 7604 27298
rect 7373 27240 7378 27296
rect 7434 27240 7604 27296
rect 7373 27238 7604 27240
rect 7373 27235 7439 27238
rect 7598 27236 7604 27238
rect 7668 27236 7674 27300
rect 24853 27298 24919 27301
rect 25540 27298 26000 27328
rect 24853 27296 26000 27298
rect 24853 27240 24858 27296
rect 24914 27240 26000 27296
rect 24853 27238 26000 27240
rect 24853 27235 24919 27238
rect 6810 27232 7126 27233
rect 6810 27168 6816 27232
rect 6880 27168 6896 27232
rect 6960 27168 6976 27232
rect 7040 27168 7056 27232
rect 7120 27168 7126 27232
rect 6810 27167 7126 27168
rect 12675 27232 12991 27233
rect 12675 27168 12681 27232
rect 12745 27168 12761 27232
rect 12825 27168 12841 27232
rect 12905 27168 12921 27232
rect 12985 27168 12991 27232
rect 12675 27167 12991 27168
rect 18540 27232 18856 27233
rect 18540 27168 18546 27232
rect 18610 27168 18626 27232
rect 18690 27168 18706 27232
rect 18770 27168 18786 27232
rect 18850 27168 18856 27232
rect 18540 27167 18856 27168
rect 24405 27232 24721 27233
rect 24405 27168 24411 27232
rect 24475 27168 24491 27232
rect 24555 27168 24571 27232
rect 24635 27168 24651 27232
rect 24715 27168 24721 27232
rect 25540 27208 26000 27238
rect 24405 27167 24721 27168
rect 4470 27100 4476 27164
rect 4540 27162 4546 27164
rect 4981 27162 5047 27165
rect 4540 27160 5047 27162
rect 4540 27104 4986 27160
rect 5042 27104 5047 27160
rect 4540 27102 5047 27104
rect 4540 27100 4546 27102
rect 4981 27099 5047 27102
rect 7414 27100 7420 27164
rect 7484 27162 7490 27164
rect 8477 27162 8543 27165
rect 7484 27160 8543 27162
rect 7484 27104 8482 27160
rect 8538 27104 8543 27160
rect 7484 27102 8543 27104
rect 7484 27100 7490 27102
rect 8477 27099 8543 27102
rect -300 27026 160 27056
rect 1301 27026 1367 27029
rect -300 27024 1367 27026
rect -300 26968 1306 27024
rect 1362 26968 1367 27024
rect -300 26966 1367 26968
rect -300 26936 160 26966
rect 1301 26963 1367 26966
rect 3734 26964 3740 27028
rect 3804 27026 3810 27028
rect 4981 27026 5047 27029
rect 10174 27026 10180 27028
rect 3804 26966 4906 27026
rect 3804 26964 3810 26966
rect 2497 26890 2563 26893
rect 4654 26890 4660 26892
rect 2497 26888 4660 26890
rect 2497 26832 2502 26888
rect 2558 26832 4660 26888
rect 2497 26830 4660 26832
rect 2497 26827 2563 26830
rect 4654 26828 4660 26830
rect 4724 26828 4730 26892
rect 4846 26890 4906 26966
rect 4981 27024 10180 27026
rect 4981 26968 4986 27024
rect 5042 26968 10180 27024
rect 4981 26966 10180 26968
rect 4981 26963 5047 26966
rect 10174 26964 10180 26966
rect 10244 26964 10250 27028
rect 11053 27026 11119 27029
rect 15193 27026 15259 27029
rect 11053 27024 15259 27026
rect 11053 26968 11058 27024
rect 11114 26968 15198 27024
rect 15254 26968 15259 27024
rect 11053 26966 15259 26968
rect 11053 26963 11119 26966
rect 15193 26963 15259 26966
rect 6126 26890 6132 26892
rect 4846 26830 6132 26890
rect 6126 26828 6132 26830
rect 6196 26828 6202 26892
rect 6310 26828 6316 26892
rect 6380 26890 6386 26892
rect 10358 26890 10364 26892
rect 6380 26830 10364 26890
rect 6380 26828 6386 26830
rect 10358 26828 10364 26830
rect 10428 26828 10434 26892
rect 10726 26828 10732 26892
rect 10796 26890 10802 26892
rect 11973 26890 12039 26893
rect 10796 26888 12039 26890
rect 10796 26832 11978 26888
rect 12034 26832 12039 26888
rect 10796 26830 12039 26832
rect 10796 26828 10802 26830
rect 11973 26827 12039 26830
rect -300 26754 160 26784
rect 1209 26754 1275 26757
rect -300 26752 1275 26754
rect -300 26696 1214 26752
rect 1270 26696 1275 26752
rect -300 26694 1275 26696
rect -300 26664 160 26694
rect 1209 26691 1275 26694
rect 7465 26754 7531 26757
rect 8477 26754 8543 26757
rect 7465 26752 8543 26754
rect 7465 26696 7470 26752
rect 7526 26696 8482 26752
rect 8538 26696 8543 26752
rect 7465 26694 8543 26696
rect 7465 26691 7531 26694
rect 8477 26691 8543 26694
rect 24117 26754 24183 26757
rect 25540 26754 26000 26784
rect 24117 26752 26000 26754
rect 24117 26696 24122 26752
rect 24178 26696 26000 26752
rect 24117 26694 26000 26696
rect 24117 26691 24183 26694
rect 3878 26688 4194 26689
rect 3878 26624 3884 26688
rect 3948 26624 3964 26688
rect 4028 26624 4044 26688
rect 4108 26624 4124 26688
rect 4188 26624 4194 26688
rect 3878 26623 4194 26624
rect 9743 26688 10059 26689
rect 9743 26624 9749 26688
rect 9813 26624 9829 26688
rect 9893 26624 9909 26688
rect 9973 26624 9989 26688
rect 10053 26624 10059 26688
rect 9743 26623 10059 26624
rect 15608 26688 15924 26689
rect 15608 26624 15614 26688
rect 15678 26624 15694 26688
rect 15758 26624 15774 26688
rect 15838 26624 15854 26688
rect 15918 26624 15924 26688
rect 15608 26623 15924 26624
rect 21473 26688 21789 26689
rect 21473 26624 21479 26688
rect 21543 26624 21559 26688
rect 21623 26624 21639 26688
rect 21703 26624 21719 26688
rect 21783 26624 21789 26688
rect 25540 26664 26000 26694
rect 21473 26623 21789 26624
rect 4337 26618 4403 26621
rect 5758 26618 5764 26620
rect 4337 26616 5764 26618
rect 4337 26560 4342 26616
rect 4398 26560 5764 26616
rect 4337 26558 5764 26560
rect 4337 26555 4403 26558
rect 5758 26556 5764 26558
rect 5828 26556 5834 26620
rect 7373 26618 7439 26621
rect 8661 26618 8727 26621
rect 7373 26616 8727 26618
rect 7373 26560 7378 26616
rect 7434 26560 8666 26616
rect 8722 26560 8727 26616
rect 7373 26558 8727 26560
rect 7373 26555 7439 26558
rect 8661 26555 8727 26558
rect 10961 26618 11027 26621
rect 11278 26618 11284 26620
rect 10961 26616 11284 26618
rect 10961 26560 10966 26616
rect 11022 26560 11284 26616
rect 10961 26558 11284 26560
rect 10961 26555 11027 26558
rect 11278 26556 11284 26558
rect 11348 26556 11354 26620
rect 14038 26556 14044 26620
rect 14108 26618 14114 26620
rect 14181 26618 14247 26621
rect 14774 26618 14780 26620
rect 14108 26616 14780 26618
rect 14108 26560 14186 26616
rect 14242 26560 14780 26616
rect 14108 26558 14780 26560
rect 14108 26556 14114 26558
rect 14181 26555 14247 26558
rect 14774 26556 14780 26558
rect 14844 26556 14850 26620
rect -300 26482 160 26512
rect 1301 26482 1367 26485
rect -300 26480 1367 26482
rect -300 26424 1306 26480
rect 1362 26424 1367 26480
rect -300 26422 1367 26424
rect -300 26392 160 26422
rect 1301 26419 1367 26422
rect 2037 26482 2103 26485
rect 7465 26482 7531 26485
rect 2037 26480 7531 26482
rect 2037 26424 2042 26480
rect 2098 26424 7470 26480
rect 7526 26424 7531 26480
rect 2037 26422 7531 26424
rect 2037 26419 2103 26422
rect 7465 26419 7531 26422
rect 9305 26482 9371 26485
rect 11973 26482 12039 26485
rect 9305 26480 12039 26482
rect 9305 26424 9310 26480
rect 9366 26424 11978 26480
rect 12034 26424 12039 26480
rect 9305 26422 12039 26424
rect 9305 26419 9371 26422
rect 11973 26419 12039 26422
rect 4153 26346 4219 26349
rect 5809 26346 5875 26349
rect 4153 26344 5875 26346
rect 4153 26288 4158 26344
rect 4214 26288 5814 26344
rect 5870 26288 5875 26344
rect 4153 26286 5875 26288
rect 4153 26283 4219 26286
rect 5809 26283 5875 26286
rect 10174 26284 10180 26348
rect 10244 26346 10250 26348
rect 12249 26346 12315 26349
rect 10244 26344 12315 26346
rect 10244 26288 12254 26344
rect 12310 26288 12315 26344
rect 10244 26286 12315 26288
rect 10244 26284 10250 26286
rect 12249 26283 12315 26286
rect -300 26210 160 26240
rect 2865 26210 2931 26213
rect 5165 26212 5231 26213
rect 5165 26210 5212 26212
rect -300 26208 2931 26210
rect -300 26152 2870 26208
rect 2926 26152 2931 26208
rect -300 26150 2931 26152
rect -300 26120 160 26150
rect 2865 26147 2931 26150
rect 3006 26208 5212 26210
rect 3006 26152 5170 26208
rect 3006 26150 5212 26152
rect 2262 26012 2268 26076
rect 2332 26074 2338 26076
rect 2405 26074 2471 26077
rect 3006 26074 3066 26150
rect 5165 26148 5212 26150
rect 5276 26148 5282 26212
rect 7966 26148 7972 26212
rect 8036 26210 8042 26212
rect 9857 26210 9923 26213
rect 8036 26208 9923 26210
rect 8036 26152 9862 26208
rect 9918 26152 9923 26208
rect 8036 26150 9923 26152
rect 8036 26148 8042 26150
rect 5165 26147 5231 26148
rect 9857 26147 9923 26150
rect 24853 26210 24919 26213
rect 25540 26210 26000 26240
rect 24853 26208 26000 26210
rect 24853 26152 24858 26208
rect 24914 26152 26000 26208
rect 24853 26150 26000 26152
rect 24853 26147 24919 26150
rect 6810 26144 7126 26145
rect 6810 26080 6816 26144
rect 6880 26080 6896 26144
rect 6960 26080 6976 26144
rect 7040 26080 7056 26144
rect 7120 26080 7126 26144
rect 6810 26079 7126 26080
rect 12675 26144 12991 26145
rect 12675 26080 12681 26144
rect 12745 26080 12761 26144
rect 12825 26080 12841 26144
rect 12905 26080 12921 26144
rect 12985 26080 12991 26144
rect 12675 26079 12991 26080
rect 18540 26144 18856 26145
rect 18540 26080 18546 26144
rect 18610 26080 18626 26144
rect 18690 26080 18706 26144
rect 18770 26080 18786 26144
rect 18850 26080 18856 26144
rect 18540 26079 18856 26080
rect 24405 26144 24721 26145
rect 24405 26080 24411 26144
rect 24475 26080 24491 26144
rect 24555 26080 24571 26144
rect 24635 26080 24651 26144
rect 24715 26080 24721 26144
rect 25540 26120 26000 26150
rect 24405 26079 24721 26080
rect 2332 26072 3066 26074
rect 2332 26016 2410 26072
rect 2466 26016 3066 26072
rect 2332 26014 3066 26016
rect 2332 26012 2338 26014
rect 2405 26011 2471 26014
rect 5206 26012 5212 26076
rect 5276 26012 5282 26076
rect -300 25938 160 25968
rect 2773 25938 2839 25941
rect -300 25936 2839 25938
rect -300 25880 2778 25936
rect 2834 25880 2839 25936
rect -300 25878 2839 25880
rect 5214 25938 5274 26012
rect 7649 25938 7715 25941
rect 5214 25936 7715 25938
rect 5214 25880 7654 25936
rect 7710 25880 7715 25936
rect 5214 25878 7715 25880
rect -300 25848 160 25878
rect 2773 25875 2839 25878
rect 7649 25875 7715 25878
rect 10777 25938 10843 25941
rect 20110 25938 20116 25940
rect 10777 25936 20116 25938
rect 10777 25880 10782 25936
rect 10838 25880 20116 25936
rect 10777 25878 20116 25880
rect 10777 25875 10843 25878
rect 20110 25876 20116 25878
rect 20180 25876 20186 25940
rect 4429 25802 4495 25805
rect 16573 25802 16639 25805
rect 4429 25800 16639 25802
rect 4429 25744 4434 25800
rect 4490 25744 16578 25800
rect 16634 25744 16639 25800
rect 4429 25742 16639 25744
rect 4429 25739 4495 25742
rect 16573 25739 16639 25742
rect -300 25666 160 25696
rect 1301 25666 1367 25669
rect -300 25664 1367 25666
rect -300 25608 1306 25664
rect 1362 25608 1367 25664
rect -300 25606 1367 25608
rect -300 25576 160 25606
rect 1301 25603 1367 25606
rect 2814 25604 2820 25668
rect 2884 25666 2890 25668
rect 3693 25666 3759 25669
rect 2884 25664 3759 25666
rect 2884 25608 3698 25664
rect 3754 25608 3759 25664
rect 2884 25606 3759 25608
rect 2884 25604 2890 25606
rect 3693 25603 3759 25606
rect 5942 25604 5948 25668
rect 6012 25666 6018 25668
rect 6545 25666 6611 25669
rect 6012 25664 6611 25666
rect 6012 25608 6550 25664
rect 6606 25608 6611 25664
rect 6012 25606 6611 25608
rect 6012 25604 6018 25606
rect 6545 25603 6611 25606
rect 23749 25666 23815 25669
rect 25540 25666 26000 25696
rect 23749 25664 26000 25666
rect 23749 25608 23754 25664
rect 23810 25608 26000 25664
rect 23749 25606 26000 25608
rect 23749 25603 23815 25606
rect 3878 25600 4194 25601
rect 3878 25536 3884 25600
rect 3948 25536 3964 25600
rect 4028 25536 4044 25600
rect 4108 25536 4124 25600
rect 4188 25536 4194 25600
rect 3878 25535 4194 25536
rect 9743 25600 10059 25601
rect 9743 25536 9749 25600
rect 9813 25536 9829 25600
rect 9893 25536 9909 25600
rect 9973 25536 9989 25600
rect 10053 25536 10059 25600
rect 9743 25535 10059 25536
rect 15608 25600 15924 25601
rect 15608 25536 15614 25600
rect 15678 25536 15694 25600
rect 15758 25536 15774 25600
rect 15838 25536 15854 25600
rect 15918 25536 15924 25600
rect 15608 25535 15924 25536
rect 21473 25600 21789 25601
rect 21473 25536 21479 25600
rect 21543 25536 21559 25600
rect 21623 25536 21639 25600
rect 21703 25536 21719 25600
rect 21783 25536 21789 25600
rect 25540 25576 26000 25606
rect 21473 25535 21789 25536
rect -300 25394 160 25424
rect 841 25394 907 25397
rect -300 25392 907 25394
rect -300 25336 846 25392
rect 902 25336 907 25392
rect -300 25334 907 25336
rect -300 25304 160 25334
rect 841 25331 907 25334
rect 5390 25332 5396 25396
rect 5460 25394 5466 25396
rect 10225 25394 10291 25397
rect 5460 25392 10291 25394
rect 5460 25336 10230 25392
rect 10286 25336 10291 25392
rect 5460 25334 10291 25336
rect 5460 25332 5466 25334
rect 10225 25331 10291 25334
rect 12065 25394 12131 25397
rect 12525 25394 12591 25397
rect 12065 25392 12591 25394
rect 12065 25336 12070 25392
rect 12126 25336 12530 25392
rect 12586 25336 12591 25392
rect 12065 25334 12591 25336
rect 12065 25331 12131 25334
rect 12525 25331 12591 25334
rect 1669 25258 1735 25261
rect 798 25256 1735 25258
rect 798 25200 1674 25256
rect 1730 25200 1735 25256
rect 798 25198 1735 25200
rect -300 25122 160 25152
rect 798 25122 858 25198
rect 1669 25195 1735 25198
rect 2865 25258 2931 25261
rect 13997 25258 14063 25261
rect 2865 25256 14063 25258
rect 2865 25200 2870 25256
rect 2926 25200 14002 25256
rect 14058 25200 14063 25256
rect 2865 25198 14063 25200
rect 2865 25195 2931 25198
rect 13997 25195 14063 25198
rect 6545 25122 6611 25125
rect -300 25062 858 25122
rect 5950 25120 6611 25122
rect 5950 25064 6550 25120
rect 6606 25064 6611 25120
rect 5950 25062 6611 25064
rect -300 25032 160 25062
rect 2630 24924 2636 24988
rect 2700 24986 2706 24988
rect 4245 24986 4311 24989
rect 2700 24984 4311 24986
rect 2700 24928 4250 24984
rect 4306 24928 4311 24984
rect 2700 24926 4311 24928
rect 2700 24924 2706 24926
rect 4245 24923 4311 24926
rect 5625 24986 5691 24989
rect 5758 24986 5764 24988
rect 5625 24984 5764 24986
rect 5625 24928 5630 24984
rect 5686 24928 5764 24984
rect 5625 24926 5764 24928
rect 5625 24923 5691 24926
rect 5758 24924 5764 24926
rect 5828 24924 5834 24988
rect -300 24850 160 24880
rect 1301 24850 1367 24853
rect -300 24848 1367 24850
rect -300 24792 1306 24848
rect 1362 24792 1367 24848
rect -300 24790 1367 24792
rect -300 24760 160 24790
rect 1301 24787 1367 24790
rect 1669 24850 1735 24853
rect 5950 24850 6010 25062
rect 6545 25059 6611 25062
rect 24853 25122 24919 25125
rect 25540 25122 26000 25152
rect 24853 25120 26000 25122
rect 24853 25064 24858 25120
rect 24914 25064 26000 25120
rect 24853 25062 26000 25064
rect 24853 25059 24919 25062
rect 6810 25056 7126 25057
rect 6810 24992 6816 25056
rect 6880 24992 6896 25056
rect 6960 24992 6976 25056
rect 7040 24992 7056 25056
rect 7120 24992 7126 25056
rect 6810 24991 7126 24992
rect 12675 25056 12991 25057
rect 12675 24992 12681 25056
rect 12745 24992 12761 25056
rect 12825 24992 12841 25056
rect 12905 24992 12921 25056
rect 12985 24992 12991 25056
rect 12675 24991 12991 24992
rect 18540 25056 18856 25057
rect 18540 24992 18546 25056
rect 18610 24992 18626 25056
rect 18690 24992 18706 25056
rect 18770 24992 18786 25056
rect 18850 24992 18856 25056
rect 18540 24991 18856 24992
rect 24405 25056 24721 25057
rect 24405 24992 24411 25056
rect 24475 24992 24491 25056
rect 24555 24992 24571 25056
rect 24635 24992 24651 25056
rect 24715 24992 24721 25056
rect 25540 25032 26000 25062
rect 24405 24991 24721 24992
rect 1669 24848 6010 24850
rect 1669 24792 1674 24848
rect 1730 24792 6010 24848
rect 1669 24790 6010 24792
rect 6085 24850 6151 24853
rect 8753 24850 8819 24853
rect 6085 24848 8819 24850
rect 6085 24792 6090 24848
rect 6146 24792 8758 24848
rect 8814 24792 8819 24848
rect 6085 24790 8819 24792
rect 1669 24787 1735 24790
rect 6085 24787 6151 24790
rect 8753 24787 8819 24790
rect 10593 24850 10659 24853
rect 11329 24850 11395 24853
rect 10593 24848 11395 24850
rect 10593 24792 10598 24848
rect 10654 24792 11334 24848
rect 11390 24792 11395 24848
rect 10593 24790 11395 24792
rect 10593 24787 10659 24790
rect 11329 24787 11395 24790
rect 1577 24714 1643 24717
rect 3417 24714 3483 24717
rect 4797 24714 4863 24717
rect 1577 24712 3483 24714
rect 1577 24656 1582 24712
rect 1638 24656 3422 24712
rect 3478 24656 3483 24712
rect 1577 24654 3483 24656
rect 1577 24651 1643 24654
rect 3417 24651 3483 24654
rect 3742 24712 4863 24714
rect 3742 24656 4802 24712
rect 4858 24656 4863 24712
rect 3742 24654 4863 24656
rect -300 24578 160 24608
rect 1209 24578 1275 24581
rect -300 24576 1275 24578
rect -300 24520 1214 24576
rect 1270 24520 1275 24576
rect -300 24518 1275 24520
rect -300 24488 160 24518
rect 1209 24515 1275 24518
rect 2814 24516 2820 24580
rect 2884 24578 2890 24580
rect 3742 24578 3802 24654
rect 4797 24651 4863 24654
rect 7833 24714 7899 24717
rect 21081 24714 21147 24717
rect 7833 24712 21147 24714
rect 7833 24656 7838 24712
rect 7894 24656 21086 24712
rect 21142 24656 21147 24712
rect 7833 24654 21147 24656
rect 7833 24651 7899 24654
rect 21081 24651 21147 24654
rect 2884 24518 3802 24578
rect 10225 24578 10291 24581
rect 14549 24578 14615 24581
rect 10225 24576 14615 24578
rect 10225 24520 10230 24576
rect 10286 24520 14554 24576
rect 14610 24520 14615 24576
rect 10225 24518 14615 24520
rect 2884 24516 2890 24518
rect 10225 24515 10291 24518
rect 14549 24515 14615 24518
rect 23841 24578 23907 24581
rect 25540 24578 26000 24608
rect 23841 24576 26000 24578
rect 23841 24520 23846 24576
rect 23902 24520 26000 24576
rect 23841 24518 26000 24520
rect 23841 24515 23907 24518
rect 3878 24512 4194 24513
rect 3878 24448 3884 24512
rect 3948 24448 3964 24512
rect 4028 24448 4044 24512
rect 4108 24448 4124 24512
rect 4188 24448 4194 24512
rect 3878 24447 4194 24448
rect 9743 24512 10059 24513
rect 9743 24448 9749 24512
rect 9813 24448 9829 24512
rect 9893 24448 9909 24512
rect 9973 24448 9989 24512
rect 10053 24448 10059 24512
rect 9743 24447 10059 24448
rect 15608 24512 15924 24513
rect 15608 24448 15614 24512
rect 15678 24448 15694 24512
rect 15758 24448 15774 24512
rect 15838 24448 15854 24512
rect 15918 24448 15924 24512
rect 15608 24447 15924 24448
rect 21473 24512 21789 24513
rect 21473 24448 21479 24512
rect 21543 24448 21559 24512
rect 21623 24448 21639 24512
rect 21703 24448 21719 24512
rect 21783 24448 21789 24512
rect 25540 24488 26000 24518
rect 21473 24447 21789 24448
rect 10409 24442 10475 24445
rect 10409 24440 10794 24442
rect 10409 24384 10414 24440
rect 10470 24384 10794 24440
rect 10409 24382 10794 24384
rect 10409 24379 10475 24382
rect -300 24306 160 24336
rect 10734 24309 10794 24382
rect 749 24306 815 24309
rect -300 24304 815 24306
rect -300 24248 754 24304
rect 810 24248 815 24304
rect -300 24246 815 24248
rect -300 24216 160 24246
rect 749 24243 815 24246
rect 3417 24306 3483 24309
rect 6453 24306 6519 24309
rect 3417 24304 6519 24306
rect 3417 24248 3422 24304
rect 3478 24248 6458 24304
rect 6514 24248 6519 24304
rect 3417 24246 6519 24248
rect 10734 24304 10843 24309
rect 10734 24248 10782 24304
rect 10838 24248 10843 24304
rect 10734 24246 10843 24248
rect 3417 24243 3483 24246
rect 6453 24243 6519 24246
rect 10777 24243 10843 24246
rect 4153 24170 4219 24173
rect 5022 24170 5028 24172
rect 4153 24168 5028 24170
rect 4153 24112 4158 24168
rect 4214 24112 5028 24168
rect 4153 24110 5028 24112
rect 4153 24107 4219 24110
rect 5022 24108 5028 24110
rect 5092 24108 5098 24172
rect 21950 24108 21956 24172
rect 22020 24170 22026 24172
rect 22553 24170 22619 24173
rect 22020 24168 22619 24170
rect 22020 24112 22558 24168
rect 22614 24112 22619 24168
rect 22020 24110 22619 24112
rect 22020 24108 22026 24110
rect 22553 24107 22619 24110
rect -300 24034 160 24064
rect 1301 24034 1367 24037
rect -300 24032 1367 24034
rect -300 23976 1306 24032
rect 1362 23976 1367 24032
rect -300 23974 1367 23976
rect -300 23944 160 23974
rect 1301 23971 1367 23974
rect 7649 24034 7715 24037
rect 8753 24034 8819 24037
rect 7649 24032 8819 24034
rect 7649 23976 7654 24032
rect 7710 23976 8758 24032
rect 8814 23976 8819 24032
rect 7649 23974 8819 23976
rect 7649 23971 7715 23974
rect 8753 23971 8819 23974
rect 24853 24034 24919 24037
rect 25540 24034 26000 24064
rect 24853 24032 26000 24034
rect 24853 23976 24858 24032
rect 24914 23976 26000 24032
rect 24853 23974 26000 23976
rect 24853 23971 24919 23974
rect 6810 23968 7126 23969
rect 6810 23904 6816 23968
rect 6880 23904 6896 23968
rect 6960 23904 6976 23968
rect 7040 23904 7056 23968
rect 7120 23904 7126 23968
rect 6810 23903 7126 23904
rect 12675 23968 12991 23969
rect 12675 23904 12681 23968
rect 12745 23904 12761 23968
rect 12825 23904 12841 23968
rect 12905 23904 12921 23968
rect 12985 23904 12991 23968
rect 12675 23903 12991 23904
rect 18540 23968 18856 23969
rect 18540 23904 18546 23968
rect 18610 23904 18626 23968
rect 18690 23904 18706 23968
rect 18770 23904 18786 23968
rect 18850 23904 18856 23968
rect 18540 23903 18856 23904
rect 24405 23968 24721 23969
rect 24405 23904 24411 23968
rect 24475 23904 24491 23968
rect 24555 23904 24571 23968
rect 24635 23904 24651 23968
rect 24715 23904 24721 23968
rect 25540 23944 26000 23974
rect 24405 23903 24721 23904
rect 9673 23898 9739 23901
rect 10593 23898 10659 23901
rect 9673 23896 10659 23898
rect 9673 23840 9678 23896
rect 9734 23840 10598 23896
rect 10654 23840 10659 23896
rect 9673 23838 10659 23840
rect 9673 23835 9739 23838
rect 10593 23835 10659 23838
rect -300 23762 160 23792
rect 841 23762 907 23765
rect -300 23760 907 23762
rect -300 23704 846 23760
rect 902 23704 907 23760
rect -300 23702 907 23704
rect -300 23672 160 23702
rect 841 23699 907 23702
rect 2497 23762 2563 23765
rect 8201 23762 8267 23765
rect 2497 23760 8267 23762
rect 2497 23704 2502 23760
rect 2558 23704 8206 23760
rect 8262 23704 8267 23760
rect 2497 23702 8267 23704
rect 2497 23699 2563 23702
rect 8201 23699 8267 23702
rect 8385 23762 8451 23765
rect 11881 23762 11947 23765
rect 8385 23760 11947 23762
rect 8385 23704 8390 23760
rect 8446 23704 11886 23760
rect 11942 23704 11947 23760
rect 8385 23702 11947 23704
rect 8385 23699 8451 23702
rect 11881 23699 11947 23702
rect 2773 23626 2839 23629
rect 9581 23626 9647 23629
rect 2773 23624 9647 23626
rect 2773 23568 2778 23624
rect 2834 23568 9586 23624
rect 9642 23568 9647 23624
rect 2773 23566 9647 23568
rect 2773 23563 2839 23566
rect 9581 23563 9647 23566
rect 10041 23626 10107 23629
rect 10501 23626 10567 23629
rect 10041 23624 10567 23626
rect 10041 23568 10046 23624
rect 10102 23568 10506 23624
rect 10562 23568 10567 23624
rect 10041 23566 10567 23568
rect 10041 23563 10107 23566
rect 10501 23563 10567 23566
rect 11278 23564 11284 23628
rect 11348 23626 11354 23628
rect 18413 23626 18479 23629
rect 11348 23624 18479 23626
rect 11348 23568 18418 23624
rect 18474 23568 18479 23624
rect 11348 23566 18479 23568
rect 11348 23564 11354 23566
rect 18413 23563 18479 23566
rect -300 23490 160 23520
rect 749 23490 815 23493
rect 1669 23490 1735 23493
rect 2497 23492 2563 23493
rect -300 23488 815 23490
rect -300 23432 754 23488
rect 810 23432 815 23488
rect -300 23430 815 23432
rect -300 23400 160 23430
rect 749 23427 815 23430
rect 936 23488 1735 23490
rect 936 23432 1674 23488
rect 1730 23432 1735 23488
rect 936 23430 1735 23432
rect -300 23218 160 23248
rect 936 23218 996 23430
rect 1669 23427 1735 23430
rect 2446 23428 2452 23492
rect 2516 23490 2563 23492
rect 4705 23490 4771 23493
rect 5022 23490 5028 23492
rect 2516 23488 2608 23490
rect 2558 23432 2608 23488
rect 2516 23430 2608 23432
rect 4705 23488 5028 23490
rect 4705 23432 4710 23488
rect 4766 23432 5028 23488
rect 4705 23430 5028 23432
rect 2516 23428 2563 23430
rect 2497 23427 2563 23428
rect 4705 23427 4771 23430
rect 5022 23428 5028 23430
rect 5092 23428 5098 23492
rect 13261 23490 13327 23493
rect 14222 23490 14228 23492
rect 13261 23488 14228 23490
rect 13261 23432 13266 23488
rect 13322 23432 14228 23488
rect 13261 23430 14228 23432
rect 13261 23427 13327 23430
rect 14222 23428 14228 23430
rect 14292 23428 14298 23492
rect 24117 23490 24183 23493
rect 25540 23490 26000 23520
rect 24117 23488 26000 23490
rect 24117 23432 24122 23488
rect 24178 23432 26000 23488
rect 24117 23430 26000 23432
rect 24117 23427 24183 23430
rect 3878 23424 4194 23425
rect 3878 23360 3884 23424
rect 3948 23360 3964 23424
rect 4028 23360 4044 23424
rect 4108 23360 4124 23424
rect 4188 23360 4194 23424
rect 3878 23359 4194 23360
rect 9743 23424 10059 23425
rect 9743 23360 9749 23424
rect 9813 23360 9829 23424
rect 9893 23360 9909 23424
rect 9973 23360 9989 23424
rect 10053 23360 10059 23424
rect 9743 23359 10059 23360
rect 15608 23424 15924 23425
rect 15608 23360 15614 23424
rect 15678 23360 15694 23424
rect 15758 23360 15774 23424
rect 15838 23360 15854 23424
rect 15918 23360 15924 23424
rect 15608 23359 15924 23360
rect 21473 23424 21789 23425
rect 21473 23360 21479 23424
rect 21543 23360 21559 23424
rect 21623 23360 21639 23424
rect 21703 23360 21719 23424
rect 21783 23360 21789 23424
rect 25540 23400 26000 23430
rect 21473 23359 21789 23360
rect 2681 23354 2747 23357
rect 3550 23354 3556 23356
rect 2681 23352 3556 23354
rect 2681 23296 2686 23352
rect 2742 23296 3556 23352
rect 2681 23294 3556 23296
rect 2681 23291 2747 23294
rect 3550 23292 3556 23294
rect 3620 23292 3626 23356
rect -300 23158 996 23218
rect -300 23128 160 23158
rect 2037 23082 2103 23085
rect 2865 23082 2931 23085
rect 2037 23080 2931 23082
rect 2037 23024 2042 23080
rect 2098 23024 2870 23080
rect 2926 23024 2931 23080
rect 2037 23022 2931 23024
rect 2037 23019 2103 23022
rect 2865 23019 2931 23022
rect 7649 23082 7715 23085
rect 10910 23082 10916 23084
rect 7649 23080 10916 23082
rect 7649 23024 7654 23080
rect 7710 23024 10916 23080
rect 7649 23022 10916 23024
rect 7649 23019 7715 23022
rect 10910 23020 10916 23022
rect 10980 23020 10986 23084
rect -300 22946 160 22976
rect 749 22946 815 22949
rect -300 22944 815 22946
rect -300 22888 754 22944
rect 810 22888 815 22944
rect -300 22886 815 22888
rect -300 22856 160 22886
rect 749 22883 815 22886
rect 24853 22946 24919 22949
rect 25540 22946 26000 22976
rect 24853 22944 26000 22946
rect 24853 22888 24858 22944
rect 24914 22888 26000 22944
rect 24853 22886 26000 22888
rect 24853 22883 24919 22886
rect 6810 22880 7126 22881
rect 6810 22816 6816 22880
rect 6880 22816 6896 22880
rect 6960 22816 6976 22880
rect 7040 22816 7056 22880
rect 7120 22816 7126 22880
rect 6810 22815 7126 22816
rect 12675 22880 12991 22881
rect 12675 22816 12681 22880
rect 12745 22816 12761 22880
rect 12825 22816 12841 22880
rect 12905 22816 12921 22880
rect 12985 22816 12991 22880
rect 12675 22815 12991 22816
rect 18540 22880 18856 22881
rect 18540 22816 18546 22880
rect 18610 22816 18626 22880
rect 18690 22816 18706 22880
rect 18770 22816 18786 22880
rect 18850 22816 18856 22880
rect 18540 22815 18856 22816
rect 24405 22880 24721 22881
rect 24405 22816 24411 22880
rect 24475 22816 24491 22880
rect 24555 22816 24571 22880
rect 24635 22816 24651 22880
rect 24715 22816 24721 22880
rect 25540 22856 26000 22886
rect 24405 22815 24721 22816
rect -300 22674 160 22704
rect 841 22674 907 22677
rect -300 22672 907 22674
rect -300 22616 846 22672
rect 902 22616 907 22672
rect -300 22614 907 22616
rect -300 22584 160 22614
rect 841 22611 907 22614
rect 6269 22674 6335 22677
rect 7741 22674 7807 22677
rect 6269 22672 7807 22674
rect 6269 22616 6274 22672
rect 6330 22616 7746 22672
rect 7802 22616 7807 22672
rect 6269 22614 7807 22616
rect 6269 22611 6335 22614
rect 7741 22611 7807 22614
rect 10593 22674 10659 22677
rect 13445 22674 13511 22677
rect 14457 22676 14523 22677
rect 14406 22674 14412 22676
rect 10593 22672 13511 22674
rect 10593 22616 10598 22672
rect 10654 22616 13450 22672
rect 13506 22616 13511 22672
rect 10593 22614 13511 22616
rect 14366 22614 14412 22674
rect 14476 22672 14523 22676
rect 14518 22616 14523 22672
rect 10593 22611 10659 22614
rect 13445 22611 13511 22614
rect 14406 22612 14412 22614
rect 14476 22612 14523 22616
rect 14457 22611 14523 22612
rect -300 22402 160 22432
rect 1301 22402 1367 22405
rect -300 22400 1367 22402
rect -300 22344 1306 22400
rect 1362 22344 1367 22400
rect -300 22342 1367 22344
rect -300 22312 160 22342
rect 1301 22339 1367 22342
rect 23749 22402 23815 22405
rect 25540 22402 26000 22432
rect 23749 22400 26000 22402
rect 23749 22344 23754 22400
rect 23810 22344 26000 22400
rect 23749 22342 26000 22344
rect 23749 22339 23815 22342
rect 3878 22336 4194 22337
rect 3878 22272 3884 22336
rect 3948 22272 3964 22336
rect 4028 22272 4044 22336
rect 4108 22272 4124 22336
rect 4188 22272 4194 22336
rect 3878 22271 4194 22272
rect 9743 22336 10059 22337
rect 9743 22272 9749 22336
rect 9813 22272 9829 22336
rect 9893 22272 9909 22336
rect 9973 22272 9989 22336
rect 10053 22272 10059 22336
rect 9743 22271 10059 22272
rect 15608 22336 15924 22337
rect 15608 22272 15614 22336
rect 15678 22272 15694 22336
rect 15758 22272 15774 22336
rect 15838 22272 15854 22336
rect 15918 22272 15924 22336
rect 15608 22271 15924 22272
rect 21473 22336 21789 22337
rect 21473 22272 21479 22336
rect 21543 22272 21559 22336
rect 21623 22272 21639 22336
rect 21703 22272 21719 22336
rect 21783 22272 21789 22336
rect 25540 22312 26000 22342
rect 21473 22271 21789 22272
rect 10542 22204 10548 22268
rect 10612 22266 10618 22268
rect 13302 22266 13308 22268
rect 10612 22206 13308 22266
rect 10612 22204 10618 22206
rect 13302 22204 13308 22206
rect 13372 22204 13378 22268
rect -300 22130 160 22160
rect 1945 22130 2011 22133
rect 2405 22130 2471 22133
rect -300 22128 2011 22130
rect -300 22072 1950 22128
rect 2006 22072 2011 22128
rect -300 22070 2011 22072
rect -300 22040 160 22070
rect 1945 22067 2011 22070
rect 2086 22128 2471 22130
rect 2086 22072 2410 22128
rect 2466 22072 2471 22128
rect 2086 22070 2471 22072
rect 2086 21994 2146 22070
rect 2405 22067 2471 22070
rect 2589 22130 2655 22133
rect 4429 22130 4495 22133
rect 6269 22130 6335 22133
rect 2589 22128 6335 22130
rect 2589 22072 2594 22128
rect 2650 22072 4434 22128
rect 4490 22072 6274 22128
rect 6330 22072 6335 22128
rect 2589 22070 6335 22072
rect 2589 22067 2655 22070
rect 4429 22067 4495 22070
rect 6269 22067 6335 22070
rect 12382 22068 12388 22132
rect 12452 22130 12458 22132
rect 13118 22130 13124 22132
rect 12452 22070 13124 22130
rect 12452 22068 12458 22070
rect 13118 22068 13124 22070
rect 13188 22068 13194 22132
rect 13261 22130 13327 22133
rect 13486 22130 13492 22132
rect 13261 22128 13492 22130
rect 13261 22072 13266 22128
rect 13322 22072 13492 22128
rect 13261 22070 13492 22072
rect 13261 22067 13327 22070
rect 13486 22068 13492 22070
rect 13556 22068 13562 22132
rect 4429 21996 4495 21997
rect 4429 21994 4476 21996
rect 1902 21934 2146 21994
rect 4384 21992 4476 21994
rect 4540 21994 4546 21996
rect 11697 21994 11763 21997
rect 4540 21992 11763 21994
rect 4384 21936 4434 21992
rect 4540 21936 11702 21992
rect 11758 21936 11763 21992
rect 4384 21934 4476 21936
rect -300 21858 160 21888
rect 933 21858 999 21861
rect 1902 21860 1962 21934
rect 4429 21932 4476 21934
rect 4540 21934 11763 21936
rect 4540 21932 4546 21934
rect 4429 21931 4495 21932
rect 11697 21931 11763 21934
rect 12382 21932 12388 21996
rect 12452 21994 12458 21996
rect 13118 21994 13124 21996
rect 12452 21934 13124 21994
rect 12452 21932 12458 21934
rect 13118 21932 13124 21934
rect 13188 21932 13194 21996
rect 21214 21932 21220 21996
rect 21284 21994 21290 21996
rect 21357 21994 21423 21997
rect 21284 21992 21423 21994
rect 21284 21936 21362 21992
rect 21418 21936 21423 21992
rect 21284 21934 21423 21936
rect 21284 21932 21290 21934
rect 21357 21931 21423 21934
rect -300 21856 999 21858
rect -300 21800 938 21856
rect 994 21800 999 21856
rect -300 21798 999 21800
rect -300 21768 160 21798
rect 933 21795 999 21798
rect 1894 21796 1900 21860
rect 1964 21796 1970 21860
rect 7598 21796 7604 21860
rect 7668 21858 7674 21860
rect 7741 21858 7807 21861
rect 12157 21858 12223 21861
rect 7668 21856 7807 21858
rect 7668 21800 7746 21856
rect 7802 21800 7807 21856
rect 7668 21798 7807 21800
rect 7668 21796 7674 21798
rect 7741 21795 7807 21798
rect 11838 21856 12223 21858
rect 11838 21800 12162 21856
rect 12218 21800 12223 21856
rect 11838 21798 12223 21800
rect 6810 21792 7126 21793
rect 6810 21728 6816 21792
rect 6880 21728 6896 21792
rect 6960 21728 6976 21792
rect 7040 21728 7056 21792
rect 7120 21728 7126 21792
rect 6810 21727 7126 21728
rect 11838 21725 11898 21798
rect 12157 21795 12223 21798
rect 24853 21858 24919 21861
rect 25540 21858 26000 21888
rect 24853 21856 26000 21858
rect 24853 21800 24858 21856
rect 24914 21800 26000 21856
rect 24853 21798 26000 21800
rect 24853 21795 24919 21798
rect 12675 21792 12991 21793
rect 12675 21728 12681 21792
rect 12745 21728 12761 21792
rect 12825 21728 12841 21792
rect 12905 21728 12921 21792
rect 12985 21728 12991 21792
rect 12675 21727 12991 21728
rect 18540 21792 18856 21793
rect 18540 21728 18546 21792
rect 18610 21728 18626 21792
rect 18690 21728 18706 21792
rect 18770 21728 18786 21792
rect 18850 21728 18856 21792
rect 18540 21727 18856 21728
rect 24405 21792 24721 21793
rect 24405 21728 24411 21792
rect 24475 21728 24491 21792
rect 24555 21728 24571 21792
rect 24635 21728 24651 21792
rect 24715 21728 24721 21792
rect 25540 21768 26000 21798
rect 24405 21727 24721 21728
rect 11789 21720 11898 21725
rect 11789 21664 11794 21720
rect 11850 21664 11898 21720
rect 11789 21662 11898 21664
rect 11789 21659 11855 21662
rect -300 21586 160 21616
rect 749 21586 815 21589
rect -300 21584 815 21586
rect -300 21528 754 21584
rect 810 21528 815 21584
rect -300 21526 815 21528
rect -300 21496 160 21526
rect 749 21523 815 21526
rect 3969 21586 4035 21589
rect 4337 21586 4403 21589
rect 3969 21584 4403 21586
rect 3969 21528 3974 21584
rect 4030 21528 4342 21584
rect 4398 21528 4403 21584
rect 3969 21526 4403 21528
rect 3969 21523 4035 21526
rect 4337 21523 4403 21526
rect 5441 21586 5507 21589
rect 5901 21586 5967 21589
rect 5441 21584 5967 21586
rect 5441 21528 5446 21584
rect 5502 21528 5906 21584
rect 5962 21528 5967 21584
rect 5441 21526 5967 21528
rect 5441 21523 5507 21526
rect 5901 21523 5967 21526
rect 6269 21586 6335 21589
rect 8518 21586 8524 21588
rect 6269 21584 8524 21586
rect 6269 21528 6274 21584
rect 6330 21528 8524 21584
rect 6269 21526 8524 21528
rect 6269 21523 6335 21526
rect 8518 21524 8524 21526
rect 8588 21524 8594 21588
rect 10409 21586 10475 21589
rect 14181 21586 14247 21589
rect 10409 21584 14247 21586
rect 10409 21528 10414 21584
rect 10470 21528 14186 21584
rect 14242 21528 14247 21584
rect 10409 21526 14247 21528
rect 10409 21523 10475 21526
rect 14181 21523 14247 21526
rect 4153 21450 4219 21453
rect 10961 21450 11027 21453
rect 14549 21450 14615 21453
rect 4153 21448 4354 21450
rect 4153 21392 4158 21448
rect 4214 21392 4354 21448
rect 4153 21390 4354 21392
rect 4153 21387 4219 21390
rect -300 21314 160 21344
rect 1117 21314 1183 21317
rect -300 21312 1183 21314
rect -300 21256 1122 21312
rect 1178 21256 1183 21312
rect -300 21254 1183 21256
rect -300 21224 160 21254
rect 1117 21251 1183 21254
rect 3878 21248 4194 21249
rect 3878 21184 3884 21248
rect 3948 21184 3964 21248
rect 4028 21184 4044 21248
rect 4108 21184 4124 21248
rect 4188 21184 4194 21248
rect 3878 21183 4194 21184
rect -300 21042 160 21072
rect 4294 21045 4354 21390
rect 10961 21448 14615 21450
rect 10961 21392 10966 21448
rect 11022 21392 14554 21448
rect 14610 21392 14615 21448
rect 10961 21390 14615 21392
rect 10961 21387 11027 21390
rect 14549 21387 14615 21390
rect 24117 21314 24183 21317
rect 25540 21314 26000 21344
rect 24117 21312 26000 21314
rect 24117 21256 24122 21312
rect 24178 21256 26000 21312
rect 24117 21254 26000 21256
rect 24117 21251 24183 21254
rect 9743 21248 10059 21249
rect 9743 21184 9749 21248
rect 9813 21184 9829 21248
rect 9893 21184 9909 21248
rect 9973 21184 9989 21248
rect 10053 21184 10059 21248
rect 9743 21183 10059 21184
rect 15608 21248 15924 21249
rect 15608 21184 15614 21248
rect 15678 21184 15694 21248
rect 15758 21184 15774 21248
rect 15838 21184 15854 21248
rect 15918 21184 15924 21248
rect 15608 21183 15924 21184
rect 21473 21248 21789 21249
rect 21473 21184 21479 21248
rect 21543 21184 21559 21248
rect 21623 21184 21639 21248
rect 21703 21184 21719 21248
rect 21783 21184 21789 21248
rect 25540 21224 26000 21254
rect 21473 21183 21789 21184
rect 1301 21042 1367 21045
rect -300 21040 1367 21042
rect -300 20984 1306 21040
rect 1362 20984 1367 21040
rect -300 20982 1367 20984
rect -300 20952 160 20982
rect 1301 20979 1367 20982
rect 4245 21040 4354 21045
rect 4245 20984 4250 21040
rect 4306 20984 4354 21040
rect 4245 20982 4354 20984
rect 8569 21042 8635 21045
rect 8702 21042 8708 21044
rect 8569 21040 8708 21042
rect 8569 20984 8574 21040
rect 8630 20984 8708 21040
rect 8569 20982 8708 20984
rect 4245 20979 4311 20982
rect 8569 20979 8635 20982
rect 8702 20980 8708 20982
rect 8772 20980 8778 21044
rect 9857 21042 9923 21045
rect 11237 21044 11303 21045
rect 11237 21042 11284 21044
rect 9857 21040 11284 21042
rect 9857 20984 9862 21040
rect 9918 20984 11242 21040
rect 9857 20982 11284 20984
rect 9857 20979 9923 20982
rect 11237 20980 11284 20982
rect 11348 20980 11354 21044
rect 11237 20979 11303 20980
rect 1485 20906 1551 20909
rect 3233 20908 3299 20909
rect 3182 20906 3188 20908
rect 1485 20904 3188 20906
rect 3252 20906 3299 20908
rect 4613 20906 4679 20909
rect 11145 20906 11211 20909
rect 3252 20904 3380 20906
rect 1485 20848 1490 20904
rect 1546 20848 3188 20904
rect 3294 20848 3380 20904
rect 1485 20846 3188 20848
rect 1485 20843 1551 20846
rect 3182 20844 3188 20846
rect 3252 20846 3380 20848
rect 4613 20904 11211 20906
rect 4613 20848 4618 20904
rect 4674 20848 11150 20904
rect 11206 20848 11211 20904
rect 4613 20846 11211 20848
rect 3252 20844 3299 20846
rect 3233 20843 3299 20844
rect 4613 20843 4679 20846
rect 11145 20843 11211 20846
rect -300 20770 160 20800
rect 1485 20770 1551 20773
rect -300 20768 1551 20770
rect -300 20712 1490 20768
rect 1546 20712 1551 20768
rect -300 20710 1551 20712
rect -300 20680 160 20710
rect 1485 20707 1551 20710
rect 2129 20770 2195 20773
rect 5165 20770 5231 20773
rect 2129 20768 5231 20770
rect 2129 20712 2134 20768
rect 2190 20712 5170 20768
rect 5226 20712 5231 20768
rect 2129 20710 5231 20712
rect 2129 20707 2195 20710
rect 5165 20707 5231 20710
rect 8385 20770 8451 20773
rect 9438 20770 9444 20772
rect 8385 20768 9444 20770
rect 8385 20712 8390 20768
rect 8446 20712 9444 20768
rect 8385 20710 9444 20712
rect 8385 20707 8451 20710
rect 9438 20708 9444 20710
rect 9508 20708 9514 20772
rect 13302 20708 13308 20772
rect 13372 20770 13378 20772
rect 13537 20770 13603 20773
rect 13372 20768 13603 20770
rect 13372 20712 13542 20768
rect 13598 20712 13603 20768
rect 13372 20710 13603 20712
rect 13372 20708 13378 20710
rect 13537 20707 13603 20710
rect 13670 20708 13676 20772
rect 13740 20770 13746 20772
rect 14590 20770 14596 20772
rect 13740 20710 14596 20770
rect 13740 20708 13746 20710
rect 14590 20708 14596 20710
rect 14660 20708 14666 20772
rect 24853 20770 24919 20773
rect 25540 20770 26000 20800
rect 24853 20768 26000 20770
rect 24853 20712 24858 20768
rect 24914 20712 26000 20768
rect 24853 20710 26000 20712
rect 24853 20707 24919 20710
rect 6810 20704 7126 20705
rect 6810 20640 6816 20704
rect 6880 20640 6896 20704
rect 6960 20640 6976 20704
rect 7040 20640 7056 20704
rect 7120 20640 7126 20704
rect 6810 20639 7126 20640
rect 12675 20704 12991 20705
rect 12675 20640 12681 20704
rect 12745 20640 12761 20704
rect 12825 20640 12841 20704
rect 12905 20640 12921 20704
rect 12985 20640 12991 20704
rect 12675 20639 12991 20640
rect 18540 20704 18856 20705
rect 18540 20640 18546 20704
rect 18610 20640 18626 20704
rect 18690 20640 18706 20704
rect 18770 20640 18786 20704
rect 18850 20640 18856 20704
rect 18540 20639 18856 20640
rect 24405 20704 24721 20705
rect 24405 20640 24411 20704
rect 24475 20640 24491 20704
rect 24555 20640 24571 20704
rect 24635 20640 24651 20704
rect 24715 20640 24721 20704
rect 25540 20680 26000 20710
rect 24405 20639 24721 20640
rect 2037 20636 2103 20637
rect 2037 20634 2084 20636
rect 1992 20632 2084 20634
rect 1992 20576 2042 20632
rect 1992 20574 2084 20576
rect 2037 20572 2084 20574
rect 2148 20572 2154 20636
rect 4337 20634 4403 20637
rect 5390 20634 5396 20636
rect 4337 20632 5396 20634
rect 4337 20576 4342 20632
rect 4398 20576 5396 20632
rect 4337 20574 5396 20576
rect 2037 20571 2103 20572
rect 4337 20571 4403 20574
rect 5390 20572 5396 20574
rect 5460 20572 5466 20636
rect 9489 20634 9555 20637
rect 7238 20632 9555 20634
rect 7238 20576 9494 20632
rect 9550 20576 9555 20632
rect 7238 20574 9555 20576
rect -300 20498 160 20528
rect 933 20498 999 20501
rect -300 20496 999 20498
rect -300 20440 938 20496
rect 994 20440 999 20496
rect -300 20438 999 20440
rect -300 20408 160 20438
rect 933 20435 999 20438
rect 1577 20498 1643 20501
rect 3417 20498 3483 20501
rect 7238 20498 7298 20574
rect 9489 20571 9555 20574
rect 14181 20634 14247 20637
rect 14406 20634 14412 20636
rect 14181 20632 14412 20634
rect 14181 20576 14186 20632
rect 14242 20576 14412 20632
rect 14181 20574 14412 20576
rect 14181 20571 14247 20574
rect 14406 20572 14412 20574
rect 14476 20572 14482 20636
rect 1577 20496 2790 20498
rect 1577 20440 1582 20496
rect 1638 20440 2790 20496
rect 1577 20438 2790 20440
rect 1577 20435 1643 20438
rect 2730 20362 2790 20438
rect 3417 20496 7298 20498
rect 3417 20440 3422 20496
rect 3478 20440 7298 20496
rect 3417 20438 7298 20440
rect 7373 20498 7439 20501
rect 12341 20498 12407 20501
rect 14958 20498 14964 20500
rect 7373 20496 14964 20498
rect 7373 20440 7378 20496
rect 7434 20440 12346 20496
rect 12402 20440 14964 20496
rect 7373 20438 14964 20440
rect 3417 20435 3483 20438
rect 7373 20435 7439 20438
rect 12341 20435 12407 20438
rect 14958 20436 14964 20438
rect 15028 20436 15034 20500
rect 10133 20362 10199 20365
rect 2730 20360 10199 20362
rect 2730 20304 10138 20360
rect 10194 20304 10199 20360
rect 2730 20302 10199 20304
rect 10133 20299 10199 20302
rect 11513 20362 11579 20365
rect 13813 20362 13879 20365
rect 11513 20360 13879 20362
rect 11513 20304 11518 20360
rect 11574 20304 13818 20360
rect 13874 20304 13879 20360
rect 11513 20302 13879 20304
rect 11513 20299 11579 20302
rect 13813 20299 13879 20302
rect -300 20226 160 20256
rect 749 20226 815 20229
rect -300 20224 815 20226
rect -300 20168 754 20224
rect 810 20168 815 20224
rect -300 20166 815 20168
rect -300 20136 160 20166
rect 749 20163 815 20166
rect 10174 20164 10180 20228
rect 10244 20226 10250 20228
rect 14958 20226 14964 20228
rect 10244 20166 14964 20226
rect 10244 20164 10250 20166
rect 14958 20164 14964 20166
rect 15028 20164 15034 20228
rect 23749 20226 23815 20229
rect 25540 20226 26000 20256
rect 23749 20224 26000 20226
rect 23749 20168 23754 20224
rect 23810 20168 26000 20224
rect 23749 20166 26000 20168
rect 23749 20163 23815 20166
rect 3878 20160 4194 20161
rect 3878 20096 3884 20160
rect 3948 20096 3964 20160
rect 4028 20096 4044 20160
rect 4108 20096 4124 20160
rect 4188 20096 4194 20160
rect 3878 20095 4194 20096
rect 9743 20160 10059 20161
rect 9743 20096 9749 20160
rect 9813 20096 9829 20160
rect 9893 20096 9909 20160
rect 9973 20096 9989 20160
rect 10053 20096 10059 20160
rect 9743 20095 10059 20096
rect 15608 20160 15924 20161
rect 15608 20096 15614 20160
rect 15678 20096 15694 20160
rect 15758 20096 15774 20160
rect 15838 20096 15854 20160
rect 15918 20096 15924 20160
rect 15608 20095 15924 20096
rect 21473 20160 21789 20161
rect 21473 20096 21479 20160
rect 21543 20096 21559 20160
rect 21623 20096 21639 20160
rect 21703 20096 21719 20160
rect 21783 20096 21789 20160
rect 25540 20136 26000 20166
rect 21473 20095 21789 20096
rect 1669 20092 1735 20093
rect 1669 20090 1716 20092
rect 1624 20088 1716 20090
rect 1624 20032 1674 20088
rect 1624 20030 1716 20032
rect 1669 20028 1716 20030
rect 1780 20028 1786 20092
rect 1669 20027 1735 20028
rect -300 19954 160 19984
rect 1393 19954 1459 19957
rect -300 19952 1459 19954
rect -300 19896 1398 19952
rect 1454 19896 1459 19952
rect -300 19894 1459 19896
rect -300 19864 160 19894
rect 1393 19891 1459 19894
rect 3509 19954 3575 19957
rect 3734 19954 3740 19956
rect 3509 19952 3740 19954
rect 3509 19896 3514 19952
rect 3570 19896 3740 19952
rect 3509 19894 3740 19896
rect 3509 19891 3575 19894
rect 3734 19892 3740 19894
rect 3804 19954 3810 19956
rect 5390 19954 5396 19956
rect 3804 19894 5396 19954
rect 3804 19892 3810 19894
rect 5390 19892 5396 19894
rect 5460 19892 5466 19956
rect 5533 19954 5599 19957
rect 10358 19954 10364 19956
rect 5533 19952 10364 19954
rect 5533 19896 5538 19952
rect 5594 19896 10364 19952
rect 5533 19894 10364 19896
rect 5533 19891 5599 19894
rect 10358 19892 10364 19894
rect 10428 19954 10434 19956
rect 10501 19954 10567 19957
rect 10428 19952 10567 19954
rect 10428 19896 10506 19952
rect 10562 19896 10567 19952
rect 10428 19894 10567 19896
rect 10428 19892 10434 19894
rect 10501 19891 10567 19894
rect 2037 19818 2103 19821
rect 4061 19818 4127 19821
rect 13905 19818 13971 19821
rect 18413 19818 18479 19821
rect 2037 19816 3618 19818
rect 2037 19760 2042 19816
rect 2098 19760 3618 19816
rect 2037 19758 3618 19760
rect 2037 19755 2103 19758
rect -300 19682 160 19712
rect 1301 19682 1367 19685
rect -300 19680 1367 19682
rect -300 19624 1306 19680
rect 1362 19624 1367 19680
rect -300 19622 1367 19624
rect -300 19592 160 19622
rect 1301 19619 1367 19622
rect 2129 19682 2195 19685
rect 3417 19684 3483 19685
rect 3366 19682 3372 19684
rect 2129 19680 3250 19682
rect 2129 19624 2134 19680
rect 2190 19624 3250 19680
rect 2129 19622 3250 19624
rect 3326 19622 3372 19682
rect 3436 19680 3483 19684
rect 3478 19624 3483 19680
rect 2129 19619 2195 19622
rect 2221 19548 2287 19549
rect 2221 19546 2268 19548
rect 2176 19544 2268 19546
rect 2176 19488 2226 19544
rect 2176 19486 2268 19488
rect 2221 19484 2268 19486
rect 2332 19484 2338 19548
rect 3190 19546 3250 19622
rect 3366 19620 3372 19622
rect 3436 19620 3483 19624
rect 3558 19682 3618 19758
rect 4061 19816 7666 19818
rect 4061 19760 4066 19816
rect 4122 19760 7666 19816
rect 4061 19758 7666 19760
rect 4061 19755 4127 19758
rect 5574 19682 5580 19684
rect 3558 19622 5580 19682
rect 5574 19620 5580 19622
rect 5644 19620 5650 19684
rect 5901 19682 5967 19685
rect 6361 19682 6427 19685
rect 5901 19680 6427 19682
rect 5901 19624 5906 19680
rect 5962 19624 6366 19680
rect 6422 19624 6427 19680
rect 5901 19622 6427 19624
rect 3417 19619 3483 19620
rect 5901 19619 5967 19622
rect 6361 19619 6427 19622
rect 6810 19616 7126 19617
rect 6810 19552 6816 19616
rect 6880 19552 6896 19616
rect 6960 19552 6976 19616
rect 7040 19552 7056 19616
rect 7120 19552 7126 19616
rect 6810 19551 7126 19552
rect 3190 19486 6746 19546
rect 2221 19483 2287 19484
rect -300 19410 160 19440
rect 1117 19410 1183 19413
rect -300 19408 1183 19410
rect -300 19352 1122 19408
rect 1178 19352 1183 19408
rect -300 19350 1183 19352
rect -300 19320 160 19350
rect 1117 19347 1183 19350
rect 1526 19348 1532 19412
rect 1596 19410 1602 19412
rect 3785 19410 3851 19413
rect 1596 19408 3851 19410
rect 1596 19352 3790 19408
rect 3846 19352 3851 19408
rect 1596 19350 3851 19352
rect 6686 19410 6746 19486
rect 7373 19444 7439 19447
rect 7192 19442 7439 19444
rect 7192 19410 7378 19442
rect 6686 19386 7378 19410
rect 7434 19386 7439 19442
rect 6686 19384 7439 19386
rect 6686 19350 7252 19384
rect 7373 19381 7439 19384
rect 7606 19353 7666 19758
rect 13905 19816 18479 19818
rect 13905 19760 13910 19816
rect 13966 19760 18418 19816
rect 18474 19760 18479 19816
rect 13905 19758 18479 19760
rect 13905 19755 13971 19758
rect 18413 19755 18479 19758
rect 13169 19682 13235 19685
rect 17493 19682 17559 19685
rect 13169 19680 17559 19682
rect 13169 19624 13174 19680
rect 13230 19624 17498 19680
rect 17554 19624 17559 19680
rect 13169 19622 17559 19624
rect 13169 19619 13235 19622
rect 17493 19619 17559 19622
rect 25129 19682 25195 19685
rect 25540 19682 26000 19712
rect 25129 19680 26000 19682
rect 25129 19624 25134 19680
rect 25190 19624 26000 19680
rect 25129 19622 26000 19624
rect 25129 19619 25195 19622
rect 12675 19616 12991 19617
rect 12675 19552 12681 19616
rect 12745 19552 12761 19616
rect 12825 19552 12841 19616
rect 12905 19552 12921 19616
rect 12985 19552 12991 19616
rect 12675 19551 12991 19552
rect 18540 19616 18856 19617
rect 18540 19552 18546 19616
rect 18610 19552 18626 19616
rect 18690 19552 18706 19616
rect 18770 19552 18786 19616
rect 18850 19552 18856 19616
rect 18540 19551 18856 19552
rect 24405 19616 24721 19617
rect 24405 19552 24411 19616
rect 24475 19552 24491 19616
rect 24555 19552 24571 19616
rect 24635 19552 24651 19616
rect 24715 19552 24721 19616
rect 25540 19592 26000 19622
rect 24405 19551 24721 19552
rect 15193 19546 15259 19549
rect 18137 19546 18203 19549
rect 15193 19544 18203 19546
rect 15193 19488 15198 19544
rect 15254 19488 18142 19544
rect 18198 19488 18203 19544
rect 15193 19486 18203 19488
rect 15193 19483 15259 19486
rect 18137 19483 18203 19486
rect 1596 19348 1602 19350
rect 3785 19347 3851 19350
rect 7557 19348 7666 19353
rect 7557 19292 7562 19348
rect 7618 19292 7666 19348
rect 12065 19410 12131 19413
rect 13353 19410 13419 19413
rect 12065 19408 13419 19410
rect 12065 19352 12070 19408
rect 12126 19352 13358 19408
rect 13414 19352 13419 19408
rect 12065 19350 13419 19352
rect 12065 19347 12131 19350
rect 13353 19347 13419 19350
rect 14273 19410 14339 19413
rect 15142 19410 15148 19412
rect 14273 19408 15148 19410
rect 14273 19352 14278 19408
rect 14334 19352 15148 19408
rect 14273 19350 15148 19352
rect 14273 19347 14339 19350
rect 15142 19348 15148 19350
rect 15212 19348 15218 19412
rect 16430 19348 16436 19412
rect 16500 19410 16506 19412
rect 16665 19410 16731 19413
rect 16500 19408 16731 19410
rect 16500 19352 16670 19408
rect 16726 19352 16731 19408
rect 16500 19350 16731 19352
rect 16500 19348 16506 19350
rect 16665 19347 16731 19350
rect 17769 19410 17835 19413
rect 18086 19410 18092 19412
rect 17769 19408 18092 19410
rect 17769 19352 17774 19408
rect 17830 19352 18092 19408
rect 17769 19350 18092 19352
rect 17769 19347 17835 19350
rect 18086 19348 18092 19350
rect 18156 19348 18162 19412
rect 7557 19290 7666 19292
rect 7557 19287 7623 19290
rect 2589 19274 2655 19277
rect 5441 19274 5507 19277
rect 2589 19272 5507 19274
rect 2589 19216 2594 19272
rect 2650 19216 5446 19272
rect 5502 19216 5507 19272
rect 2589 19214 5507 19216
rect 2589 19211 2655 19214
rect 5441 19211 5507 19214
rect -300 19138 160 19168
rect 749 19138 815 19141
rect -300 19136 815 19138
rect -300 19080 754 19136
rect 810 19080 815 19136
rect -300 19078 815 19080
rect -300 19048 160 19078
rect 749 19075 815 19078
rect 4286 19076 4292 19140
rect 4356 19138 4362 19140
rect 6453 19138 6519 19141
rect 4356 19136 6519 19138
rect 4356 19080 6458 19136
rect 6514 19080 6519 19136
rect 4356 19078 6519 19080
rect 4356 19076 4362 19078
rect 6453 19075 6519 19078
rect 8753 19138 8819 19141
rect 23933 19138 23999 19141
rect 25540 19138 26000 19168
rect 8753 19136 9322 19138
rect 8753 19080 8758 19136
rect 8814 19080 9322 19136
rect 8753 19078 9322 19080
rect 8753 19075 8819 19078
rect 3878 19072 4194 19073
rect 3878 19008 3884 19072
rect 3948 19008 3964 19072
rect 4028 19008 4044 19072
rect 4108 19008 4124 19072
rect 4188 19008 4194 19072
rect 3878 19007 4194 19008
rect 4521 19002 4587 19005
rect 7741 19002 7807 19005
rect 9121 19002 9187 19005
rect 4521 19000 9187 19002
rect 4521 18944 4526 19000
rect 4582 18944 7746 19000
rect 7802 18944 9126 19000
rect 9182 18944 9187 19000
rect 4521 18942 9187 18944
rect 4521 18939 4587 18942
rect 7741 18939 7807 18942
rect 9121 18939 9187 18942
rect -300 18866 160 18896
rect 2773 18866 2839 18869
rect 8753 18866 8819 18869
rect -300 18864 2839 18866
rect -300 18808 2778 18864
rect 2834 18808 2839 18864
rect -300 18806 2839 18808
rect -300 18776 160 18806
rect 2773 18803 2839 18806
rect 5030 18864 8819 18866
rect 5030 18808 8758 18864
rect 8814 18808 8819 18864
rect 5030 18806 8819 18808
rect 9262 18866 9322 19078
rect 23933 19136 26000 19138
rect 23933 19080 23938 19136
rect 23994 19080 26000 19136
rect 23933 19078 26000 19080
rect 23933 19075 23999 19078
rect 9743 19072 10059 19073
rect 9743 19008 9749 19072
rect 9813 19008 9829 19072
rect 9893 19008 9909 19072
rect 9973 19008 9989 19072
rect 10053 19008 10059 19072
rect 9743 19007 10059 19008
rect 15608 19072 15924 19073
rect 15608 19008 15614 19072
rect 15678 19008 15694 19072
rect 15758 19008 15774 19072
rect 15838 19008 15854 19072
rect 15918 19008 15924 19072
rect 15608 19007 15924 19008
rect 21473 19072 21789 19073
rect 21473 19008 21479 19072
rect 21543 19008 21559 19072
rect 21623 19008 21639 19072
rect 21703 19008 21719 19072
rect 21783 19008 21789 19072
rect 25540 19048 26000 19078
rect 21473 19007 21789 19008
rect 9949 18866 10015 18869
rect 9262 18864 10015 18866
rect 9262 18808 9954 18864
rect 10010 18808 10015 18864
rect 9262 18806 10015 18808
rect 1761 18730 1827 18733
rect 2630 18730 2636 18732
rect 1761 18728 2636 18730
rect 1761 18672 1766 18728
rect 1822 18672 2636 18728
rect 1761 18670 2636 18672
rect 1761 18667 1827 18670
rect 2630 18668 2636 18670
rect 2700 18730 2706 18732
rect 5030 18730 5090 18806
rect 8753 18803 8819 18806
rect 9949 18803 10015 18806
rect 2700 18670 5090 18730
rect 5349 18730 5415 18733
rect 11145 18730 11211 18733
rect 5349 18728 11211 18730
rect 5349 18672 5354 18728
rect 5410 18672 11150 18728
rect 11206 18672 11211 18728
rect 5349 18670 11211 18672
rect 2700 18668 2706 18670
rect 5349 18667 5415 18670
rect 11145 18667 11211 18670
rect -300 18594 160 18624
rect 3785 18594 3851 18597
rect -300 18592 3851 18594
rect -300 18536 3790 18592
rect 3846 18536 3851 18592
rect -300 18534 3851 18536
rect -300 18504 160 18534
rect 3785 18531 3851 18534
rect 8569 18594 8635 18597
rect 10225 18594 10291 18597
rect 8569 18592 10291 18594
rect 8569 18536 8574 18592
rect 8630 18536 10230 18592
rect 10286 18536 10291 18592
rect 8569 18534 10291 18536
rect 8569 18531 8635 18534
rect 10225 18531 10291 18534
rect 24853 18594 24919 18597
rect 25540 18594 26000 18624
rect 24853 18592 26000 18594
rect 24853 18536 24858 18592
rect 24914 18536 26000 18592
rect 24853 18534 26000 18536
rect 24853 18531 24919 18534
rect 6810 18528 7126 18529
rect 6810 18464 6816 18528
rect 6880 18464 6896 18528
rect 6960 18464 6976 18528
rect 7040 18464 7056 18528
rect 7120 18464 7126 18528
rect 6810 18463 7126 18464
rect 12675 18528 12991 18529
rect 12675 18464 12681 18528
rect 12745 18464 12761 18528
rect 12825 18464 12841 18528
rect 12905 18464 12921 18528
rect 12985 18464 12991 18528
rect 12675 18463 12991 18464
rect 18540 18528 18856 18529
rect 18540 18464 18546 18528
rect 18610 18464 18626 18528
rect 18690 18464 18706 18528
rect 18770 18464 18786 18528
rect 18850 18464 18856 18528
rect 18540 18463 18856 18464
rect 24405 18528 24721 18529
rect 24405 18464 24411 18528
rect 24475 18464 24491 18528
rect 24555 18464 24571 18528
rect 24635 18464 24651 18528
rect 24715 18464 24721 18528
rect 25540 18504 26000 18534
rect 24405 18463 24721 18464
rect 2129 18458 2195 18461
rect 6453 18458 6519 18461
rect 2129 18456 6519 18458
rect 2129 18400 2134 18456
rect 2190 18400 6458 18456
rect 6514 18400 6519 18456
rect 2129 18398 6519 18400
rect 2129 18395 2195 18398
rect 6453 18395 6519 18398
rect 8702 18396 8708 18460
rect 8772 18458 8778 18460
rect 9397 18458 9463 18461
rect 8772 18456 9463 18458
rect 8772 18400 9402 18456
rect 9458 18400 9463 18456
rect 8772 18398 9463 18400
rect 8772 18396 8778 18398
rect 9397 18395 9463 18398
rect -300 18322 160 18352
rect 2773 18322 2839 18325
rect -300 18320 2839 18322
rect -300 18264 2778 18320
rect 2834 18264 2839 18320
rect -300 18262 2839 18264
rect -300 18232 160 18262
rect 2773 18259 2839 18262
rect 2957 18322 3023 18325
rect 11237 18322 11303 18325
rect 2957 18320 11303 18322
rect 2957 18264 2962 18320
rect 3018 18264 11242 18320
rect 11298 18264 11303 18320
rect 2957 18262 11303 18264
rect 2957 18259 3023 18262
rect 11237 18259 11303 18262
rect 6269 18186 6335 18189
rect 9489 18186 9555 18189
rect 6269 18184 9555 18186
rect 6269 18128 6274 18184
rect 6330 18128 9494 18184
rect 9550 18128 9555 18184
rect 6269 18126 9555 18128
rect 6269 18123 6335 18126
rect 9489 18123 9555 18126
rect -300 18050 160 18080
rect 3601 18050 3667 18053
rect -300 18048 3667 18050
rect -300 17992 3606 18048
rect 3662 17992 3667 18048
rect -300 17990 3667 17992
rect -300 17960 160 17990
rect 3601 17987 3667 17990
rect 5993 18050 6059 18053
rect 6310 18050 6316 18052
rect 5993 18048 6316 18050
rect 5993 17992 5998 18048
rect 6054 17992 6316 18048
rect 5993 17990 6316 17992
rect 5993 17987 6059 17990
rect 6310 17988 6316 17990
rect 6380 17988 6386 18052
rect 23565 18050 23631 18053
rect 25540 18050 26000 18080
rect 23565 18048 26000 18050
rect 23565 17992 23570 18048
rect 23626 17992 26000 18048
rect 23565 17990 26000 17992
rect 23565 17987 23631 17990
rect 3878 17984 4194 17985
rect 3878 17920 3884 17984
rect 3948 17920 3964 17984
rect 4028 17920 4044 17984
rect 4108 17920 4124 17984
rect 4188 17920 4194 17984
rect 3878 17919 4194 17920
rect 9743 17984 10059 17985
rect 9743 17920 9749 17984
rect 9813 17920 9829 17984
rect 9893 17920 9909 17984
rect 9973 17920 9989 17984
rect 10053 17920 10059 17984
rect 9743 17919 10059 17920
rect 15608 17984 15924 17985
rect 15608 17920 15614 17984
rect 15678 17920 15694 17984
rect 15758 17920 15774 17984
rect 15838 17920 15854 17984
rect 15918 17920 15924 17984
rect 15608 17919 15924 17920
rect 21473 17984 21789 17985
rect 21473 17920 21479 17984
rect 21543 17920 21559 17984
rect 21623 17920 21639 17984
rect 21703 17920 21719 17984
rect 21783 17920 21789 17984
rect 25540 17960 26000 17990
rect 21473 17919 21789 17920
rect 5625 17914 5691 17917
rect 5758 17914 5764 17916
rect 5625 17912 5764 17914
rect 5625 17856 5630 17912
rect 5686 17856 5764 17912
rect 5625 17854 5764 17856
rect 5625 17851 5691 17854
rect 5758 17852 5764 17854
rect 5828 17852 5834 17916
rect -300 17778 160 17808
rect 3233 17778 3299 17781
rect -300 17776 3299 17778
rect -300 17720 3238 17776
rect 3294 17720 3299 17776
rect -300 17718 3299 17720
rect -300 17688 160 17718
rect 3233 17715 3299 17718
rect 13854 17716 13860 17780
rect 13924 17778 13930 17780
rect 14733 17778 14799 17781
rect 16246 17778 16252 17780
rect 13924 17776 16252 17778
rect 13924 17720 14738 17776
rect 14794 17720 16252 17776
rect 13924 17718 16252 17720
rect 13924 17716 13930 17718
rect 14733 17715 14799 17718
rect 16246 17716 16252 17718
rect 16316 17716 16322 17780
rect -300 17506 160 17536
rect 1301 17506 1367 17509
rect -300 17504 1367 17506
rect -300 17448 1306 17504
rect 1362 17448 1367 17504
rect -300 17446 1367 17448
rect -300 17416 160 17446
rect 1301 17443 1367 17446
rect 2589 17506 2655 17509
rect 2998 17506 3004 17508
rect 2589 17504 3004 17506
rect 2589 17448 2594 17504
rect 2650 17448 3004 17504
rect 2589 17446 3004 17448
rect 2589 17443 2655 17446
rect 2998 17444 3004 17446
rect 3068 17444 3074 17508
rect 24853 17506 24919 17509
rect 25540 17506 26000 17536
rect 24853 17504 26000 17506
rect 24853 17448 24858 17504
rect 24914 17448 26000 17504
rect 24853 17446 26000 17448
rect 24853 17443 24919 17446
rect 6810 17440 7126 17441
rect 6810 17376 6816 17440
rect 6880 17376 6896 17440
rect 6960 17376 6976 17440
rect 7040 17376 7056 17440
rect 7120 17376 7126 17440
rect 6810 17375 7126 17376
rect 12675 17440 12991 17441
rect 12675 17376 12681 17440
rect 12745 17376 12761 17440
rect 12825 17376 12841 17440
rect 12905 17376 12921 17440
rect 12985 17376 12991 17440
rect 12675 17375 12991 17376
rect 18540 17440 18856 17441
rect 18540 17376 18546 17440
rect 18610 17376 18626 17440
rect 18690 17376 18706 17440
rect 18770 17376 18786 17440
rect 18850 17376 18856 17440
rect 18540 17375 18856 17376
rect 24405 17440 24721 17441
rect 24405 17376 24411 17440
rect 24475 17376 24491 17440
rect 24555 17376 24571 17440
rect 24635 17376 24651 17440
rect 24715 17376 24721 17440
rect 25540 17416 26000 17446
rect 24405 17375 24721 17376
rect 1710 17308 1716 17372
rect 1780 17370 1786 17372
rect 2221 17370 2287 17373
rect 6637 17370 6703 17373
rect 1780 17368 6703 17370
rect 1780 17312 2226 17368
rect 2282 17312 6642 17368
rect 6698 17312 6703 17368
rect 1780 17310 6703 17312
rect 1780 17308 1786 17310
rect 2221 17307 2287 17310
rect 6637 17307 6703 17310
rect -300 17234 160 17264
rect 3417 17234 3483 17237
rect -300 17232 3483 17234
rect -300 17176 3422 17232
rect 3478 17176 3483 17232
rect -300 17174 3483 17176
rect -300 17144 160 17174
rect 3417 17171 3483 17174
rect 4061 17234 4127 17237
rect 6494 17234 6500 17236
rect 4061 17232 6500 17234
rect 4061 17176 4066 17232
rect 4122 17176 6500 17232
rect 4061 17174 6500 17176
rect 4061 17171 4127 17174
rect 6494 17172 6500 17174
rect 6564 17234 6570 17236
rect 6821 17234 6887 17237
rect 6564 17232 6887 17234
rect 6564 17176 6826 17232
rect 6882 17176 6887 17232
rect 6564 17174 6887 17176
rect 6564 17172 6570 17174
rect 6821 17171 6887 17174
rect 7281 17234 7347 17237
rect 9305 17234 9371 17237
rect 7281 17232 9371 17234
rect 7281 17176 7286 17232
rect 7342 17176 9310 17232
rect 9366 17176 9371 17232
rect 7281 17174 9371 17176
rect 7281 17171 7347 17174
rect 9305 17171 9371 17174
rect 13813 17234 13879 17237
rect 16481 17234 16547 17237
rect 13813 17232 16547 17234
rect 13813 17176 13818 17232
rect 13874 17176 16486 17232
rect 16542 17176 16547 17232
rect 13813 17174 16547 17176
rect 13813 17171 13879 17174
rect 16481 17171 16547 17174
rect 5165 17098 5231 17101
rect 6453 17098 6519 17101
rect 8017 17098 8083 17101
rect 16573 17098 16639 17101
rect 5165 17096 8083 17098
rect 5165 17040 5170 17096
rect 5226 17040 6458 17096
rect 6514 17040 8022 17096
rect 8078 17040 8083 17096
rect 5165 17038 8083 17040
rect 5165 17035 5231 17038
rect 6453 17035 6519 17038
rect 8017 17035 8083 17038
rect 10182 17096 16639 17098
rect 10182 17040 16578 17096
rect 16634 17040 16639 17096
rect 10182 17038 16639 17040
rect -300 16962 160 16992
rect 841 16962 907 16965
rect -300 16960 907 16962
rect -300 16904 846 16960
rect 902 16904 907 16960
rect -300 16902 907 16904
rect -300 16872 160 16902
rect 841 16899 907 16902
rect 3878 16896 4194 16897
rect 3878 16832 3884 16896
rect 3948 16832 3964 16896
rect 4028 16832 4044 16896
rect 4108 16832 4124 16896
rect 4188 16832 4194 16896
rect 3878 16831 4194 16832
rect 9743 16896 10059 16897
rect 9743 16832 9749 16896
rect 9813 16832 9829 16896
rect 9893 16832 9909 16896
rect 9973 16832 9989 16896
rect 10053 16832 10059 16896
rect 9743 16831 10059 16832
rect -300 16690 160 16720
rect 3693 16690 3759 16693
rect -300 16688 3759 16690
rect -300 16632 3698 16688
rect 3754 16632 3759 16688
rect -300 16630 3759 16632
rect -300 16600 160 16630
rect 3693 16627 3759 16630
rect 4613 16690 4679 16693
rect 8017 16690 8083 16693
rect 4613 16688 8083 16690
rect 4613 16632 4618 16688
rect 4674 16632 8022 16688
rect 8078 16632 8083 16688
rect 4613 16630 8083 16632
rect 4613 16627 4679 16630
rect 8017 16627 8083 16630
rect 10041 16690 10107 16693
rect 10182 16690 10242 17038
rect 16573 17035 16639 17038
rect 23565 16962 23631 16965
rect 25540 16962 26000 16992
rect 23565 16960 26000 16962
rect 23565 16904 23570 16960
rect 23626 16904 26000 16960
rect 23565 16902 26000 16904
rect 23565 16899 23631 16902
rect 15608 16896 15924 16897
rect 15608 16832 15614 16896
rect 15678 16832 15694 16896
rect 15758 16832 15774 16896
rect 15838 16832 15854 16896
rect 15918 16832 15924 16896
rect 15608 16831 15924 16832
rect 21473 16896 21789 16897
rect 21473 16832 21479 16896
rect 21543 16832 21559 16896
rect 21623 16832 21639 16896
rect 21703 16832 21719 16896
rect 21783 16832 21789 16896
rect 25540 16872 26000 16902
rect 21473 16831 21789 16832
rect 10317 16826 10383 16829
rect 10869 16826 10935 16829
rect 10317 16824 10935 16826
rect 10317 16768 10322 16824
rect 10378 16768 10874 16824
rect 10930 16768 10935 16824
rect 10317 16766 10935 16768
rect 10317 16763 10383 16766
rect 10869 16763 10935 16766
rect 10041 16688 10242 16690
rect 10041 16632 10046 16688
rect 10102 16632 10242 16688
rect 10041 16630 10242 16632
rect 11605 16690 11671 16693
rect 13353 16690 13419 16693
rect 11605 16688 13419 16690
rect 11605 16632 11610 16688
rect 11666 16632 13358 16688
rect 13414 16632 13419 16688
rect 11605 16630 13419 16632
rect 10041 16627 10107 16630
rect 11605 16627 11671 16630
rect 13353 16627 13419 16630
rect 4245 16554 4311 16557
rect 7465 16554 7531 16557
rect 4245 16552 7531 16554
rect 4245 16496 4250 16552
rect 4306 16496 7470 16552
rect 7526 16496 7531 16552
rect 4245 16494 7531 16496
rect 4245 16491 4311 16494
rect 7465 16491 7531 16494
rect 8109 16554 8175 16557
rect 9070 16554 9076 16556
rect 8109 16552 9076 16554
rect 8109 16496 8114 16552
rect 8170 16496 9076 16552
rect 8109 16494 9076 16496
rect 8109 16491 8175 16494
rect 9070 16492 9076 16494
rect 9140 16492 9146 16556
rect 10910 16492 10916 16556
rect 10980 16554 10986 16556
rect 20846 16554 20852 16556
rect 10980 16494 20852 16554
rect 10980 16492 10986 16494
rect 20846 16492 20852 16494
rect 20916 16492 20922 16556
rect -300 16418 160 16448
rect 3325 16418 3391 16421
rect -300 16416 3391 16418
rect -300 16360 3330 16416
rect 3386 16360 3391 16416
rect -300 16358 3391 16360
rect -300 16328 160 16358
rect 3325 16355 3391 16358
rect 24853 16418 24919 16421
rect 25540 16418 26000 16448
rect 24853 16416 26000 16418
rect 24853 16360 24858 16416
rect 24914 16360 26000 16416
rect 24853 16358 26000 16360
rect 24853 16355 24919 16358
rect 6810 16352 7126 16353
rect 6810 16288 6816 16352
rect 6880 16288 6896 16352
rect 6960 16288 6976 16352
rect 7040 16288 7056 16352
rect 7120 16288 7126 16352
rect 6810 16287 7126 16288
rect 12675 16352 12991 16353
rect 12675 16288 12681 16352
rect 12745 16288 12761 16352
rect 12825 16288 12841 16352
rect 12905 16288 12921 16352
rect 12985 16288 12991 16352
rect 12675 16287 12991 16288
rect 18540 16352 18856 16353
rect 18540 16288 18546 16352
rect 18610 16288 18626 16352
rect 18690 16288 18706 16352
rect 18770 16288 18786 16352
rect 18850 16288 18856 16352
rect 18540 16287 18856 16288
rect 24405 16352 24721 16353
rect 24405 16288 24411 16352
rect 24475 16288 24491 16352
rect 24555 16288 24571 16352
rect 24635 16288 24651 16352
rect 24715 16288 24721 16352
rect 25540 16328 26000 16358
rect 24405 16287 24721 16288
rect 4153 16282 4219 16285
rect 6453 16282 6519 16285
rect 4153 16280 6519 16282
rect 4153 16224 4158 16280
rect 4214 16224 6458 16280
rect 6514 16224 6519 16280
rect 4153 16222 6519 16224
rect 4153 16219 4219 16222
rect 6453 16219 6519 16222
rect -300 16146 160 16176
rect 1577 16146 1643 16149
rect -300 16144 1643 16146
rect -300 16088 1582 16144
rect 1638 16088 1643 16144
rect -300 16086 1643 16088
rect -300 16056 160 16086
rect 1577 16083 1643 16086
rect 5390 16084 5396 16148
rect 5460 16146 5466 16148
rect 8293 16146 8359 16149
rect 5460 16144 8359 16146
rect 5460 16088 8298 16144
rect 8354 16088 8359 16144
rect 5460 16086 8359 16088
rect 5460 16084 5466 16086
rect 8293 16083 8359 16086
rect 14958 16084 14964 16148
rect 15028 16146 15034 16148
rect 15285 16146 15351 16149
rect 15028 16144 15351 16146
rect 15028 16088 15290 16144
rect 15346 16088 15351 16144
rect 15028 16086 15351 16088
rect 15028 16084 15034 16086
rect 15285 16083 15351 16086
rect 1485 16010 1551 16013
rect 13169 16010 13235 16013
rect 1485 16008 13235 16010
rect 1485 15952 1490 16008
rect 1546 15952 13174 16008
rect 13230 15952 13235 16008
rect 1485 15950 13235 15952
rect 1485 15947 1551 15950
rect 13169 15947 13235 15950
rect -300 15874 160 15904
rect 1117 15874 1183 15877
rect -300 15872 1183 15874
rect -300 15816 1122 15872
rect 1178 15816 1183 15872
rect -300 15814 1183 15816
rect -300 15784 160 15814
rect 1117 15811 1183 15814
rect 5206 15812 5212 15876
rect 5276 15874 5282 15876
rect 6085 15874 6151 15877
rect 5276 15872 6151 15874
rect 5276 15816 6090 15872
rect 6146 15816 6151 15872
rect 5276 15814 6151 15816
rect 5276 15812 5282 15814
rect 6085 15811 6151 15814
rect 23749 15874 23815 15877
rect 25540 15874 26000 15904
rect 23749 15872 26000 15874
rect 23749 15816 23754 15872
rect 23810 15816 26000 15872
rect 23749 15814 26000 15816
rect 23749 15811 23815 15814
rect 3878 15808 4194 15809
rect 3878 15744 3884 15808
rect 3948 15744 3964 15808
rect 4028 15744 4044 15808
rect 4108 15744 4124 15808
rect 4188 15744 4194 15808
rect 3878 15743 4194 15744
rect 9743 15808 10059 15809
rect 9743 15744 9749 15808
rect 9813 15744 9829 15808
rect 9893 15744 9909 15808
rect 9973 15744 9989 15808
rect 10053 15744 10059 15808
rect 9743 15743 10059 15744
rect 15608 15808 15924 15809
rect 15608 15744 15614 15808
rect 15678 15744 15694 15808
rect 15758 15744 15774 15808
rect 15838 15744 15854 15808
rect 15918 15744 15924 15808
rect 15608 15743 15924 15744
rect 21473 15808 21789 15809
rect 21473 15744 21479 15808
rect 21543 15744 21559 15808
rect 21623 15744 21639 15808
rect 21703 15744 21719 15808
rect 21783 15744 21789 15808
rect 25540 15784 26000 15814
rect 21473 15743 21789 15744
rect 1894 15676 1900 15740
rect 1964 15738 1970 15740
rect 3233 15738 3299 15741
rect 1964 15736 3299 15738
rect 1964 15680 3238 15736
rect 3294 15680 3299 15736
rect 1964 15678 3299 15680
rect 1964 15676 1970 15678
rect 3233 15675 3299 15678
rect -300 15602 160 15632
rect 1301 15602 1367 15605
rect -300 15600 1367 15602
rect -300 15544 1306 15600
rect 1362 15544 1367 15600
rect -300 15542 1367 15544
rect -300 15512 160 15542
rect 1301 15539 1367 15542
rect 3877 15602 3943 15605
rect 8569 15602 8635 15605
rect 3877 15600 8635 15602
rect 3877 15544 3882 15600
rect 3938 15544 8574 15600
rect 8630 15544 8635 15600
rect 3877 15542 8635 15544
rect 3877 15539 3943 15542
rect 8569 15539 8635 15542
rect 8293 15466 8359 15469
rect 12525 15466 12591 15469
rect 8293 15464 12591 15466
rect 8293 15408 8298 15464
rect 8354 15408 12530 15464
rect 12586 15408 12591 15464
rect 8293 15406 12591 15408
rect 8293 15403 8359 15406
rect 12525 15403 12591 15406
rect 14733 15468 14799 15469
rect 14733 15464 14780 15468
rect 14844 15466 14850 15468
rect 14733 15408 14738 15464
rect 14733 15404 14780 15408
rect 14844 15406 14890 15466
rect 14844 15404 14850 15406
rect 14733 15403 14799 15404
rect -300 15330 160 15360
rect 1209 15330 1275 15333
rect -300 15328 1275 15330
rect -300 15272 1214 15328
rect 1270 15272 1275 15328
rect -300 15270 1275 15272
rect -300 15240 160 15270
rect 1209 15267 1275 15270
rect 2630 15268 2636 15332
rect 2700 15330 2706 15332
rect 3049 15330 3115 15333
rect 2700 15328 3115 15330
rect 2700 15272 3054 15328
rect 3110 15272 3115 15328
rect 2700 15270 3115 15272
rect 2700 15268 2706 15270
rect 3049 15267 3115 15270
rect 24853 15330 24919 15333
rect 25540 15330 26000 15360
rect 24853 15328 26000 15330
rect 24853 15272 24858 15328
rect 24914 15272 26000 15328
rect 24853 15270 26000 15272
rect 24853 15267 24919 15270
rect 6810 15264 7126 15265
rect 6810 15200 6816 15264
rect 6880 15200 6896 15264
rect 6960 15200 6976 15264
rect 7040 15200 7056 15264
rect 7120 15200 7126 15264
rect 6810 15199 7126 15200
rect 12675 15264 12991 15265
rect 12675 15200 12681 15264
rect 12745 15200 12761 15264
rect 12825 15200 12841 15264
rect 12905 15200 12921 15264
rect 12985 15200 12991 15264
rect 12675 15199 12991 15200
rect 18540 15264 18856 15265
rect 18540 15200 18546 15264
rect 18610 15200 18626 15264
rect 18690 15200 18706 15264
rect 18770 15200 18786 15264
rect 18850 15200 18856 15264
rect 18540 15199 18856 15200
rect 24405 15264 24721 15265
rect 24405 15200 24411 15264
rect 24475 15200 24491 15264
rect 24555 15200 24571 15264
rect 24635 15200 24651 15264
rect 24715 15200 24721 15264
rect 25540 15240 26000 15270
rect 24405 15199 24721 15200
rect 933 15194 999 15197
rect 5349 15194 5415 15197
rect 933 15192 5415 15194
rect 933 15136 938 15192
rect 994 15136 5354 15192
rect 5410 15136 5415 15192
rect 933 15134 5415 15136
rect 933 15131 999 15134
rect 5349 15131 5415 15134
rect 8201 15194 8267 15197
rect 8334 15194 8340 15196
rect 8201 15192 8340 15194
rect 8201 15136 8206 15192
rect 8262 15136 8340 15192
rect 8201 15134 8340 15136
rect 8201 15131 8267 15134
rect 8334 15132 8340 15134
rect 8404 15132 8410 15196
rect 13905 15194 13971 15197
rect 17718 15194 17724 15196
rect 13905 15192 17724 15194
rect 13905 15136 13910 15192
rect 13966 15136 17724 15192
rect 13905 15134 17724 15136
rect 13905 15131 13971 15134
rect 17718 15132 17724 15134
rect 17788 15132 17794 15196
rect 22645 15194 22711 15197
rect 23013 15194 23079 15197
rect 22645 15192 23079 15194
rect 22645 15136 22650 15192
rect 22706 15136 23018 15192
rect 23074 15136 23079 15192
rect 22645 15134 23079 15136
rect 22645 15131 22711 15134
rect 23013 15131 23079 15134
rect -300 15058 160 15088
rect 1117 15058 1183 15061
rect 7465 15058 7531 15061
rect 21725 15058 21791 15061
rect 22829 15058 22895 15061
rect -300 15056 1183 15058
rect -300 15000 1122 15056
rect 1178 15000 1183 15056
rect -300 14998 1183 15000
rect -300 14968 160 14998
rect 1117 14995 1183 14998
rect 2730 15056 22895 15058
rect 2730 15000 7470 15056
rect 7526 15000 21730 15056
rect 21786 15000 22834 15056
rect 22890 15000 22895 15056
rect 2730 14998 22895 15000
rect 2262 14860 2268 14924
rect 2332 14922 2338 14924
rect 2730 14922 2790 14998
rect 7465 14995 7531 14998
rect 21725 14995 21791 14998
rect 22829 14995 22895 14998
rect 2332 14862 2790 14922
rect 4153 14922 4219 14925
rect 4981 14922 5047 14925
rect 4153 14920 5047 14922
rect 4153 14864 4158 14920
rect 4214 14864 4986 14920
rect 5042 14864 5047 14920
rect 4153 14862 5047 14864
rect 2332 14860 2338 14862
rect 4153 14859 4219 14862
rect 4981 14859 5047 14862
rect 5574 14860 5580 14924
rect 5644 14922 5650 14924
rect 8293 14922 8359 14925
rect 11513 14922 11579 14925
rect 19701 14922 19767 14925
rect 5644 14920 8359 14922
rect 5644 14864 8298 14920
rect 8354 14864 8359 14920
rect 5644 14862 8359 14864
rect 5644 14860 5650 14862
rect 8293 14859 8359 14862
rect 8526 14920 19767 14922
rect 8526 14864 11518 14920
rect 11574 14864 19706 14920
rect 19762 14864 19767 14920
rect 8526 14862 19767 14864
rect -300 14786 160 14816
rect 1301 14786 1367 14789
rect -300 14784 1367 14786
rect -300 14728 1306 14784
rect 1362 14728 1367 14784
rect -300 14726 1367 14728
rect -300 14696 160 14726
rect 1301 14723 1367 14726
rect 5165 14786 5231 14789
rect 8526 14786 8586 14862
rect 11513 14859 11579 14862
rect 19701 14859 19767 14862
rect 5165 14784 8586 14786
rect 5165 14728 5170 14784
rect 5226 14728 8586 14784
rect 5165 14726 8586 14728
rect 24117 14786 24183 14789
rect 25540 14786 26000 14816
rect 24117 14784 26000 14786
rect 24117 14728 24122 14784
rect 24178 14728 26000 14784
rect 24117 14726 26000 14728
rect 5165 14723 5231 14726
rect 24117 14723 24183 14726
rect 3878 14720 4194 14721
rect 3878 14656 3884 14720
rect 3948 14656 3964 14720
rect 4028 14656 4044 14720
rect 4108 14656 4124 14720
rect 4188 14656 4194 14720
rect 3878 14655 4194 14656
rect 9743 14720 10059 14721
rect 9743 14656 9749 14720
rect 9813 14656 9829 14720
rect 9893 14656 9909 14720
rect 9973 14656 9989 14720
rect 10053 14656 10059 14720
rect 9743 14655 10059 14656
rect 15608 14720 15924 14721
rect 15608 14656 15614 14720
rect 15678 14656 15694 14720
rect 15758 14656 15774 14720
rect 15838 14656 15854 14720
rect 15918 14656 15924 14720
rect 15608 14655 15924 14656
rect 21473 14720 21789 14721
rect 21473 14656 21479 14720
rect 21543 14656 21559 14720
rect 21623 14656 21639 14720
rect 21703 14656 21719 14720
rect 21783 14656 21789 14720
rect 25540 14696 26000 14726
rect 21473 14655 21789 14656
rect -300 14514 160 14544
rect 3969 14514 4035 14517
rect -300 14512 4035 14514
rect -300 14456 3974 14512
rect 4030 14456 4035 14512
rect -300 14454 4035 14456
rect -300 14424 160 14454
rect 3969 14451 4035 14454
rect 8753 14514 8819 14517
rect 16205 14514 16271 14517
rect 16849 14514 16915 14517
rect 8753 14512 16915 14514
rect 8753 14456 8758 14512
rect 8814 14456 16210 14512
rect 16266 14456 16854 14512
rect 16910 14456 16915 14512
rect 8753 14454 16915 14456
rect 8753 14451 8819 14454
rect 16205 14451 16271 14454
rect 16849 14451 16915 14454
rect 1761 14378 1827 14381
rect 2313 14378 2379 14381
rect 4153 14378 4219 14381
rect 1761 14376 4219 14378
rect 1761 14320 1766 14376
rect 1822 14320 2318 14376
rect 2374 14320 4158 14376
rect 4214 14320 4219 14376
rect 1761 14318 4219 14320
rect 1761 14315 1827 14318
rect 2313 14315 2379 14318
rect 4153 14315 4219 14318
rect 6126 14316 6132 14380
rect 6196 14378 6202 14380
rect 10317 14378 10383 14381
rect 6196 14376 10383 14378
rect 6196 14320 10322 14376
rect 10378 14320 10383 14376
rect 6196 14318 10383 14320
rect 6196 14316 6202 14318
rect 10317 14315 10383 14318
rect -300 14242 160 14272
rect 24853 14242 24919 14245
rect 25540 14242 26000 14272
rect -300 14182 1226 14242
rect -300 14152 160 14182
rect -300 13970 160 14000
rect 1166 13970 1226 14182
rect 24853 14240 26000 14242
rect 24853 14184 24858 14240
rect 24914 14184 26000 14240
rect 24853 14182 26000 14184
rect 24853 14179 24919 14182
rect 6810 14176 7126 14177
rect 6810 14112 6816 14176
rect 6880 14112 6896 14176
rect 6960 14112 6976 14176
rect 7040 14112 7056 14176
rect 7120 14112 7126 14176
rect 6810 14111 7126 14112
rect 12675 14176 12991 14177
rect 12675 14112 12681 14176
rect 12745 14112 12761 14176
rect 12825 14112 12841 14176
rect 12905 14112 12921 14176
rect 12985 14112 12991 14176
rect 12675 14111 12991 14112
rect 18540 14176 18856 14177
rect 18540 14112 18546 14176
rect 18610 14112 18626 14176
rect 18690 14112 18706 14176
rect 18770 14112 18786 14176
rect 18850 14112 18856 14176
rect 18540 14111 18856 14112
rect 24405 14176 24721 14177
rect 24405 14112 24411 14176
rect 24475 14112 24491 14176
rect 24555 14112 24571 14176
rect 24635 14112 24651 14176
rect 24715 14112 24721 14176
rect 25540 14152 26000 14182
rect 24405 14111 24721 14112
rect 1577 13970 1643 13973
rect -300 13910 1042 13970
rect 1166 13968 1643 13970
rect 1166 13912 1582 13968
rect 1638 13912 1643 13968
rect 1166 13910 1643 13912
rect -300 13880 160 13910
rect 982 13834 1042 13910
rect 1577 13907 1643 13910
rect 2957 13970 3023 13973
rect 12341 13970 12407 13973
rect 2957 13968 12407 13970
rect 2957 13912 2962 13968
rect 3018 13912 12346 13968
rect 12402 13912 12407 13968
rect 2957 13910 12407 13912
rect 2957 13907 3023 13910
rect 12341 13907 12407 13910
rect 1301 13834 1367 13837
rect 982 13832 1367 13834
rect 982 13776 1306 13832
rect 1362 13776 1367 13832
rect 982 13774 1367 13776
rect 1301 13771 1367 13774
rect 5349 13834 5415 13837
rect 8017 13834 8083 13837
rect 5349 13832 8083 13834
rect 5349 13776 5354 13832
rect 5410 13776 8022 13832
rect 8078 13776 8083 13832
rect 5349 13774 8083 13776
rect 5349 13771 5415 13774
rect 8017 13771 8083 13774
rect 10685 13834 10751 13837
rect 12433 13834 12499 13837
rect 10685 13832 12499 13834
rect 10685 13776 10690 13832
rect 10746 13776 12438 13832
rect 12494 13776 12499 13832
rect 10685 13774 12499 13776
rect 10685 13771 10751 13774
rect 12433 13771 12499 13774
rect 21214 13772 21220 13836
rect 21284 13834 21290 13836
rect 22645 13834 22711 13837
rect 21284 13832 22711 13834
rect 21284 13776 22650 13832
rect 22706 13776 22711 13832
rect 21284 13774 22711 13776
rect 21284 13772 21290 13774
rect 22645 13771 22711 13774
rect -300 13698 160 13728
rect 3601 13698 3667 13701
rect -300 13696 3667 13698
rect -300 13640 3606 13696
rect 3662 13640 3667 13696
rect -300 13638 3667 13640
rect -300 13608 160 13638
rect 3601 13635 3667 13638
rect 24117 13698 24183 13701
rect 25540 13698 26000 13728
rect 24117 13696 26000 13698
rect 24117 13640 24122 13696
rect 24178 13640 26000 13696
rect 24117 13638 26000 13640
rect 24117 13635 24183 13638
rect 3878 13632 4194 13633
rect 3878 13568 3884 13632
rect 3948 13568 3964 13632
rect 4028 13568 4044 13632
rect 4108 13568 4124 13632
rect 4188 13568 4194 13632
rect 3878 13567 4194 13568
rect 9743 13632 10059 13633
rect 9743 13568 9749 13632
rect 9813 13568 9829 13632
rect 9893 13568 9909 13632
rect 9973 13568 9989 13632
rect 10053 13568 10059 13632
rect 9743 13567 10059 13568
rect 15608 13632 15924 13633
rect 15608 13568 15614 13632
rect 15678 13568 15694 13632
rect 15758 13568 15774 13632
rect 15838 13568 15854 13632
rect 15918 13568 15924 13632
rect 15608 13567 15924 13568
rect 21473 13632 21789 13633
rect 21473 13568 21479 13632
rect 21543 13568 21559 13632
rect 21623 13568 21639 13632
rect 21703 13568 21719 13632
rect 21783 13568 21789 13632
rect 25540 13608 26000 13638
rect 21473 13567 21789 13568
rect -300 13426 160 13456
rect 657 13426 723 13429
rect -300 13424 723 13426
rect -300 13368 662 13424
rect 718 13368 723 13424
rect -300 13366 723 13368
rect -300 13336 160 13366
rect 657 13363 723 13366
rect 10501 13426 10567 13429
rect 11605 13426 11671 13429
rect 10501 13424 11671 13426
rect 10501 13368 10506 13424
rect 10562 13368 11610 13424
rect 11666 13368 11671 13424
rect 10501 13366 11671 13368
rect 10501 13363 10567 13366
rect -300 13154 160 13184
rect 10734 13157 10794 13366
rect 11605 13363 11671 13366
rect 20805 13426 20871 13429
rect 22829 13426 22895 13429
rect 20805 13424 22895 13426
rect 20805 13368 20810 13424
rect 20866 13368 22834 13424
rect 22890 13368 22895 13424
rect 20805 13366 22895 13368
rect 20805 13363 20871 13366
rect 22829 13363 22895 13366
rect 1209 13154 1275 13157
rect -300 13152 1275 13154
rect -300 13096 1214 13152
rect 1270 13096 1275 13152
rect -300 13094 1275 13096
rect -300 13064 160 13094
rect 1209 13091 1275 13094
rect 8518 13092 8524 13156
rect 8588 13154 8594 13156
rect 8753 13154 8819 13157
rect 8588 13152 8819 13154
rect 8588 13096 8758 13152
rect 8814 13096 8819 13152
rect 8588 13094 8819 13096
rect 10734 13152 10843 13157
rect 10734 13096 10782 13152
rect 10838 13096 10843 13152
rect 10734 13094 10843 13096
rect 8588 13092 8594 13094
rect 8753 13091 8819 13094
rect 10777 13091 10843 13094
rect 24853 13154 24919 13157
rect 25540 13154 26000 13184
rect 24853 13152 26000 13154
rect 24853 13096 24858 13152
rect 24914 13096 26000 13152
rect 24853 13094 26000 13096
rect 24853 13091 24919 13094
rect 6810 13088 7126 13089
rect 6810 13024 6816 13088
rect 6880 13024 6896 13088
rect 6960 13024 6976 13088
rect 7040 13024 7056 13088
rect 7120 13024 7126 13088
rect 6810 13023 7126 13024
rect 12675 13088 12991 13089
rect 12675 13024 12681 13088
rect 12745 13024 12761 13088
rect 12825 13024 12841 13088
rect 12905 13024 12921 13088
rect 12985 13024 12991 13088
rect 12675 13023 12991 13024
rect 18540 13088 18856 13089
rect 18540 13024 18546 13088
rect 18610 13024 18626 13088
rect 18690 13024 18706 13088
rect 18770 13024 18786 13088
rect 18850 13024 18856 13088
rect 18540 13023 18856 13024
rect 24405 13088 24721 13089
rect 24405 13024 24411 13088
rect 24475 13024 24491 13088
rect 24555 13024 24571 13088
rect 24635 13024 24651 13088
rect 24715 13024 24721 13088
rect 25540 13064 26000 13094
rect 24405 13023 24721 13024
rect -300 12882 160 12912
rect 3601 12882 3667 12885
rect -300 12880 3667 12882
rect -300 12824 3606 12880
rect 3662 12824 3667 12880
rect -300 12822 3667 12824
rect -300 12792 160 12822
rect 3601 12819 3667 12822
rect 9489 12882 9555 12885
rect 21030 12882 21036 12884
rect 9489 12880 21036 12882
rect 9489 12824 9494 12880
rect 9550 12824 21036 12880
rect 9489 12822 21036 12824
rect 9489 12819 9555 12822
rect 21030 12820 21036 12822
rect 21100 12820 21106 12884
rect 12382 12684 12388 12748
rect 12452 12746 12458 12748
rect 13118 12746 13124 12748
rect 12452 12686 13124 12746
rect 12452 12684 12458 12686
rect 13118 12684 13124 12686
rect 13188 12684 13194 12748
rect 19333 12746 19399 12749
rect 22185 12746 22251 12749
rect 19333 12744 22251 12746
rect 19333 12688 19338 12744
rect 19394 12688 22190 12744
rect 22246 12688 22251 12744
rect 19333 12686 22251 12688
rect 19333 12683 19399 12686
rect 22185 12683 22251 12686
rect -300 12610 160 12640
rect 1761 12610 1827 12613
rect 4429 12612 4495 12613
rect 4429 12610 4476 12612
rect -300 12608 1827 12610
rect -300 12552 1766 12608
rect 1822 12552 1827 12608
rect -300 12550 1827 12552
rect 4384 12608 4476 12610
rect 4384 12552 4434 12608
rect 4384 12550 4476 12552
rect -300 12520 160 12550
rect 1761 12547 1827 12550
rect 4429 12548 4476 12550
rect 4540 12548 4546 12612
rect 23933 12610 23999 12613
rect 25540 12610 26000 12640
rect 23933 12608 26000 12610
rect 23933 12552 23938 12608
rect 23994 12552 26000 12608
rect 23933 12550 26000 12552
rect 4429 12547 4495 12548
rect 23933 12547 23999 12550
rect 3878 12544 4194 12545
rect 3878 12480 3884 12544
rect 3948 12480 3964 12544
rect 4028 12480 4044 12544
rect 4108 12480 4124 12544
rect 4188 12480 4194 12544
rect 3878 12479 4194 12480
rect 9743 12544 10059 12545
rect 9743 12480 9749 12544
rect 9813 12480 9829 12544
rect 9893 12480 9909 12544
rect 9973 12480 9989 12544
rect 10053 12480 10059 12544
rect 9743 12479 10059 12480
rect 15608 12544 15924 12545
rect 15608 12480 15614 12544
rect 15678 12480 15694 12544
rect 15758 12480 15774 12544
rect 15838 12480 15854 12544
rect 15918 12480 15924 12544
rect 15608 12479 15924 12480
rect 21473 12544 21789 12545
rect 21473 12480 21479 12544
rect 21543 12480 21559 12544
rect 21623 12480 21639 12544
rect 21703 12480 21719 12544
rect 21783 12480 21789 12544
rect 25540 12520 26000 12550
rect 21473 12479 21789 12480
rect 19425 12474 19491 12477
rect 19558 12474 19564 12476
rect 19425 12472 19564 12474
rect 19425 12416 19430 12472
rect 19486 12416 19564 12472
rect 19425 12414 19564 12416
rect 19425 12411 19491 12414
rect 19558 12412 19564 12414
rect 19628 12412 19634 12476
rect -300 12338 160 12368
rect 3693 12338 3759 12341
rect -300 12336 3759 12338
rect -300 12280 3698 12336
rect 3754 12280 3759 12336
rect -300 12278 3759 12280
rect -300 12248 160 12278
rect 3693 12275 3759 12278
rect 5901 12338 5967 12341
rect 6545 12338 6611 12341
rect 5901 12336 6611 12338
rect 5901 12280 5906 12336
rect 5962 12280 6550 12336
rect 6606 12280 6611 12336
rect 5901 12278 6611 12280
rect 5901 12275 5967 12278
rect 6545 12275 6611 12278
rect 7281 12338 7347 12341
rect 7281 12336 13370 12338
rect 7281 12280 7286 12336
rect 7342 12280 13370 12336
rect 7281 12278 13370 12280
rect 7281 12275 7347 12278
rect 1485 12204 1551 12205
rect 1485 12200 1532 12204
rect 1596 12202 1602 12204
rect 1485 12144 1490 12200
rect 1485 12140 1532 12144
rect 1596 12142 1642 12202
rect 1596 12140 1602 12142
rect 2078 12140 2084 12204
rect 2148 12202 2154 12204
rect 7414 12202 7420 12204
rect 2148 12142 7420 12202
rect 2148 12140 2154 12142
rect 7414 12140 7420 12142
rect 7484 12140 7490 12204
rect 12382 12140 12388 12204
rect 12452 12202 12458 12204
rect 13118 12202 13124 12204
rect 12452 12142 13124 12202
rect 12452 12140 12458 12142
rect 13118 12140 13124 12142
rect 13188 12140 13194 12204
rect 1485 12139 1551 12140
rect -300 12066 160 12096
rect 1301 12066 1367 12069
rect -300 12064 1367 12066
rect -300 12008 1306 12064
rect 1362 12008 1367 12064
rect -300 12006 1367 12008
rect 13310 12066 13370 12278
rect 13854 12276 13860 12340
rect 13924 12338 13930 12340
rect 19977 12338 20043 12341
rect 13924 12336 20043 12338
rect 13924 12280 19982 12336
rect 20038 12280 20043 12336
rect 13924 12278 20043 12280
rect 13924 12276 13930 12278
rect 19977 12275 20043 12278
rect 13537 12202 13603 12205
rect 20161 12202 20227 12205
rect 13537 12200 20227 12202
rect 13537 12144 13542 12200
rect 13598 12144 20166 12200
rect 20222 12144 20227 12200
rect 13537 12142 20227 12144
rect 13537 12139 13603 12142
rect 20161 12139 20227 12142
rect 15653 12066 15719 12069
rect 13310 12064 15719 12066
rect 13310 12008 15658 12064
rect 15714 12008 15719 12064
rect 13310 12006 15719 12008
rect -300 11976 160 12006
rect 1301 12003 1367 12006
rect 15653 12003 15719 12006
rect 19333 12066 19399 12069
rect 19558 12066 19564 12068
rect 19333 12064 19564 12066
rect 19333 12008 19338 12064
rect 19394 12008 19564 12064
rect 19333 12006 19564 12008
rect 19333 12003 19399 12006
rect 19558 12004 19564 12006
rect 19628 12004 19634 12068
rect 24853 12066 24919 12069
rect 25540 12066 26000 12096
rect 24853 12064 26000 12066
rect 24853 12008 24858 12064
rect 24914 12008 26000 12064
rect 24853 12006 26000 12008
rect 24853 12003 24919 12006
rect 6810 12000 7126 12001
rect 6810 11936 6816 12000
rect 6880 11936 6896 12000
rect 6960 11936 6976 12000
rect 7040 11936 7056 12000
rect 7120 11936 7126 12000
rect 6810 11935 7126 11936
rect 12675 12000 12991 12001
rect 12675 11936 12681 12000
rect 12745 11936 12761 12000
rect 12825 11936 12841 12000
rect 12905 11936 12921 12000
rect 12985 11936 12991 12000
rect 12675 11935 12991 11936
rect 18540 12000 18856 12001
rect 18540 11936 18546 12000
rect 18610 11936 18626 12000
rect 18690 11936 18706 12000
rect 18770 11936 18786 12000
rect 18850 11936 18856 12000
rect 18540 11935 18856 11936
rect 24405 12000 24721 12001
rect 24405 11936 24411 12000
rect 24475 11936 24491 12000
rect 24555 11936 24571 12000
rect 24635 11936 24651 12000
rect 24715 11936 24721 12000
rect 25540 11976 26000 12006
rect 24405 11935 24721 11936
rect 381 11930 447 11933
rect 4470 11930 4476 11932
rect 381 11928 4476 11930
rect 381 11872 386 11928
rect 442 11872 4476 11928
rect 381 11870 4476 11872
rect 381 11867 447 11870
rect 4470 11868 4476 11870
rect 4540 11868 4546 11932
rect 11973 11930 12039 11933
rect 11973 11928 12450 11930
rect 11973 11872 11978 11928
rect 12034 11872 12450 11928
rect 11973 11870 12450 11872
rect 11973 11867 12039 11870
rect -300 11794 160 11824
rect 12390 11797 12450 11870
rect 3417 11794 3483 11797
rect -300 11792 3483 11794
rect -300 11736 3422 11792
rect 3478 11736 3483 11792
rect -300 11734 3483 11736
rect 12390 11794 12499 11797
rect 14273 11794 14339 11797
rect 19149 11794 19215 11797
rect 12390 11792 12534 11794
rect 12390 11736 12438 11792
rect 12494 11736 12534 11792
rect 12390 11734 12534 11736
rect 14273 11792 19215 11794
rect 14273 11736 14278 11792
rect 14334 11736 19154 11792
rect 19210 11736 19215 11792
rect 14273 11734 19215 11736
rect -300 11704 160 11734
rect 3417 11731 3483 11734
rect 12433 11731 12499 11734
rect 14273 11731 14339 11734
rect 19149 11731 19215 11734
rect 2313 11658 2379 11661
rect 6821 11658 6887 11661
rect 13854 11658 13860 11660
rect 2313 11656 13860 11658
rect 2313 11600 2318 11656
rect 2374 11600 6826 11656
rect 6882 11600 13860 11656
rect 2313 11598 13860 11600
rect 2313 11595 2379 11598
rect 6821 11595 6887 11598
rect 13854 11596 13860 11598
rect 13924 11596 13930 11660
rect -300 11522 160 11552
rect 1577 11522 1643 11525
rect -300 11520 1643 11522
rect -300 11464 1582 11520
rect 1638 11464 1643 11520
rect -300 11462 1643 11464
rect -300 11432 160 11462
rect 1577 11459 1643 11462
rect 10726 11460 10732 11524
rect 10796 11460 10802 11524
rect 24025 11522 24091 11525
rect 25540 11522 26000 11552
rect 24025 11520 26000 11522
rect 24025 11464 24030 11520
rect 24086 11464 26000 11520
rect 24025 11462 26000 11464
rect 3878 11456 4194 11457
rect 3878 11392 3884 11456
rect 3948 11392 3964 11456
rect 4028 11392 4044 11456
rect 4108 11392 4124 11456
rect 4188 11392 4194 11456
rect 3878 11391 4194 11392
rect 9743 11456 10059 11457
rect 9743 11392 9749 11456
rect 9813 11392 9829 11456
rect 9893 11392 9909 11456
rect 9973 11392 9989 11456
rect 10053 11392 10059 11456
rect 9743 11391 10059 11392
rect 7833 11388 7899 11389
rect 7782 11386 7788 11388
rect 7742 11326 7788 11386
rect 7852 11384 7899 11388
rect 7894 11328 7899 11384
rect 7782 11324 7788 11326
rect 7852 11324 7899 11328
rect 7833 11323 7899 11324
rect -300 11250 160 11280
rect 2957 11250 3023 11253
rect 10734 11250 10794 11460
rect 24025 11459 24091 11462
rect 15608 11456 15924 11457
rect 15608 11392 15614 11456
rect 15678 11392 15694 11456
rect 15758 11392 15774 11456
rect 15838 11392 15854 11456
rect 15918 11392 15924 11456
rect 15608 11391 15924 11392
rect 21473 11456 21789 11457
rect 21473 11392 21479 11456
rect 21543 11392 21559 11456
rect 21623 11392 21639 11456
rect 21703 11392 21719 11456
rect 21783 11392 21789 11456
rect 25540 11432 26000 11462
rect 21473 11391 21789 11392
rect -300 11248 3023 11250
rect -300 11192 2962 11248
rect 3018 11192 3023 11248
rect -300 11190 3023 11192
rect -300 11160 160 11190
rect 2957 11187 3023 11190
rect 5214 11190 10794 11250
rect 12341 11250 12407 11253
rect 13997 11250 14063 11253
rect 12341 11248 14063 11250
rect 12341 11192 12346 11248
rect 12402 11192 14002 11248
rect 14058 11192 14063 11248
rect 12341 11190 14063 11192
rect 2589 11114 2655 11117
rect 5214 11114 5274 11190
rect 12341 11187 12407 11190
rect 13997 11187 14063 11190
rect 2589 11112 5274 11114
rect 2589 11056 2594 11112
rect 2650 11056 5274 11112
rect 2589 11054 5274 11056
rect 2589 11051 2655 11054
rect 5390 11052 5396 11116
rect 5460 11114 5466 11116
rect 5993 11114 6059 11117
rect 5460 11112 6059 11114
rect 5460 11056 5998 11112
rect 6054 11056 6059 11112
rect 5460 11054 6059 11056
rect 5460 11052 5466 11054
rect 5993 11051 6059 11054
rect 7414 11052 7420 11116
rect 7484 11114 7490 11116
rect 8385 11114 8451 11117
rect 7484 11112 8451 11114
rect 7484 11056 8390 11112
rect 8446 11056 8451 11112
rect 7484 11054 8451 11056
rect 7484 11052 7490 11054
rect 8385 11051 8451 11054
rect 10358 11052 10364 11116
rect 10428 11114 10434 11116
rect 11830 11114 11836 11116
rect 10428 11054 11836 11114
rect 10428 11052 10434 11054
rect 11830 11052 11836 11054
rect 11900 11052 11906 11116
rect 13721 11114 13787 11117
rect 14406 11114 14412 11116
rect 13721 11112 14412 11114
rect 13721 11056 13726 11112
rect 13782 11056 14412 11112
rect 13721 11054 14412 11056
rect 13721 11051 13787 11054
rect 14406 11052 14412 11054
rect 14476 11052 14482 11116
rect -300 10978 160 11008
rect 3969 10978 4035 10981
rect -300 10976 4035 10978
rect -300 10920 3974 10976
rect 4030 10920 4035 10976
rect -300 10918 4035 10920
rect -300 10888 160 10918
rect 3969 10915 4035 10918
rect 4153 10978 4219 10981
rect 4286 10978 4292 10980
rect 4153 10976 4292 10978
rect 4153 10920 4158 10976
rect 4214 10920 4292 10976
rect 4153 10918 4292 10920
rect 4153 10915 4219 10918
rect 4286 10916 4292 10918
rect 4356 10916 4362 10980
rect 24853 10978 24919 10981
rect 25540 10978 26000 11008
rect 24853 10976 26000 10978
rect 24853 10920 24858 10976
rect 24914 10920 26000 10976
rect 24853 10918 26000 10920
rect 24853 10915 24919 10918
rect 6810 10912 7126 10913
rect 6810 10848 6816 10912
rect 6880 10848 6896 10912
rect 6960 10848 6976 10912
rect 7040 10848 7056 10912
rect 7120 10848 7126 10912
rect 6810 10847 7126 10848
rect 12675 10912 12991 10913
rect 12675 10848 12681 10912
rect 12745 10848 12761 10912
rect 12825 10848 12841 10912
rect 12905 10848 12921 10912
rect 12985 10848 12991 10912
rect 12675 10847 12991 10848
rect 18540 10912 18856 10913
rect 18540 10848 18546 10912
rect 18610 10848 18626 10912
rect 18690 10848 18706 10912
rect 18770 10848 18786 10912
rect 18850 10848 18856 10912
rect 18540 10847 18856 10848
rect 24405 10912 24721 10913
rect 24405 10848 24411 10912
rect 24475 10848 24491 10912
rect 24555 10848 24571 10912
rect 24635 10848 24651 10912
rect 24715 10848 24721 10912
rect 25540 10888 26000 10918
rect 24405 10847 24721 10848
rect 2865 10842 2931 10845
rect 4889 10842 4955 10845
rect 2865 10840 4955 10842
rect 2865 10784 2870 10840
rect 2926 10784 4894 10840
rect 4950 10784 4955 10840
rect 2865 10782 4955 10784
rect 2865 10779 2931 10782
rect 4889 10779 4955 10782
rect -300 10706 160 10736
rect 3693 10706 3759 10709
rect -300 10704 3759 10706
rect -300 10648 3698 10704
rect 3754 10648 3759 10704
rect -300 10646 3759 10648
rect -300 10616 160 10646
rect 3693 10643 3759 10646
rect 6545 10706 6611 10709
rect 17401 10706 17467 10709
rect 6545 10704 17467 10706
rect 6545 10648 6550 10704
rect 6606 10648 17406 10704
rect 17462 10648 17467 10704
rect 6545 10646 17467 10648
rect 6545 10643 6611 10646
rect 17401 10643 17467 10646
rect 2773 10570 2839 10573
rect 2998 10570 3004 10572
rect 2773 10568 3004 10570
rect 2773 10512 2778 10568
rect 2834 10512 3004 10568
rect 2773 10510 3004 10512
rect 2773 10507 2839 10510
rect 2998 10508 3004 10510
rect 3068 10570 3074 10572
rect 4521 10570 4587 10573
rect 20161 10570 20227 10573
rect 3068 10568 4587 10570
rect 3068 10512 4526 10568
rect 4582 10512 4587 10568
rect 3068 10510 4587 10512
rect 3068 10508 3074 10510
rect 4521 10507 4587 10510
rect 12390 10568 20227 10570
rect 12390 10512 20166 10568
rect 20222 10512 20227 10568
rect 12390 10510 20227 10512
rect -300 10434 160 10464
rect 3601 10434 3667 10437
rect -300 10432 3667 10434
rect -300 10376 3606 10432
rect 3662 10376 3667 10432
rect -300 10374 3667 10376
rect -300 10344 160 10374
rect 3601 10371 3667 10374
rect 3878 10368 4194 10369
rect 3878 10304 3884 10368
rect 3948 10304 3964 10368
rect 4028 10304 4044 10368
rect 4108 10304 4124 10368
rect 4188 10304 4194 10368
rect 3878 10303 4194 10304
rect 9743 10368 10059 10369
rect 9743 10304 9749 10368
rect 9813 10304 9829 10368
rect 9893 10304 9909 10368
rect 9973 10304 9989 10368
rect 10053 10304 10059 10368
rect 9743 10303 10059 10304
rect -300 10162 160 10192
rect 4061 10162 4127 10165
rect -300 10160 4127 10162
rect -300 10104 4066 10160
rect 4122 10104 4127 10160
rect -300 10102 4127 10104
rect -300 10072 160 10102
rect 4061 10099 4127 10102
rect 1853 10026 1919 10029
rect 12390 10026 12450 10510
rect 20161 10507 20227 10510
rect 25129 10434 25195 10437
rect 25540 10434 26000 10464
rect 25129 10432 26000 10434
rect 25129 10376 25134 10432
rect 25190 10376 26000 10432
rect 25129 10374 26000 10376
rect 25129 10371 25195 10374
rect 15608 10368 15924 10369
rect 15608 10304 15614 10368
rect 15678 10304 15694 10368
rect 15758 10304 15774 10368
rect 15838 10304 15854 10368
rect 15918 10304 15924 10368
rect 15608 10303 15924 10304
rect 21473 10368 21789 10369
rect 21473 10304 21479 10368
rect 21543 10304 21559 10368
rect 21623 10304 21639 10368
rect 21703 10304 21719 10368
rect 21783 10304 21789 10368
rect 25540 10344 26000 10374
rect 21473 10303 21789 10304
rect 14733 10162 14799 10165
rect 15193 10162 15259 10165
rect 14733 10160 15259 10162
rect 14733 10104 14738 10160
rect 14794 10104 15198 10160
rect 15254 10104 15259 10160
rect 14733 10102 15259 10104
rect 14733 10099 14799 10102
rect 15193 10099 15259 10102
rect 17033 10162 17099 10165
rect 22686 10162 22692 10164
rect 17033 10160 22692 10162
rect 17033 10104 17038 10160
rect 17094 10104 22692 10160
rect 17033 10102 22692 10104
rect 17033 10099 17099 10102
rect 22686 10100 22692 10102
rect 22756 10100 22762 10164
rect 14365 10026 14431 10029
rect 1853 10024 12450 10026
rect 1853 9968 1858 10024
rect 1914 9968 12450 10024
rect 1853 9966 12450 9968
rect 12528 10024 14431 10026
rect 12528 9968 14370 10024
rect 14426 9968 14431 10024
rect 12528 9966 14431 9968
rect 1853 9963 1919 9966
rect -300 9890 160 9920
rect 2865 9890 2931 9893
rect -300 9888 2931 9890
rect -300 9832 2870 9888
rect 2926 9832 2931 9888
rect -300 9830 2931 9832
rect -300 9800 160 9830
rect 2865 9827 2931 9830
rect 3693 9890 3759 9893
rect 5022 9890 5028 9892
rect 3693 9888 5028 9890
rect 3693 9832 3698 9888
rect 3754 9832 5028 9888
rect 3693 9830 5028 9832
rect 3693 9827 3759 9830
rect 5022 9828 5028 9830
rect 5092 9828 5098 9892
rect 11789 9890 11855 9893
rect 12528 9890 12588 9966
rect 14365 9963 14431 9966
rect 14641 10026 14707 10029
rect 15745 10026 15811 10029
rect 14641 10024 15811 10026
rect 14641 9968 14646 10024
rect 14702 9968 15750 10024
rect 15806 9968 15811 10024
rect 14641 9966 15811 9968
rect 14641 9963 14707 9966
rect 15745 9963 15811 9966
rect 11789 9888 12588 9890
rect 11789 9832 11794 9888
rect 11850 9832 12588 9888
rect 11789 9830 12588 9832
rect 24853 9890 24919 9893
rect 25540 9890 26000 9920
rect 24853 9888 26000 9890
rect 24853 9832 24858 9888
rect 24914 9832 26000 9888
rect 24853 9830 26000 9832
rect 11789 9827 11855 9830
rect 24853 9827 24919 9830
rect 6810 9824 7126 9825
rect 6810 9760 6816 9824
rect 6880 9760 6896 9824
rect 6960 9760 6976 9824
rect 7040 9760 7056 9824
rect 7120 9760 7126 9824
rect 6810 9759 7126 9760
rect 12675 9824 12991 9825
rect 12675 9760 12681 9824
rect 12745 9760 12761 9824
rect 12825 9760 12841 9824
rect 12905 9760 12921 9824
rect 12985 9760 12991 9824
rect 12675 9759 12991 9760
rect 18540 9824 18856 9825
rect 18540 9760 18546 9824
rect 18610 9760 18626 9824
rect 18690 9760 18706 9824
rect 18770 9760 18786 9824
rect 18850 9760 18856 9824
rect 18540 9759 18856 9760
rect 24405 9824 24721 9825
rect 24405 9760 24411 9824
rect 24475 9760 24491 9824
rect 24555 9760 24571 9824
rect 24635 9760 24651 9824
rect 24715 9760 24721 9824
rect 25540 9800 26000 9830
rect 24405 9759 24721 9760
rect 8150 9692 8156 9756
rect 8220 9754 8226 9756
rect 9254 9754 9260 9756
rect 8220 9694 9260 9754
rect 8220 9692 8226 9694
rect 9254 9692 9260 9694
rect 9324 9692 9330 9756
rect 14549 9754 14615 9757
rect 15837 9754 15903 9757
rect 14549 9752 15903 9754
rect 14549 9696 14554 9752
rect 14610 9696 15842 9752
rect 15898 9696 15903 9752
rect 14549 9694 15903 9696
rect 14549 9691 14615 9694
rect 15837 9691 15903 9694
rect -300 9618 160 9648
rect 4061 9618 4127 9621
rect 4337 9620 4403 9621
rect 4286 9618 4292 9620
rect -300 9616 4127 9618
rect -300 9560 4066 9616
rect 4122 9560 4127 9616
rect -300 9558 4127 9560
rect 4246 9558 4292 9618
rect 4356 9616 4403 9620
rect 4398 9560 4403 9616
rect -300 9528 160 9558
rect 4061 9555 4127 9558
rect 4286 9556 4292 9558
rect 4356 9556 4403 9560
rect 4337 9555 4403 9556
rect 12157 9618 12223 9621
rect 17309 9618 17375 9621
rect 12157 9616 17375 9618
rect 12157 9560 12162 9616
rect 12218 9560 17314 9616
rect 17370 9560 17375 9616
rect 12157 9558 17375 9560
rect 12157 9555 12223 9558
rect 17309 9555 17375 9558
rect 4797 9482 4863 9485
rect 2730 9480 4863 9482
rect 2730 9424 4802 9480
rect 4858 9424 4863 9480
rect 2730 9422 4863 9424
rect -300 9346 160 9376
rect 2730 9346 2790 9422
rect 4797 9419 4863 9422
rect 11053 9482 11119 9485
rect 18505 9482 18571 9485
rect 11053 9480 18571 9482
rect 11053 9424 11058 9480
rect 11114 9424 18510 9480
rect 18566 9424 18571 9480
rect 11053 9422 18571 9424
rect 11053 9419 11119 9422
rect 18505 9419 18571 9422
rect -300 9286 2790 9346
rect 24117 9346 24183 9349
rect 25540 9346 26000 9376
rect 24117 9344 26000 9346
rect 24117 9288 24122 9344
rect 24178 9288 26000 9344
rect 24117 9286 26000 9288
rect -300 9256 160 9286
rect 24117 9283 24183 9286
rect 3878 9280 4194 9281
rect 3878 9216 3884 9280
rect 3948 9216 3964 9280
rect 4028 9216 4044 9280
rect 4108 9216 4124 9280
rect 4188 9216 4194 9280
rect 3878 9215 4194 9216
rect 9743 9280 10059 9281
rect 9743 9216 9749 9280
rect 9813 9216 9829 9280
rect 9893 9216 9909 9280
rect 9973 9216 9989 9280
rect 10053 9216 10059 9280
rect 9743 9215 10059 9216
rect 15608 9280 15924 9281
rect 15608 9216 15614 9280
rect 15678 9216 15694 9280
rect 15758 9216 15774 9280
rect 15838 9216 15854 9280
rect 15918 9216 15924 9280
rect 15608 9215 15924 9216
rect 21473 9280 21789 9281
rect 21473 9216 21479 9280
rect 21543 9216 21559 9280
rect 21623 9216 21639 9280
rect 21703 9216 21719 9280
rect 21783 9216 21789 9280
rect 25540 9256 26000 9286
rect 21473 9215 21789 9216
rect -300 9074 160 9104
rect 4286 9074 4292 9076
rect -300 9014 4292 9074
rect -300 8984 160 9014
rect 4286 9012 4292 9014
rect 4356 9012 4362 9076
rect 11237 9074 11303 9077
rect 15101 9074 15167 9077
rect 11237 9072 15167 9074
rect 11237 9016 11242 9072
rect 11298 9016 15106 9072
rect 15162 9016 15167 9072
rect 11237 9014 15167 9016
rect 11237 9011 11303 9014
rect 15101 9011 15167 9014
rect 19333 9074 19399 9077
rect 20253 9074 20319 9077
rect 19333 9072 20319 9074
rect 19333 9016 19338 9072
rect 19394 9016 20258 9072
rect 20314 9016 20319 9072
rect 19333 9014 20319 9016
rect 19333 9011 19399 9014
rect 20253 9011 20319 9014
rect 3417 8938 3483 8941
rect 5441 8938 5507 8941
rect 3417 8936 5507 8938
rect 3417 8880 3422 8936
rect 3478 8880 5446 8936
rect 5502 8880 5507 8936
rect 3417 8878 5507 8880
rect 3417 8875 3483 8878
rect 5441 8875 5507 8878
rect 8702 8876 8708 8940
rect 8772 8938 8778 8940
rect 11145 8938 11211 8941
rect 8772 8936 11211 8938
rect 8772 8880 11150 8936
rect 11206 8880 11211 8936
rect 8772 8878 11211 8880
rect 8772 8876 8778 8878
rect 11145 8875 11211 8878
rect 18045 8938 18111 8941
rect 18965 8938 19031 8941
rect 18045 8936 19031 8938
rect 18045 8880 18050 8936
rect 18106 8880 18970 8936
rect 19026 8880 19031 8936
rect 18045 8878 19031 8880
rect 18045 8875 18111 8878
rect 18965 8875 19031 8878
rect 23565 8938 23631 8941
rect 23565 8936 24962 8938
rect 23565 8880 23570 8936
rect 23626 8880 24962 8936
rect 23565 8878 24962 8880
rect 23565 8875 23631 8878
rect -300 8802 160 8832
rect 3509 8802 3575 8805
rect -300 8800 3575 8802
rect -300 8744 3514 8800
rect 3570 8744 3575 8800
rect -300 8742 3575 8744
rect -300 8712 160 8742
rect 3509 8739 3575 8742
rect 20713 8802 20779 8805
rect 23381 8802 23447 8805
rect 20713 8800 23447 8802
rect 20713 8744 20718 8800
rect 20774 8744 23386 8800
rect 23442 8744 23447 8800
rect 20713 8742 23447 8744
rect 24902 8802 24962 8878
rect 25540 8802 26000 8832
rect 24902 8742 26000 8802
rect 20713 8739 20779 8742
rect 23381 8739 23447 8742
rect 6810 8736 7126 8737
rect 6810 8672 6816 8736
rect 6880 8672 6896 8736
rect 6960 8672 6976 8736
rect 7040 8672 7056 8736
rect 7120 8672 7126 8736
rect 6810 8671 7126 8672
rect 12675 8736 12991 8737
rect 12675 8672 12681 8736
rect 12745 8672 12761 8736
rect 12825 8672 12841 8736
rect 12905 8672 12921 8736
rect 12985 8672 12991 8736
rect 12675 8671 12991 8672
rect 18540 8736 18856 8737
rect 18540 8672 18546 8736
rect 18610 8672 18626 8736
rect 18690 8672 18706 8736
rect 18770 8672 18786 8736
rect 18850 8672 18856 8736
rect 18540 8671 18856 8672
rect 24405 8736 24721 8737
rect 24405 8672 24411 8736
rect 24475 8672 24491 8736
rect 24555 8672 24571 8736
rect 24635 8672 24651 8736
rect 24715 8672 24721 8736
rect 25540 8712 26000 8742
rect 24405 8671 24721 8672
rect 2129 8666 2195 8669
rect 5165 8666 5231 8669
rect 2129 8664 5231 8666
rect 2129 8608 2134 8664
rect 2190 8608 5170 8664
rect 5226 8608 5231 8664
rect 2129 8606 5231 8608
rect 2129 8603 2195 8606
rect 5165 8603 5231 8606
rect -300 8530 160 8560
rect 1945 8530 2011 8533
rect -300 8528 2011 8530
rect -300 8472 1950 8528
rect 2006 8472 2011 8528
rect -300 8470 2011 8472
rect -300 8440 160 8470
rect 1945 8467 2011 8470
rect 2814 8468 2820 8532
rect 2884 8530 2890 8532
rect 3233 8530 3299 8533
rect 2884 8528 3299 8530
rect 2884 8472 3238 8528
rect 3294 8472 3299 8528
rect 2884 8470 3299 8472
rect 2884 8468 2890 8470
rect 3233 8467 3299 8470
rect 5993 8530 6059 8533
rect 7649 8530 7715 8533
rect 5993 8528 7715 8530
rect 5993 8472 5998 8528
rect 6054 8472 7654 8528
rect 7710 8472 7715 8528
rect 5993 8470 7715 8472
rect 5993 8467 6059 8470
rect 7649 8467 7715 8470
rect 18965 8530 19031 8533
rect 19742 8530 19748 8532
rect 18965 8528 19748 8530
rect 18965 8472 18970 8528
rect 19026 8472 19748 8528
rect 18965 8470 19748 8472
rect 18965 8467 19031 8470
rect 19742 8468 19748 8470
rect 19812 8468 19818 8532
rect 1485 8394 1551 8397
rect 3182 8394 3188 8396
rect 1485 8392 3188 8394
rect 1485 8336 1490 8392
rect 1546 8336 3188 8392
rect 1485 8334 3188 8336
rect 1485 8331 1551 8334
rect 3182 8332 3188 8334
rect 3252 8394 3258 8396
rect 3734 8394 3740 8396
rect 3252 8334 3740 8394
rect 3252 8332 3258 8334
rect 3734 8332 3740 8334
rect 3804 8394 3810 8396
rect 3877 8394 3943 8397
rect 3804 8392 3943 8394
rect 3804 8336 3882 8392
rect 3938 8336 3943 8392
rect 3804 8334 3943 8336
rect 3804 8332 3810 8334
rect 3877 8331 3943 8334
rect 14365 8394 14431 8397
rect 19517 8396 19583 8397
rect 17902 8394 17908 8396
rect 14365 8392 17908 8394
rect 14365 8336 14370 8392
rect 14426 8336 17908 8392
rect 14365 8334 17908 8336
rect 14365 8331 14431 8334
rect 17902 8332 17908 8334
rect 17972 8332 17978 8396
rect 19517 8394 19564 8396
rect 19472 8392 19564 8394
rect 19472 8336 19522 8392
rect 19472 8334 19564 8336
rect 19517 8332 19564 8334
rect 19628 8332 19634 8396
rect 19926 8332 19932 8396
rect 19996 8394 20002 8396
rect 20846 8394 20852 8396
rect 19996 8334 20852 8394
rect 19996 8332 20002 8334
rect 20846 8332 20852 8334
rect 20916 8332 20922 8396
rect 19517 8331 19583 8332
rect -300 8258 160 8288
rect 3049 8258 3115 8261
rect -300 8256 3115 8258
rect -300 8200 3054 8256
rect 3110 8200 3115 8256
rect -300 8198 3115 8200
rect -300 8168 160 8198
rect 3049 8195 3115 8198
rect 24209 8258 24275 8261
rect 25540 8258 26000 8288
rect 24209 8256 26000 8258
rect 24209 8200 24214 8256
rect 24270 8200 26000 8256
rect 24209 8198 26000 8200
rect 24209 8195 24275 8198
rect 3878 8192 4194 8193
rect 3878 8128 3884 8192
rect 3948 8128 3964 8192
rect 4028 8128 4044 8192
rect 4108 8128 4124 8192
rect 4188 8128 4194 8192
rect 3878 8127 4194 8128
rect 9743 8192 10059 8193
rect 9743 8128 9749 8192
rect 9813 8128 9829 8192
rect 9893 8128 9909 8192
rect 9973 8128 9989 8192
rect 10053 8128 10059 8192
rect 9743 8127 10059 8128
rect 15608 8192 15924 8193
rect 15608 8128 15614 8192
rect 15678 8128 15694 8192
rect 15758 8128 15774 8192
rect 15838 8128 15854 8192
rect 15918 8128 15924 8192
rect 15608 8127 15924 8128
rect 21473 8192 21789 8193
rect 21473 8128 21479 8192
rect 21543 8128 21559 8192
rect 21623 8128 21639 8192
rect 21703 8128 21719 8192
rect 21783 8128 21789 8192
rect 25540 8168 26000 8198
rect 21473 8127 21789 8128
rect -300 7986 160 8016
rect 1853 7986 1919 7989
rect -300 7984 1919 7986
rect -300 7928 1858 7984
rect 1914 7928 1919 7984
rect -300 7926 1919 7928
rect -300 7896 160 7926
rect 1853 7923 1919 7926
rect 3601 7986 3667 7989
rect 5717 7986 5783 7989
rect 3601 7984 5783 7986
rect 3601 7928 3606 7984
rect 3662 7928 5722 7984
rect 5778 7928 5783 7984
rect 3601 7926 5783 7928
rect 3601 7923 3667 7926
rect 5717 7923 5783 7926
rect 7649 7986 7715 7989
rect 9765 7986 9831 7989
rect 7649 7984 9831 7986
rect 7649 7928 7654 7984
rect 7710 7928 9770 7984
rect 9826 7928 9831 7984
rect 7649 7926 9831 7928
rect 7649 7923 7715 7926
rect 9765 7923 9831 7926
rect 2865 7850 2931 7853
rect 3366 7850 3372 7852
rect 2865 7848 3372 7850
rect 2865 7792 2870 7848
rect 2926 7792 3372 7848
rect 2865 7790 3372 7792
rect 2865 7787 2931 7790
rect 3366 7788 3372 7790
rect 3436 7850 3442 7852
rect 4061 7850 4127 7853
rect 3436 7848 4127 7850
rect 3436 7792 4066 7848
rect 4122 7792 4127 7848
rect 3436 7790 4127 7792
rect 3436 7788 3442 7790
rect 4061 7787 4127 7790
rect 24025 7850 24091 7853
rect 24025 7848 24962 7850
rect 24025 7792 24030 7848
rect 24086 7792 24962 7848
rect 24025 7790 24962 7792
rect 24025 7787 24091 7790
rect -300 7714 160 7744
rect 4061 7714 4127 7717
rect -300 7712 4127 7714
rect -300 7656 4066 7712
rect 4122 7656 4127 7712
rect -300 7654 4127 7656
rect 24902 7714 24962 7790
rect 25540 7714 26000 7744
rect 24902 7654 26000 7714
rect -300 7624 160 7654
rect 4061 7651 4127 7654
rect 6810 7648 7126 7649
rect 6810 7584 6816 7648
rect 6880 7584 6896 7648
rect 6960 7584 6976 7648
rect 7040 7584 7056 7648
rect 7120 7584 7126 7648
rect 6810 7583 7126 7584
rect 12675 7648 12991 7649
rect 12675 7584 12681 7648
rect 12745 7584 12761 7648
rect 12825 7584 12841 7648
rect 12905 7584 12921 7648
rect 12985 7584 12991 7648
rect 12675 7583 12991 7584
rect 18540 7648 18856 7649
rect 18540 7584 18546 7648
rect 18610 7584 18626 7648
rect 18690 7584 18706 7648
rect 18770 7584 18786 7648
rect 18850 7584 18856 7648
rect 18540 7583 18856 7584
rect 24405 7648 24721 7649
rect 24405 7584 24411 7648
rect 24475 7584 24491 7648
rect 24555 7584 24571 7648
rect 24635 7584 24651 7648
rect 24715 7584 24721 7648
rect 25540 7624 26000 7654
rect 24405 7583 24721 7584
rect 20713 7578 20779 7581
rect 24025 7578 24091 7581
rect 20713 7576 24091 7578
rect 20713 7520 20718 7576
rect 20774 7520 24030 7576
rect 24086 7520 24091 7576
rect 20713 7518 24091 7520
rect 20713 7515 20779 7518
rect 24025 7515 24091 7518
rect -300 7442 160 7472
rect 4061 7442 4127 7445
rect -300 7440 4127 7442
rect -300 7384 4066 7440
rect 4122 7384 4127 7440
rect -300 7382 4127 7384
rect -300 7352 160 7382
rect 4061 7379 4127 7382
rect 3141 7306 3207 7309
rect 7557 7306 7623 7309
rect 3141 7304 7623 7306
rect 3141 7248 3146 7304
rect 3202 7248 7562 7304
rect 7618 7248 7623 7304
rect 3141 7246 7623 7248
rect 3141 7243 3207 7246
rect 7557 7243 7623 7246
rect -300 7170 160 7200
rect 3509 7170 3575 7173
rect -300 7168 3575 7170
rect -300 7112 3514 7168
rect 3570 7112 3575 7168
rect -300 7110 3575 7112
rect -300 7080 160 7110
rect 3509 7107 3575 7110
rect 24025 7170 24091 7173
rect 25540 7170 26000 7200
rect 24025 7168 26000 7170
rect 24025 7112 24030 7168
rect 24086 7112 26000 7168
rect 24025 7110 26000 7112
rect 24025 7107 24091 7110
rect 3878 7104 4194 7105
rect 3878 7040 3884 7104
rect 3948 7040 3964 7104
rect 4028 7040 4044 7104
rect 4108 7040 4124 7104
rect 4188 7040 4194 7104
rect 3878 7039 4194 7040
rect 9743 7104 10059 7105
rect 9743 7040 9749 7104
rect 9813 7040 9829 7104
rect 9893 7040 9909 7104
rect 9973 7040 9989 7104
rect 10053 7040 10059 7104
rect 9743 7039 10059 7040
rect 15608 7104 15924 7105
rect 15608 7040 15614 7104
rect 15678 7040 15694 7104
rect 15758 7040 15774 7104
rect 15838 7040 15854 7104
rect 15918 7040 15924 7104
rect 15608 7039 15924 7040
rect 21473 7104 21789 7105
rect 21473 7040 21479 7104
rect 21543 7040 21559 7104
rect 21623 7040 21639 7104
rect 21703 7040 21719 7104
rect 21783 7040 21789 7104
rect 25540 7080 26000 7110
rect 21473 7039 21789 7040
rect -300 6898 160 6928
rect 4705 6898 4771 6901
rect 15929 6898 15995 6901
rect -300 6896 4771 6898
rect -300 6840 4710 6896
rect 4766 6840 4771 6896
rect -300 6838 4771 6840
rect -300 6808 160 6838
rect 4705 6835 4771 6838
rect 7606 6896 15995 6898
rect 7606 6840 15934 6896
rect 15990 6840 15995 6896
rect 7606 6838 15995 6840
rect 1485 6762 1551 6765
rect 7606 6762 7666 6838
rect 15929 6835 15995 6838
rect 23841 6898 23907 6901
rect 23841 6896 24226 6898
rect 23841 6840 23846 6896
rect 23902 6840 24226 6896
rect 23841 6838 24226 6840
rect 23841 6835 23907 6838
rect 1485 6760 7666 6762
rect 1485 6704 1490 6760
rect 1546 6704 7666 6760
rect 1485 6702 7666 6704
rect 9673 6762 9739 6765
rect 12801 6762 12867 6765
rect 9673 6760 12867 6762
rect 9673 6704 9678 6760
rect 9734 6704 12806 6760
rect 12862 6704 12867 6760
rect 9673 6702 12867 6704
rect 1485 6699 1551 6702
rect 9673 6699 9739 6702
rect 12801 6699 12867 6702
rect -300 6626 160 6656
rect 2865 6626 2931 6629
rect -300 6624 2931 6626
rect -300 6568 2870 6624
rect 2926 6568 2931 6624
rect -300 6566 2931 6568
rect -300 6536 160 6566
rect 2865 6563 2931 6566
rect 10225 6626 10291 6629
rect 12433 6626 12499 6629
rect 10225 6624 12499 6626
rect 10225 6568 10230 6624
rect 10286 6568 12438 6624
rect 12494 6568 12499 6624
rect 10225 6566 12499 6568
rect 10225 6563 10291 6566
rect 12433 6563 12499 6566
rect 20805 6626 20871 6629
rect 21081 6626 21147 6629
rect 20805 6624 21147 6626
rect 20805 6568 20810 6624
rect 20866 6568 21086 6624
rect 21142 6568 21147 6624
rect 20805 6566 21147 6568
rect 20805 6563 20871 6566
rect 21081 6563 21147 6566
rect 6810 6560 7126 6561
rect 6810 6496 6816 6560
rect 6880 6496 6896 6560
rect 6960 6496 6976 6560
rect 7040 6496 7056 6560
rect 7120 6496 7126 6560
rect 6810 6495 7126 6496
rect 12675 6560 12991 6561
rect 12675 6496 12681 6560
rect 12745 6496 12761 6560
rect 12825 6496 12841 6560
rect 12905 6496 12921 6560
rect 12985 6496 12991 6560
rect 12675 6495 12991 6496
rect 18540 6560 18856 6561
rect 18540 6496 18546 6560
rect 18610 6496 18626 6560
rect 18690 6496 18706 6560
rect 18770 6496 18786 6560
rect 18850 6496 18856 6560
rect 18540 6495 18856 6496
rect 2262 6428 2268 6492
rect 2332 6490 2338 6492
rect 2589 6490 2655 6493
rect 2332 6488 2655 6490
rect 2332 6432 2594 6488
rect 2650 6432 2655 6488
rect 2332 6430 2655 6432
rect 2332 6428 2338 6430
rect 2589 6427 2655 6430
rect -300 6354 160 6384
rect 2589 6354 2655 6357
rect -300 6352 2655 6354
rect -300 6296 2594 6352
rect 2650 6296 2655 6352
rect -300 6294 2655 6296
rect -300 6264 160 6294
rect 2589 6291 2655 6294
rect 9121 6354 9187 6357
rect 13353 6354 13419 6357
rect 9121 6352 13419 6354
rect 9121 6296 9126 6352
rect 9182 6296 13358 6352
rect 13414 6296 13419 6352
rect 9121 6294 13419 6296
rect 9121 6291 9187 6294
rect 13353 6291 13419 6294
rect 3233 6218 3299 6221
rect 3417 6218 3483 6221
rect 9121 6218 9187 6221
rect 3233 6216 9187 6218
rect 3233 6160 3238 6216
rect 3294 6160 3422 6216
rect 3478 6160 9126 6216
rect 9182 6160 9187 6216
rect 3233 6158 9187 6160
rect 3233 6155 3299 6158
rect 3417 6155 3483 6158
rect 9121 6155 9187 6158
rect 19241 6218 19307 6221
rect 21541 6218 21607 6221
rect 19241 6216 21607 6218
rect 19241 6160 19246 6216
rect 19302 6160 21546 6216
rect 21602 6160 21607 6216
rect 19241 6158 21607 6160
rect 19241 6155 19307 6158
rect 21541 6155 21607 6158
rect -300 6082 160 6112
rect 3233 6082 3299 6085
rect -300 6080 3299 6082
rect -300 6024 3238 6080
rect 3294 6024 3299 6080
rect -300 6022 3299 6024
rect 24166 6082 24226 6838
rect 24853 6626 24919 6629
rect 25540 6626 26000 6656
rect 24853 6624 26000 6626
rect 24853 6568 24858 6624
rect 24914 6568 26000 6624
rect 24853 6566 26000 6568
rect 24853 6563 24919 6566
rect 24405 6560 24721 6561
rect 24405 6496 24411 6560
rect 24475 6496 24491 6560
rect 24555 6496 24571 6560
rect 24635 6496 24651 6560
rect 24715 6496 24721 6560
rect 25540 6536 26000 6566
rect 24405 6495 24721 6496
rect 25540 6082 26000 6112
rect 24166 6022 26000 6082
rect -300 5992 160 6022
rect 3233 6019 3299 6022
rect 3878 6016 4194 6017
rect 3878 5952 3884 6016
rect 3948 5952 3964 6016
rect 4028 5952 4044 6016
rect 4108 5952 4124 6016
rect 4188 5952 4194 6016
rect 3878 5951 4194 5952
rect 9743 6016 10059 6017
rect 9743 5952 9749 6016
rect 9813 5952 9829 6016
rect 9893 5952 9909 6016
rect 9973 5952 9989 6016
rect 10053 5952 10059 6016
rect 9743 5951 10059 5952
rect 15608 6016 15924 6017
rect 15608 5952 15614 6016
rect 15678 5952 15694 6016
rect 15758 5952 15774 6016
rect 15838 5952 15854 6016
rect 15918 5952 15924 6016
rect 15608 5951 15924 5952
rect 21473 6016 21789 6017
rect 21473 5952 21479 6016
rect 21543 5952 21559 6016
rect 21623 5952 21639 6016
rect 21703 5952 21719 6016
rect 21783 5952 21789 6016
rect 25540 5992 26000 6022
rect 21473 5951 21789 5952
rect -300 5810 160 5840
rect 2773 5810 2839 5813
rect -300 5808 2839 5810
rect -300 5752 2778 5808
rect 2834 5752 2839 5808
rect -300 5750 2839 5752
rect -300 5720 160 5750
rect 2773 5747 2839 5750
rect 17493 5810 17559 5813
rect 22461 5810 22527 5813
rect 17493 5808 22527 5810
rect 17493 5752 17498 5808
rect 17554 5752 22466 5808
rect 22522 5752 22527 5808
rect 17493 5750 22527 5752
rect 17493 5747 17559 5750
rect 22461 5747 22527 5750
rect 3734 5612 3740 5676
rect 3804 5674 3810 5676
rect 4061 5674 4127 5677
rect 23841 5674 23907 5677
rect 3804 5672 23907 5674
rect 3804 5616 4066 5672
rect 4122 5616 23846 5672
rect 23902 5616 23907 5672
rect 3804 5614 23907 5616
rect 3804 5612 3810 5614
rect 4061 5611 4127 5614
rect 23841 5611 23907 5614
rect -300 5538 160 5568
rect 1669 5538 1735 5541
rect 11605 5540 11671 5541
rect 1894 5538 1900 5540
rect -300 5478 1042 5538
rect -300 5448 160 5478
rect 982 5402 1042 5478
rect 1669 5536 1900 5538
rect 1669 5480 1674 5536
rect 1730 5480 1900 5536
rect 1669 5478 1900 5480
rect 1669 5475 1735 5478
rect 1894 5476 1900 5478
rect 1964 5476 1970 5540
rect 11605 5536 11652 5540
rect 11716 5538 11722 5540
rect 17401 5538 17467 5541
rect 18270 5538 18276 5540
rect 11605 5480 11610 5536
rect 11605 5476 11652 5480
rect 11716 5478 11762 5538
rect 17401 5536 18276 5538
rect 17401 5480 17406 5536
rect 17462 5480 18276 5536
rect 17401 5478 18276 5480
rect 11716 5476 11722 5478
rect 11605 5475 11671 5476
rect 17401 5475 17467 5478
rect 18270 5476 18276 5478
rect 18340 5476 18346 5540
rect 23105 5538 23171 5541
rect 23381 5538 23447 5541
rect 25540 5538 26000 5568
rect 23105 5536 23306 5538
rect 23105 5480 23110 5536
rect 23166 5480 23306 5536
rect 23105 5478 23306 5480
rect 23105 5475 23171 5478
rect 6810 5472 7126 5473
rect 6810 5408 6816 5472
rect 6880 5408 6896 5472
rect 6960 5408 6976 5472
rect 7040 5408 7056 5472
rect 7120 5408 7126 5472
rect 6810 5407 7126 5408
rect 12675 5472 12991 5473
rect 12675 5408 12681 5472
rect 12745 5408 12761 5472
rect 12825 5408 12841 5472
rect 12905 5408 12921 5472
rect 12985 5408 12991 5472
rect 12675 5407 12991 5408
rect 18540 5472 18856 5473
rect 18540 5408 18546 5472
rect 18610 5408 18626 5472
rect 18690 5408 18706 5472
rect 18770 5408 18786 5472
rect 18850 5408 18856 5472
rect 18540 5407 18856 5408
rect 1761 5402 1827 5405
rect 982 5400 1827 5402
rect 982 5344 1766 5400
rect 1822 5344 1827 5400
rect 982 5342 1827 5344
rect 1761 5339 1827 5342
rect 19517 5402 19583 5405
rect 20345 5402 20411 5405
rect 19517 5400 20411 5402
rect 19517 5344 19522 5400
rect 19578 5344 20350 5400
rect 20406 5344 20411 5400
rect 19517 5342 20411 5344
rect 19517 5339 19583 5342
rect 20345 5339 20411 5342
rect 22185 5402 22251 5405
rect 22318 5402 22324 5404
rect 22185 5400 22324 5402
rect 22185 5344 22190 5400
rect 22246 5344 22324 5400
rect 22185 5342 22324 5344
rect 22185 5339 22251 5342
rect 22318 5340 22324 5342
rect 22388 5340 22394 5404
rect -300 5266 160 5296
rect 3693 5266 3759 5269
rect 8937 5266 9003 5269
rect -300 5264 3759 5266
rect -300 5208 3698 5264
rect 3754 5208 3759 5264
rect -300 5206 3759 5208
rect -300 5176 160 5206
rect 3693 5203 3759 5206
rect 4892 5264 9003 5266
rect 4892 5208 8942 5264
rect 8998 5208 9003 5264
rect 4892 5206 9003 5208
rect 2405 5130 2471 5133
rect 4892 5130 4952 5206
rect 8937 5203 9003 5206
rect 19425 5266 19491 5269
rect 19793 5266 19859 5269
rect 19425 5264 19859 5266
rect 19425 5208 19430 5264
rect 19486 5208 19798 5264
rect 19854 5208 19859 5264
rect 19425 5206 19859 5208
rect 19425 5203 19491 5206
rect 19793 5203 19859 5206
rect 2405 5128 4952 5130
rect 2405 5072 2410 5128
rect 2466 5072 4952 5128
rect 2405 5070 4952 5072
rect 5073 5130 5139 5133
rect 16614 5130 16620 5132
rect 5073 5128 16620 5130
rect 5073 5072 5078 5128
rect 5134 5072 16620 5128
rect 5073 5070 16620 5072
rect 2405 5067 2471 5070
rect 5073 5067 5139 5070
rect 16614 5068 16620 5070
rect 16684 5068 16690 5132
rect -300 4994 160 5024
rect 1301 4994 1367 4997
rect -300 4992 1367 4994
rect -300 4936 1306 4992
rect 1362 4936 1367 4992
rect -300 4934 1367 4936
rect -300 4904 160 4934
rect 1301 4931 1367 4934
rect 11421 4994 11487 4997
rect 13629 4994 13695 4997
rect 14917 4994 14983 4997
rect 11421 4992 14983 4994
rect 11421 4936 11426 4992
rect 11482 4936 13634 4992
rect 13690 4936 14922 4992
rect 14978 4936 14983 4992
rect 11421 4934 14983 4936
rect 11421 4931 11487 4934
rect 13629 4931 13695 4934
rect 14917 4931 14983 4934
rect 3878 4928 4194 4929
rect 3878 4864 3884 4928
rect 3948 4864 3964 4928
rect 4028 4864 4044 4928
rect 4108 4864 4124 4928
rect 4188 4864 4194 4928
rect 3878 4863 4194 4864
rect 9743 4928 10059 4929
rect 9743 4864 9749 4928
rect 9813 4864 9829 4928
rect 9893 4864 9909 4928
rect 9973 4864 9989 4928
rect 10053 4864 10059 4928
rect 9743 4863 10059 4864
rect 15608 4928 15924 4929
rect 15608 4864 15614 4928
rect 15678 4864 15694 4928
rect 15758 4864 15774 4928
rect 15838 4864 15854 4928
rect 15918 4864 15924 4928
rect 15608 4863 15924 4864
rect 21473 4928 21789 4929
rect 21473 4864 21479 4928
rect 21543 4864 21559 4928
rect 21623 4864 21639 4928
rect 21703 4864 21719 4928
rect 21783 4864 21789 4928
rect 21473 4863 21789 4864
rect 1669 4724 1735 4725
rect 1669 4722 1716 4724
rect 1588 4720 1716 4722
rect 1780 4722 1786 4724
rect 17585 4722 17651 4725
rect 1780 4720 17651 4722
rect 1588 4664 1674 4720
rect 1780 4664 17590 4720
rect 17646 4664 17651 4720
rect 1588 4662 1716 4664
rect 1669 4660 1716 4662
rect 1780 4662 17651 4664
rect 1780 4660 1786 4662
rect 1669 4659 1735 4660
rect 17585 4659 17651 4662
rect 21633 4722 21699 4725
rect 21950 4722 21956 4724
rect 21633 4720 21956 4722
rect 21633 4664 21638 4720
rect 21694 4664 21956 4720
rect 21633 4662 21956 4664
rect 21633 4659 21699 4662
rect 21950 4660 21956 4662
rect 22020 4660 22026 4724
rect 23246 4722 23306 5478
rect 23381 5536 24226 5538
rect 23381 5480 23386 5536
rect 23442 5480 24226 5536
rect 23381 5478 24226 5480
rect 23381 5475 23447 5478
rect 24166 5266 24226 5478
rect 24902 5478 26000 5538
rect 24405 5472 24721 5473
rect 24405 5408 24411 5472
rect 24475 5408 24491 5472
rect 24555 5408 24571 5472
rect 24635 5408 24651 5472
rect 24715 5408 24721 5472
rect 24405 5407 24721 5408
rect 24902 5266 24962 5478
rect 25540 5448 26000 5478
rect 24166 5206 24962 5266
rect 24025 4994 24091 4997
rect 25540 4994 26000 5024
rect 24025 4992 26000 4994
rect 24025 4936 24030 4992
rect 24086 4936 26000 4992
rect 24025 4934 26000 4936
rect 24025 4931 24091 4934
rect 25540 4904 26000 4934
rect 23246 4662 24962 4722
rect 8017 4586 8083 4589
rect 11145 4586 11211 4589
rect 8017 4584 11211 4586
rect 8017 4528 8022 4584
rect 8078 4528 11150 4584
rect 11206 4528 11211 4584
rect 8017 4526 11211 4528
rect 8017 4523 8083 4526
rect 11145 4523 11211 4526
rect 11329 4586 11395 4589
rect 24301 4586 24367 4589
rect 11329 4584 24367 4586
rect 11329 4528 11334 4584
rect 11390 4528 24306 4584
rect 24362 4528 24367 4584
rect 11329 4526 24367 4528
rect 11329 4523 11395 4526
rect 24301 4523 24367 4526
rect 19977 4450 20043 4453
rect 21081 4450 21147 4453
rect 19977 4448 21147 4450
rect 19977 4392 19982 4448
rect 20038 4392 21086 4448
rect 21142 4392 21147 4448
rect 19977 4390 21147 4392
rect 24902 4450 24962 4662
rect 25540 4450 26000 4480
rect 24902 4390 26000 4450
rect 19977 4387 20043 4390
rect 21081 4387 21147 4390
rect 6810 4384 7126 4385
rect 6810 4320 6816 4384
rect 6880 4320 6896 4384
rect 6960 4320 6976 4384
rect 7040 4320 7056 4384
rect 7120 4320 7126 4384
rect 6810 4319 7126 4320
rect 12675 4384 12991 4385
rect 12675 4320 12681 4384
rect 12745 4320 12761 4384
rect 12825 4320 12841 4384
rect 12905 4320 12921 4384
rect 12985 4320 12991 4384
rect 12675 4319 12991 4320
rect 18540 4384 18856 4385
rect 18540 4320 18546 4384
rect 18610 4320 18626 4384
rect 18690 4320 18706 4384
rect 18770 4320 18786 4384
rect 18850 4320 18856 4384
rect 18540 4319 18856 4320
rect 24405 4384 24721 4385
rect 24405 4320 24411 4384
rect 24475 4320 24491 4384
rect 24555 4320 24571 4384
rect 24635 4320 24651 4384
rect 24715 4320 24721 4384
rect 25540 4360 26000 4390
rect 24405 4319 24721 4320
rect 2681 4314 2747 4317
rect 5717 4314 5783 4317
rect 2681 4312 5783 4314
rect 2681 4256 2686 4312
rect 2742 4256 5722 4312
rect 5778 4256 5783 4312
rect 2681 4254 5783 4256
rect 2681 4251 2747 4254
rect 5717 4251 5783 4254
rect 19425 4314 19491 4317
rect 20253 4314 20319 4317
rect 19425 4312 20319 4314
rect 19425 4256 19430 4312
rect 19486 4256 20258 4312
rect 20314 4256 20319 4312
rect 19425 4254 20319 4256
rect 19425 4251 19491 4254
rect 20253 4251 20319 4254
rect 3233 4178 3299 4181
rect 2960 4176 3299 4178
rect 2960 4120 3238 4176
rect 3294 4120 3299 4176
rect 2960 4118 3299 4120
rect 1577 4042 1643 4045
rect 2814 4042 2820 4044
rect 1577 4040 2820 4042
rect 1577 3984 1582 4040
rect 1638 3984 2820 4040
rect 1577 3982 2820 3984
rect 1577 3979 1643 3982
rect 2814 3980 2820 3982
rect 2884 3980 2890 4044
rect 2960 3909 3020 4118
rect 3233 4115 3299 4118
rect 3509 4178 3575 4181
rect 3734 4178 3740 4180
rect 3509 4176 3740 4178
rect 3509 4120 3514 4176
rect 3570 4120 3740 4176
rect 3509 4118 3740 4120
rect 3509 4115 3575 4118
rect 3734 4116 3740 4118
rect 3804 4116 3810 4180
rect 4981 4178 5047 4181
rect 5625 4178 5691 4181
rect 4981 4176 5691 4178
rect 4981 4120 4986 4176
rect 5042 4120 5630 4176
rect 5686 4120 5691 4176
rect 4981 4118 5691 4120
rect 4981 4115 5047 4118
rect 5625 4115 5691 4118
rect 7281 4178 7347 4181
rect 12985 4178 13051 4181
rect 7281 4176 13051 4178
rect 7281 4120 7286 4176
rect 7342 4120 12990 4176
rect 13046 4120 13051 4176
rect 7281 4118 13051 4120
rect 7281 4115 7347 4118
rect 12985 4115 13051 4118
rect 3233 4042 3299 4045
rect 7925 4042 7991 4045
rect 3233 4040 7991 4042
rect 3233 3984 3238 4040
rect 3294 3984 7930 4040
rect 7986 3984 7991 4040
rect 3233 3982 7991 3984
rect 3233 3979 3299 3982
rect 7925 3979 7991 3982
rect 10869 4044 10935 4045
rect 10869 4040 10916 4044
rect 10980 4042 10986 4044
rect 11605 4042 11671 4045
rect 19701 4042 19767 4045
rect 10869 3984 10874 4040
rect 10869 3980 10916 3984
rect 10980 3982 11026 4042
rect 11605 4040 19767 4042
rect 11605 3984 11610 4040
rect 11666 3984 19706 4040
rect 19762 3984 19767 4040
rect 11605 3982 19767 3984
rect 10980 3980 10986 3982
rect 10869 3979 10935 3980
rect 11605 3979 11671 3982
rect 19701 3979 19767 3982
rect 19977 4042 20043 4045
rect 20110 4042 20116 4044
rect 19977 4040 20116 4042
rect 19977 3984 19982 4040
rect 20038 3984 20116 4040
rect 19977 3982 20116 3984
rect 19977 3979 20043 3982
rect 20110 3980 20116 3982
rect 20180 3980 20186 4044
rect 20897 4042 20963 4045
rect 20897 4040 23858 4042
rect 20897 3984 20902 4040
rect 20958 3984 23858 4040
rect 20897 3982 23858 3984
rect 20897 3979 20963 3982
rect 1945 3906 2011 3909
rect 2078 3906 2084 3908
rect 1945 3904 2084 3906
rect 1945 3848 1950 3904
rect 2006 3848 2084 3904
rect 1945 3846 2084 3848
rect 1945 3843 2011 3846
rect 2078 3844 2084 3846
rect 2148 3844 2154 3908
rect 2957 3904 3023 3909
rect 2957 3848 2962 3904
rect 3018 3848 3023 3904
rect 2957 3843 3023 3848
rect 22737 3906 22803 3909
rect 23798 3906 23858 3982
rect 25540 3906 26000 3936
rect 22737 3904 23674 3906
rect 22737 3848 22742 3904
rect 22798 3848 23674 3904
rect 22737 3846 23674 3848
rect 23798 3846 26000 3906
rect 22737 3843 22803 3846
rect 3878 3840 4194 3841
rect 3878 3776 3884 3840
rect 3948 3776 3964 3840
rect 4028 3776 4044 3840
rect 4108 3776 4124 3840
rect 4188 3776 4194 3840
rect 3878 3775 4194 3776
rect 9743 3840 10059 3841
rect 9743 3776 9749 3840
rect 9813 3776 9829 3840
rect 9893 3776 9909 3840
rect 9973 3776 9989 3840
rect 10053 3776 10059 3840
rect 9743 3775 10059 3776
rect 15608 3840 15924 3841
rect 15608 3776 15614 3840
rect 15678 3776 15694 3840
rect 15758 3776 15774 3840
rect 15838 3776 15854 3840
rect 15918 3776 15924 3840
rect 15608 3775 15924 3776
rect 21473 3840 21789 3841
rect 21473 3776 21479 3840
rect 21543 3776 21559 3840
rect 21623 3776 21639 3840
rect 21703 3776 21719 3840
rect 21783 3776 21789 3840
rect 21473 3775 21789 3776
rect 4797 3770 4863 3773
rect 5257 3770 5323 3773
rect 7373 3770 7439 3773
rect 4797 3768 7439 3770
rect 4797 3712 4802 3768
rect 4858 3712 5262 3768
rect 5318 3712 7378 3768
rect 7434 3712 7439 3768
rect 4797 3710 7439 3712
rect 4797 3707 4863 3710
rect 5257 3707 5323 3710
rect 7373 3707 7439 3710
rect 16021 3770 16087 3773
rect 19425 3770 19491 3773
rect 16021 3768 19491 3770
rect 16021 3712 16026 3768
rect 16082 3712 19430 3768
rect 19486 3712 19491 3768
rect 16021 3710 19491 3712
rect 16021 3707 16130 3710
rect 19425 3707 19491 3710
rect 3877 3634 3943 3637
rect 4613 3634 4679 3637
rect 16070 3634 16130 3707
rect 3877 3632 16130 3634
rect 3877 3576 3882 3632
rect 3938 3576 4618 3632
rect 4674 3576 16130 3632
rect 3877 3574 16130 3576
rect 17217 3634 17283 3637
rect 22185 3634 22251 3637
rect 17217 3632 22251 3634
rect 17217 3576 17222 3632
rect 17278 3576 22190 3632
rect 22246 3576 22251 3632
rect 17217 3574 22251 3576
rect 3877 3571 3943 3574
rect 4613 3571 4679 3574
rect 17217 3571 17283 3574
rect 22185 3571 22251 3574
rect 197 3498 263 3501
rect 4613 3498 4679 3501
rect 197 3496 4679 3498
rect 197 3440 202 3496
rect 258 3440 4618 3496
rect 4674 3440 4679 3496
rect 197 3438 4679 3440
rect 197 3435 263 3438
rect 4613 3435 4679 3438
rect 6269 3498 6335 3501
rect 8201 3498 8267 3501
rect 22277 3498 22343 3501
rect 6269 3496 7298 3498
rect 6269 3440 6274 3496
rect 6330 3440 7298 3496
rect 6269 3438 7298 3440
rect 6269 3435 6335 3438
rect 3601 3362 3667 3365
rect 4337 3362 4403 3365
rect 4797 3362 4863 3365
rect 3601 3360 4863 3362
rect 3601 3304 3606 3360
rect 3662 3304 4342 3360
rect 4398 3304 4802 3360
rect 4858 3304 4863 3360
rect 3601 3302 4863 3304
rect 7238 3362 7298 3438
rect 8201 3496 22343 3498
rect 8201 3440 8206 3496
rect 8262 3440 22282 3496
rect 22338 3440 22343 3496
rect 8201 3438 22343 3440
rect 23614 3498 23674 3846
rect 25540 3816 26000 3846
rect 23614 3438 24962 3498
rect 8201 3435 8267 3438
rect 22277 3435 22343 3438
rect 12157 3362 12223 3365
rect 7238 3360 12223 3362
rect 7238 3304 12162 3360
rect 12218 3304 12223 3360
rect 7238 3302 12223 3304
rect 3601 3299 3667 3302
rect 4337 3299 4403 3302
rect 4797 3299 4863 3302
rect 12157 3299 12223 3302
rect 20846 3300 20852 3364
rect 20916 3362 20922 3364
rect 21633 3362 21699 3365
rect 20916 3360 21699 3362
rect 20916 3304 21638 3360
rect 21694 3304 21699 3360
rect 20916 3302 21699 3304
rect 24902 3362 24962 3438
rect 25540 3362 26000 3392
rect 24902 3302 26000 3362
rect 20916 3300 20922 3302
rect 21633 3299 21699 3302
rect 6810 3296 7126 3297
rect 6810 3232 6816 3296
rect 6880 3232 6896 3296
rect 6960 3232 6976 3296
rect 7040 3232 7056 3296
rect 7120 3232 7126 3296
rect 6810 3231 7126 3232
rect 12675 3296 12991 3297
rect 12675 3232 12681 3296
rect 12745 3232 12761 3296
rect 12825 3232 12841 3296
rect 12905 3232 12921 3296
rect 12985 3232 12991 3296
rect 12675 3231 12991 3232
rect 18540 3296 18856 3297
rect 18540 3232 18546 3296
rect 18610 3232 18626 3296
rect 18690 3232 18706 3296
rect 18770 3232 18786 3296
rect 18850 3232 18856 3296
rect 18540 3231 18856 3232
rect 24405 3296 24721 3297
rect 24405 3232 24411 3296
rect 24475 3232 24491 3296
rect 24555 3232 24571 3296
rect 24635 3232 24651 3296
rect 24715 3232 24721 3296
rect 25540 3272 26000 3302
rect 24405 3231 24721 3232
rect 7373 3226 7439 3229
rect 12525 3226 12591 3229
rect 7373 3224 12591 3226
rect 7373 3168 7378 3224
rect 7434 3168 12530 3224
rect 12586 3168 12591 3224
rect 7373 3166 12591 3168
rect 7373 3163 7439 3166
rect 12525 3163 12591 3166
rect 20345 3226 20411 3229
rect 20897 3226 20963 3229
rect 20345 3224 20963 3226
rect 20345 3168 20350 3224
rect 20406 3168 20902 3224
rect 20958 3168 20963 3224
rect 20345 3166 20963 3168
rect 20345 3163 20411 3166
rect 20897 3163 20963 3166
rect 5349 3090 5415 3093
rect 8845 3090 8911 3093
rect 5349 3088 8911 3090
rect 5349 3032 5354 3088
rect 5410 3032 8850 3088
rect 8906 3032 8911 3088
rect 5349 3030 8911 3032
rect 5349 3027 5415 3030
rect 8845 3027 8911 3030
rect 12382 3028 12388 3092
rect 12452 3090 12458 3092
rect 13118 3090 13124 3092
rect 12452 3030 13124 3090
rect 12452 3028 12458 3030
rect 13118 3028 13124 3030
rect 13188 3028 13194 3092
rect 16481 3090 16547 3093
rect 17769 3090 17835 3093
rect 20529 3090 20595 3093
rect 23749 3090 23815 3093
rect 16481 3088 17602 3090
rect 16481 3032 16486 3088
rect 16542 3032 17602 3088
rect 16481 3030 17602 3032
rect 16481 3027 16547 3030
rect 1669 2954 1735 2957
rect 11789 2954 11855 2957
rect 1669 2952 11855 2954
rect 1669 2896 1674 2952
rect 1730 2896 11794 2952
rect 11850 2896 11855 2952
rect 1669 2894 11855 2896
rect 17542 2954 17602 3030
rect 17769 3088 20595 3090
rect 17769 3032 17774 3088
rect 17830 3032 20534 3088
rect 20590 3032 20595 3088
rect 17769 3030 20595 3032
rect 17769 3027 17835 3030
rect 20529 3027 20595 3030
rect 20670 3088 23815 3090
rect 20670 3032 23754 3088
rect 23810 3032 23815 3088
rect 20670 3030 23815 3032
rect 19885 2954 19951 2957
rect 20670 2954 20730 3030
rect 23749 3027 23815 3030
rect 17542 2952 20730 2954
rect 17542 2896 19890 2952
rect 19946 2896 20730 2952
rect 17542 2894 20730 2896
rect 20989 2954 21055 2957
rect 20989 2952 22110 2954
rect 20989 2896 20994 2952
rect 21050 2896 22110 2952
rect 20989 2894 22110 2896
rect 1669 2891 1735 2894
rect 11789 2891 11855 2894
rect 19885 2891 19951 2894
rect 20989 2891 21055 2894
rect 6361 2818 6427 2821
rect 6637 2818 6703 2821
rect 7741 2818 7807 2821
rect 6361 2816 6562 2818
rect 6361 2760 6366 2816
rect 6422 2760 6562 2816
rect 6361 2758 6562 2760
rect 6361 2755 6427 2758
rect 3878 2752 4194 2753
rect 3878 2688 3884 2752
rect 3948 2688 3964 2752
rect 4028 2688 4044 2752
rect 4108 2688 4124 2752
rect 4188 2688 4194 2752
rect 3878 2687 4194 2688
rect 5349 2684 5415 2685
rect 5349 2682 5396 2684
rect 5304 2680 5396 2682
rect 5304 2624 5354 2680
rect 5304 2622 5396 2624
rect 5349 2620 5396 2622
rect 5460 2620 5466 2684
rect 6502 2682 6562 2758
rect 6637 2816 7807 2818
rect 6637 2760 6642 2816
rect 6698 2760 7746 2816
rect 7802 2760 7807 2816
rect 6637 2758 7807 2760
rect 22050 2818 22110 2894
rect 25540 2818 26000 2848
rect 22050 2758 26000 2818
rect 6637 2755 6703 2758
rect 7741 2755 7807 2758
rect 9743 2752 10059 2753
rect 9743 2688 9749 2752
rect 9813 2688 9829 2752
rect 9893 2688 9909 2752
rect 9973 2688 9989 2752
rect 10053 2688 10059 2752
rect 9743 2687 10059 2688
rect 15608 2752 15924 2753
rect 15608 2688 15614 2752
rect 15678 2688 15694 2752
rect 15758 2688 15774 2752
rect 15838 2688 15854 2752
rect 15918 2688 15924 2752
rect 15608 2687 15924 2688
rect 21473 2752 21789 2753
rect 21473 2688 21479 2752
rect 21543 2688 21559 2752
rect 21623 2688 21639 2752
rect 21703 2688 21719 2752
rect 21783 2688 21789 2752
rect 25540 2728 26000 2758
rect 21473 2687 21789 2688
rect 11789 2682 11855 2685
rect 13302 2682 13308 2684
rect 6502 2622 7804 2682
rect 5349 2619 5415 2620
rect 606 2484 612 2548
rect 676 2546 682 2548
rect 7465 2546 7531 2549
rect 676 2544 7531 2546
rect 676 2488 7470 2544
rect 7526 2488 7531 2544
rect 676 2486 7531 2488
rect 676 2484 682 2486
rect 7465 2483 7531 2486
rect 3969 2410 4035 2413
rect 6269 2410 6335 2413
rect 7744 2410 7804 2622
rect 11789 2680 13308 2682
rect 11789 2624 11794 2680
rect 11850 2624 13308 2680
rect 11789 2622 13308 2624
rect 11789 2619 11855 2622
rect 13302 2620 13308 2622
rect 13372 2620 13378 2684
rect 16849 2682 16915 2685
rect 17125 2684 17191 2685
rect 19609 2684 19675 2685
rect 22185 2684 22251 2685
rect 16982 2682 16988 2684
rect 16849 2680 16988 2682
rect 16849 2624 16854 2680
rect 16910 2624 16988 2680
rect 16849 2622 16988 2624
rect 16849 2619 16915 2622
rect 16982 2620 16988 2622
rect 17052 2620 17058 2684
rect 17125 2680 17172 2684
rect 17236 2682 17242 2684
rect 19558 2682 19564 2684
rect 17125 2624 17130 2680
rect 17125 2620 17172 2624
rect 17236 2622 17282 2682
rect 19518 2622 19564 2682
rect 19628 2680 19675 2684
rect 22134 2682 22140 2684
rect 19670 2624 19675 2680
rect 17236 2620 17242 2622
rect 19558 2620 19564 2622
rect 19628 2620 19675 2624
rect 22094 2622 22140 2682
rect 22204 2680 22251 2684
rect 22246 2624 22251 2680
rect 22134 2620 22140 2622
rect 22204 2620 22251 2624
rect 17125 2619 17191 2620
rect 19609 2619 19675 2620
rect 22185 2619 22251 2620
rect 10225 2546 10291 2549
rect 10358 2546 10364 2548
rect 10225 2544 10364 2546
rect 10225 2488 10230 2544
rect 10286 2488 10364 2544
rect 10225 2486 10364 2488
rect 10225 2483 10291 2486
rect 10358 2484 10364 2486
rect 10428 2484 10434 2548
rect 13905 2546 13971 2549
rect 15326 2546 15332 2548
rect 13862 2544 15332 2546
rect 13862 2488 13910 2544
rect 13966 2488 15332 2544
rect 13862 2486 15332 2488
rect 13862 2483 13971 2486
rect 15326 2484 15332 2486
rect 15396 2484 15402 2548
rect 16389 2546 16455 2549
rect 20621 2546 20687 2549
rect 16389 2544 20687 2546
rect 16389 2488 16394 2544
rect 16450 2488 20626 2544
rect 20682 2488 20687 2544
rect 16389 2486 20687 2488
rect 16389 2483 16455 2486
rect 20621 2483 20687 2486
rect 21817 2546 21883 2549
rect 21817 2544 24962 2546
rect 21817 2488 21822 2544
rect 21878 2488 24962 2544
rect 21817 2486 24962 2488
rect 21817 2483 21883 2486
rect 11237 2410 11303 2413
rect 3969 2408 7620 2410
rect 3969 2352 3974 2408
rect 4030 2352 6274 2408
rect 6330 2352 7620 2408
rect 3969 2350 7620 2352
rect 7744 2408 11303 2410
rect 7744 2352 11242 2408
rect 11298 2352 11303 2408
rect 7744 2350 11303 2352
rect 3969 2347 4035 2350
rect 6269 2347 6335 2350
rect 7281 2274 7347 2277
rect 7414 2274 7420 2276
rect 7281 2272 7420 2274
rect 7281 2216 7286 2272
rect 7342 2216 7420 2272
rect 7281 2214 7420 2216
rect 7281 2211 7347 2214
rect 7414 2212 7420 2214
rect 7484 2212 7490 2276
rect 6810 2208 7126 2209
rect 6810 2144 6816 2208
rect 6880 2144 6896 2208
rect 6960 2144 6976 2208
rect 7040 2144 7056 2208
rect 7120 2144 7126 2208
rect 6810 2143 7126 2144
rect 7560 2138 7620 2350
rect 11237 2347 11303 2350
rect 11881 2410 11947 2413
rect 12014 2410 12020 2412
rect 11881 2408 12020 2410
rect 11881 2352 11886 2408
rect 11942 2352 12020 2408
rect 11881 2350 12020 2352
rect 11881 2347 11947 2350
rect 12014 2348 12020 2350
rect 12084 2348 12090 2412
rect 13862 2410 13922 2483
rect 12390 2350 13922 2410
rect 15745 2410 15811 2413
rect 21081 2410 21147 2413
rect 21214 2410 21220 2412
rect 15745 2408 20914 2410
rect 15745 2352 15750 2408
rect 15806 2352 20914 2408
rect 15745 2350 20914 2352
rect 8109 2276 8175 2277
rect 8845 2276 8911 2277
rect 8109 2274 8156 2276
rect 8064 2272 8156 2274
rect 8064 2216 8114 2272
rect 8064 2214 8156 2216
rect 8109 2212 8156 2214
rect 8220 2212 8226 2276
rect 8845 2274 8892 2276
rect 8800 2272 8892 2274
rect 8800 2216 8850 2272
rect 8800 2214 8892 2216
rect 8845 2212 8892 2214
rect 8956 2212 8962 2276
rect 9673 2274 9739 2277
rect 11145 2274 11211 2277
rect 9673 2272 11211 2274
rect 9673 2216 9678 2272
rect 9734 2216 11150 2272
rect 11206 2216 11211 2272
rect 9673 2214 11211 2216
rect 8109 2211 8175 2212
rect 8845 2211 8911 2212
rect 9673 2211 9739 2214
rect 11145 2211 11211 2214
rect 11973 2274 12039 2277
rect 12390 2274 12450 2350
rect 15745 2347 15811 2350
rect 11973 2272 12450 2274
rect 11973 2216 11978 2272
rect 12034 2216 12450 2272
rect 11973 2214 12450 2216
rect 20854 2274 20914 2350
rect 21081 2408 21220 2410
rect 21081 2352 21086 2408
rect 21142 2352 21220 2408
rect 21081 2350 21220 2352
rect 21081 2347 21147 2350
rect 21214 2348 21220 2350
rect 21284 2348 21290 2412
rect 22185 2410 22251 2413
rect 22050 2408 22251 2410
rect 22050 2352 22190 2408
rect 22246 2352 22251 2408
rect 22050 2350 22251 2352
rect 22050 2274 22110 2350
rect 22185 2347 22251 2350
rect 20854 2214 22110 2274
rect 24902 2274 24962 2486
rect 25540 2274 26000 2304
rect 24902 2214 26000 2274
rect 11973 2211 12039 2214
rect 12675 2208 12991 2209
rect 12675 2144 12681 2208
rect 12745 2144 12761 2208
rect 12825 2144 12841 2208
rect 12905 2144 12921 2208
rect 12985 2144 12991 2208
rect 12675 2143 12991 2144
rect 18540 2208 18856 2209
rect 18540 2144 18546 2208
rect 18610 2144 18626 2208
rect 18690 2144 18706 2208
rect 18770 2144 18786 2208
rect 18850 2144 18856 2208
rect 18540 2143 18856 2144
rect 24405 2208 24721 2209
rect 24405 2144 24411 2208
rect 24475 2144 24491 2208
rect 24555 2144 24571 2208
rect 24635 2144 24651 2208
rect 24715 2144 24721 2208
rect 25540 2184 26000 2214
rect 24405 2143 24721 2144
rect 12249 2138 12315 2141
rect 14457 2140 14523 2141
rect 7560 2136 12315 2138
rect 7560 2080 12254 2136
rect 12310 2080 12315 2136
rect 7560 2078 12315 2080
rect 12249 2075 12315 2078
rect 14406 2076 14412 2140
rect 14476 2138 14523 2140
rect 14476 2136 14568 2138
rect 14518 2080 14568 2136
rect 14476 2078 14568 2080
rect 14476 2076 14523 2078
rect 14457 2075 14523 2076
rect 974 1940 980 2004
rect 1044 2002 1050 2004
rect 7649 2002 7715 2005
rect 1044 2000 7715 2002
rect 1044 1944 7654 2000
rect 7710 1944 7715 2000
rect 1044 1942 7715 1944
rect 1044 1940 1050 1942
rect 7649 1939 7715 1942
rect 9489 2002 9555 2005
rect 22502 2002 22508 2004
rect 9489 2000 22508 2002
rect 9489 1944 9494 2000
rect 9550 1944 22508 2000
rect 9489 1942 22508 1944
rect 9489 1939 9555 1942
rect 22502 1940 22508 1942
rect 22572 1940 22578 2004
rect 1158 1804 1164 1868
rect 1228 1866 1234 1868
rect 8385 1866 8451 1869
rect 1228 1864 8451 1866
rect 1228 1808 8390 1864
rect 8446 1808 8451 1864
rect 1228 1806 8451 1808
rect 1228 1804 1234 1806
rect 8385 1803 8451 1806
rect 9949 1866 10015 1869
rect 13077 1866 13143 1869
rect 9949 1864 13143 1866
rect 9949 1808 9954 1864
rect 10010 1808 13082 1864
rect 13138 1808 13143 1864
rect 9949 1806 13143 1808
rect 9949 1803 10015 1806
rect 13077 1803 13143 1806
rect 19977 1866 20043 1869
rect 21541 1866 21607 1869
rect 19977 1864 21607 1866
rect 19977 1808 19982 1864
rect 20038 1808 21546 1864
rect 21602 1808 21607 1864
rect 19977 1806 21607 1808
rect 19977 1803 20043 1806
rect 21541 1803 21607 1806
rect 10225 1730 10291 1733
rect 11513 1730 11579 1733
rect 10225 1728 11579 1730
rect 10225 1672 10230 1728
rect 10286 1672 11518 1728
rect 11574 1672 11579 1728
rect 10225 1670 11579 1672
rect 10225 1667 10291 1670
rect 11513 1667 11579 1670
rect 22001 1730 22067 1733
rect 25540 1730 26000 1760
rect 22001 1728 26000 1730
rect 22001 1672 22006 1728
rect 22062 1672 26000 1728
rect 22001 1670 26000 1672
rect 22001 1667 22067 1670
rect 3878 1664 4194 1665
rect 3878 1600 3884 1664
rect 3948 1600 3964 1664
rect 4028 1600 4044 1664
rect 4108 1600 4124 1664
rect 4188 1600 4194 1664
rect 3878 1599 4194 1600
rect 9743 1664 10059 1665
rect 9743 1600 9749 1664
rect 9813 1600 9829 1664
rect 9893 1600 9909 1664
rect 9973 1600 9989 1664
rect 10053 1600 10059 1664
rect 9743 1599 10059 1600
rect 15608 1664 15924 1665
rect 15608 1600 15614 1664
rect 15678 1600 15694 1664
rect 15758 1600 15774 1664
rect 15838 1600 15854 1664
rect 15918 1600 15924 1664
rect 15608 1599 15924 1600
rect 21473 1664 21789 1665
rect 21473 1600 21479 1664
rect 21543 1600 21559 1664
rect 21623 1600 21639 1664
rect 21703 1600 21719 1664
rect 21783 1600 21789 1664
rect 25540 1640 26000 1670
rect 21473 1599 21789 1600
rect 3785 1460 3851 1461
rect 3734 1458 3740 1460
rect 3658 1398 3740 1458
rect 3804 1458 3851 1460
rect 11053 1458 11119 1461
rect 3804 1456 11119 1458
rect 3846 1400 11058 1456
rect 11114 1400 11119 1456
rect 3734 1396 3740 1398
rect 3804 1398 11119 1400
rect 3804 1396 3851 1398
rect 3785 1395 3851 1396
rect 11053 1395 11119 1398
rect 4429 1324 4495 1325
rect 4429 1320 4476 1324
rect 4540 1322 4546 1324
rect 7925 1322 7991 1325
rect 8702 1322 8708 1324
rect 4429 1264 4434 1320
rect 4429 1260 4476 1264
rect 4540 1262 4586 1322
rect 7925 1320 8708 1322
rect 7925 1264 7930 1320
rect 7986 1264 8708 1320
rect 7925 1262 8708 1264
rect 4540 1260 4546 1262
rect 4429 1259 4495 1260
rect 7925 1259 7991 1262
rect 8702 1260 8708 1262
rect 8772 1260 8778 1324
rect 9627 1322 9693 1325
rect 10041 1322 10107 1325
rect 9627 1320 10107 1322
rect 9627 1264 9632 1320
rect 9688 1264 10046 1320
rect 10102 1264 10107 1320
rect 9627 1262 10107 1264
rect 9627 1259 9693 1262
rect 10041 1259 10107 1262
rect 11053 1324 11119 1325
rect 11053 1320 11100 1324
rect 11164 1322 11170 1324
rect 11053 1264 11058 1320
rect 11053 1260 11100 1264
rect 11164 1262 11210 1322
rect 11164 1260 11170 1262
rect 12382 1260 12388 1324
rect 12452 1322 12458 1324
rect 12709 1322 12775 1325
rect 12452 1320 12775 1322
rect 12452 1264 12714 1320
rect 12770 1264 12775 1320
rect 12452 1262 12775 1264
rect 12452 1260 12458 1262
rect 11053 1259 11119 1260
rect 12709 1259 12775 1262
rect 13445 1324 13511 1325
rect 13445 1320 13492 1324
rect 13556 1322 13562 1324
rect 14089 1322 14155 1325
rect 14549 1324 14615 1325
rect 15193 1324 15259 1325
rect 14222 1322 14228 1324
rect 13445 1264 13450 1320
rect 13445 1260 13492 1264
rect 13556 1262 13602 1322
rect 14089 1320 14228 1322
rect 14089 1264 14094 1320
rect 14150 1264 14228 1320
rect 14089 1262 14228 1264
rect 13556 1260 13562 1262
rect 13445 1259 13511 1260
rect 14089 1259 14155 1262
rect 14222 1260 14228 1262
rect 14292 1260 14298 1324
rect 14549 1320 14596 1324
rect 14660 1322 14666 1324
rect 14549 1264 14554 1320
rect 14549 1260 14596 1264
rect 14660 1262 14706 1322
rect 14660 1260 14666 1262
rect 15142 1260 15148 1324
rect 15212 1322 15259 1324
rect 15212 1320 15304 1322
rect 15254 1264 15304 1320
rect 15212 1262 15304 1264
rect 24166 1262 24962 1322
rect 15212 1260 15259 1262
rect 14549 1259 14615 1260
rect 15193 1259 15259 1260
rect 2129 1186 2195 1189
rect 6126 1186 6132 1188
rect 2129 1184 6132 1186
rect 2129 1128 2134 1184
rect 2190 1128 6132 1184
rect 2129 1126 6132 1128
rect 2129 1123 2195 1126
rect 6126 1124 6132 1126
rect 6196 1124 6202 1188
rect 7465 1186 7531 1189
rect 8334 1186 8340 1188
rect 7465 1184 8340 1186
rect 7465 1128 7470 1184
rect 7526 1128 8340 1184
rect 7465 1126 8340 1128
rect 7465 1123 7531 1126
rect 8334 1124 8340 1126
rect 8404 1124 8410 1188
rect 9213 1186 9279 1189
rect 11513 1186 11579 1189
rect 9213 1184 11579 1186
rect 9213 1128 9218 1184
rect 9274 1128 11518 1184
rect 11574 1128 11579 1184
rect 9213 1126 11579 1128
rect 9213 1123 9279 1126
rect 11513 1123 11579 1126
rect 20713 1186 20779 1189
rect 24166 1186 24226 1262
rect 20713 1184 24226 1186
rect 20713 1128 20718 1184
rect 20774 1128 24226 1184
rect 20713 1126 24226 1128
rect 24902 1186 24962 1262
rect 25540 1186 26000 1216
rect 24902 1126 26000 1186
rect 20713 1123 20779 1126
rect 6810 1120 7126 1121
rect 6810 1056 6816 1120
rect 6880 1056 6896 1120
rect 6960 1056 6976 1120
rect 7040 1056 7056 1120
rect 7120 1056 7126 1120
rect 6810 1055 7126 1056
rect 12675 1120 12991 1121
rect 12675 1056 12681 1120
rect 12745 1056 12761 1120
rect 12825 1056 12841 1120
rect 12905 1056 12921 1120
rect 12985 1056 12991 1120
rect 12675 1055 12991 1056
rect 18540 1120 18856 1121
rect 18540 1056 18546 1120
rect 18610 1056 18626 1120
rect 18690 1056 18706 1120
rect 18770 1056 18786 1120
rect 18850 1056 18856 1120
rect 18540 1055 18856 1056
rect 24405 1120 24721 1121
rect 24405 1056 24411 1120
rect 24475 1056 24491 1120
rect 24555 1056 24571 1120
rect 24635 1056 24651 1120
rect 24715 1056 24721 1120
rect 25540 1096 26000 1126
rect 24405 1055 24721 1056
rect 2773 914 2839 917
rect 19374 914 19380 916
rect 2773 912 19380 914
rect 2773 856 2778 912
rect 2834 856 19380 912
rect 2773 854 19380 856
rect 2773 851 2839 854
rect 19374 852 19380 854
rect 19444 852 19450 916
rect 4061 778 4127 781
rect 10542 778 10548 780
rect 4061 776 10548 778
rect 4061 720 4066 776
rect 4122 720 10548 776
rect 4061 718 10548 720
rect 4061 715 4127 718
rect 10542 716 10548 718
rect 10612 716 10618 780
rect 22369 642 22435 645
rect 25540 642 26000 672
rect 22369 640 26000 642
rect 22369 584 22374 640
rect 22430 584 26000 640
rect 22369 582 26000 584
rect 22369 579 22435 582
rect 25540 552 26000 582
rect 790 444 796 508
rect 860 506 866 508
rect 7741 506 7807 509
rect 860 504 7807 506
rect 860 448 7746 504
rect 7802 448 7807 504
rect 860 446 7807 448
rect 860 444 866 446
rect 7741 443 7807 446
<< via3 >>
rect 6816 43548 6880 43552
rect 6816 43492 6820 43548
rect 6820 43492 6876 43548
rect 6876 43492 6880 43548
rect 6816 43488 6880 43492
rect 6896 43548 6960 43552
rect 6896 43492 6900 43548
rect 6900 43492 6956 43548
rect 6956 43492 6960 43548
rect 6896 43488 6960 43492
rect 6976 43548 7040 43552
rect 6976 43492 6980 43548
rect 6980 43492 7036 43548
rect 7036 43492 7040 43548
rect 6976 43488 7040 43492
rect 7056 43548 7120 43552
rect 7056 43492 7060 43548
rect 7060 43492 7116 43548
rect 7116 43492 7120 43548
rect 7056 43488 7120 43492
rect 12681 43548 12745 43552
rect 12681 43492 12685 43548
rect 12685 43492 12741 43548
rect 12741 43492 12745 43548
rect 12681 43488 12745 43492
rect 12761 43548 12825 43552
rect 12761 43492 12765 43548
rect 12765 43492 12821 43548
rect 12821 43492 12825 43548
rect 12761 43488 12825 43492
rect 12841 43548 12905 43552
rect 12841 43492 12845 43548
rect 12845 43492 12901 43548
rect 12901 43492 12905 43548
rect 12841 43488 12905 43492
rect 12921 43548 12985 43552
rect 12921 43492 12925 43548
rect 12925 43492 12981 43548
rect 12981 43492 12985 43548
rect 12921 43488 12985 43492
rect 18546 43548 18610 43552
rect 18546 43492 18550 43548
rect 18550 43492 18606 43548
rect 18606 43492 18610 43548
rect 18546 43488 18610 43492
rect 18626 43548 18690 43552
rect 18626 43492 18630 43548
rect 18630 43492 18686 43548
rect 18686 43492 18690 43548
rect 18626 43488 18690 43492
rect 18706 43548 18770 43552
rect 18706 43492 18710 43548
rect 18710 43492 18766 43548
rect 18766 43492 18770 43548
rect 18706 43488 18770 43492
rect 18786 43548 18850 43552
rect 18786 43492 18790 43548
rect 18790 43492 18846 43548
rect 18846 43492 18850 43548
rect 18786 43488 18850 43492
rect 24411 43548 24475 43552
rect 24411 43492 24415 43548
rect 24415 43492 24471 43548
rect 24471 43492 24475 43548
rect 24411 43488 24475 43492
rect 24491 43548 24555 43552
rect 24491 43492 24495 43548
rect 24495 43492 24551 43548
rect 24551 43492 24555 43548
rect 24491 43488 24555 43492
rect 24571 43548 24635 43552
rect 24571 43492 24575 43548
rect 24575 43492 24631 43548
rect 24631 43492 24635 43548
rect 24571 43488 24635 43492
rect 24651 43548 24715 43552
rect 24651 43492 24655 43548
rect 24655 43492 24711 43548
rect 24711 43492 24715 43548
rect 24651 43488 24715 43492
rect 3884 43004 3948 43008
rect 3884 42948 3888 43004
rect 3888 42948 3944 43004
rect 3944 42948 3948 43004
rect 3884 42944 3948 42948
rect 3964 43004 4028 43008
rect 3964 42948 3968 43004
rect 3968 42948 4024 43004
rect 4024 42948 4028 43004
rect 3964 42944 4028 42948
rect 4044 43004 4108 43008
rect 4044 42948 4048 43004
rect 4048 42948 4104 43004
rect 4104 42948 4108 43004
rect 4044 42944 4108 42948
rect 4124 43004 4188 43008
rect 4124 42948 4128 43004
rect 4128 42948 4184 43004
rect 4184 42948 4188 43004
rect 4124 42944 4188 42948
rect 9749 43004 9813 43008
rect 9749 42948 9753 43004
rect 9753 42948 9809 43004
rect 9809 42948 9813 43004
rect 9749 42944 9813 42948
rect 9829 43004 9893 43008
rect 9829 42948 9833 43004
rect 9833 42948 9889 43004
rect 9889 42948 9893 43004
rect 9829 42944 9893 42948
rect 9909 43004 9973 43008
rect 9909 42948 9913 43004
rect 9913 42948 9969 43004
rect 9969 42948 9973 43004
rect 9909 42944 9973 42948
rect 9989 43004 10053 43008
rect 9989 42948 9993 43004
rect 9993 42948 10049 43004
rect 10049 42948 10053 43004
rect 9989 42944 10053 42948
rect 980 42740 1044 42804
rect 21956 43148 22020 43212
rect 11652 43012 11716 43076
rect 15614 43004 15678 43008
rect 15614 42948 15618 43004
rect 15618 42948 15674 43004
rect 15674 42948 15678 43004
rect 15614 42944 15678 42948
rect 15694 43004 15758 43008
rect 15694 42948 15698 43004
rect 15698 42948 15754 43004
rect 15754 42948 15758 43004
rect 15694 42944 15758 42948
rect 15774 43004 15838 43008
rect 15774 42948 15778 43004
rect 15778 42948 15834 43004
rect 15834 42948 15838 43004
rect 15774 42944 15838 42948
rect 15854 43004 15918 43008
rect 15854 42948 15858 43004
rect 15858 42948 15914 43004
rect 15914 42948 15918 43004
rect 15854 42944 15918 42948
rect 21479 43004 21543 43008
rect 21479 42948 21483 43004
rect 21483 42948 21539 43004
rect 21539 42948 21543 43004
rect 21479 42944 21543 42948
rect 21559 43004 21623 43008
rect 21559 42948 21563 43004
rect 21563 42948 21619 43004
rect 21619 42948 21623 43004
rect 21559 42944 21623 42948
rect 21639 43004 21703 43008
rect 21639 42948 21643 43004
rect 21643 42948 21699 43004
rect 21699 42948 21703 43004
rect 21639 42944 21703 42948
rect 21719 43004 21783 43008
rect 21719 42948 21723 43004
rect 21723 42948 21779 43004
rect 21779 42948 21783 43004
rect 21719 42944 21783 42948
rect 11836 42936 11900 42940
rect 11836 42880 11850 42936
rect 11850 42880 11900 42936
rect 11836 42876 11900 42880
rect 14964 42936 15028 42940
rect 14964 42880 15014 42936
rect 15014 42880 15028 42936
rect 14964 42876 15028 42880
rect 15332 42876 15396 42940
rect 17724 42876 17788 42940
rect 16620 42604 16684 42668
rect 22140 42604 22204 42668
rect 4844 42468 4908 42532
rect 6816 42460 6880 42464
rect 6816 42404 6820 42460
rect 6820 42404 6876 42460
rect 6876 42404 6880 42460
rect 6816 42400 6880 42404
rect 6896 42460 6960 42464
rect 6896 42404 6900 42460
rect 6900 42404 6956 42460
rect 6956 42404 6960 42460
rect 6896 42400 6960 42404
rect 6976 42460 7040 42464
rect 6976 42404 6980 42460
rect 6980 42404 7036 42460
rect 7036 42404 7040 42460
rect 6976 42400 7040 42404
rect 7056 42460 7120 42464
rect 7056 42404 7060 42460
rect 7060 42404 7116 42460
rect 7116 42404 7120 42460
rect 7056 42400 7120 42404
rect 12681 42460 12745 42464
rect 12681 42404 12685 42460
rect 12685 42404 12741 42460
rect 12741 42404 12745 42460
rect 12681 42400 12745 42404
rect 12761 42460 12825 42464
rect 12761 42404 12765 42460
rect 12765 42404 12821 42460
rect 12821 42404 12825 42460
rect 12761 42400 12825 42404
rect 12841 42460 12905 42464
rect 12841 42404 12845 42460
rect 12845 42404 12901 42460
rect 12901 42404 12905 42460
rect 12841 42400 12905 42404
rect 12921 42460 12985 42464
rect 12921 42404 12925 42460
rect 12925 42404 12981 42460
rect 12981 42404 12985 42460
rect 12921 42400 12985 42404
rect 18546 42460 18610 42464
rect 18546 42404 18550 42460
rect 18550 42404 18606 42460
rect 18606 42404 18610 42460
rect 18546 42400 18610 42404
rect 18626 42460 18690 42464
rect 18626 42404 18630 42460
rect 18630 42404 18686 42460
rect 18686 42404 18690 42460
rect 18626 42400 18690 42404
rect 18706 42460 18770 42464
rect 18706 42404 18710 42460
rect 18710 42404 18766 42460
rect 18766 42404 18770 42460
rect 18706 42400 18770 42404
rect 18786 42460 18850 42464
rect 18786 42404 18790 42460
rect 18790 42404 18846 42460
rect 18846 42404 18850 42460
rect 18786 42400 18850 42404
rect 24411 42460 24475 42464
rect 24411 42404 24415 42460
rect 24415 42404 24471 42460
rect 24471 42404 24475 42460
rect 24411 42400 24475 42404
rect 24491 42460 24555 42464
rect 24491 42404 24495 42460
rect 24495 42404 24551 42460
rect 24551 42404 24555 42460
rect 24491 42400 24555 42404
rect 24571 42460 24635 42464
rect 24571 42404 24575 42460
rect 24575 42404 24631 42460
rect 24631 42404 24635 42460
rect 24571 42400 24635 42404
rect 24651 42460 24715 42464
rect 24651 42404 24655 42460
rect 24655 42404 24711 42460
rect 24711 42404 24715 42460
rect 24651 42400 24715 42404
rect 5580 42060 5644 42124
rect 10364 42060 10428 42124
rect 16988 42060 17052 42124
rect 8892 41924 8956 41988
rect 17172 41924 17236 41988
rect 18276 41984 18340 41988
rect 18276 41928 18326 41984
rect 18326 41928 18340 41984
rect 18276 41924 18340 41928
rect 19564 41984 19628 41988
rect 19564 41928 19578 41984
rect 19578 41928 19628 41984
rect 19564 41924 19628 41928
rect 19932 41924 19996 41988
rect 3884 41916 3948 41920
rect 3884 41860 3888 41916
rect 3888 41860 3944 41916
rect 3944 41860 3948 41916
rect 3884 41856 3948 41860
rect 3964 41916 4028 41920
rect 3964 41860 3968 41916
rect 3968 41860 4024 41916
rect 4024 41860 4028 41916
rect 3964 41856 4028 41860
rect 4044 41916 4108 41920
rect 4044 41860 4048 41916
rect 4048 41860 4104 41916
rect 4104 41860 4108 41916
rect 4044 41856 4108 41860
rect 4124 41916 4188 41920
rect 4124 41860 4128 41916
rect 4128 41860 4184 41916
rect 4184 41860 4188 41916
rect 4124 41856 4188 41860
rect 9749 41916 9813 41920
rect 9749 41860 9753 41916
rect 9753 41860 9809 41916
rect 9809 41860 9813 41916
rect 9749 41856 9813 41860
rect 9829 41916 9893 41920
rect 9829 41860 9833 41916
rect 9833 41860 9889 41916
rect 9889 41860 9893 41916
rect 9829 41856 9893 41860
rect 9909 41916 9973 41920
rect 9909 41860 9913 41916
rect 9913 41860 9969 41916
rect 9969 41860 9973 41916
rect 9909 41856 9973 41860
rect 9989 41916 10053 41920
rect 9989 41860 9993 41916
rect 9993 41860 10049 41916
rect 10049 41860 10053 41916
rect 9989 41856 10053 41860
rect 15614 41916 15678 41920
rect 15614 41860 15618 41916
rect 15618 41860 15674 41916
rect 15674 41860 15678 41916
rect 15614 41856 15678 41860
rect 15694 41916 15758 41920
rect 15694 41860 15698 41916
rect 15698 41860 15754 41916
rect 15754 41860 15758 41916
rect 15694 41856 15758 41860
rect 15774 41916 15838 41920
rect 15774 41860 15778 41916
rect 15778 41860 15834 41916
rect 15834 41860 15838 41916
rect 15774 41856 15838 41860
rect 15854 41916 15918 41920
rect 15854 41860 15858 41916
rect 15858 41860 15914 41916
rect 15914 41860 15918 41916
rect 15854 41856 15918 41860
rect 21479 41916 21543 41920
rect 21479 41860 21483 41916
rect 21483 41860 21539 41916
rect 21539 41860 21543 41916
rect 21479 41856 21543 41860
rect 21559 41916 21623 41920
rect 21559 41860 21563 41916
rect 21563 41860 21619 41916
rect 21619 41860 21623 41916
rect 21559 41856 21623 41860
rect 21639 41916 21703 41920
rect 21639 41860 21643 41916
rect 21643 41860 21699 41916
rect 21699 41860 21703 41916
rect 21639 41856 21703 41860
rect 21719 41916 21783 41920
rect 21719 41860 21723 41916
rect 21723 41860 21779 41916
rect 21779 41860 21783 41916
rect 21719 41856 21783 41860
rect 9076 41848 9140 41852
rect 9076 41792 9090 41848
rect 9090 41792 9140 41848
rect 9076 41788 9140 41792
rect 3740 41516 3804 41580
rect 1532 41380 1596 41444
rect 2452 41380 2516 41444
rect 6132 41380 6196 41444
rect 6816 41372 6880 41376
rect 6816 41316 6820 41372
rect 6820 41316 6876 41372
rect 6876 41316 6880 41372
rect 6816 41312 6880 41316
rect 6896 41372 6960 41376
rect 6896 41316 6900 41372
rect 6900 41316 6956 41372
rect 6956 41316 6960 41372
rect 6896 41312 6960 41316
rect 6976 41372 7040 41376
rect 6976 41316 6980 41372
rect 6980 41316 7036 41372
rect 7036 41316 7040 41372
rect 6976 41312 7040 41316
rect 7056 41372 7120 41376
rect 7056 41316 7060 41372
rect 7060 41316 7116 41372
rect 7116 41316 7120 41372
rect 7056 41312 7120 41316
rect 9260 41516 9324 41580
rect 9444 41516 9508 41580
rect 21220 41516 21284 41580
rect 10916 41380 10980 41444
rect 12681 41372 12745 41376
rect 12681 41316 12685 41372
rect 12685 41316 12741 41372
rect 12741 41316 12745 41372
rect 12681 41312 12745 41316
rect 12761 41372 12825 41376
rect 12761 41316 12765 41372
rect 12765 41316 12821 41372
rect 12821 41316 12825 41372
rect 12761 41312 12825 41316
rect 12841 41372 12905 41376
rect 12841 41316 12845 41372
rect 12845 41316 12901 41372
rect 12901 41316 12905 41372
rect 12841 41312 12905 41316
rect 12921 41372 12985 41376
rect 12921 41316 12925 41372
rect 12925 41316 12981 41372
rect 12981 41316 12985 41372
rect 12921 41312 12985 41316
rect 18546 41372 18610 41376
rect 18546 41316 18550 41372
rect 18550 41316 18606 41372
rect 18606 41316 18610 41372
rect 18546 41312 18610 41316
rect 18626 41372 18690 41376
rect 18626 41316 18630 41372
rect 18630 41316 18686 41372
rect 18686 41316 18690 41372
rect 18626 41312 18690 41316
rect 18706 41372 18770 41376
rect 18706 41316 18710 41372
rect 18710 41316 18766 41372
rect 18766 41316 18770 41372
rect 18706 41312 18770 41316
rect 18786 41372 18850 41376
rect 18786 41316 18790 41372
rect 18790 41316 18846 41372
rect 18846 41316 18850 41372
rect 18786 41312 18850 41316
rect 24411 41372 24475 41376
rect 24411 41316 24415 41372
rect 24415 41316 24471 41372
rect 24471 41316 24475 41372
rect 24411 41312 24475 41316
rect 24491 41372 24555 41376
rect 24491 41316 24495 41372
rect 24495 41316 24551 41372
rect 24551 41316 24555 41372
rect 24491 41312 24555 41316
rect 24571 41372 24635 41376
rect 24571 41316 24575 41372
rect 24575 41316 24631 41372
rect 24631 41316 24635 41372
rect 24571 41312 24635 41316
rect 24651 41372 24715 41376
rect 24651 41316 24655 41372
rect 24655 41316 24711 41372
rect 24711 41316 24715 41372
rect 24651 41312 24715 41316
rect 3884 40828 3948 40832
rect 3884 40772 3888 40828
rect 3888 40772 3944 40828
rect 3944 40772 3948 40828
rect 3884 40768 3948 40772
rect 3964 40828 4028 40832
rect 3964 40772 3968 40828
rect 3968 40772 4024 40828
rect 4024 40772 4028 40828
rect 3964 40768 4028 40772
rect 4044 40828 4108 40832
rect 4044 40772 4048 40828
rect 4048 40772 4104 40828
rect 4104 40772 4108 40828
rect 4044 40768 4108 40772
rect 4124 40828 4188 40832
rect 4124 40772 4128 40828
rect 4128 40772 4184 40828
rect 4184 40772 4188 40828
rect 4124 40768 4188 40772
rect 9749 40828 9813 40832
rect 9749 40772 9753 40828
rect 9753 40772 9809 40828
rect 9809 40772 9813 40828
rect 9749 40768 9813 40772
rect 9829 40828 9893 40832
rect 9829 40772 9833 40828
rect 9833 40772 9889 40828
rect 9889 40772 9893 40828
rect 9829 40768 9893 40772
rect 9909 40828 9973 40832
rect 9909 40772 9913 40828
rect 9913 40772 9969 40828
rect 9969 40772 9973 40828
rect 9909 40768 9973 40772
rect 9989 40828 10053 40832
rect 9989 40772 9993 40828
rect 9993 40772 10049 40828
rect 10049 40772 10053 40828
rect 9989 40768 10053 40772
rect 15614 40828 15678 40832
rect 15614 40772 15618 40828
rect 15618 40772 15674 40828
rect 15674 40772 15678 40828
rect 15614 40768 15678 40772
rect 15694 40828 15758 40832
rect 15694 40772 15698 40828
rect 15698 40772 15754 40828
rect 15754 40772 15758 40828
rect 15694 40768 15758 40772
rect 15774 40828 15838 40832
rect 15774 40772 15778 40828
rect 15778 40772 15834 40828
rect 15834 40772 15838 40828
rect 15774 40768 15838 40772
rect 15854 40828 15918 40832
rect 15854 40772 15858 40828
rect 15858 40772 15914 40828
rect 15914 40772 15918 40828
rect 15854 40768 15918 40772
rect 21479 40828 21543 40832
rect 21479 40772 21483 40828
rect 21483 40772 21539 40828
rect 21539 40772 21543 40828
rect 21479 40768 21543 40772
rect 21559 40828 21623 40832
rect 21559 40772 21563 40828
rect 21563 40772 21619 40828
rect 21619 40772 21623 40828
rect 21559 40768 21623 40772
rect 21639 40828 21703 40832
rect 21639 40772 21643 40828
rect 21643 40772 21699 40828
rect 21699 40772 21703 40828
rect 21639 40768 21703 40772
rect 21719 40828 21783 40832
rect 21719 40772 21723 40828
rect 21723 40772 21779 40828
rect 21779 40772 21783 40828
rect 21719 40768 21783 40772
rect 2636 40292 2700 40356
rect 6816 40284 6880 40288
rect 6816 40228 6820 40284
rect 6820 40228 6876 40284
rect 6876 40228 6880 40284
rect 6816 40224 6880 40228
rect 6896 40284 6960 40288
rect 6896 40228 6900 40284
rect 6900 40228 6956 40284
rect 6956 40228 6960 40284
rect 6896 40224 6960 40228
rect 6976 40284 7040 40288
rect 6976 40228 6980 40284
rect 6980 40228 7036 40284
rect 7036 40228 7040 40284
rect 6976 40224 7040 40228
rect 7056 40284 7120 40288
rect 7056 40228 7060 40284
rect 7060 40228 7116 40284
rect 7116 40228 7120 40284
rect 7056 40224 7120 40228
rect 12681 40284 12745 40288
rect 12681 40228 12685 40284
rect 12685 40228 12741 40284
rect 12741 40228 12745 40284
rect 12681 40224 12745 40228
rect 12761 40284 12825 40288
rect 12761 40228 12765 40284
rect 12765 40228 12821 40284
rect 12821 40228 12825 40284
rect 12761 40224 12825 40228
rect 12841 40284 12905 40288
rect 12841 40228 12845 40284
rect 12845 40228 12901 40284
rect 12901 40228 12905 40284
rect 12841 40224 12905 40228
rect 12921 40284 12985 40288
rect 12921 40228 12925 40284
rect 12925 40228 12981 40284
rect 12981 40228 12985 40284
rect 12921 40224 12985 40228
rect 18546 40284 18610 40288
rect 18546 40228 18550 40284
rect 18550 40228 18606 40284
rect 18606 40228 18610 40284
rect 18546 40224 18610 40228
rect 18626 40284 18690 40288
rect 18626 40228 18630 40284
rect 18630 40228 18686 40284
rect 18686 40228 18690 40284
rect 18626 40224 18690 40228
rect 18706 40284 18770 40288
rect 18706 40228 18710 40284
rect 18710 40228 18766 40284
rect 18766 40228 18770 40284
rect 18706 40224 18770 40228
rect 18786 40284 18850 40288
rect 18786 40228 18790 40284
rect 18790 40228 18846 40284
rect 18846 40228 18850 40284
rect 18786 40224 18850 40228
rect 24411 40284 24475 40288
rect 24411 40228 24415 40284
rect 24415 40228 24471 40284
rect 24471 40228 24475 40284
rect 24411 40224 24475 40228
rect 24491 40284 24555 40288
rect 24491 40228 24495 40284
rect 24495 40228 24551 40284
rect 24551 40228 24555 40284
rect 24491 40224 24555 40228
rect 24571 40284 24635 40288
rect 24571 40228 24575 40284
rect 24575 40228 24631 40284
rect 24631 40228 24635 40284
rect 24571 40224 24635 40228
rect 24651 40284 24715 40288
rect 24651 40228 24655 40284
rect 24655 40228 24711 40284
rect 24711 40228 24715 40284
rect 24651 40224 24715 40228
rect 612 40020 676 40084
rect 4844 40020 4908 40084
rect 13308 39884 13372 39948
rect 21956 39748 22020 39812
rect 3884 39740 3948 39744
rect 3884 39684 3888 39740
rect 3888 39684 3944 39740
rect 3944 39684 3948 39740
rect 3884 39680 3948 39684
rect 3964 39740 4028 39744
rect 3964 39684 3968 39740
rect 3968 39684 4024 39740
rect 4024 39684 4028 39740
rect 3964 39680 4028 39684
rect 4044 39740 4108 39744
rect 4044 39684 4048 39740
rect 4048 39684 4104 39740
rect 4104 39684 4108 39740
rect 4044 39680 4108 39684
rect 4124 39740 4188 39744
rect 4124 39684 4128 39740
rect 4128 39684 4184 39740
rect 4184 39684 4188 39740
rect 4124 39680 4188 39684
rect 9749 39740 9813 39744
rect 9749 39684 9753 39740
rect 9753 39684 9809 39740
rect 9809 39684 9813 39740
rect 9749 39680 9813 39684
rect 9829 39740 9893 39744
rect 9829 39684 9833 39740
rect 9833 39684 9889 39740
rect 9889 39684 9893 39740
rect 9829 39680 9893 39684
rect 9909 39740 9973 39744
rect 9909 39684 9913 39740
rect 9913 39684 9969 39740
rect 9969 39684 9973 39740
rect 9909 39680 9973 39684
rect 9989 39740 10053 39744
rect 9989 39684 9993 39740
rect 9993 39684 10049 39740
rect 10049 39684 10053 39740
rect 9989 39680 10053 39684
rect 15614 39740 15678 39744
rect 15614 39684 15618 39740
rect 15618 39684 15674 39740
rect 15674 39684 15678 39740
rect 15614 39680 15678 39684
rect 15694 39740 15758 39744
rect 15694 39684 15698 39740
rect 15698 39684 15754 39740
rect 15754 39684 15758 39740
rect 15694 39680 15758 39684
rect 15774 39740 15838 39744
rect 15774 39684 15778 39740
rect 15778 39684 15834 39740
rect 15834 39684 15838 39740
rect 15774 39680 15838 39684
rect 15854 39740 15918 39744
rect 15854 39684 15858 39740
rect 15858 39684 15914 39740
rect 15914 39684 15918 39740
rect 15854 39680 15918 39684
rect 21479 39740 21543 39744
rect 21479 39684 21483 39740
rect 21483 39684 21539 39740
rect 21539 39684 21543 39740
rect 21479 39680 21543 39684
rect 21559 39740 21623 39744
rect 21559 39684 21563 39740
rect 21563 39684 21619 39740
rect 21619 39684 21623 39740
rect 21559 39680 21623 39684
rect 21639 39740 21703 39744
rect 21639 39684 21643 39740
rect 21643 39684 21699 39740
rect 21699 39684 21703 39740
rect 21639 39680 21703 39684
rect 21719 39740 21783 39744
rect 21719 39684 21723 39740
rect 21723 39684 21779 39740
rect 21779 39684 21783 39740
rect 21719 39680 21783 39684
rect 1164 39612 1228 39676
rect 19380 39476 19444 39540
rect 3740 39204 3804 39268
rect 5212 39204 5276 39268
rect 21036 39340 21100 39404
rect 6816 39196 6880 39200
rect 6816 39140 6820 39196
rect 6820 39140 6876 39196
rect 6876 39140 6880 39196
rect 6816 39136 6880 39140
rect 6896 39196 6960 39200
rect 6896 39140 6900 39196
rect 6900 39140 6956 39196
rect 6956 39140 6960 39196
rect 6896 39136 6960 39140
rect 6976 39196 7040 39200
rect 6976 39140 6980 39196
rect 6980 39140 7036 39196
rect 7036 39140 7040 39196
rect 6976 39136 7040 39140
rect 7056 39196 7120 39200
rect 7056 39140 7060 39196
rect 7060 39140 7116 39196
rect 7116 39140 7120 39196
rect 7056 39136 7120 39140
rect 12681 39196 12745 39200
rect 12681 39140 12685 39196
rect 12685 39140 12741 39196
rect 12741 39140 12745 39196
rect 12681 39136 12745 39140
rect 12761 39196 12825 39200
rect 12761 39140 12765 39196
rect 12765 39140 12821 39196
rect 12821 39140 12825 39196
rect 12761 39136 12825 39140
rect 12841 39196 12905 39200
rect 12841 39140 12845 39196
rect 12845 39140 12901 39196
rect 12901 39140 12905 39196
rect 12841 39136 12905 39140
rect 12921 39196 12985 39200
rect 12921 39140 12925 39196
rect 12925 39140 12981 39196
rect 12981 39140 12985 39196
rect 12921 39136 12985 39140
rect 18546 39196 18610 39200
rect 18546 39140 18550 39196
rect 18550 39140 18606 39196
rect 18606 39140 18610 39196
rect 18546 39136 18610 39140
rect 18626 39196 18690 39200
rect 18626 39140 18630 39196
rect 18630 39140 18686 39196
rect 18686 39140 18690 39196
rect 18626 39136 18690 39140
rect 18706 39196 18770 39200
rect 18706 39140 18710 39196
rect 18710 39140 18766 39196
rect 18766 39140 18770 39196
rect 18706 39136 18770 39140
rect 18786 39196 18850 39200
rect 18786 39140 18790 39196
rect 18790 39140 18846 39196
rect 18846 39140 18850 39196
rect 18786 39136 18850 39140
rect 24411 39196 24475 39200
rect 24411 39140 24415 39196
rect 24415 39140 24471 39196
rect 24471 39140 24475 39196
rect 24411 39136 24475 39140
rect 24491 39196 24555 39200
rect 24491 39140 24495 39196
rect 24495 39140 24551 39196
rect 24551 39140 24555 39196
rect 24491 39136 24555 39140
rect 24571 39196 24635 39200
rect 24571 39140 24575 39196
rect 24575 39140 24631 39196
rect 24631 39140 24635 39196
rect 24571 39136 24635 39140
rect 24651 39196 24715 39200
rect 24651 39140 24655 39196
rect 24655 39140 24711 39196
rect 24711 39140 24715 39196
rect 24651 39136 24715 39140
rect 6316 39068 6380 39132
rect 3740 38932 3804 38996
rect 796 38796 860 38860
rect 11468 38660 11532 38724
rect 3884 38652 3948 38656
rect 3884 38596 3888 38652
rect 3888 38596 3944 38652
rect 3944 38596 3948 38652
rect 3884 38592 3948 38596
rect 3964 38652 4028 38656
rect 3964 38596 3968 38652
rect 3968 38596 4024 38652
rect 4024 38596 4028 38652
rect 3964 38592 4028 38596
rect 4044 38652 4108 38656
rect 4044 38596 4048 38652
rect 4048 38596 4104 38652
rect 4104 38596 4108 38652
rect 4044 38592 4108 38596
rect 4124 38652 4188 38656
rect 4124 38596 4128 38652
rect 4128 38596 4184 38652
rect 4184 38596 4188 38652
rect 4124 38592 4188 38596
rect 9749 38652 9813 38656
rect 9749 38596 9753 38652
rect 9753 38596 9809 38652
rect 9809 38596 9813 38652
rect 9749 38592 9813 38596
rect 9829 38652 9893 38656
rect 9829 38596 9833 38652
rect 9833 38596 9889 38652
rect 9889 38596 9893 38652
rect 9829 38592 9893 38596
rect 9909 38652 9973 38656
rect 9909 38596 9913 38652
rect 9913 38596 9969 38652
rect 9969 38596 9973 38652
rect 9909 38592 9973 38596
rect 9989 38652 10053 38656
rect 9989 38596 9993 38652
rect 9993 38596 10049 38652
rect 10049 38596 10053 38652
rect 9989 38592 10053 38596
rect 15614 38652 15678 38656
rect 15614 38596 15618 38652
rect 15618 38596 15674 38652
rect 15674 38596 15678 38652
rect 15614 38592 15678 38596
rect 15694 38652 15758 38656
rect 15694 38596 15698 38652
rect 15698 38596 15754 38652
rect 15754 38596 15758 38652
rect 15694 38592 15758 38596
rect 15774 38652 15838 38656
rect 15774 38596 15778 38652
rect 15778 38596 15834 38652
rect 15834 38596 15838 38652
rect 15774 38592 15838 38596
rect 15854 38652 15918 38656
rect 15854 38596 15858 38652
rect 15858 38596 15914 38652
rect 15914 38596 15918 38652
rect 15854 38592 15918 38596
rect 21479 38652 21543 38656
rect 21479 38596 21483 38652
rect 21483 38596 21539 38652
rect 21539 38596 21543 38652
rect 21479 38592 21543 38596
rect 21559 38652 21623 38656
rect 21559 38596 21563 38652
rect 21563 38596 21619 38652
rect 21619 38596 21623 38652
rect 21559 38592 21623 38596
rect 21639 38652 21703 38656
rect 21639 38596 21643 38652
rect 21643 38596 21699 38652
rect 21699 38596 21703 38652
rect 21639 38592 21703 38596
rect 21719 38652 21783 38656
rect 21719 38596 21723 38652
rect 21723 38596 21779 38652
rect 21779 38596 21783 38652
rect 21719 38592 21783 38596
rect 3556 38388 3620 38452
rect 2452 38252 2516 38316
rect 3372 38116 3436 38180
rect 4292 38116 4356 38180
rect 6816 38108 6880 38112
rect 6816 38052 6820 38108
rect 6820 38052 6876 38108
rect 6876 38052 6880 38108
rect 6816 38048 6880 38052
rect 6896 38108 6960 38112
rect 6896 38052 6900 38108
rect 6900 38052 6956 38108
rect 6956 38052 6960 38108
rect 6896 38048 6960 38052
rect 6976 38108 7040 38112
rect 6976 38052 6980 38108
rect 6980 38052 7036 38108
rect 7036 38052 7040 38108
rect 6976 38048 7040 38052
rect 7056 38108 7120 38112
rect 7056 38052 7060 38108
rect 7060 38052 7116 38108
rect 7116 38052 7120 38108
rect 7056 38048 7120 38052
rect 12681 38108 12745 38112
rect 12681 38052 12685 38108
rect 12685 38052 12741 38108
rect 12741 38052 12745 38108
rect 12681 38048 12745 38052
rect 12761 38108 12825 38112
rect 12761 38052 12765 38108
rect 12765 38052 12821 38108
rect 12821 38052 12825 38108
rect 12761 38048 12825 38052
rect 12841 38108 12905 38112
rect 12841 38052 12845 38108
rect 12845 38052 12901 38108
rect 12901 38052 12905 38108
rect 12841 38048 12905 38052
rect 12921 38108 12985 38112
rect 12921 38052 12925 38108
rect 12925 38052 12981 38108
rect 12981 38052 12985 38108
rect 12921 38048 12985 38052
rect 18546 38108 18610 38112
rect 18546 38052 18550 38108
rect 18550 38052 18606 38108
rect 18606 38052 18610 38108
rect 18546 38048 18610 38052
rect 18626 38108 18690 38112
rect 18626 38052 18630 38108
rect 18630 38052 18686 38108
rect 18686 38052 18690 38108
rect 18626 38048 18690 38052
rect 18706 38108 18770 38112
rect 18706 38052 18710 38108
rect 18710 38052 18766 38108
rect 18766 38052 18770 38108
rect 18706 38048 18770 38052
rect 18786 38108 18850 38112
rect 18786 38052 18790 38108
rect 18790 38052 18846 38108
rect 18846 38052 18850 38108
rect 18786 38048 18850 38052
rect 24411 38108 24475 38112
rect 24411 38052 24415 38108
rect 24415 38052 24471 38108
rect 24471 38052 24475 38108
rect 24411 38048 24475 38052
rect 24491 38108 24555 38112
rect 24491 38052 24495 38108
rect 24495 38052 24551 38108
rect 24551 38052 24555 38108
rect 24491 38048 24555 38052
rect 24571 38108 24635 38112
rect 24571 38052 24575 38108
rect 24575 38052 24631 38108
rect 24631 38052 24635 38108
rect 24571 38048 24635 38052
rect 24651 38108 24715 38112
rect 24651 38052 24655 38108
rect 24655 38052 24711 38108
rect 24711 38052 24715 38108
rect 24651 38048 24715 38052
rect 3884 37564 3948 37568
rect 3884 37508 3888 37564
rect 3888 37508 3944 37564
rect 3944 37508 3948 37564
rect 3884 37504 3948 37508
rect 3964 37564 4028 37568
rect 3964 37508 3968 37564
rect 3968 37508 4024 37564
rect 4024 37508 4028 37564
rect 3964 37504 4028 37508
rect 4044 37564 4108 37568
rect 4044 37508 4048 37564
rect 4048 37508 4104 37564
rect 4104 37508 4108 37564
rect 4044 37504 4108 37508
rect 4124 37564 4188 37568
rect 4124 37508 4128 37564
rect 4128 37508 4184 37564
rect 4184 37508 4188 37564
rect 4124 37504 4188 37508
rect 9749 37564 9813 37568
rect 9749 37508 9753 37564
rect 9753 37508 9809 37564
rect 9809 37508 9813 37564
rect 9749 37504 9813 37508
rect 9829 37564 9893 37568
rect 9829 37508 9833 37564
rect 9833 37508 9889 37564
rect 9889 37508 9893 37564
rect 9829 37504 9893 37508
rect 9909 37564 9973 37568
rect 9909 37508 9913 37564
rect 9913 37508 9969 37564
rect 9969 37508 9973 37564
rect 9909 37504 9973 37508
rect 9989 37564 10053 37568
rect 9989 37508 9993 37564
rect 9993 37508 10049 37564
rect 10049 37508 10053 37564
rect 9989 37504 10053 37508
rect 15614 37564 15678 37568
rect 15614 37508 15618 37564
rect 15618 37508 15674 37564
rect 15674 37508 15678 37564
rect 15614 37504 15678 37508
rect 15694 37564 15758 37568
rect 15694 37508 15698 37564
rect 15698 37508 15754 37564
rect 15754 37508 15758 37564
rect 15694 37504 15758 37508
rect 15774 37564 15838 37568
rect 15774 37508 15778 37564
rect 15778 37508 15834 37564
rect 15834 37508 15838 37564
rect 15774 37504 15838 37508
rect 15854 37564 15918 37568
rect 15854 37508 15858 37564
rect 15858 37508 15914 37564
rect 15914 37508 15918 37564
rect 15854 37504 15918 37508
rect 21479 37564 21543 37568
rect 21479 37508 21483 37564
rect 21483 37508 21539 37564
rect 21539 37508 21543 37564
rect 21479 37504 21543 37508
rect 21559 37564 21623 37568
rect 21559 37508 21563 37564
rect 21563 37508 21619 37564
rect 21619 37508 21623 37564
rect 21559 37504 21623 37508
rect 21639 37564 21703 37568
rect 21639 37508 21643 37564
rect 21643 37508 21699 37564
rect 21699 37508 21703 37564
rect 21639 37504 21703 37508
rect 21719 37564 21783 37568
rect 21719 37508 21723 37564
rect 21723 37508 21779 37564
rect 21779 37508 21783 37564
rect 21719 37504 21783 37508
rect 5396 37436 5460 37500
rect 13676 37300 13740 37364
rect 4660 37028 4724 37092
rect 6816 37020 6880 37024
rect 6816 36964 6820 37020
rect 6820 36964 6876 37020
rect 6876 36964 6880 37020
rect 6816 36960 6880 36964
rect 6896 37020 6960 37024
rect 6896 36964 6900 37020
rect 6900 36964 6956 37020
rect 6956 36964 6960 37020
rect 6896 36960 6960 36964
rect 6976 37020 7040 37024
rect 6976 36964 6980 37020
rect 6980 36964 7036 37020
rect 7036 36964 7040 37020
rect 6976 36960 7040 36964
rect 7056 37020 7120 37024
rect 7056 36964 7060 37020
rect 7060 36964 7116 37020
rect 7116 36964 7120 37020
rect 7056 36960 7120 36964
rect 12681 37020 12745 37024
rect 12681 36964 12685 37020
rect 12685 36964 12741 37020
rect 12741 36964 12745 37020
rect 12681 36960 12745 36964
rect 12761 37020 12825 37024
rect 12761 36964 12765 37020
rect 12765 36964 12821 37020
rect 12821 36964 12825 37020
rect 12761 36960 12825 36964
rect 12841 37020 12905 37024
rect 12841 36964 12845 37020
rect 12845 36964 12901 37020
rect 12901 36964 12905 37020
rect 12841 36960 12905 36964
rect 12921 37020 12985 37024
rect 12921 36964 12925 37020
rect 12925 36964 12981 37020
rect 12981 36964 12985 37020
rect 12921 36960 12985 36964
rect 18546 37020 18610 37024
rect 18546 36964 18550 37020
rect 18550 36964 18606 37020
rect 18606 36964 18610 37020
rect 18546 36960 18610 36964
rect 18626 37020 18690 37024
rect 18626 36964 18630 37020
rect 18630 36964 18686 37020
rect 18686 36964 18690 37020
rect 18626 36960 18690 36964
rect 18706 37020 18770 37024
rect 18706 36964 18710 37020
rect 18710 36964 18766 37020
rect 18766 36964 18770 37020
rect 18706 36960 18770 36964
rect 18786 37020 18850 37024
rect 18786 36964 18790 37020
rect 18790 36964 18846 37020
rect 18846 36964 18850 37020
rect 18786 36960 18850 36964
rect 24411 37020 24475 37024
rect 24411 36964 24415 37020
rect 24415 36964 24471 37020
rect 24471 36964 24475 37020
rect 24411 36960 24475 36964
rect 24491 37020 24555 37024
rect 24491 36964 24495 37020
rect 24495 36964 24551 37020
rect 24551 36964 24555 37020
rect 24491 36960 24555 36964
rect 24571 37020 24635 37024
rect 24571 36964 24575 37020
rect 24575 36964 24631 37020
rect 24631 36964 24635 37020
rect 24571 36960 24635 36964
rect 24651 37020 24715 37024
rect 24651 36964 24655 37020
rect 24655 36964 24711 37020
rect 24711 36964 24715 37020
rect 24651 36960 24715 36964
rect 3740 36756 3804 36820
rect 4476 36484 4540 36548
rect 3884 36476 3948 36480
rect 3884 36420 3888 36476
rect 3888 36420 3944 36476
rect 3944 36420 3948 36476
rect 3884 36416 3948 36420
rect 3964 36476 4028 36480
rect 3964 36420 3968 36476
rect 3968 36420 4024 36476
rect 4024 36420 4028 36476
rect 3964 36416 4028 36420
rect 4044 36476 4108 36480
rect 4044 36420 4048 36476
rect 4048 36420 4104 36476
rect 4104 36420 4108 36476
rect 4044 36416 4108 36420
rect 4124 36476 4188 36480
rect 4124 36420 4128 36476
rect 4128 36420 4184 36476
rect 4184 36420 4188 36476
rect 4124 36416 4188 36420
rect 9749 36476 9813 36480
rect 9749 36420 9753 36476
rect 9753 36420 9809 36476
rect 9809 36420 9813 36476
rect 9749 36416 9813 36420
rect 9829 36476 9893 36480
rect 9829 36420 9833 36476
rect 9833 36420 9889 36476
rect 9889 36420 9893 36476
rect 9829 36416 9893 36420
rect 9909 36476 9973 36480
rect 9909 36420 9913 36476
rect 9913 36420 9969 36476
rect 9969 36420 9973 36476
rect 9909 36416 9973 36420
rect 9989 36476 10053 36480
rect 9989 36420 9993 36476
rect 9993 36420 10049 36476
rect 10049 36420 10053 36476
rect 9989 36416 10053 36420
rect 15614 36476 15678 36480
rect 15614 36420 15618 36476
rect 15618 36420 15674 36476
rect 15674 36420 15678 36476
rect 15614 36416 15678 36420
rect 15694 36476 15758 36480
rect 15694 36420 15698 36476
rect 15698 36420 15754 36476
rect 15754 36420 15758 36476
rect 15694 36416 15758 36420
rect 15774 36476 15838 36480
rect 15774 36420 15778 36476
rect 15778 36420 15834 36476
rect 15834 36420 15838 36476
rect 15774 36416 15838 36420
rect 15854 36476 15918 36480
rect 15854 36420 15858 36476
rect 15858 36420 15914 36476
rect 15914 36420 15918 36476
rect 15854 36416 15918 36420
rect 21479 36476 21543 36480
rect 21479 36420 21483 36476
rect 21483 36420 21539 36476
rect 21539 36420 21543 36476
rect 21479 36416 21543 36420
rect 21559 36476 21623 36480
rect 21559 36420 21563 36476
rect 21563 36420 21619 36476
rect 21619 36420 21623 36476
rect 21559 36416 21623 36420
rect 21639 36476 21703 36480
rect 21639 36420 21643 36476
rect 21643 36420 21699 36476
rect 21699 36420 21703 36476
rect 21639 36416 21703 36420
rect 21719 36476 21783 36480
rect 21719 36420 21723 36476
rect 21723 36420 21779 36476
rect 21779 36420 21783 36476
rect 21719 36416 21783 36420
rect 3556 36212 3620 36276
rect 3556 36076 3620 36140
rect 10180 36076 10244 36140
rect 6816 35932 6880 35936
rect 6816 35876 6820 35932
rect 6820 35876 6876 35932
rect 6876 35876 6880 35932
rect 6816 35872 6880 35876
rect 6896 35932 6960 35936
rect 6896 35876 6900 35932
rect 6900 35876 6956 35932
rect 6956 35876 6960 35932
rect 6896 35872 6960 35876
rect 6976 35932 7040 35936
rect 6976 35876 6980 35932
rect 6980 35876 7036 35932
rect 7036 35876 7040 35932
rect 6976 35872 7040 35876
rect 7056 35932 7120 35936
rect 7056 35876 7060 35932
rect 7060 35876 7116 35932
rect 7116 35876 7120 35932
rect 7056 35872 7120 35876
rect 12681 35932 12745 35936
rect 12681 35876 12685 35932
rect 12685 35876 12741 35932
rect 12741 35876 12745 35932
rect 12681 35872 12745 35876
rect 12761 35932 12825 35936
rect 12761 35876 12765 35932
rect 12765 35876 12821 35932
rect 12821 35876 12825 35932
rect 12761 35872 12825 35876
rect 12841 35932 12905 35936
rect 12841 35876 12845 35932
rect 12845 35876 12901 35932
rect 12901 35876 12905 35932
rect 12841 35872 12905 35876
rect 12921 35932 12985 35936
rect 12921 35876 12925 35932
rect 12925 35876 12981 35932
rect 12981 35876 12985 35932
rect 12921 35872 12985 35876
rect 18546 35932 18610 35936
rect 18546 35876 18550 35932
rect 18550 35876 18606 35932
rect 18606 35876 18610 35932
rect 18546 35872 18610 35876
rect 18626 35932 18690 35936
rect 18626 35876 18630 35932
rect 18630 35876 18686 35932
rect 18686 35876 18690 35932
rect 18626 35872 18690 35876
rect 18706 35932 18770 35936
rect 18706 35876 18710 35932
rect 18710 35876 18766 35932
rect 18766 35876 18770 35932
rect 18706 35872 18770 35876
rect 18786 35932 18850 35936
rect 18786 35876 18790 35932
rect 18790 35876 18846 35932
rect 18846 35876 18850 35932
rect 18786 35872 18850 35876
rect 24411 35932 24475 35936
rect 24411 35876 24415 35932
rect 24415 35876 24471 35932
rect 24471 35876 24475 35932
rect 24411 35872 24475 35876
rect 24491 35932 24555 35936
rect 24491 35876 24495 35932
rect 24495 35876 24551 35932
rect 24551 35876 24555 35932
rect 24491 35872 24555 35876
rect 24571 35932 24635 35936
rect 24571 35876 24575 35932
rect 24575 35876 24631 35932
rect 24631 35876 24635 35932
rect 24571 35872 24635 35876
rect 24651 35932 24715 35936
rect 24651 35876 24655 35932
rect 24655 35876 24711 35932
rect 24711 35876 24715 35932
rect 24651 35872 24715 35876
rect 5212 35728 5276 35732
rect 5212 35672 5262 35728
rect 5262 35672 5276 35728
rect 5212 35668 5276 35672
rect 5948 35668 6012 35732
rect 22508 35532 22572 35596
rect 3884 35388 3948 35392
rect 3884 35332 3888 35388
rect 3888 35332 3944 35388
rect 3944 35332 3948 35388
rect 3884 35328 3948 35332
rect 3964 35388 4028 35392
rect 3964 35332 3968 35388
rect 3968 35332 4024 35388
rect 4024 35332 4028 35388
rect 3964 35328 4028 35332
rect 4044 35388 4108 35392
rect 4044 35332 4048 35388
rect 4048 35332 4104 35388
rect 4104 35332 4108 35388
rect 4044 35328 4108 35332
rect 4124 35388 4188 35392
rect 4124 35332 4128 35388
rect 4128 35332 4184 35388
rect 4184 35332 4188 35388
rect 4124 35328 4188 35332
rect 9749 35388 9813 35392
rect 9749 35332 9753 35388
rect 9753 35332 9809 35388
rect 9809 35332 9813 35388
rect 9749 35328 9813 35332
rect 9829 35388 9893 35392
rect 9829 35332 9833 35388
rect 9833 35332 9889 35388
rect 9889 35332 9893 35388
rect 9829 35328 9893 35332
rect 9909 35388 9973 35392
rect 9909 35332 9913 35388
rect 9913 35332 9969 35388
rect 9969 35332 9973 35388
rect 9909 35328 9973 35332
rect 9989 35388 10053 35392
rect 9989 35332 9993 35388
rect 9993 35332 10049 35388
rect 10049 35332 10053 35388
rect 9989 35328 10053 35332
rect 15614 35388 15678 35392
rect 15614 35332 15618 35388
rect 15618 35332 15674 35388
rect 15674 35332 15678 35388
rect 15614 35328 15678 35332
rect 15694 35388 15758 35392
rect 15694 35332 15698 35388
rect 15698 35332 15754 35388
rect 15754 35332 15758 35388
rect 15694 35328 15758 35332
rect 15774 35388 15838 35392
rect 15774 35332 15778 35388
rect 15778 35332 15834 35388
rect 15834 35332 15838 35388
rect 15774 35328 15838 35332
rect 15854 35388 15918 35392
rect 15854 35332 15858 35388
rect 15858 35332 15914 35388
rect 15914 35332 15918 35388
rect 15854 35328 15918 35332
rect 21479 35388 21543 35392
rect 21479 35332 21483 35388
rect 21483 35332 21539 35388
rect 21539 35332 21543 35388
rect 21479 35328 21543 35332
rect 21559 35388 21623 35392
rect 21559 35332 21563 35388
rect 21563 35332 21619 35388
rect 21619 35332 21623 35388
rect 21559 35328 21623 35332
rect 21639 35388 21703 35392
rect 21639 35332 21643 35388
rect 21643 35332 21699 35388
rect 21699 35332 21703 35388
rect 21639 35328 21703 35332
rect 21719 35388 21783 35392
rect 21719 35332 21723 35388
rect 21723 35332 21779 35388
rect 21779 35332 21783 35388
rect 21719 35328 21783 35332
rect 17908 34988 17972 35052
rect 6816 34844 6880 34848
rect 6816 34788 6820 34844
rect 6820 34788 6876 34844
rect 6876 34788 6880 34844
rect 6816 34784 6880 34788
rect 6896 34844 6960 34848
rect 6896 34788 6900 34844
rect 6900 34788 6956 34844
rect 6956 34788 6960 34844
rect 6896 34784 6960 34788
rect 6976 34844 7040 34848
rect 6976 34788 6980 34844
rect 6980 34788 7036 34844
rect 7036 34788 7040 34844
rect 6976 34784 7040 34788
rect 7056 34844 7120 34848
rect 7056 34788 7060 34844
rect 7060 34788 7116 34844
rect 7116 34788 7120 34844
rect 7056 34784 7120 34788
rect 12681 34844 12745 34848
rect 12681 34788 12685 34844
rect 12685 34788 12741 34844
rect 12741 34788 12745 34844
rect 12681 34784 12745 34788
rect 12761 34844 12825 34848
rect 12761 34788 12765 34844
rect 12765 34788 12821 34844
rect 12821 34788 12825 34844
rect 12761 34784 12825 34788
rect 12841 34844 12905 34848
rect 12841 34788 12845 34844
rect 12845 34788 12901 34844
rect 12901 34788 12905 34844
rect 12841 34784 12905 34788
rect 12921 34844 12985 34848
rect 12921 34788 12925 34844
rect 12925 34788 12981 34844
rect 12981 34788 12985 34844
rect 12921 34784 12985 34788
rect 18546 34844 18610 34848
rect 18546 34788 18550 34844
rect 18550 34788 18606 34844
rect 18606 34788 18610 34844
rect 18546 34784 18610 34788
rect 18626 34844 18690 34848
rect 18626 34788 18630 34844
rect 18630 34788 18686 34844
rect 18686 34788 18690 34844
rect 18626 34784 18690 34788
rect 18706 34844 18770 34848
rect 18706 34788 18710 34844
rect 18710 34788 18766 34844
rect 18766 34788 18770 34844
rect 18706 34784 18770 34788
rect 18786 34844 18850 34848
rect 18786 34788 18790 34844
rect 18790 34788 18846 34844
rect 18846 34788 18850 34844
rect 18786 34784 18850 34788
rect 24411 34844 24475 34848
rect 24411 34788 24415 34844
rect 24415 34788 24471 34844
rect 24471 34788 24475 34844
rect 24411 34784 24475 34788
rect 24491 34844 24555 34848
rect 24491 34788 24495 34844
rect 24495 34788 24551 34844
rect 24551 34788 24555 34844
rect 24491 34784 24555 34788
rect 24571 34844 24635 34848
rect 24571 34788 24575 34844
rect 24575 34788 24631 34844
rect 24631 34788 24635 34844
rect 24571 34784 24635 34788
rect 24651 34844 24715 34848
rect 24651 34788 24655 34844
rect 24655 34788 24711 34844
rect 24711 34788 24715 34844
rect 24651 34784 24715 34788
rect 22324 34580 22388 34644
rect 6132 34444 6196 34508
rect 7972 34444 8036 34508
rect 3884 34300 3948 34304
rect 3884 34244 3888 34300
rect 3888 34244 3944 34300
rect 3944 34244 3948 34300
rect 3884 34240 3948 34244
rect 3964 34300 4028 34304
rect 3964 34244 3968 34300
rect 3968 34244 4024 34300
rect 4024 34244 4028 34300
rect 3964 34240 4028 34244
rect 4044 34300 4108 34304
rect 4044 34244 4048 34300
rect 4048 34244 4104 34300
rect 4104 34244 4108 34300
rect 4044 34240 4108 34244
rect 4124 34300 4188 34304
rect 4124 34244 4128 34300
rect 4128 34244 4184 34300
rect 4184 34244 4188 34300
rect 4124 34240 4188 34244
rect 9749 34300 9813 34304
rect 9749 34244 9753 34300
rect 9753 34244 9809 34300
rect 9809 34244 9813 34300
rect 9749 34240 9813 34244
rect 9829 34300 9893 34304
rect 9829 34244 9833 34300
rect 9833 34244 9889 34300
rect 9889 34244 9893 34300
rect 9829 34240 9893 34244
rect 9909 34300 9973 34304
rect 9909 34244 9913 34300
rect 9913 34244 9969 34300
rect 9969 34244 9973 34300
rect 9909 34240 9973 34244
rect 9989 34300 10053 34304
rect 9989 34244 9993 34300
rect 9993 34244 10049 34300
rect 10049 34244 10053 34300
rect 9989 34240 10053 34244
rect 5212 34172 5276 34236
rect 7604 34036 7668 34100
rect 15614 34300 15678 34304
rect 15614 34244 15618 34300
rect 15618 34244 15674 34300
rect 15674 34244 15678 34300
rect 15614 34240 15678 34244
rect 15694 34300 15758 34304
rect 15694 34244 15698 34300
rect 15698 34244 15754 34300
rect 15754 34244 15758 34300
rect 15694 34240 15758 34244
rect 15774 34300 15838 34304
rect 15774 34244 15778 34300
rect 15778 34244 15834 34300
rect 15834 34244 15838 34300
rect 15774 34240 15838 34244
rect 15854 34300 15918 34304
rect 15854 34244 15858 34300
rect 15858 34244 15914 34300
rect 15914 34244 15918 34300
rect 15854 34240 15918 34244
rect 21479 34300 21543 34304
rect 21479 34244 21483 34300
rect 21483 34244 21539 34300
rect 21539 34244 21543 34300
rect 21479 34240 21543 34244
rect 21559 34300 21623 34304
rect 21559 34244 21563 34300
rect 21563 34244 21619 34300
rect 21619 34244 21623 34300
rect 21559 34240 21623 34244
rect 21639 34300 21703 34304
rect 21639 34244 21643 34300
rect 21643 34244 21699 34300
rect 21699 34244 21703 34300
rect 21639 34240 21703 34244
rect 21719 34300 21783 34304
rect 21719 34244 21723 34300
rect 21723 34244 21779 34300
rect 21779 34244 21783 34300
rect 21719 34240 21783 34244
rect 4476 33900 4540 33964
rect 6816 33756 6880 33760
rect 6816 33700 6820 33756
rect 6820 33700 6876 33756
rect 6876 33700 6880 33756
rect 6816 33696 6880 33700
rect 6896 33756 6960 33760
rect 6896 33700 6900 33756
rect 6900 33700 6956 33756
rect 6956 33700 6960 33756
rect 6896 33696 6960 33700
rect 6976 33756 7040 33760
rect 6976 33700 6980 33756
rect 6980 33700 7036 33756
rect 7036 33700 7040 33756
rect 6976 33696 7040 33700
rect 7056 33756 7120 33760
rect 7056 33700 7060 33756
rect 7060 33700 7116 33756
rect 7116 33700 7120 33756
rect 7056 33696 7120 33700
rect 12681 33756 12745 33760
rect 12681 33700 12685 33756
rect 12685 33700 12741 33756
rect 12741 33700 12745 33756
rect 12681 33696 12745 33700
rect 12761 33756 12825 33760
rect 12761 33700 12765 33756
rect 12765 33700 12821 33756
rect 12821 33700 12825 33756
rect 12761 33696 12825 33700
rect 12841 33756 12905 33760
rect 12841 33700 12845 33756
rect 12845 33700 12901 33756
rect 12901 33700 12905 33756
rect 12841 33696 12905 33700
rect 12921 33756 12985 33760
rect 12921 33700 12925 33756
rect 12925 33700 12981 33756
rect 12981 33700 12985 33756
rect 12921 33696 12985 33700
rect 18546 33756 18610 33760
rect 18546 33700 18550 33756
rect 18550 33700 18606 33756
rect 18606 33700 18610 33756
rect 18546 33696 18610 33700
rect 18626 33756 18690 33760
rect 18626 33700 18630 33756
rect 18630 33700 18686 33756
rect 18686 33700 18690 33756
rect 18626 33696 18690 33700
rect 18706 33756 18770 33760
rect 18706 33700 18710 33756
rect 18710 33700 18766 33756
rect 18766 33700 18770 33756
rect 18706 33696 18770 33700
rect 18786 33756 18850 33760
rect 18786 33700 18790 33756
rect 18790 33700 18846 33756
rect 18846 33700 18850 33756
rect 18786 33696 18850 33700
rect 24411 33756 24475 33760
rect 24411 33700 24415 33756
rect 24415 33700 24471 33756
rect 24471 33700 24475 33756
rect 24411 33696 24475 33700
rect 24491 33756 24555 33760
rect 24491 33700 24495 33756
rect 24495 33700 24551 33756
rect 24551 33700 24555 33756
rect 24491 33696 24555 33700
rect 24571 33756 24635 33760
rect 24571 33700 24575 33756
rect 24575 33700 24631 33756
rect 24631 33700 24635 33756
rect 24571 33696 24635 33700
rect 24651 33756 24715 33760
rect 24651 33700 24655 33756
rect 24655 33700 24711 33756
rect 24711 33700 24715 33756
rect 24651 33696 24715 33700
rect 3372 33492 3436 33556
rect 6500 33492 6564 33556
rect 3884 33212 3948 33216
rect 3884 33156 3888 33212
rect 3888 33156 3944 33212
rect 3944 33156 3948 33212
rect 3884 33152 3948 33156
rect 3964 33212 4028 33216
rect 3964 33156 3968 33212
rect 3968 33156 4024 33212
rect 4024 33156 4028 33212
rect 3964 33152 4028 33156
rect 4044 33212 4108 33216
rect 4044 33156 4048 33212
rect 4048 33156 4104 33212
rect 4104 33156 4108 33212
rect 4044 33152 4108 33156
rect 4124 33212 4188 33216
rect 4124 33156 4128 33212
rect 4128 33156 4184 33212
rect 4184 33156 4188 33212
rect 4124 33152 4188 33156
rect 9749 33212 9813 33216
rect 9749 33156 9753 33212
rect 9753 33156 9809 33212
rect 9809 33156 9813 33212
rect 9749 33152 9813 33156
rect 9829 33212 9893 33216
rect 9829 33156 9833 33212
rect 9833 33156 9889 33212
rect 9889 33156 9893 33212
rect 9829 33152 9893 33156
rect 9909 33212 9973 33216
rect 9909 33156 9913 33212
rect 9913 33156 9969 33212
rect 9969 33156 9973 33212
rect 9909 33152 9973 33156
rect 9989 33212 10053 33216
rect 9989 33156 9993 33212
rect 9993 33156 10049 33212
rect 10049 33156 10053 33212
rect 9989 33152 10053 33156
rect 15614 33212 15678 33216
rect 15614 33156 15618 33212
rect 15618 33156 15674 33212
rect 15674 33156 15678 33212
rect 15614 33152 15678 33156
rect 15694 33212 15758 33216
rect 15694 33156 15698 33212
rect 15698 33156 15754 33212
rect 15754 33156 15758 33212
rect 15694 33152 15758 33156
rect 15774 33212 15838 33216
rect 15774 33156 15778 33212
rect 15778 33156 15834 33212
rect 15834 33156 15838 33212
rect 15774 33152 15838 33156
rect 15854 33212 15918 33216
rect 15854 33156 15858 33212
rect 15858 33156 15914 33212
rect 15914 33156 15918 33212
rect 15854 33152 15918 33156
rect 21479 33212 21543 33216
rect 21479 33156 21483 33212
rect 21483 33156 21539 33212
rect 21539 33156 21543 33212
rect 21479 33152 21543 33156
rect 21559 33212 21623 33216
rect 21559 33156 21563 33212
rect 21563 33156 21619 33212
rect 21619 33156 21623 33212
rect 21559 33152 21623 33156
rect 21639 33212 21703 33216
rect 21639 33156 21643 33212
rect 21643 33156 21699 33212
rect 21699 33156 21703 33212
rect 21639 33152 21703 33156
rect 21719 33212 21783 33216
rect 21719 33156 21723 33212
rect 21723 33156 21779 33212
rect 21779 33156 21783 33212
rect 21719 33152 21783 33156
rect 3740 33084 3804 33148
rect 4292 33084 4356 33148
rect 6132 33084 6196 33148
rect 2084 32812 2148 32876
rect 6816 32668 6880 32672
rect 6816 32612 6820 32668
rect 6820 32612 6876 32668
rect 6876 32612 6880 32668
rect 6816 32608 6880 32612
rect 6896 32668 6960 32672
rect 6896 32612 6900 32668
rect 6900 32612 6956 32668
rect 6956 32612 6960 32668
rect 6896 32608 6960 32612
rect 6976 32668 7040 32672
rect 6976 32612 6980 32668
rect 6980 32612 7036 32668
rect 7036 32612 7040 32668
rect 6976 32608 7040 32612
rect 7056 32668 7120 32672
rect 7056 32612 7060 32668
rect 7060 32612 7116 32668
rect 7116 32612 7120 32668
rect 7056 32608 7120 32612
rect 12681 32668 12745 32672
rect 12681 32612 12685 32668
rect 12685 32612 12741 32668
rect 12741 32612 12745 32668
rect 12681 32608 12745 32612
rect 12761 32668 12825 32672
rect 12761 32612 12765 32668
rect 12765 32612 12821 32668
rect 12821 32612 12825 32668
rect 12761 32608 12825 32612
rect 12841 32668 12905 32672
rect 12841 32612 12845 32668
rect 12845 32612 12901 32668
rect 12901 32612 12905 32668
rect 12841 32608 12905 32612
rect 12921 32668 12985 32672
rect 12921 32612 12925 32668
rect 12925 32612 12981 32668
rect 12981 32612 12985 32668
rect 12921 32608 12985 32612
rect 18546 32668 18610 32672
rect 18546 32612 18550 32668
rect 18550 32612 18606 32668
rect 18606 32612 18610 32668
rect 18546 32608 18610 32612
rect 18626 32668 18690 32672
rect 18626 32612 18630 32668
rect 18630 32612 18686 32668
rect 18686 32612 18690 32668
rect 18626 32608 18690 32612
rect 18706 32668 18770 32672
rect 18706 32612 18710 32668
rect 18710 32612 18766 32668
rect 18766 32612 18770 32668
rect 18706 32608 18770 32612
rect 18786 32668 18850 32672
rect 18786 32612 18790 32668
rect 18790 32612 18846 32668
rect 18846 32612 18850 32668
rect 18786 32608 18850 32612
rect 24411 32668 24475 32672
rect 24411 32612 24415 32668
rect 24415 32612 24471 32668
rect 24471 32612 24475 32668
rect 24411 32608 24475 32612
rect 24491 32668 24555 32672
rect 24491 32612 24495 32668
rect 24495 32612 24551 32668
rect 24551 32612 24555 32668
rect 24491 32608 24555 32612
rect 24571 32668 24635 32672
rect 24571 32612 24575 32668
rect 24575 32612 24631 32668
rect 24631 32612 24635 32668
rect 24571 32608 24635 32612
rect 24651 32668 24715 32672
rect 24651 32612 24655 32668
rect 24655 32612 24711 32668
rect 24711 32612 24715 32668
rect 24651 32608 24715 32612
rect 10180 32540 10244 32604
rect 7788 32464 7852 32468
rect 7788 32408 7802 32464
rect 7802 32408 7852 32464
rect 7788 32404 7852 32408
rect 2452 32268 2516 32332
rect 8156 32268 8220 32332
rect 5948 32132 6012 32196
rect 3884 32124 3948 32128
rect 3884 32068 3888 32124
rect 3888 32068 3944 32124
rect 3944 32068 3948 32124
rect 3884 32064 3948 32068
rect 3964 32124 4028 32128
rect 3964 32068 3968 32124
rect 3968 32068 4024 32124
rect 4024 32068 4028 32124
rect 3964 32064 4028 32068
rect 4044 32124 4108 32128
rect 4044 32068 4048 32124
rect 4048 32068 4104 32124
rect 4104 32068 4108 32124
rect 4044 32064 4108 32068
rect 4124 32124 4188 32128
rect 4124 32068 4128 32124
rect 4128 32068 4184 32124
rect 4184 32068 4188 32124
rect 4124 32064 4188 32068
rect 9749 32124 9813 32128
rect 9749 32068 9753 32124
rect 9753 32068 9809 32124
rect 9809 32068 9813 32124
rect 9749 32064 9813 32068
rect 9829 32124 9893 32128
rect 9829 32068 9833 32124
rect 9833 32068 9889 32124
rect 9889 32068 9893 32124
rect 9829 32064 9893 32068
rect 9909 32124 9973 32128
rect 9909 32068 9913 32124
rect 9913 32068 9969 32124
rect 9969 32068 9973 32124
rect 9909 32064 9973 32068
rect 9989 32124 10053 32128
rect 9989 32068 9993 32124
rect 9993 32068 10049 32124
rect 10049 32068 10053 32124
rect 9989 32064 10053 32068
rect 11100 32268 11164 32332
rect 15614 32124 15678 32128
rect 15614 32068 15618 32124
rect 15618 32068 15674 32124
rect 15674 32068 15678 32124
rect 15614 32064 15678 32068
rect 15694 32124 15758 32128
rect 15694 32068 15698 32124
rect 15698 32068 15754 32124
rect 15754 32068 15758 32124
rect 15694 32064 15758 32068
rect 15774 32124 15838 32128
rect 15774 32068 15778 32124
rect 15778 32068 15834 32124
rect 15834 32068 15838 32124
rect 15774 32064 15838 32068
rect 15854 32124 15918 32128
rect 15854 32068 15858 32124
rect 15858 32068 15914 32124
rect 15914 32068 15918 32124
rect 15854 32064 15918 32068
rect 21479 32124 21543 32128
rect 21479 32068 21483 32124
rect 21483 32068 21539 32124
rect 21539 32068 21543 32124
rect 21479 32064 21543 32068
rect 21559 32124 21623 32128
rect 21559 32068 21563 32124
rect 21563 32068 21619 32124
rect 21619 32068 21623 32124
rect 21559 32064 21623 32068
rect 21639 32124 21703 32128
rect 21639 32068 21643 32124
rect 21643 32068 21699 32124
rect 21699 32068 21703 32124
rect 21639 32064 21703 32068
rect 21719 32124 21783 32128
rect 21719 32068 21723 32124
rect 21723 32068 21779 32124
rect 21779 32068 21783 32124
rect 21719 32064 21783 32068
rect 2820 31724 2884 31788
rect 5580 31724 5644 31788
rect 15148 31860 15212 31924
rect 7604 31648 7668 31652
rect 7604 31592 7654 31648
rect 7654 31592 7668 31648
rect 7604 31588 7668 31592
rect 6816 31580 6880 31584
rect 6816 31524 6820 31580
rect 6820 31524 6876 31580
rect 6876 31524 6880 31580
rect 6816 31520 6880 31524
rect 6896 31580 6960 31584
rect 6896 31524 6900 31580
rect 6900 31524 6956 31580
rect 6956 31524 6960 31580
rect 6896 31520 6960 31524
rect 6976 31580 7040 31584
rect 6976 31524 6980 31580
rect 6980 31524 7036 31580
rect 7036 31524 7040 31580
rect 6976 31520 7040 31524
rect 7056 31580 7120 31584
rect 7056 31524 7060 31580
rect 7060 31524 7116 31580
rect 7116 31524 7120 31580
rect 7056 31520 7120 31524
rect 12681 31580 12745 31584
rect 12681 31524 12685 31580
rect 12685 31524 12741 31580
rect 12741 31524 12745 31580
rect 12681 31520 12745 31524
rect 12761 31580 12825 31584
rect 12761 31524 12765 31580
rect 12765 31524 12821 31580
rect 12821 31524 12825 31580
rect 12761 31520 12825 31524
rect 12841 31580 12905 31584
rect 12841 31524 12845 31580
rect 12845 31524 12901 31580
rect 12901 31524 12905 31580
rect 12841 31520 12905 31524
rect 12921 31580 12985 31584
rect 12921 31524 12925 31580
rect 12925 31524 12981 31580
rect 12981 31524 12985 31580
rect 12921 31520 12985 31524
rect 18546 31580 18610 31584
rect 18546 31524 18550 31580
rect 18550 31524 18606 31580
rect 18606 31524 18610 31580
rect 18546 31520 18610 31524
rect 18626 31580 18690 31584
rect 18626 31524 18630 31580
rect 18630 31524 18686 31580
rect 18686 31524 18690 31580
rect 18626 31520 18690 31524
rect 18706 31580 18770 31584
rect 18706 31524 18710 31580
rect 18710 31524 18766 31580
rect 18766 31524 18770 31580
rect 18706 31520 18770 31524
rect 18786 31580 18850 31584
rect 18786 31524 18790 31580
rect 18790 31524 18846 31580
rect 18846 31524 18850 31580
rect 18786 31520 18850 31524
rect 24411 31580 24475 31584
rect 24411 31524 24415 31580
rect 24415 31524 24471 31580
rect 24471 31524 24475 31580
rect 24411 31520 24475 31524
rect 24491 31580 24555 31584
rect 24491 31524 24495 31580
rect 24495 31524 24551 31580
rect 24551 31524 24555 31580
rect 24491 31520 24555 31524
rect 24571 31580 24635 31584
rect 24571 31524 24575 31580
rect 24575 31524 24631 31580
rect 24631 31524 24635 31580
rect 24571 31520 24635 31524
rect 24651 31580 24715 31584
rect 24651 31524 24655 31580
rect 24655 31524 24711 31580
rect 24711 31524 24715 31580
rect 24651 31520 24715 31524
rect 2636 31452 2700 31516
rect 5580 31512 5644 31516
rect 5580 31456 5594 31512
rect 5594 31456 5644 31512
rect 5580 31452 5644 31456
rect 2636 31316 2700 31380
rect 10180 31180 10244 31244
rect 3884 31036 3948 31040
rect 3884 30980 3888 31036
rect 3888 30980 3944 31036
rect 3944 30980 3948 31036
rect 3884 30976 3948 30980
rect 3964 31036 4028 31040
rect 3964 30980 3968 31036
rect 3968 30980 4024 31036
rect 4024 30980 4028 31036
rect 3964 30976 4028 30980
rect 4044 31036 4108 31040
rect 4044 30980 4048 31036
rect 4048 30980 4104 31036
rect 4104 30980 4108 31036
rect 4044 30976 4108 30980
rect 4124 31036 4188 31040
rect 4124 30980 4128 31036
rect 4128 30980 4184 31036
rect 4184 30980 4188 31036
rect 4124 30976 4188 30980
rect 9749 31036 9813 31040
rect 9749 30980 9753 31036
rect 9753 30980 9809 31036
rect 9809 30980 9813 31036
rect 9749 30976 9813 30980
rect 9829 31036 9893 31040
rect 9829 30980 9833 31036
rect 9833 30980 9889 31036
rect 9889 30980 9893 31036
rect 9829 30976 9893 30980
rect 9909 31036 9973 31040
rect 9909 30980 9913 31036
rect 9913 30980 9969 31036
rect 9969 30980 9973 31036
rect 9909 30976 9973 30980
rect 9989 31036 10053 31040
rect 9989 30980 9993 31036
rect 9993 30980 10049 31036
rect 10049 30980 10053 31036
rect 9989 30976 10053 30980
rect 15614 31036 15678 31040
rect 15614 30980 15618 31036
rect 15618 30980 15674 31036
rect 15674 30980 15678 31036
rect 15614 30976 15678 30980
rect 15694 31036 15758 31040
rect 15694 30980 15698 31036
rect 15698 30980 15754 31036
rect 15754 30980 15758 31036
rect 15694 30976 15758 30980
rect 15774 31036 15838 31040
rect 15774 30980 15778 31036
rect 15778 30980 15834 31036
rect 15834 30980 15838 31036
rect 15774 30976 15838 30980
rect 15854 31036 15918 31040
rect 15854 30980 15858 31036
rect 15858 30980 15914 31036
rect 15914 30980 15918 31036
rect 15854 30976 15918 30980
rect 21479 31036 21543 31040
rect 21479 30980 21483 31036
rect 21483 30980 21539 31036
rect 21539 30980 21543 31036
rect 21479 30976 21543 30980
rect 21559 31036 21623 31040
rect 21559 30980 21563 31036
rect 21563 30980 21619 31036
rect 21619 30980 21623 31036
rect 21559 30976 21623 30980
rect 21639 31036 21703 31040
rect 21639 30980 21643 31036
rect 21643 30980 21699 31036
rect 21699 30980 21703 31036
rect 21639 30976 21703 30980
rect 21719 31036 21783 31040
rect 21719 30980 21723 31036
rect 21723 30980 21779 31036
rect 21779 30980 21783 31036
rect 21719 30976 21783 30980
rect 6816 30492 6880 30496
rect 6816 30436 6820 30492
rect 6820 30436 6876 30492
rect 6876 30436 6880 30492
rect 6816 30432 6880 30436
rect 6896 30492 6960 30496
rect 6896 30436 6900 30492
rect 6900 30436 6956 30492
rect 6956 30436 6960 30492
rect 6896 30432 6960 30436
rect 6976 30492 7040 30496
rect 6976 30436 6980 30492
rect 6980 30436 7036 30492
rect 7036 30436 7040 30492
rect 6976 30432 7040 30436
rect 7056 30492 7120 30496
rect 7056 30436 7060 30492
rect 7060 30436 7116 30492
rect 7116 30436 7120 30492
rect 7056 30432 7120 30436
rect 12681 30492 12745 30496
rect 12681 30436 12685 30492
rect 12685 30436 12741 30492
rect 12741 30436 12745 30492
rect 12681 30432 12745 30436
rect 12761 30492 12825 30496
rect 12761 30436 12765 30492
rect 12765 30436 12821 30492
rect 12821 30436 12825 30492
rect 12761 30432 12825 30436
rect 12841 30492 12905 30496
rect 12841 30436 12845 30492
rect 12845 30436 12901 30492
rect 12901 30436 12905 30492
rect 12841 30432 12905 30436
rect 12921 30492 12985 30496
rect 12921 30436 12925 30492
rect 12925 30436 12981 30492
rect 12981 30436 12985 30492
rect 12921 30432 12985 30436
rect 18546 30492 18610 30496
rect 18546 30436 18550 30492
rect 18550 30436 18606 30492
rect 18606 30436 18610 30492
rect 18546 30432 18610 30436
rect 18626 30492 18690 30496
rect 18626 30436 18630 30492
rect 18630 30436 18686 30492
rect 18686 30436 18690 30492
rect 18626 30432 18690 30436
rect 18706 30492 18770 30496
rect 18706 30436 18710 30492
rect 18710 30436 18766 30492
rect 18766 30436 18770 30492
rect 18706 30432 18770 30436
rect 18786 30492 18850 30496
rect 18786 30436 18790 30492
rect 18790 30436 18846 30492
rect 18846 30436 18850 30492
rect 18786 30432 18850 30436
rect 24411 30492 24475 30496
rect 24411 30436 24415 30492
rect 24415 30436 24471 30492
rect 24471 30436 24475 30492
rect 24411 30432 24475 30436
rect 24491 30492 24555 30496
rect 24491 30436 24495 30492
rect 24495 30436 24551 30492
rect 24551 30436 24555 30492
rect 24491 30432 24555 30436
rect 24571 30492 24635 30496
rect 24571 30436 24575 30492
rect 24575 30436 24631 30492
rect 24631 30436 24635 30492
rect 24571 30432 24635 30436
rect 24651 30492 24715 30496
rect 24651 30436 24655 30492
rect 24655 30436 24711 30492
rect 24711 30436 24715 30492
rect 24651 30432 24715 30436
rect 10180 30364 10244 30428
rect 11468 30364 11532 30428
rect 12020 30364 12084 30428
rect 5212 30228 5276 30292
rect 1532 30092 1596 30156
rect 7972 29956 8036 30020
rect 3884 29948 3948 29952
rect 3884 29892 3888 29948
rect 3888 29892 3944 29948
rect 3944 29892 3948 29948
rect 3884 29888 3948 29892
rect 3964 29948 4028 29952
rect 3964 29892 3968 29948
rect 3968 29892 4024 29948
rect 4024 29892 4028 29948
rect 3964 29888 4028 29892
rect 4044 29948 4108 29952
rect 4044 29892 4048 29948
rect 4048 29892 4104 29948
rect 4104 29892 4108 29948
rect 4044 29888 4108 29892
rect 4124 29948 4188 29952
rect 4124 29892 4128 29948
rect 4128 29892 4184 29948
rect 4184 29892 4188 29948
rect 4124 29888 4188 29892
rect 9749 29948 9813 29952
rect 9749 29892 9753 29948
rect 9753 29892 9809 29948
rect 9809 29892 9813 29948
rect 9749 29888 9813 29892
rect 9829 29948 9893 29952
rect 9829 29892 9833 29948
rect 9833 29892 9889 29948
rect 9889 29892 9893 29948
rect 9829 29888 9893 29892
rect 9909 29948 9973 29952
rect 9909 29892 9913 29948
rect 9913 29892 9969 29948
rect 9969 29892 9973 29948
rect 9909 29888 9973 29892
rect 9989 29948 10053 29952
rect 9989 29892 9993 29948
rect 9993 29892 10049 29948
rect 10049 29892 10053 29948
rect 9989 29888 10053 29892
rect 15614 29948 15678 29952
rect 15614 29892 15618 29948
rect 15618 29892 15674 29948
rect 15674 29892 15678 29948
rect 15614 29888 15678 29892
rect 15694 29948 15758 29952
rect 15694 29892 15698 29948
rect 15698 29892 15754 29948
rect 15754 29892 15758 29948
rect 15694 29888 15758 29892
rect 15774 29948 15838 29952
rect 15774 29892 15778 29948
rect 15778 29892 15834 29948
rect 15834 29892 15838 29948
rect 15774 29888 15838 29892
rect 15854 29948 15918 29952
rect 15854 29892 15858 29948
rect 15858 29892 15914 29948
rect 15914 29892 15918 29948
rect 15854 29888 15918 29892
rect 21479 29948 21543 29952
rect 21479 29892 21483 29948
rect 21483 29892 21539 29948
rect 21539 29892 21543 29948
rect 21479 29888 21543 29892
rect 21559 29948 21623 29952
rect 21559 29892 21563 29948
rect 21563 29892 21619 29948
rect 21619 29892 21623 29948
rect 21559 29888 21623 29892
rect 21639 29948 21703 29952
rect 21639 29892 21643 29948
rect 21643 29892 21699 29948
rect 21699 29892 21703 29948
rect 21639 29888 21703 29892
rect 21719 29948 21783 29952
rect 21719 29892 21723 29948
rect 21723 29892 21779 29948
rect 21779 29892 21783 29948
rect 21719 29888 21783 29892
rect 5028 29820 5092 29884
rect 8708 29820 8772 29884
rect 16436 29548 16500 29612
rect 1716 29412 1780 29476
rect 6816 29404 6880 29408
rect 6816 29348 6820 29404
rect 6820 29348 6876 29404
rect 6876 29348 6880 29404
rect 6816 29344 6880 29348
rect 6896 29404 6960 29408
rect 6896 29348 6900 29404
rect 6900 29348 6956 29404
rect 6956 29348 6960 29404
rect 6896 29344 6960 29348
rect 6976 29404 7040 29408
rect 6976 29348 6980 29404
rect 6980 29348 7036 29404
rect 7036 29348 7040 29404
rect 6976 29344 7040 29348
rect 7056 29404 7120 29408
rect 7056 29348 7060 29404
rect 7060 29348 7116 29404
rect 7116 29348 7120 29404
rect 7056 29344 7120 29348
rect 12681 29404 12745 29408
rect 12681 29348 12685 29404
rect 12685 29348 12741 29404
rect 12741 29348 12745 29404
rect 12681 29344 12745 29348
rect 12761 29404 12825 29408
rect 12761 29348 12765 29404
rect 12765 29348 12821 29404
rect 12821 29348 12825 29404
rect 12761 29344 12825 29348
rect 12841 29404 12905 29408
rect 12841 29348 12845 29404
rect 12845 29348 12901 29404
rect 12901 29348 12905 29404
rect 12841 29344 12905 29348
rect 12921 29404 12985 29408
rect 12921 29348 12925 29404
rect 12925 29348 12981 29404
rect 12981 29348 12985 29404
rect 12921 29344 12985 29348
rect 18546 29404 18610 29408
rect 18546 29348 18550 29404
rect 18550 29348 18606 29404
rect 18606 29348 18610 29404
rect 18546 29344 18610 29348
rect 18626 29404 18690 29408
rect 18626 29348 18630 29404
rect 18630 29348 18686 29404
rect 18686 29348 18690 29404
rect 18626 29344 18690 29348
rect 18706 29404 18770 29408
rect 18706 29348 18710 29404
rect 18710 29348 18766 29404
rect 18766 29348 18770 29404
rect 18706 29344 18770 29348
rect 18786 29404 18850 29408
rect 18786 29348 18790 29404
rect 18790 29348 18846 29404
rect 18846 29348 18850 29404
rect 18786 29344 18850 29348
rect 24411 29404 24475 29408
rect 24411 29348 24415 29404
rect 24415 29348 24471 29404
rect 24471 29348 24475 29404
rect 24411 29344 24475 29348
rect 24491 29404 24555 29408
rect 24491 29348 24495 29404
rect 24495 29348 24551 29404
rect 24551 29348 24555 29404
rect 24491 29344 24555 29348
rect 24571 29404 24635 29408
rect 24571 29348 24575 29404
rect 24575 29348 24631 29404
rect 24631 29348 24635 29404
rect 24571 29344 24635 29348
rect 24651 29404 24715 29408
rect 24651 29348 24655 29404
rect 24655 29348 24711 29404
rect 24711 29348 24715 29404
rect 24651 29344 24715 29348
rect 18092 29140 18156 29204
rect 5580 29004 5644 29068
rect 6500 29004 6564 29068
rect 13124 29004 13188 29068
rect 20852 29004 20916 29068
rect 3884 28860 3948 28864
rect 3884 28804 3888 28860
rect 3888 28804 3944 28860
rect 3944 28804 3948 28860
rect 3884 28800 3948 28804
rect 3964 28860 4028 28864
rect 3964 28804 3968 28860
rect 3968 28804 4024 28860
rect 4024 28804 4028 28860
rect 3964 28800 4028 28804
rect 4044 28860 4108 28864
rect 4044 28804 4048 28860
rect 4048 28804 4104 28860
rect 4104 28804 4108 28860
rect 4044 28800 4108 28804
rect 4124 28860 4188 28864
rect 4124 28804 4128 28860
rect 4128 28804 4184 28860
rect 4184 28804 4188 28860
rect 4124 28800 4188 28804
rect 9749 28860 9813 28864
rect 9749 28804 9753 28860
rect 9753 28804 9809 28860
rect 9809 28804 9813 28860
rect 9749 28800 9813 28804
rect 9829 28860 9893 28864
rect 9829 28804 9833 28860
rect 9833 28804 9889 28860
rect 9889 28804 9893 28860
rect 9829 28800 9893 28804
rect 9909 28860 9973 28864
rect 9909 28804 9913 28860
rect 9913 28804 9969 28860
rect 9969 28804 9973 28860
rect 9909 28800 9973 28804
rect 9989 28860 10053 28864
rect 9989 28804 9993 28860
rect 9993 28804 10049 28860
rect 10049 28804 10053 28860
rect 9989 28800 10053 28804
rect 15614 28860 15678 28864
rect 15614 28804 15618 28860
rect 15618 28804 15674 28860
rect 15674 28804 15678 28860
rect 15614 28800 15678 28804
rect 15694 28860 15758 28864
rect 15694 28804 15698 28860
rect 15698 28804 15754 28860
rect 15754 28804 15758 28860
rect 15694 28800 15758 28804
rect 15774 28860 15838 28864
rect 15774 28804 15778 28860
rect 15778 28804 15834 28860
rect 15834 28804 15838 28860
rect 15774 28800 15838 28804
rect 15854 28860 15918 28864
rect 15854 28804 15858 28860
rect 15858 28804 15914 28860
rect 15914 28804 15918 28860
rect 15854 28800 15918 28804
rect 21479 28860 21543 28864
rect 21479 28804 21483 28860
rect 21483 28804 21539 28860
rect 21539 28804 21543 28860
rect 21479 28800 21543 28804
rect 21559 28860 21623 28864
rect 21559 28804 21563 28860
rect 21563 28804 21619 28860
rect 21619 28804 21623 28860
rect 21559 28800 21623 28804
rect 21639 28860 21703 28864
rect 21639 28804 21643 28860
rect 21643 28804 21699 28860
rect 21699 28804 21703 28860
rect 21639 28800 21703 28804
rect 21719 28860 21783 28864
rect 21719 28804 21723 28860
rect 21723 28804 21779 28860
rect 21779 28804 21783 28860
rect 21719 28800 21783 28804
rect 6316 28460 6380 28524
rect 8708 28460 8772 28524
rect 14044 28460 14108 28524
rect 6816 28316 6880 28320
rect 6816 28260 6820 28316
rect 6820 28260 6876 28316
rect 6876 28260 6880 28316
rect 6816 28256 6880 28260
rect 6896 28316 6960 28320
rect 6896 28260 6900 28316
rect 6900 28260 6956 28316
rect 6956 28260 6960 28316
rect 6896 28256 6960 28260
rect 6976 28316 7040 28320
rect 6976 28260 6980 28316
rect 6980 28260 7036 28316
rect 7036 28260 7040 28316
rect 6976 28256 7040 28260
rect 7056 28316 7120 28320
rect 7056 28260 7060 28316
rect 7060 28260 7116 28316
rect 7116 28260 7120 28316
rect 7056 28256 7120 28260
rect 12681 28316 12745 28320
rect 12681 28260 12685 28316
rect 12685 28260 12741 28316
rect 12741 28260 12745 28316
rect 12681 28256 12745 28260
rect 12761 28316 12825 28320
rect 12761 28260 12765 28316
rect 12765 28260 12821 28316
rect 12821 28260 12825 28316
rect 12761 28256 12825 28260
rect 12841 28316 12905 28320
rect 12841 28260 12845 28316
rect 12845 28260 12901 28316
rect 12901 28260 12905 28316
rect 12841 28256 12905 28260
rect 12921 28316 12985 28320
rect 12921 28260 12925 28316
rect 12925 28260 12981 28316
rect 12981 28260 12985 28316
rect 12921 28256 12985 28260
rect 18546 28316 18610 28320
rect 18546 28260 18550 28316
rect 18550 28260 18606 28316
rect 18606 28260 18610 28316
rect 18546 28256 18610 28260
rect 18626 28316 18690 28320
rect 18626 28260 18630 28316
rect 18630 28260 18686 28316
rect 18686 28260 18690 28316
rect 18626 28256 18690 28260
rect 18706 28316 18770 28320
rect 18706 28260 18710 28316
rect 18710 28260 18766 28316
rect 18766 28260 18770 28316
rect 18706 28256 18770 28260
rect 18786 28316 18850 28320
rect 18786 28260 18790 28316
rect 18790 28260 18846 28316
rect 18846 28260 18850 28316
rect 18786 28256 18850 28260
rect 24411 28316 24475 28320
rect 24411 28260 24415 28316
rect 24415 28260 24471 28316
rect 24471 28260 24475 28316
rect 24411 28256 24475 28260
rect 24491 28316 24555 28320
rect 24491 28260 24495 28316
rect 24495 28260 24551 28316
rect 24551 28260 24555 28316
rect 24491 28256 24555 28260
rect 24571 28316 24635 28320
rect 24571 28260 24575 28316
rect 24575 28260 24631 28316
rect 24631 28260 24635 28316
rect 24571 28256 24635 28260
rect 24651 28316 24715 28320
rect 24651 28260 24655 28316
rect 24655 28260 24711 28316
rect 24711 28260 24715 28316
rect 24651 28256 24715 28260
rect 15148 28052 15212 28116
rect 16252 28052 16316 28116
rect 22692 27916 22756 27980
rect 3884 27772 3948 27776
rect 3884 27716 3888 27772
rect 3888 27716 3944 27772
rect 3944 27716 3948 27772
rect 3884 27712 3948 27716
rect 3964 27772 4028 27776
rect 3964 27716 3968 27772
rect 3968 27716 4024 27772
rect 4024 27716 4028 27772
rect 3964 27712 4028 27716
rect 4044 27772 4108 27776
rect 4044 27716 4048 27772
rect 4048 27716 4104 27772
rect 4104 27716 4108 27772
rect 4044 27712 4108 27716
rect 4124 27772 4188 27776
rect 4124 27716 4128 27772
rect 4128 27716 4184 27772
rect 4184 27716 4188 27772
rect 4124 27712 4188 27716
rect 9749 27772 9813 27776
rect 9749 27716 9753 27772
rect 9753 27716 9809 27772
rect 9809 27716 9813 27772
rect 9749 27712 9813 27716
rect 9829 27772 9893 27776
rect 9829 27716 9833 27772
rect 9833 27716 9889 27772
rect 9889 27716 9893 27772
rect 9829 27712 9893 27716
rect 9909 27772 9973 27776
rect 9909 27716 9913 27772
rect 9913 27716 9969 27772
rect 9969 27716 9973 27772
rect 9909 27712 9973 27716
rect 9989 27772 10053 27776
rect 9989 27716 9993 27772
rect 9993 27716 10049 27772
rect 10049 27716 10053 27772
rect 9989 27712 10053 27716
rect 5764 27644 5828 27708
rect 6132 27644 6196 27708
rect 4292 27508 4356 27572
rect 15614 27772 15678 27776
rect 15614 27716 15618 27772
rect 15618 27716 15674 27772
rect 15674 27716 15678 27772
rect 15614 27712 15678 27716
rect 15694 27772 15758 27776
rect 15694 27716 15698 27772
rect 15698 27716 15754 27772
rect 15754 27716 15758 27772
rect 15694 27712 15758 27716
rect 15774 27772 15838 27776
rect 15774 27716 15778 27772
rect 15778 27716 15834 27772
rect 15834 27716 15838 27772
rect 15774 27712 15838 27716
rect 15854 27772 15918 27776
rect 15854 27716 15858 27772
rect 15858 27716 15914 27772
rect 15914 27716 15918 27772
rect 15854 27712 15918 27716
rect 21479 27772 21543 27776
rect 21479 27716 21483 27772
rect 21483 27716 21539 27772
rect 21539 27716 21543 27772
rect 21479 27712 21543 27716
rect 21559 27772 21623 27776
rect 21559 27716 21563 27772
rect 21563 27716 21619 27772
rect 21619 27716 21623 27772
rect 21559 27712 21623 27716
rect 21639 27772 21703 27776
rect 21639 27716 21643 27772
rect 21643 27716 21699 27772
rect 21699 27716 21703 27772
rect 21639 27712 21703 27716
rect 21719 27772 21783 27776
rect 21719 27716 21723 27772
rect 21723 27716 21779 27772
rect 21779 27716 21783 27772
rect 21719 27712 21783 27716
rect 10548 27508 10612 27572
rect 4660 27236 4724 27300
rect 7604 27236 7668 27300
rect 6816 27228 6880 27232
rect 6816 27172 6820 27228
rect 6820 27172 6876 27228
rect 6876 27172 6880 27228
rect 6816 27168 6880 27172
rect 6896 27228 6960 27232
rect 6896 27172 6900 27228
rect 6900 27172 6956 27228
rect 6956 27172 6960 27228
rect 6896 27168 6960 27172
rect 6976 27228 7040 27232
rect 6976 27172 6980 27228
rect 6980 27172 7036 27228
rect 7036 27172 7040 27228
rect 6976 27168 7040 27172
rect 7056 27228 7120 27232
rect 7056 27172 7060 27228
rect 7060 27172 7116 27228
rect 7116 27172 7120 27228
rect 7056 27168 7120 27172
rect 12681 27228 12745 27232
rect 12681 27172 12685 27228
rect 12685 27172 12741 27228
rect 12741 27172 12745 27228
rect 12681 27168 12745 27172
rect 12761 27228 12825 27232
rect 12761 27172 12765 27228
rect 12765 27172 12821 27228
rect 12821 27172 12825 27228
rect 12761 27168 12825 27172
rect 12841 27228 12905 27232
rect 12841 27172 12845 27228
rect 12845 27172 12901 27228
rect 12901 27172 12905 27228
rect 12841 27168 12905 27172
rect 12921 27228 12985 27232
rect 12921 27172 12925 27228
rect 12925 27172 12981 27228
rect 12981 27172 12985 27228
rect 12921 27168 12985 27172
rect 18546 27228 18610 27232
rect 18546 27172 18550 27228
rect 18550 27172 18606 27228
rect 18606 27172 18610 27228
rect 18546 27168 18610 27172
rect 18626 27228 18690 27232
rect 18626 27172 18630 27228
rect 18630 27172 18686 27228
rect 18686 27172 18690 27228
rect 18626 27168 18690 27172
rect 18706 27228 18770 27232
rect 18706 27172 18710 27228
rect 18710 27172 18766 27228
rect 18766 27172 18770 27228
rect 18706 27168 18770 27172
rect 18786 27228 18850 27232
rect 18786 27172 18790 27228
rect 18790 27172 18846 27228
rect 18846 27172 18850 27228
rect 18786 27168 18850 27172
rect 24411 27228 24475 27232
rect 24411 27172 24415 27228
rect 24415 27172 24471 27228
rect 24471 27172 24475 27228
rect 24411 27168 24475 27172
rect 24491 27228 24555 27232
rect 24491 27172 24495 27228
rect 24495 27172 24551 27228
rect 24551 27172 24555 27228
rect 24491 27168 24555 27172
rect 24571 27228 24635 27232
rect 24571 27172 24575 27228
rect 24575 27172 24631 27228
rect 24631 27172 24635 27228
rect 24571 27168 24635 27172
rect 24651 27228 24715 27232
rect 24651 27172 24655 27228
rect 24655 27172 24711 27228
rect 24711 27172 24715 27228
rect 24651 27168 24715 27172
rect 4476 27100 4540 27164
rect 7420 27100 7484 27164
rect 3740 26964 3804 27028
rect 4660 26828 4724 26892
rect 10180 26964 10244 27028
rect 6132 26828 6196 26892
rect 6316 26828 6380 26892
rect 10364 26828 10428 26892
rect 10732 26828 10796 26892
rect 3884 26684 3948 26688
rect 3884 26628 3888 26684
rect 3888 26628 3944 26684
rect 3944 26628 3948 26684
rect 3884 26624 3948 26628
rect 3964 26684 4028 26688
rect 3964 26628 3968 26684
rect 3968 26628 4024 26684
rect 4024 26628 4028 26684
rect 3964 26624 4028 26628
rect 4044 26684 4108 26688
rect 4044 26628 4048 26684
rect 4048 26628 4104 26684
rect 4104 26628 4108 26684
rect 4044 26624 4108 26628
rect 4124 26684 4188 26688
rect 4124 26628 4128 26684
rect 4128 26628 4184 26684
rect 4184 26628 4188 26684
rect 4124 26624 4188 26628
rect 9749 26684 9813 26688
rect 9749 26628 9753 26684
rect 9753 26628 9809 26684
rect 9809 26628 9813 26684
rect 9749 26624 9813 26628
rect 9829 26684 9893 26688
rect 9829 26628 9833 26684
rect 9833 26628 9889 26684
rect 9889 26628 9893 26684
rect 9829 26624 9893 26628
rect 9909 26684 9973 26688
rect 9909 26628 9913 26684
rect 9913 26628 9969 26684
rect 9969 26628 9973 26684
rect 9909 26624 9973 26628
rect 9989 26684 10053 26688
rect 9989 26628 9993 26684
rect 9993 26628 10049 26684
rect 10049 26628 10053 26684
rect 9989 26624 10053 26628
rect 15614 26684 15678 26688
rect 15614 26628 15618 26684
rect 15618 26628 15674 26684
rect 15674 26628 15678 26684
rect 15614 26624 15678 26628
rect 15694 26684 15758 26688
rect 15694 26628 15698 26684
rect 15698 26628 15754 26684
rect 15754 26628 15758 26684
rect 15694 26624 15758 26628
rect 15774 26684 15838 26688
rect 15774 26628 15778 26684
rect 15778 26628 15834 26684
rect 15834 26628 15838 26684
rect 15774 26624 15838 26628
rect 15854 26684 15918 26688
rect 15854 26628 15858 26684
rect 15858 26628 15914 26684
rect 15914 26628 15918 26684
rect 15854 26624 15918 26628
rect 21479 26684 21543 26688
rect 21479 26628 21483 26684
rect 21483 26628 21539 26684
rect 21539 26628 21543 26684
rect 21479 26624 21543 26628
rect 21559 26684 21623 26688
rect 21559 26628 21563 26684
rect 21563 26628 21619 26684
rect 21619 26628 21623 26684
rect 21559 26624 21623 26628
rect 21639 26684 21703 26688
rect 21639 26628 21643 26684
rect 21643 26628 21699 26684
rect 21699 26628 21703 26684
rect 21639 26624 21703 26628
rect 21719 26684 21783 26688
rect 21719 26628 21723 26684
rect 21723 26628 21779 26684
rect 21779 26628 21783 26684
rect 21719 26624 21783 26628
rect 5764 26556 5828 26620
rect 11284 26556 11348 26620
rect 14044 26556 14108 26620
rect 14780 26556 14844 26620
rect 10180 26284 10244 26348
rect 5212 26208 5276 26212
rect 5212 26152 5226 26208
rect 5226 26152 5276 26208
rect 2268 26012 2332 26076
rect 5212 26148 5276 26152
rect 7972 26148 8036 26212
rect 6816 26140 6880 26144
rect 6816 26084 6820 26140
rect 6820 26084 6876 26140
rect 6876 26084 6880 26140
rect 6816 26080 6880 26084
rect 6896 26140 6960 26144
rect 6896 26084 6900 26140
rect 6900 26084 6956 26140
rect 6956 26084 6960 26140
rect 6896 26080 6960 26084
rect 6976 26140 7040 26144
rect 6976 26084 6980 26140
rect 6980 26084 7036 26140
rect 7036 26084 7040 26140
rect 6976 26080 7040 26084
rect 7056 26140 7120 26144
rect 7056 26084 7060 26140
rect 7060 26084 7116 26140
rect 7116 26084 7120 26140
rect 7056 26080 7120 26084
rect 12681 26140 12745 26144
rect 12681 26084 12685 26140
rect 12685 26084 12741 26140
rect 12741 26084 12745 26140
rect 12681 26080 12745 26084
rect 12761 26140 12825 26144
rect 12761 26084 12765 26140
rect 12765 26084 12821 26140
rect 12821 26084 12825 26140
rect 12761 26080 12825 26084
rect 12841 26140 12905 26144
rect 12841 26084 12845 26140
rect 12845 26084 12901 26140
rect 12901 26084 12905 26140
rect 12841 26080 12905 26084
rect 12921 26140 12985 26144
rect 12921 26084 12925 26140
rect 12925 26084 12981 26140
rect 12981 26084 12985 26140
rect 12921 26080 12985 26084
rect 18546 26140 18610 26144
rect 18546 26084 18550 26140
rect 18550 26084 18606 26140
rect 18606 26084 18610 26140
rect 18546 26080 18610 26084
rect 18626 26140 18690 26144
rect 18626 26084 18630 26140
rect 18630 26084 18686 26140
rect 18686 26084 18690 26140
rect 18626 26080 18690 26084
rect 18706 26140 18770 26144
rect 18706 26084 18710 26140
rect 18710 26084 18766 26140
rect 18766 26084 18770 26140
rect 18706 26080 18770 26084
rect 18786 26140 18850 26144
rect 18786 26084 18790 26140
rect 18790 26084 18846 26140
rect 18846 26084 18850 26140
rect 18786 26080 18850 26084
rect 24411 26140 24475 26144
rect 24411 26084 24415 26140
rect 24415 26084 24471 26140
rect 24471 26084 24475 26140
rect 24411 26080 24475 26084
rect 24491 26140 24555 26144
rect 24491 26084 24495 26140
rect 24495 26084 24551 26140
rect 24551 26084 24555 26140
rect 24491 26080 24555 26084
rect 24571 26140 24635 26144
rect 24571 26084 24575 26140
rect 24575 26084 24631 26140
rect 24631 26084 24635 26140
rect 24571 26080 24635 26084
rect 24651 26140 24715 26144
rect 24651 26084 24655 26140
rect 24655 26084 24711 26140
rect 24711 26084 24715 26140
rect 24651 26080 24715 26084
rect 5212 26012 5276 26076
rect 20116 25876 20180 25940
rect 2820 25604 2884 25668
rect 5948 25604 6012 25668
rect 3884 25596 3948 25600
rect 3884 25540 3888 25596
rect 3888 25540 3944 25596
rect 3944 25540 3948 25596
rect 3884 25536 3948 25540
rect 3964 25596 4028 25600
rect 3964 25540 3968 25596
rect 3968 25540 4024 25596
rect 4024 25540 4028 25596
rect 3964 25536 4028 25540
rect 4044 25596 4108 25600
rect 4044 25540 4048 25596
rect 4048 25540 4104 25596
rect 4104 25540 4108 25596
rect 4044 25536 4108 25540
rect 4124 25596 4188 25600
rect 4124 25540 4128 25596
rect 4128 25540 4184 25596
rect 4184 25540 4188 25596
rect 4124 25536 4188 25540
rect 9749 25596 9813 25600
rect 9749 25540 9753 25596
rect 9753 25540 9809 25596
rect 9809 25540 9813 25596
rect 9749 25536 9813 25540
rect 9829 25596 9893 25600
rect 9829 25540 9833 25596
rect 9833 25540 9889 25596
rect 9889 25540 9893 25596
rect 9829 25536 9893 25540
rect 9909 25596 9973 25600
rect 9909 25540 9913 25596
rect 9913 25540 9969 25596
rect 9969 25540 9973 25596
rect 9909 25536 9973 25540
rect 9989 25596 10053 25600
rect 9989 25540 9993 25596
rect 9993 25540 10049 25596
rect 10049 25540 10053 25596
rect 9989 25536 10053 25540
rect 15614 25596 15678 25600
rect 15614 25540 15618 25596
rect 15618 25540 15674 25596
rect 15674 25540 15678 25596
rect 15614 25536 15678 25540
rect 15694 25596 15758 25600
rect 15694 25540 15698 25596
rect 15698 25540 15754 25596
rect 15754 25540 15758 25596
rect 15694 25536 15758 25540
rect 15774 25596 15838 25600
rect 15774 25540 15778 25596
rect 15778 25540 15834 25596
rect 15834 25540 15838 25596
rect 15774 25536 15838 25540
rect 15854 25596 15918 25600
rect 15854 25540 15858 25596
rect 15858 25540 15914 25596
rect 15914 25540 15918 25596
rect 15854 25536 15918 25540
rect 21479 25596 21543 25600
rect 21479 25540 21483 25596
rect 21483 25540 21539 25596
rect 21539 25540 21543 25596
rect 21479 25536 21543 25540
rect 21559 25596 21623 25600
rect 21559 25540 21563 25596
rect 21563 25540 21619 25596
rect 21619 25540 21623 25596
rect 21559 25536 21623 25540
rect 21639 25596 21703 25600
rect 21639 25540 21643 25596
rect 21643 25540 21699 25596
rect 21699 25540 21703 25596
rect 21639 25536 21703 25540
rect 21719 25596 21783 25600
rect 21719 25540 21723 25596
rect 21723 25540 21779 25596
rect 21779 25540 21783 25596
rect 21719 25536 21783 25540
rect 5396 25332 5460 25396
rect 2636 24924 2700 24988
rect 5764 24924 5828 24988
rect 6816 25052 6880 25056
rect 6816 24996 6820 25052
rect 6820 24996 6876 25052
rect 6876 24996 6880 25052
rect 6816 24992 6880 24996
rect 6896 25052 6960 25056
rect 6896 24996 6900 25052
rect 6900 24996 6956 25052
rect 6956 24996 6960 25052
rect 6896 24992 6960 24996
rect 6976 25052 7040 25056
rect 6976 24996 6980 25052
rect 6980 24996 7036 25052
rect 7036 24996 7040 25052
rect 6976 24992 7040 24996
rect 7056 25052 7120 25056
rect 7056 24996 7060 25052
rect 7060 24996 7116 25052
rect 7116 24996 7120 25052
rect 7056 24992 7120 24996
rect 12681 25052 12745 25056
rect 12681 24996 12685 25052
rect 12685 24996 12741 25052
rect 12741 24996 12745 25052
rect 12681 24992 12745 24996
rect 12761 25052 12825 25056
rect 12761 24996 12765 25052
rect 12765 24996 12821 25052
rect 12821 24996 12825 25052
rect 12761 24992 12825 24996
rect 12841 25052 12905 25056
rect 12841 24996 12845 25052
rect 12845 24996 12901 25052
rect 12901 24996 12905 25052
rect 12841 24992 12905 24996
rect 12921 25052 12985 25056
rect 12921 24996 12925 25052
rect 12925 24996 12981 25052
rect 12981 24996 12985 25052
rect 12921 24992 12985 24996
rect 18546 25052 18610 25056
rect 18546 24996 18550 25052
rect 18550 24996 18606 25052
rect 18606 24996 18610 25052
rect 18546 24992 18610 24996
rect 18626 25052 18690 25056
rect 18626 24996 18630 25052
rect 18630 24996 18686 25052
rect 18686 24996 18690 25052
rect 18626 24992 18690 24996
rect 18706 25052 18770 25056
rect 18706 24996 18710 25052
rect 18710 24996 18766 25052
rect 18766 24996 18770 25052
rect 18706 24992 18770 24996
rect 18786 25052 18850 25056
rect 18786 24996 18790 25052
rect 18790 24996 18846 25052
rect 18846 24996 18850 25052
rect 18786 24992 18850 24996
rect 24411 25052 24475 25056
rect 24411 24996 24415 25052
rect 24415 24996 24471 25052
rect 24471 24996 24475 25052
rect 24411 24992 24475 24996
rect 24491 25052 24555 25056
rect 24491 24996 24495 25052
rect 24495 24996 24551 25052
rect 24551 24996 24555 25052
rect 24491 24992 24555 24996
rect 24571 25052 24635 25056
rect 24571 24996 24575 25052
rect 24575 24996 24631 25052
rect 24631 24996 24635 25052
rect 24571 24992 24635 24996
rect 24651 25052 24715 25056
rect 24651 24996 24655 25052
rect 24655 24996 24711 25052
rect 24711 24996 24715 25052
rect 24651 24992 24715 24996
rect 2820 24516 2884 24580
rect 3884 24508 3948 24512
rect 3884 24452 3888 24508
rect 3888 24452 3944 24508
rect 3944 24452 3948 24508
rect 3884 24448 3948 24452
rect 3964 24508 4028 24512
rect 3964 24452 3968 24508
rect 3968 24452 4024 24508
rect 4024 24452 4028 24508
rect 3964 24448 4028 24452
rect 4044 24508 4108 24512
rect 4044 24452 4048 24508
rect 4048 24452 4104 24508
rect 4104 24452 4108 24508
rect 4044 24448 4108 24452
rect 4124 24508 4188 24512
rect 4124 24452 4128 24508
rect 4128 24452 4184 24508
rect 4184 24452 4188 24508
rect 4124 24448 4188 24452
rect 9749 24508 9813 24512
rect 9749 24452 9753 24508
rect 9753 24452 9809 24508
rect 9809 24452 9813 24508
rect 9749 24448 9813 24452
rect 9829 24508 9893 24512
rect 9829 24452 9833 24508
rect 9833 24452 9889 24508
rect 9889 24452 9893 24508
rect 9829 24448 9893 24452
rect 9909 24508 9973 24512
rect 9909 24452 9913 24508
rect 9913 24452 9969 24508
rect 9969 24452 9973 24508
rect 9909 24448 9973 24452
rect 9989 24508 10053 24512
rect 9989 24452 9993 24508
rect 9993 24452 10049 24508
rect 10049 24452 10053 24508
rect 9989 24448 10053 24452
rect 15614 24508 15678 24512
rect 15614 24452 15618 24508
rect 15618 24452 15674 24508
rect 15674 24452 15678 24508
rect 15614 24448 15678 24452
rect 15694 24508 15758 24512
rect 15694 24452 15698 24508
rect 15698 24452 15754 24508
rect 15754 24452 15758 24508
rect 15694 24448 15758 24452
rect 15774 24508 15838 24512
rect 15774 24452 15778 24508
rect 15778 24452 15834 24508
rect 15834 24452 15838 24508
rect 15774 24448 15838 24452
rect 15854 24508 15918 24512
rect 15854 24452 15858 24508
rect 15858 24452 15914 24508
rect 15914 24452 15918 24508
rect 15854 24448 15918 24452
rect 21479 24508 21543 24512
rect 21479 24452 21483 24508
rect 21483 24452 21539 24508
rect 21539 24452 21543 24508
rect 21479 24448 21543 24452
rect 21559 24508 21623 24512
rect 21559 24452 21563 24508
rect 21563 24452 21619 24508
rect 21619 24452 21623 24508
rect 21559 24448 21623 24452
rect 21639 24508 21703 24512
rect 21639 24452 21643 24508
rect 21643 24452 21699 24508
rect 21699 24452 21703 24508
rect 21639 24448 21703 24452
rect 21719 24508 21783 24512
rect 21719 24452 21723 24508
rect 21723 24452 21779 24508
rect 21779 24452 21783 24508
rect 21719 24448 21783 24452
rect 5028 24108 5092 24172
rect 21956 24108 22020 24172
rect 6816 23964 6880 23968
rect 6816 23908 6820 23964
rect 6820 23908 6876 23964
rect 6876 23908 6880 23964
rect 6816 23904 6880 23908
rect 6896 23964 6960 23968
rect 6896 23908 6900 23964
rect 6900 23908 6956 23964
rect 6956 23908 6960 23964
rect 6896 23904 6960 23908
rect 6976 23964 7040 23968
rect 6976 23908 6980 23964
rect 6980 23908 7036 23964
rect 7036 23908 7040 23964
rect 6976 23904 7040 23908
rect 7056 23964 7120 23968
rect 7056 23908 7060 23964
rect 7060 23908 7116 23964
rect 7116 23908 7120 23964
rect 7056 23904 7120 23908
rect 12681 23964 12745 23968
rect 12681 23908 12685 23964
rect 12685 23908 12741 23964
rect 12741 23908 12745 23964
rect 12681 23904 12745 23908
rect 12761 23964 12825 23968
rect 12761 23908 12765 23964
rect 12765 23908 12821 23964
rect 12821 23908 12825 23964
rect 12761 23904 12825 23908
rect 12841 23964 12905 23968
rect 12841 23908 12845 23964
rect 12845 23908 12901 23964
rect 12901 23908 12905 23964
rect 12841 23904 12905 23908
rect 12921 23964 12985 23968
rect 12921 23908 12925 23964
rect 12925 23908 12981 23964
rect 12981 23908 12985 23964
rect 12921 23904 12985 23908
rect 18546 23964 18610 23968
rect 18546 23908 18550 23964
rect 18550 23908 18606 23964
rect 18606 23908 18610 23964
rect 18546 23904 18610 23908
rect 18626 23964 18690 23968
rect 18626 23908 18630 23964
rect 18630 23908 18686 23964
rect 18686 23908 18690 23964
rect 18626 23904 18690 23908
rect 18706 23964 18770 23968
rect 18706 23908 18710 23964
rect 18710 23908 18766 23964
rect 18766 23908 18770 23964
rect 18706 23904 18770 23908
rect 18786 23964 18850 23968
rect 18786 23908 18790 23964
rect 18790 23908 18846 23964
rect 18846 23908 18850 23964
rect 18786 23904 18850 23908
rect 24411 23964 24475 23968
rect 24411 23908 24415 23964
rect 24415 23908 24471 23964
rect 24471 23908 24475 23964
rect 24411 23904 24475 23908
rect 24491 23964 24555 23968
rect 24491 23908 24495 23964
rect 24495 23908 24551 23964
rect 24551 23908 24555 23964
rect 24491 23904 24555 23908
rect 24571 23964 24635 23968
rect 24571 23908 24575 23964
rect 24575 23908 24631 23964
rect 24631 23908 24635 23964
rect 24571 23904 24635 23908
rect 24651 23964 24715 23968
rect 24651 23908 24655 23964
rect 24655 23908 24711 23964
rect 24711 23908 24715 23964
rect 24651 23904 24715 23908
rect 11284 23564 11348 23628
rect 2452 23488 2516 23492
rect 2452 23432 2502 23488
rect 2502 23432 2516 23488
rect 2452 23428 2516 23432
rect 5028 23428 5092 23492
rect 14228 23428 14292 23492
rect 3884 23420 3948 23424
rect 3884 23364 3888 23420
rect 3888 23364 3944 23420
rect 3944 23364 3948 23420
rect 3884 23360 3948 23364
rect 3964 23420 4028 23424
rect 3964 23364 3968 23420
rect 3968 23364 4024 23420
rect 4024 23364 4028 23420
rect 3964 23360 4028 23364
rect 4044 23420 4108 23424
rect 4044 23364 4048 23420
rect 4048 23364 4104 23420
rect 4104 23364 4108 23420
rect 4044 23360 4108 23364
rect 4124 23420 4188 23424
rect 4124 23364 4128 23420
rect 4128 23364 4184 23420
rect 4184 23364 4188 23420
rect 4124 23360 4188 23364
rect 9749 23420 9813 23424
rect 9749 23364 9753 23420
rect 9753 23364 9809 23420
rect 9809 23364 9813 23420
rect 9749 23360 9813 23364
rect 9829 23420 9893 23424
rect 9829 23364 9833 23420
rect 9833 23364 9889 23420
rect 9889 23364 9893 23420
rect 9829 23360 9893 23364
rect 9909 23420 9973 23424
rect 9909 23364 9913 23420
rect 9913 23364 9969 23420
rect 9969 23364 9973 23420
rect 9909 23360 9973 23364
rect 9989 23420 10053 23424
rect 9989 23364 9993 23420
rect 9993 23364 10049 23420
rect 10049 23364 10053 23420
rect 9989 23360 10053 23364
rect 15614 23420 15678 23424
rect 15614 23364 15618 23420
rect 15618 23364 15674 23420
rect 15674 23364 15678 23420
rect 15614 23360 15678 23364
rect 15694 23420 15758 23424
rect 15694 23364 15698 23420
rect 15698 23364 15754 23420
rect 15754 23364 15758 23420
rect 15694 23360 15758 23364
rect 15774 23420 15838 23424
rect 15774 23364 15778 23420
rect 15778 23364 15834 23420
rect 15834 23364 15838 23420
rect 15774 23360 15838 23364
rect 15854 23420 15918 23424
rect 15854 23364 15858 23420
rect 15858 23364 15914 23420
rect 15914 23364 15918 23420
rect 15854 23360 15918 23364
rect 21479 23420 21543 23424
rect 21479 23364 21483 23420
rect 21483 23364 21539 23420
rect 21539 23364 21543 23420
rect 21479 23360 21543 23364
rect 21559 23420 21623 23424
rect 21559 23364 21563 23420
rect 21563 23364 21619 23420
rect 21619 23364 21623 23420
rect 21559 23360 21623 23364
rect 21639 23420 21703 23424
rect 21639 23364 21643 23420
rect 21643 23364 21699 23420
rect 21699 23364 21703 23420
rect 21639 23360 21703 23364
rect 21719 23420 21783 23424
rect 21719 23364 21723 23420
rect 21723 23364 21779 23420
rect 21779 23364 21783 23420
rect 21719 23360 21783 23364
rect 3556 23292 3620 23356
rect 10916 23020 10980 23084
rect 6816 22876 6880 22880
rect 6816 22820 6820 22876
rect 6820 22820 6876 22876
rect 6876 22820 6880 22876
rect 6816 22816 6880 22820
rect 6896 22876 6960 22880
rect 6896 22820 6900 22876
rect 6900 22820 6956 22876
rect 6956 22820 6960 22876
rect 6896 22816 6960 22820
rect 6976 22876 7040 22880
rect 6976 22820 6980 22876
rect 6980 22820 7036 22876
rect 7036 22820 7040 22876
rect 6976 22816 7040 22820
rect 7056 22876 7120 22880
rect 7056 22820 7060 22876
rect 7060 22820 7116 22876
rect 7116 22820 7120 22876
rect 7056 22816 7120 22820
rect 12681 22876 12745 22880
rect 12681 22820 12685 22876
rect 12685 22820 12741 22876
rect 12741 22820 12745 22876
rect 12681 22816 12745 22820
rect 12761 22876 12825 22880
rect 12761 22820 12765 22876
rect 12765 22820 12821 22876
rect 12821 22820 12825 22876
rect 12761 22816 12825 22820
rect 12841 22876 12905 22880
rect 12841 22820 12845 22876
rect 12845 22820 12901 22876
rect 12901 22820 12905 22876
rect 12841 22816 12905 22820
rect 12921 22876 12985 22880
rect 12921 22820 12925 22876
rect 12925 22820 12981 22876
rect 12981 22820 12985 22876
rect 12921 22816 12985 22820
rect 18546 22876 18610 22880
rect 18546 22820 18550 22876
rect 18550 22820 18606 22876
rect 18606 22820 18610 22876
rect 18546 22816 18610 22820
rect 18626 22876 18690 22880
rect 18626 22820 18630 22876
rect 18630 22820 18686 22876
rect 18686 22820 18690 22876
rect 18626 22816 18690 22820
rect 18706 22876 18770 22880
rect 18706 22820 18710 22876
rect 18710 22820 18766 22876
rect 18766 22820 18770 22876
rect 18706 22816 18770 22820
rect 18786 22876 18850 22880
rect 18786 22820 18790 22876
rect 18790 22820 18846 22876
rect 18846 22820 18850 22876
rect 18786 22816 18850 22820
rect 24411 22876 24475 22880
rect 24411 22820 24415 22876
rect 24415 22820 24471 22876
rect 24471 22820 24475 22876
rect 24411 22816 24475 22820
rect 24491 22876 24555 22880
rect 24491 22820 24495 22876
rect 24495 22820 24551 22876
rect 24551 22820 24555 22876
rect 24491 22816 24555 22820
rect 24571 22876 24635 22880
rect 24571 22820 24575 22876
rect 24575 22820 24631 22876
rect 24631 22820 24635 22876
rect 24571 22816 24635 22820
rect 24651 22876 24715 22880
rect 24651 22820 24655 22876
rect 24655 22820 24711 22876
rect 24711 22820 24715 22876
rect 24651 22816 24715 22820
rect 14412 22672 14476 22676
rect 14412 22616 14462 22672
rect 14462 22616 14476 22672
rect 14412 22612 14476 22616
rect 3884 22332 3948 22336
rect 3884 22276 3888 22332
rect 3888 22276 3944 22332
rect 3944 22276 3948 22332
rect 3884 22272 3948 22276
rect 3964 22332 4028 22336
rect 3964 22276 3968 22332
rect 3968 22276 4024 22332
rect 4024 22276 4028 22332
rect 3964 22272 4028 22276
rect 4044 22332 4108 22336
rect 4044 22276 4048 22332
rect 4048 22276 4104 22332
rect 4104 22276 4108 22332
rect 4044 22272 4108 22276
rect 4124 22332 4188 22336
rect 4124 22276 4128 22332
rect 4128 22276 4184 22332
rect 4184 22276 4188 22332
rect 4124 22272 4188 22276
rect 9749 22332 9813 22336
rect 9749 22276 9753 22332
rect 9753 22276 9809 22332
rect 9809 22276 9813 22332
rect 9749 22272 9813 22276
rect 9829 22332 9893 22336
rect 9829 22276 9833 22332
rect 9833 22276 9889 22332
rect 9889 22276 9893 22332
rect 9829 22272 9893 22276
rect 9909 22332 9973 22336
rect 9909 22276 9913 22332
rect 9913 22276 9969 22332
rect 9969 22276 9973 22332
rect 9909 22272 9973 22276
rect 9989 22332 10053 22336
rect 9989 22276 9993 22332
rect 9993 22276 10049 22332
rect 10049 22276 10053 22332
rect 9989 22272 10053 22276
rect 15614 22332 15678 22336
rect 15614 22276 15618 22332
rect 15618 22276 15674 22332
rect 15674 22276 15678 22332
rect 15614 22272 15678 22276
rect 15694 22332 15758 22336
rect 15694 22276 15698 22332
rect 15698 22276 15754 22332
rect 15754 22276 15758 22332
rect 15694 22272 15758 22276
rect 15774 22332 15838 22336
rect 15774 22276 15778 22332
rect 15778 22276 15834 22332
rect 15834 22276 15838 22332
rect 15774 22272 15838 22276
rect 15854 22332 15918 22336
rect 15854 22276 15858 22332
rect 15858 22276 15914 22332
rect 15914 22276 15918 22332
rect 15854 22272 15918 22276
rect 21479 22332 21543 22336
rect 21479 22276 21483 22332
rect 21483 22276 21539 22332
rect 21539 22276 21543 22332
rect 21479 22272 21543 22276
rect 21559 22332 21623 22336
rect 21559 22276 21563 22332
rect 21563 22276 21619 22332
rect 21619 22276 21623 22332
rect 21559 22272 21623 22276
rect 21639 22332 21703 22336
rect 21639 22276 21643 22332
rect 21643 22276 21699 22332
rect 21699 22276 21703 22332
rect 21639 22272 21703 22276
rect 21719 22332 21783 22336
rect 21719 22276 21723 22332
rect 21723 22276 21779 22332
rect 21779 22276 21783 22332
rect 21719 22272 21783 22276
rect 10548 22204 10612 22268
rect 13308 22204 13372 22268
rect 12388 22068 12452 22132
rect 13124 22068 13188 22132
rect 13492 22068 13556 22132
rect 4476 21992 4540 21996
rect 4476 21936 4490 21992
rect 4490 21936 4540 21992
rect 4476 21932 4540 21936
rect 12388 21932 12452 21996
rect 13124 21932 13188 21996
rect 21220 21932 21284 21996
rect 1900 21796 1964 21860
rect 7604 21796 7668 21860
rect 6816 21788 6880 21792
rect 6816 21732 6820 21788
rect 6820 21732 6876 21788
rect 6876 21732 6880 21788
rect 6816 21728 6880 21732
rect 6896 21788 6960 21792
rect 6896 21732 6900 21788
rect 6900 21732 6956 21788
rect 6956 21732 6960 21788
rect 6896 21728 6960 21732
rect 6976 21788 7040 21792
rect 6976 21732 6980 21788
rect 6980 21732 7036 21788
rect 7036 21732 7040 21788
rect 6976 21728 7040 21732
rect 7056 21788 7120 21792
rect 7056 21732 7060 21788
rect 7060 21732 7116 21788
rect 7116 21732 7120 21788
rect 7056 21728 7120 21732
rect 12681 21788 12745 21792
rect 12681 21732 12685 21788
rect 12685 21732 12741 21788
rect 12741 21732 12745 21788
rect 12681 21728 12745 21732
rect 12761 21788 12825 21792
rect 12761 21732 12765 21788
rect 12765 21732 12821 21788
rect 12821 21732 12825 21788
rect 12761 21728 12825 21732
rect 12841 21788 12905 21792
rect 12841 21732 12845 21788
rect 12845 21732 12901 21788
rect 12901 21732 12905 21788
rect 12841 21728 12905 21732
rect 12921 21788 12985 21792
rect 12921 21732 12925 21788
rect 12925 21732 12981 21788
rect 12981 21732 12985 21788
rect 12921 21728 12985 21732
rect 18546 21788 18610 21792
rect 18546 21732 18550 21788
rect 18550 21732 18606 21788
rect 18606 21732 18610 21788
rect 18546 21728 18610 21732
rect 18626 21788 18690 21792
rect 18626 21732 18630 21788
rect 18630 21732 18686 21788
rect 18686 21732 18690 21788
rect 18626 21728 18690 21732
rect 18706 21788 18770 21792
rect 18706 21732 18710 21788
rect 18710 21732 18766 21788
rect 18766 21732 18770 21788
rect 18706 21728 18770 21732
rect 18786 21788 18850 21792
rect 18786 21732 18790 21788
rect 18790 21732 18846 21788
rect 18846 21732 18850 21788
rect 18786 21728 18850 21732
rect 24411 21788 24475 21792
rect 24411 21732 24415 21788
rect 24415 21732 24471 21788
rect 24471 21732 24475 21788
rect 24411 21728 24475 21732
rect 24491 21788 24555 21792
rect 24491 21732 24495 21788
rect 24495 21732 24551 21788
rect 24551 21732 24555 21788
rect 24491 21728 24555 21732
rect 24571 21788 24635 21792
rect 24571 21732 24575 21788
rect 24575 21732 24631 21788
rect 24631 21732 24635 21788
rect 24571 21728 24635 21732
rect 24651 21788 24715 21792
rect 24651 21732 24655 21788
rect 24655 21732 24711 21788
rect 24711 21732 24715 21788
rect 24651 21728 24715 21732
rect 8524 21524 8588 21588
rect 3884 21244 3948 21248
rect 3884 21188 3888 21244
rect 3888 21188 3944 21244
rect 3944 21188 3948 21244
rect 3884 21184 3948 21188
rect 3964 21244 4028 21248
rect 3964 21188 3968 21244
rect 3968 21188 4024 21244
rect 4024 21188 4028 21244
rect 3964 21184 4028 21188
rect 4044 21244 4108 21248
rect 4044 21188 4048 21244
rect 4048 21188 4104 21244
rect 4104 21188 4108 21244
rect 4044 21184 4108 21188
rect 4124 21244 4188 21248
rect 4124 21188 4128 21244
rect 4128 21188 4184 21244
rect 4184 21188 4188 21244
rect 4124 21184 4188 21188
rect 9749 21244 9813 21248
rect 9749 21188 9753 21244
rect 9753 21188 9809 21244
rect 9809 21188 9813 21244
rect 9749 21184 9813 21188
rect 9829 21244 9893 21248
rect 9829 21188 9833 21244
rect 9833 21188 9889 21244
rect 9889 21188 9893 21244
rect 9829 21184 9893 21188
rect 9909 21244 9973 21248
rect 9909 21188 9913 21244
rect 9913 21188 9969 21244
rect 9969 21188 9973 21244
rect 9909 21184 9973 21188
rect 9989 21244 10053 21248
rect 9989 21188 9993 21244
rect 9993 21188 10049 21244
rect 10049 21188 10053 21244
rect 9989 21184 10053 21188
rect 15614 21244 15678 21248
rect 15614 21188 15618 21244
rect 15618 21188 15674 21244
rect 15674 21188 15678 21244
rect 15614 21184 15678 21188
rect 15694 21244 15758 21248
rect 15694 21188 15698 21244
rect 15698 21188 15754 21244
rect 15754 21188 15758 21244
rect 15694 21184 15758 21188
rect 15774 21244 15838 21248
rect 15774 21188 15778 21244
rect 15778 21188 15834 21244
rect 15834 21188 15838 21244
rect 15774 21184 15838 21188
rect 15854 21244 15918 21248
rect 15854 21188 15858 21244
rect 15858 21188 15914 21244
rect 15914 21188 15918 21244
rect 15854 21184 15918 21188
rect 21479 21244 21543 21248
rect 21479 21188 21483 21244
rect 21483 21188 21539 21244
rect 21539 21188 21543 21244
rect 21479 21184 21543 21188
rect 21559 21244 21623 21248
rect 21559 21188 21563 21244
rect 21563 21188 21619 21244
rect 21619 21188 21623 21244
rect 21559 21184 21623 21188
rect 21639 21244 21703 21248
rect 21639 21188 21643 21244
rect 21643 21188 21699 21244
rect 21699 21188 21703 21244
rect 21639 21184 21703 21188
rect 21719 21244 21783 21248
rect 21719 21188 21723 21244
rect 21723 21188 21779 21244
rect 21779 21188 21783 21244
rect 21719 21184 21783 21188
rect 8708 20980 8772 21044
rect 11284 21040 11348 21044
rect 11284 20984 11298 21040
rect 11298 20984 11348 21040
rect 11284 20980 11348 20984
rect 3188 20904 3252 20908
rect 3188 20848 3238 20904
rect 3238 20848 3252 20904
rect 3188 20844 3252 20848
rect 9444 20708 9508 20772
rect 13308 20708 13372 20772
rect 13676 20708 13740 20772
rect 14596 20708 14660 20772
rect 6816 20700 6880 20704
rect 6816 20644 6820 20700
rect 6820 20644 6876 20700
rect 6876 20644 6880 20700
rect 6816 20640 6880 20644
rect 6896 20700 6960 20704
rect 6896 20644 6900 20700
rect 6900 20644 6956 20700
rect 6956 20644 6960 20700
rect 6896 20640 6960 20644
rect 6976 20700 7040 20704
rect 6976 20644 6980 20700
rect 6980 20644 7036 20700
rect 7036 20644 7040 20700
rect 6976 20640 7040 20644
rect 7056 20700 7120 20704
rect 7056 20644 7060 20700
rect 7060 20644 7116 20700
rect 7116 20644 7120 20700
rect 7056 20640 7120 20644
rect 12681 20700 12745 20704
rect 12681 20644 12685 20700
rect 12685 20644 12741 20700
rect 12741 20644 12745 20700
rect 12681 20640 12745 20644
rect 12761 20700 12825 20704
rect 12761 20644 12765 20700
rect 12765 20644 12821 20700
rect 12821 20644 12825 20700
rect 12761 20640 12825 20644
rect 12841 20700 12905 20704
rect 12841 20644 12845 20700
rect 12845 20644 12901 20700
rect 12901 20644 12905 20700
rect 12841 20640 12905 20644
rect 12921 20700 12985 20704
rect 12921 20644 12925 20700
rect 12925 20644 12981 20700
rect 12981 20644 12985 20700
rect 12921 20640 12985 20644
rect 18546 20700 18610 20704
rect 18546 20644 18550 20700
rect 18550 20644 18606 20700
rect 18606 20644 18610 20700
rect 18546 20640 18610 20644
rect 18626 20700 18690 20704
rect 18626 20644 18630 20700
rect 18630 20644 18686 20700
rect 18686 20644 18690 20700
rect 18626 20640 18690 20644
rect 18706 20700 18770 20704
rect 18706 20644 18710 20700
rect 18710 20644 18766 20700
rect 18766 20644 18770 20700
rect 18706 20640 18770 20644
rect 18786 20700 18850 20704
rect 18786 20644 18790 20700
rect 18790 20644 18846 20700
rect 18846 20644 18850 20700
rect 18786 20640 18850 20644
rect 24411 20700 24475 20704
rect 24411 20644 24415 20700
rect 24415 20644 24471 20700
rect 24471 20644 24475 20700
rect 24411 20640 24475 20644
rect 24491 20700 24555 20704
rect 24491 20644 24495 20700
rect 24495 20644 24551 20700
rect 24551 20644 24555 20700
rect 24491 20640 24555 20644
rect 24571 20700 24635 20704
rect 24571 20644 24575 20700
rect 24575 20644 24631 20700
rect 24631 20644 24635 20700
rect 24571 20640 24635 20644
rect 24651 20700 24715 20704
rect 24651 20644 24655 20700
rect 24655 20644 24711 20700
rect 24711 20644 24715 20700
rect 24651 20640 24715 20644
rect 2084 20632 2148 20636
rect 2084 20576 2098 20632
rect 2098 20576 2148 20632
rect 2084 20572 2148 20576
rect 5396 20572 5460 20636
rect 14412 20572 14476 20636
rect 14964 20436 15028 20500
rect 10180 20164 10244 20228
rect 14964 20164 15028 20228
rect 3884 20156 3948 20160
rect 3884 20100 3888 20156
rect 3888 20100 3944 20156
rect 3944 20100 3948 20156
rect 3884 20096 3948 20100
rect 3964 20156 4028 20160
rect 3964 20100 3968 20156
rect 3968 20100 4024 20156
rect 4024 20100 4028 20156
rect 3964 20096 4028 20100
rect 4044 20156 4108 20160
rect 4044 20100 4048 20156
rect 4048 20100 4104 20156
rect 4104 20100 4108 20156
rect 4044 20096 4108 20100
rect 4124 20156 4188 20160
rect 4124 20100 4128 20156
rect 4128 20100 4184 20156
rect 4184 20100 4188 20156
rect 4124 20096 4188 20100
rect 9749 20156 9813 20160
rect 9749 20100 9753 20156
rect 9753 20100 9809 20156
rect 9809 20100 9813 20156
rect 9749 20096 9813 20100
rect 9829 20156 9893 20160
rect 9829 20100 9833 20156
rect 9833 20100 9889 20156
rect 9889 20100 9893 20156
rect 9829 20096 9893 20100
rect 9909 20156 9973 20160
rect 9909 20100 9913 20156
rect 9913 20100 9969 20156
rect 9969 20100 9973 20156
rect 9909 20096 9973 20100
rect 9989 20156 10053 20160
rect 9989 20100 9993 20156
rect 9993 20100 10049 20156
rect 10049 20100 10053 20156
rect 9989 20096 10053 20100
rect 15614 20156 15678 20160
rect 15614 20100 15618 20156
rect 15618 20100 15674 20156
rect 15674 20100 15678 20156
rect 15614 20096 15678 20100
rect 15694 20156 15758 20160
rect 15694 20100 15698 20156
rect 15698 20100 15754 20156
rect 15754 20100 15758 20156
rect 15694 20096 15758 20100
rect 15774 20156 15838 20160
rect 15774 20100 15778 20156
rect 15778 20100 15834 20156
rect 15834 20100 15838 20156
rect 15774 20096 15838 20100
rect 15854 20156 15918 20160
rect 15854 20100 15858 20156
rect 15858 20100 15914 20156
rect 15914 20100 15918 20156
rect 15854 20096 15918 20100
rect 21479 20156 21543 20160
rect 21479 20100 21483 20156
rect 21483 20100 21539 20156
rect 21539 20100 21543 20156
rect 21479 20096 21543 20100
rect 21559 20156 21623 20160
rect 21559 20100 21563 20156
rect 21563 20100 21619 20156
rect 21619 20100 21623 20156
rect 21559 20096 21623 20100
rect 21639 20156 21703 20160
rect 21639 20100 21643 20156
rect 21643 20100 21699 20156
rect 21699 20100 21703 20156
rect 21639 20096 21703 20100
rect 21719 20156 21783 20160
rect 21719 20100 21723 20156
rect 21723 20100 21779 20156
rect 21779 20100 21783 20156
rect 21719 20096 21783 20100
rect 1716 20088 1780 20092
rect 1716 20032 1730 20088
rect 1730 20032 1780 20088
rect 1716 20028 1780 20032
rect 3740 19892 3804 19956
rect 5396 19892 5460 19956
rect 10364 19892 10428 19956
rect 3372 19680 3436 19684
rect 3372 19624 3422 19680
rect 3422 19624 3436 19680
rect 2268 19544 2332 19548
rect 2268 19488 2282 19544
rect 2282 19488 2332 19544
rect 2268 19484 2332 19488
rect 3372 19620 3436 19624
rect 5580 19620 5644 19684
rect 6816 19612 6880 19616
rect 6816 19556 6820 19612
rect 6820 19556 6876 19612
rect 6876 19556 6880 19612
rect 6816 19552 6880 19556
rect 6896 19612 6960 19616
rect 6896 19556 6900 19612
rect 6900 19556 6956 19612
rect 6956 19556 6960 19612
rect 6896 19552 6960 19556
rect 6976 19612 7040 19616
rect 6976 19556 6980 19612
rect 6980 19556 7036 19612
rect 7036 19556 7040 19612
rect 6976 19552 7040 19556
rect 7056 19612 7120 19616
rect 7056 19556 7060 19612
rect 7060 19556 7116 19612
rect 7116 19556 7120 19612
rect 7056 19552 7120 19556
rect 1532 19348 1596 19412
rect 12681 19612 12745 19616
rect 12681 19556 12685 19612
rect 12685 19556 12741 19612
rect 12741 19556 12745 19612
rect 12681 19552 12745 19556
rect 12761 19612 12825 19616
rect 12761 19556 12765 19612
rect 12765 19556 12821 19612
rect 12821 19556 12825 19612
rect 12761 19552 12825 19556
rect 12841 19612 12905 19616
rect 12841 19556 12845 19612
rect 12845 19556 12901 19612
rect 12901 19556 12905 19612
rect 12841 19552 12905 19556
rect 12921 19612 12985 19616
rect 12921 19556 12925 19612
rect 12925 19556 12981 19612
rect 12981 19556 12985 19612
rect 12921 19552 12985 19556
rect 18546 19612 18610 19616
rect 18546 19556 18550 19612
rect 18550 19556 18606 19612
rect 18606 19556 18610 19612
rect 18546 19552 18610 19556
rect 18626 19612 18690 19616
rect 18626 19556 18630 19612
rect 18630 19556 18686 19612
rect 18686 19556 18690 19612
rect 18626 19552 18690 19556
rect 18706 19612 18770 19616
rect 18706 19556 18710 19612
rect 18710 19556 18766 19612
rect 18766 19556 18770 19612
rect 18706 19552 18770 19556
rect 18786 19612 18850 19616
rect 18786 19556 18790 19612
rect 18790 19556 18846 19612
rect 18846 19556 18850 19612
rect 18786 19552 18850 19556
rect 24411 19612 24475 19616
rect 24411 19556 24415 19612
rect 24415 19556 24471 19612
rect 24471 19556 24475 19612
rect 24411 19552 24475 19556
rect 24491 19612 24555 19616
rect 24491 19556 24495 19612
rect 24495 19556 24551 19612
rect 24551 19556 24555 19612
rect 24491 19552 24555 19556
rect 24571 19612 24635 19616
rect 24571 19556 24575 19612
rect 24575 19556 24631 19612
rect 24631 19556 24635 19612
rect 24571 19552 24635 19556
rect 24651 19612 24715 19616
rect 24651 19556 24655 19612
rect 24655 19556 24711 19612
rect 24711 19556 24715 19612
rect 24651 19552 24715 19556
rect 15148 19348 15212 19412
rect 16436 19348 16500 19412
rect 18092 19348 18156 19412
rect 4292 19076 4356 19140
rect 3884 19068 3948 19072
rect 3884 19012 3888 19068
rect 3888 19012 3944 19068
rect 3944 19012 3948 19068
rect 3884 19008 3948 19012
rect 3964 19068 4028 19072
rect 3964 19012 3968 19068
rect 3968 19012 4024 19068
rect 4024 19012 4028 19068
rect 3964 19008 4028 19012
rect 4044 19068 4108 19072
rect 4044 19012 4048 19068
rect 4048 19012 4104 19068
rect 4104 19012 4108 19068
rect 4044 19008 4108 19012
rect 4124 19068 4188 19072
rect 4124 19012 4128 19068
rect 4128 19012 4184 19068
rect 4184 19012 4188 19068
rect 4124 19008 4188 19012
rect 9749 19068 9813 19072
rect 9749 19012 9753 19068
rect 9753 19012 9809 19068
rect 9809 19012 9813 19068
rect 9749 19008 9813 19012
rect 9829 19068 9893 19072
rect 9829 19012 9833 19068
rect 9833 19012 9889 19068
rect 9889 19012 9893 19068
rect 9829 19008 9893 19012
rect 9909 19068 9973 19072
rect 9909 19012 9913 19068
rect 9913 19012 9969 19068
rect 9969 19012 9973 19068
rect 9909 19008 9973 19012
rect 9989 19068 10053 19072
rect 9989 19012 9993 19068
rect 9993 19012 10049 19068
rect 10049 19012 10053 19068
rect 9989 19008 10053 19012
rect 15614 19068 15678 19072
rect 15614 19012 15618 19068
rect 15618 19012 15674 19068
rect 15674 19012 15678 19068
rect 15614 19008 15678 19012
rect 15694 19068 15758 19072
rect 15694 19012 15698 19068
rect 15698 19012 15754 19068
rect 15754 19012 15758 19068
rect 15694 19008 15758 19012
rect 15774 19068 15838 19072
rect 15774 19012 15778 19068
rect 15778 19012 15834 19068
rect 15834 19012 15838 19068
rect 15774 19008 15838 19012
rect 15854 19068 15918 19072
rect 15854 19012 15858 19068
rect 15858 19012 15914 19068
rect 15914 19012 15918 19068
rect 15854 19008 15918 19012
rect 21479 19068 21543 19072
rect 21479 19012 21483 19068
rect 21483 19012 21539 19068
rect 21539 19012 21543 19068
rect 21479 19008 21543 19012
rect 21559 19068 21623 19072
rect 21559 19012 21563 19068
rect 21563 19012 21619 19068
rect 21619 19012 21623 19068
rect 21559 19008 21623 19012
rect 21639 19068 21703 19072
rect 21639 19012 21643 19068
rect 21643 19012 21699 19068
rect 21699 19012 21703 19068
rect 21639 19008 21703 19012
rect 21719 19068 21783 19072
rect 21719 19012 21723 19068
rect 21723 19012 21779 19068
rect 21779 19012 21783 19068
rect 21719 19008 21783 19012
rect 2636 18668 2700 18732
rect 6816 18524 6880 18528
rect 6816 18468 6820 18524
rect 6820 18468 6876 18524
rect 6876 18468 6880 18524
rect 6816 18464 6880 18468
rect 6896 18524 6960 18528
rect 6896 18468 6900 18524
rect 6900 18468 6956 18524
rect 6956 18468 6960 18524
rect 6896 18464 6960 18468
rect 6976 18524 7040 18528
rect 6976 18468 6980 18524
rect 6980 18468 7036 18524
rect 7036 18468 7040 18524
rect 6976 18464 7040 18468
rect 7056 18524 7120 18528
rect 7056 18468 7060 18524
rect 7060 18468 7116 18524
rect 7116 18468 7120 18524
rect 7056 18464 7120 18468
rect 12681 18524 12745 18528
rect 12681 18468 12685 18524
rect 12685 18468 12741 18524
rect 12741 18468 12745 18524
rect 12681 18464 12745 18468
rect 12761 18524 12825 18528
rect 12761 18468 12765 18524
rect 12765 18468 12821 18524
rect 12821 18468 12825 18524
rect 12761 18464 12825 18468
rect 12841 18524 12905 18528
rect 12841 18468 12845 18524
rect 12845 18468 12901 18524
rect 12901 18468 12905 18524
rect 12841 18464 12905 18468
rect 12921 18524 12985 18528
rect 12921 18468 12925 18524
rect 12925 18468 12981 18524
rect 12981 18468 12985 18524
rect 12921 18464 12985 18468
rect 18546 18524 18610 18528
rect 18546 18468 18550 18524
rect 18550 18468 18606 18524
rect 18606 18468 18610 18524
rect 18546 18464 18610 18468
rect 18626 18524 18690 18528
rect 18626 18468 18630 18524
rect 18630 18468 18686 18524
rect 18686 18468 18690 18524
rect 18626 18464 18690 18468
rect 18706 18524 18770 18528
rect 18706 18468 18710 18524
rect 18710 18468 18766 18524
rect 18766 18468 18770 18524
rect 18706 18464 18770 18468
rect 18786 18524 18850 18528
rect 18786 18468 18790 18524
rect 18790 18468 18846 18524
rect 18846 18468 18850 18524
rect 18786 18464 18850 18468
rect 24411 18524 24475 18528
rect 24411 18468 24415 18524
rect 24415 18468 24471 18524
rect 24471 18468 24475 18524
rect 24411 18464 24475 18468
rect 24491 18524 24555 18528
rect 24491 18468 24495 18524
rect 24495 18468 24551 18524
rect 24551 18468 24555 18524
rect 24491 18464 24555 18468
rect 24571 18524 24635 18528
rect 24571 18468 24575 18524
rect 24575 18468 24631 18524
rect 24631 18468 24635 18524
rect 24571 18464 24635 18468
rect 24651 18524 24715 18528
rect 24651 18468 24655 18524
rect 24655 18468 24711 18524
rect 24711 18468 24715 18524
rect 24651 18464 24715 18468
rect 8708 18396 8772 18460
rect 6316 17988 6380 18052
rect 3884 17980 3948 17984
rect 3884 17924 3888 17980
rect 3888 17924 3944 17980
rect 3944 17924 3948 17980
rect 3884 17920 3948 17924
rect 3964 17980 4028 17984
rect 3964 17924 3968 17980
rect 3968 17924 4024 17980
rect 4024 17924 4028 17980
rect 3964 17920 4028 17924
rect 4044 17980 4108 17984
rect 4044 17924 4048 17980
rect 4048 17924 4104 17980
rect 4104 17924 4108 17980
rect 4044 17920 4108 17924
rect 4124 17980 4188 17984
rect 4124 17924 4128 17980
rect 4128 17924 4184 17980
rect 4184 17924 4188 17980
rect 4124 17920 4188 17924
rect 9749 17980 9813 17984
rect 9749 17924 9753 17980
rect 9753 17924 9809 17980
rect 9809 17924 9813 17980
rect 9749 17920 9813 17924
rect 9829 17980 9893 17984
rect 9829 17924 9833 17980
rect 9833 17924 9889 17980
rect 9889 17924 9893 17980
rect 9829 17920 9893 17924
rect 9909 17980 9973 17984
rect 9909 17924 9913 17980
rect 9913 17924 9969 17980
rect 9969 17924 9973 17980
rect 9909 17920 9973 17924
rect 9989 17980 10053 17984
rect 9989 17924 9993 17980
rect 9993 17924 10049 17980
rect 10049 17924 10053 17980
rect 9989 17920 10053 17924
rect 15614 17980 15678 17984
rect 15614 17924 15618 17980
rect 15618 17924 15674 17980
rect 15674 17924 15678 17980
rect 15614 17920 15678 17924
rect 15694 17980 15758 17984
rect 15694 17924 15698 17980
rect 15698 17924 15754 17980
rect 15754 17924 15758 17980
rect 15694 17920 15758 17924
rect 15774 17980 15838 17984
rect 15774 17924 15778 17980
rect 15778 17924 15834 17980
rect 15834 17924 15838 17980
rect 15774 17920 15838 17924
rect 15854 17980 15918 17984
rect 15854 17924 15858 17980
rect 15858 17924 15914 17980
rect 15914 17924 15918 17980
rect 15854 17920 15918 17924
rect 21479 17980 21543 17984
rect 21479 17924 21483 17980
rect 21483 17924 21539 17980
rect 21539 17924 21543 17980
rect 21479 17920 21543 17924
rect 21559 17980 21623 17984
rect 21559 17924 21563 17980
rect 21563 17924 21619 17980
rect 21619 17924 21623 17980
rect 21559 17920 21623 17924
rect 21639 17980 21703 17984
rect 21639 17924 21643 17980
rect 21643 17924 21699 17980
rect 21699 17924 21703 17980
rect 21639 17920 21703 17924
rect 21719 17980 21783 17984
rect 21719 17924 21723 17980
rect 21723 17924 21779 17980
rect 21779 17924 21783 17980
rect 21719 17920 21783 17924
rect 5764 17852 5828 17916
rect 13860 17716 13924 17780
rect 16252 17716 16316 17780
rect 3004 17444 3068 17508
rect 6816 17436 6880 17440
rect 6816 17380 6820 17436
rect 6820 17380 6876 17436
rect 6876 17380 6880 17436
rect 6816 17376 6880 17380
rect 6896 17436 6960 17440
rect 6896 17380 6900 17436
rect 6900 17380 6956 17436
rect 6956 17380 6960 17436
rect 6896 17376 6960 17380
rect 6976 17436 7040 17440
rect 6976 17380 6980 17436
rect 6980 17380 7036 17436
rect 7036 17380 7040 17436
rect 6976 17376 7040 17380
rect 7056 17436 7120 17440
rect 7056 17380 7060 17436
rect 7060 17380 7116 17436
rect 7116 17380 7120 17436
rect 7056 17376 7120 17380
rect 12681 17436 12745 17440
rect 12681 17380 12685 17436
rect 12685 17380 12741 17436
rect 12741 17380 12745 17436
rect 12681 17376 12745 17380
rect 12761 17436 12825 17440
rect 12761 17380 12765 17436
rect 12765 17380 12821 17436
rect 12821 17380 12825 17436
rect 12761 17376 12825 17380
rect 12841 17436 12905 17440
rect 12841 17380 12845 17436
rect 12845 17380 12901 17436
rect 12901 17380 12905 17436
rect 12841 17376 12905 17380
rect 12921 17436 12985 17440
rect 12921 17380 12925 17436
rect 12925 17380 12981 17436
rect 12981 17380 12985 17436
rect 12921 17376 12985 17380
rect 18546 17436 18610 17440
rect 18546 17380 18550 17436
rect 18550 17380 18606 17436
rect 18606 17380 18610 17436
rect 18546 17376 18610 17380
rect 18626 17436 18690 17440
rect 18626 17380 18630 17436
rect 18630 17380 18686 17436
rect 18686 17380 18690 17436
rect 18626 17376 18690 17380
rect 18706 17436 18770 17440
rect 18706 17380 18710 17436
rect 18710 17380 18766 17436
rect 18766 17380 18770 17436
rect 18706 17376 18770 17380
rect 18786 17436 18850 17440
rect 18786 17380 18790 17436
rect 18790 17380 18846 17436
rect 18846 17380 18850 17436
rect 18786 17376 18850 17380
rect 24411 17436 24475 17440
rect 24411 17380 24415 17436
rect 24415 17380 24471 17436
rect 24471 17380 24475 17436
rect 24411 17376 24475 17380
rect 24491 17436 24555 17440
rect 24491 17380 24495 17436
rect 24495 17380 24551 17436
rect 24551 17380 24555 17436
rect 24491 17376 24555 17380
rect 24571 17436 24635 17440
rect 24571 17380 24575 17436
rect 24575 17380 24631 17436
rect 24631 17380 24635 17436
rect 24571 17376 24635 17380
rect 24651 17436 24715 17440
rect 24651 17380 24655 17436
rect 24655 17380 24711 17436
rect 24711 17380 24715 17436
rect 24651 17376 24715 17380
rect 1716 17308 1780 17372
rect 6500 17172 6564 17236
rect 3884 16892 3948 16896
rect 3884 16836 3888 16892
rect 3888 16836 3944 16892
rect 3944 16836 3948 16892
rect 3884 16832 3948 16836
rect 3964 16892 4028 16896
rect 3964 16836 3968 16892
rect 3968 16836 4024 16892
rect 4024 16836 4028 16892
rect 3964 16832 4028 16836
rect 4044 16892 4108 16896
rect 4044 16836 4048 16892
rect 4048 16836 4104 16892
rect 4104 16836 4108 16892
rect 4044 16832 4108 16836
rect 4124 16892 4188 16896
rect 4124 16836 4128 16892
rect 4128 16836 4184 16892
rect 4184 16836 4188 16892
rect 4124 16832 4188 16836
rect 9749 16892 9813 16896
rect 9749 16836 9753 16892
rect 9753 16836 9809 16892
rect 9809 16836 9813 16892
rect 9749 16832 9813 16836
rect 9829 16892 9893 16896
rect 9829 16836 9833 16892
rect 9833 16836 9889 16892
rect 9889 16836 9893 16892
rect 9829 16832 9893 16836
rect 9909 16892 9973 16896
rect 9909 16836 9913 16892
rect 9913 16836 9969 16892
rect 9969 16836 9973 16892
rect 9909 16832 9973 16836
rect 9989 16892 10053 16896
rect 9989 16836 9993 16892
rect 9993 16836 10049 16892
rect 10049 16836 10053 16892
rect 9989 16832 10053 16836
rect 15614 16892 15678 16896
rect 15614 16836 15618 16892
rect 15618 16836 15674 16892
rect 15674 16836 15678 16892
rect 15614 16832 15678 16836
rect 15694 16892 15758 16896
rect 15694 16836 15698 16892
rect 15698 16836 15754 16892
rect 15754 16836 15758 16892
rect 15694 16832 15758 16836
rect 15774 16892 15838 16896
rect 15774 16836 15778 16892
rect 15778 16836 15834 16892
rect 15834 16836 15838 16892
rect 15774 16832 15838 16836
rect 15854 16892 15918 16896
rect 15854 16836 15858 16892
rect 15858 16836 15914 16892
rect 15914 16836 15918 16892
rect 15854 16832 15918 16836
rect 21479 16892 21543 16896
rect 21479 16836 21483 16892
rect 21483 16836 21539 16892
rect 21539 16836 21543 16892
rect 21479 16832 21543 16836
rect 21559 16892 21623 16896
rect 21559 16836 21563 16892
rect 21563 16836 21619 16892
rect 21619 16836 21623 16892
rect 21559 16832 21623 16836
rect 21639 16892 21703 16896
rect 21639 16836 21643 16892
rect 21643 16836 21699 16892
rect 21699 16836 21703 16892
rect 21639 16832 21703 16836
rect 21719 16892 21783 16896
rect 21719 16836 21723 16892
rect 21723 16836 21779 16892
rect 21779 16836 21783 16892
rect 21719 16832 21783 16836
rect 9076 16492 9140 16556
rect 10916 16492 10980 16556
rect 20852 16492 20916 16556
rect 6816 16348 6880 16352
rect 6816 16292 6820 16348
rect 6820 16292 6876 16348
rect 6876 16292 6880 16348
rect 6816 16288 6880 16292
rect 6896 16348 6960 16352
rect 6896 16292 6900 16348
rect 6900 16292 6956 16348
rect 6956 16292 6960 16348
rect 6896 16288 6960 16292
rect 6976 16348 7040 16352
rect 6976 16292 6980 16348
rect 6980 16292 7036 16348
rect 7036 16292 7040 16348
rect 6976 16288 7040 16292
rect 7056 16348 7120 16352
rect 7056 16292 7060 16348
rect 7060 16292 7116 16348
rect 7116 16292 7120 16348
rect 7056 16288 7120 16292
rect 12681 16348 12745 16352
rect 12681 16292 12685 16348
rect 12685 16292 12741 16348
rect 12741 16292 12745 16348
rect 12681 16288 12745 16292
rect 12761 16348 12825 16352
rect 12761 16292 12765 16348
rect 12765 16292 12821 16348
rect 12821 16292 12825 16348
rect 12761 16288 12825 16292
rect 12841 16348 12905 16352
rect 12841 16292 12845 16348
rect 12845 16292 12901 16348
rect 12901 16292 12905 16348
rect 12841 16288 12905 16292
rect 12921 16348 12985 16352
rect 12921 16292 12925 16348
rect 12925 16292 12981 16348
rect 12981 16292 12985 16348
rect 12921 16288 12985 16292
rect 18546 16348 18610 16352
rect 18546 16292 18550 16348
rect 18550 16292 18606 16348
rect 18606 16292 18610 16348
rect 18546 16288 18610 16292
rect 18626 16348 18690 16352
rect 18626 16292 18630 16348
rect 18630 16292 18686 16348
rect 18686 16292 18690 16348
rect 18626 16288 18690 16292
rect 18706 16348 18770 16352
rect 18706 16292 18710 16348
rect 18710 16292 18766 16348
rect 18766 16292 18770 16348
rect 18706 16288 18770 16292
rect 18786 16348 18850 16352
rect 18786 16292 18790 16348
rect 18790 16292 18846 16348
rect 18846 16292 18850 16348
rect 18786 16288 18850 16292
rect 24411 16348 24475 16352
rect 24411 16292 24415 16348
rect 24415 16292 24471 16348
rect 24471 16292 24475 16348
rect 24411 16288 24475 16292
rect 24491 16348 24555 16352
rect 24491 16292 24495 16348
rect 24495 16292 24551 16348
rect 24551 16292 24555 16348
rect 24491 16288 24555 16292
rect 24571 16348 24635 16352
rect 24571 16292 24575 16348
rect 24575 16292 24631 16348
rect 24631 16292 24635 16348
rect 24571 16288 24635 16292
rect 24651 16348 24715 16352
rect 24651 16292 24655 16348
rect 24655 16292 24711 16348
rect 24711 16292 24715 16348
rect 24651 16288 24715 16292
rect 5396 16084 5460 16148
rect 14964 16084 15028 16148
rect 5212 15812 5276 15876
rect 3884 15804 3948 15808
rect 3884 15748 3888 15804
rect 3888 15748 3944 15804
rect 3944 15748 3948 15804
rect 3884 15744 3948 15748
rect 3964 15804 4028 15808
rect 3964 15748 3968 15804
rect 3968 15748 4024 15804
rect 4024 15748 4028 15804
rect 3964 15744 4028 15748
rect 4044 15804 4108 15808
rect 4044 15748 4048 15804
rect 4048 15748 4104 15804
rect 4104 15748 4108 15804
rect 4044 15744 4108 15748
rect 4124 15804 4188 15808
rect 4124 15748 4128 15804
rect 4128 15748 4184 15804
rect 4184 15748 4188 15804
rect 4124 15744 4188 15748
rect 9749 15804 9813 15808
rect 9749 15748 9753 15804
rect 9753 15748 9809 15804
rect 9809 15748 9813 15804
rect 9749 15744 9813 15748
rect 9829 15804 9893 15808
rect 9829 15748 9833 15804
rect 9833 15748 9889 15804
rect 9889 15748 9893 15804
rect 9829 15744 9893 15748
rect 9909 15804 9973 15808
rect 9909 15748 9913 15804
rect 9913 15748 9969 15804
rect 9969 15748 9973 15804
rect 9909 15744 9973 15748
rect 9989 15804 10053 15808
rect 9989 15748 9993 15804
rect 9993 15748 10049 15804
rect 10049 15748 10053 15804
rect 9989 15744 10053 15748
rect 15614 15804 15678 15808
rect 15614 15748 15618 15804
rect 15618 15748 15674 15804
rect 15674 15748 15678 15804
rect 15614 15744 15678 15748
rect 15694 15804 15758 15808
rect 15694 15748 15698 15804
rect 15698 15748 15754 15804
rect 15754 15748 15758 15804
rect 15694 15744 15758 15748
rect 15774 15804 15838 15808
rect 15774 15748 15778 15804
rect 15778 15748 15834 15804
rect 15834 15748 15838 15804
rect 15774 15744 15838 15748
rect 15854 15804 15918 15808
rect 15854 15748 15858 15804
rect 15858 15748 15914 15804
rect 15914 15748 15918 15804
rect 15854 15744 15918 15748
rect 21479 15804 21543 15808
rect 21479 15748 21483 15804
rect 21483 15748 21539 15804
rect 21539 15748 21543 15804
rect 21479 15744 21543 15748
rect 21559 15804 21623 15808
rect 21559 15748 21563 15804
rect 21563 15748 21619 15804
rect 21619 15748 21623 15804
rect 21559 15744 21623 15748
rect 21639 15804 21703 15808
rect 21639 15748 21643 15804
rect 21643 15748 21699 15804
rect 21699 15748 21703 15804
rect 21639 15744 21703 15748
rect 21719 15804 21783 15808
rect 21719 15748 21723 15804
rect 21723 15748 21779 15804
rect 21779 15748 21783 15804
rect 21719 15744 21783 15748
rect 1900 15676 1964 15740
rect 14780 15464 14844 15468
rect 14780 15408 14794 15464
rect 14794 15408 14844 15464
rect 14780 15404 14844 15408
rect 2636 15268 2700 15332
rect 6816 15260 6880 15264
rect 6816 15204 6820 15260
rect 6820 15204 6876 15260
rect 6876 15204 6880 15260
rect 6816 15200 6880 15204
rect 6896 15260 6960 15264
rect 6896 15204 6900 15260
rect 6900 15204 6956 15260
rect 6956 15204 6960 15260
rect 6896 15200 6960 15204
rect 6976 15260 7040 15264
rect 6976 15204 6980 15260
rect 6980 15204 7036 15260
rect 7036 15204 7040 15260
rect 6976 15200 7040 15204
rect 7056 15260 7120 15264
rect 7056 15204 7060 15260
rect 7060 15204 7116 15260
rect 7116 15204 7120 15260
rect 7056 15200 7120 15204
rect 12681 15260 12745 15264
rect 12681 15204 12685 15260
rect 12685 15204 12741 15260
rect 12741 15204 12745 15260
rect 12681 15200 12745 15204
rect 12761 15260 12825 15264
rect 12761 15204 12765 15260
rect 12765 15204 12821 15260
rect 12821 15204 12825 15260
rect 12761 15200 12825 15204
rect 12841 15260 12905 15264
rect 12841 15204 12845 15260
rect 12845 15204 12901 15260
rect 12901 15204 12905 15260
rect 12841 15200 12905 15204
rect 12921 15260 12985 15264
rect 12921 15204 12925 15260
rect 12925 15204 12981 15260
rect 12981 15204 12985 15260
rect 12921 15200 12985 15204
rect 18546 15260 18610 15264
rect 18546 15204 18550 15260
rect 18550 15204 18606 15260
rect 18606 15204 18610 15260
rect 18546 15200 18610 15204
rect 18626 15260 18690 15264
rect 18626 15204 18630 15260
rect 18630 15204 18686 15260
rect 18686 15204 18690 15260
rect 18626 15200 18690 15204
rect 18706 15260 18770 15264
rect 18706 15204 18710 15260
rect 18710 15204 18766 15260
rect 18766 15204 18770 15260
rect 18706 15200 18770 15204
rect 18786 15260 18850 15264
rect 18786 15204 18790 15260
rect 18790 15204 18846 15260
rect 18846 15204 18850 15260
rect 18786 15200 18850 15204
rect 24411 15260 24475 15264
rect 24411 15204 24415 15260
rect 24415 15204 24471 15260
rect 24471 15204 24475 15260
rect 24411 15200 24475 15204
rect 24491 15260 24555 15264
rect 24491 15204 24495 15260
rect 24495 15204 24551 15260
rect 24551 15204 24555 15260
rect 24491 15200 24555 15204
rect 24571 15260 24635 15264
rect 24571 15204 24575 15260
rect 24575 15204 24631 15260
rect 24631 15204 24635 15260
rect 24571 15200 24635 15204
rect 24651 15260 24715 15264
rect 24651 15204 24655 15260
rect 24655 15204 24711 15260
rect 24711 15204 24715 15260
rect 24651 15200 24715 15204
rect 8340 15132 8404 15196
rect 17724 15132 17788 15196
rect 2268 14860 2332 14924
rect 5580 14860 5644 14924
rect 3884 14716 3948 14720
rect 3884 14660 3888 14716
rect 3888 14660 3944 14716
rect 3944 14660 3948 14716
rect 3884 14656 3948 14660
rect 3964 14716 4028 14720
rect 3964 14660 3968 14716
rect 3968 14660 4024 14716
rect 4024 14660 4028 14716
rect 3964 14656 4028 14660
rect 4044 14716 4108 14720
rect 4044 14660 4048 14716
rect 4048 14660 4104 14716
rect 4104 14660 4108 14716
rect 4044 14656 4108 14660
rect 4124 14716 4188 14720
rect 4124 14660 4128 14716
rect 4128 14660 4184 14716
rect 4184 14660 4188 14716
rect 4124 14656 4188 14660
rect 9749 14716 9813 14720
rect 9749 14660 9753 14716
rect 9753 14660 9809 14716
rect 9809 14660 9813 14716
rect 9749 14656 9813 14660
rect 9829 14716 9893 14720
rect 9829 14660 9833 14716
rect 9833 14660 9889 14716
rect 9889 14660 9893 14716
rect 9829 14656 9893 14660
rect 9909 14716 9973 14720
rect 9909 14660 9913 14716
rect 9913 14660 9969 14716
rect 9969 14660 9973 14716
rect 9909 14656 9973 14660
rect 9989 14716 10053 14720
rect 9989 14660 9993 14716
rect 9993 14660 10049 14716
rect 10049 14660 10053 14716
rect 9989 14656 10053 14660
rect 15614 14716 15678 14720
rect 15614 14660 15618 14716
rect 15618 14660 15674 14716
rect 15674 14660 15678 14716
rect 15614 14656 15678 14660
rect 15694 14716 15758 14720
rect 15694 14660 15698 14716
rect 15698 14660 15754 14716
rect 15754 14660 15758 14716
rect 15694 14656 15758 14660
rect 15774 14716 15838 14720
rect 15774 14660 15778 14716
rect 15778 14660 15834 14716
rect 15834 14660 15838 14716
rect 15774 14656 15838 14660
rect 15854 14716 15918 14720
rect 15854 14660 15858 14716
rect 15858 14660 15914 14716
rect 15914 14660 15918 14716
rect 15854 14656 15918 14660
rect 21479 14716 21543 14720
rect 21479 14660 21483 14716
rect 21483 14660 21539 14716
rect 21539 14660 21543 14716
rect 21479 14656 21543 14660
rect 21559 14716 21623 14720
rect 21559 14660 21563 14716
rect 21563 14660 21619 14716
rect 21619 14660 21623 14716
rect 21559 14656 21623 14660
rect 21639 14716 21703 14720
rect 21639 14660 21643 14716
rect 21643 14660 21699 14716
rect 21699 14660 21703 14716
rect 21639 14656 21703 14660
rect 21719 14716 21783 14720
rect 21719 14660 21723 14716
rect 21723 14660 21779 14716
rect 21779 14660 21783 14716
rect 21719 14656 21783 14660
rect 6132 14316 6196 14380
rect 6816 14172 6880 14176
rect 6816 14116 6820 14172
rect 6820 14116 6876 14172
rect 6876 14116 6880 14172
rect 6816 14112 6880 14116
rect 6896 14172 6960 14176
rect 6896 14116 6900 14172
rect 6900 14116 6956 14172
rect 6956 14116 6960 14172
rect 6896 14112 6960 14116
rect 6976 14172 7040 14176
rect 6976 14116 6980 14172
rect 6980 14116 7036 14172
rect 7036 14116 7040 14172
rect 6976 14112 7040 14116
rect 7056 14172 7120 14176
rect 7056 14116 7060 14172
rect 7060 14116 7116 14172
rect 7116 14116 7120 14172
rect 7056 14112 7120 14116
rect 12681 14172 12745 14176
rect 12681 14116 12685 14172
rect 12685 14116 12741 14172
rect 12741 14116 12745 14172
rect 12681 14112 12745 14116
rect 12761 14172 12825 14176
rect 12761 14116 12765 14172
rect 12765 14116 12821 14172
rect 12821 14116 12825 14172
rect 12761 14112 12825 14116
rect 12841 14172 12905 14176
rect 12841 14116 12845 14172
rect 12845 14116 12901 14172
rect 12901 14116 12905 14172
rect 12841 14112 12905 14116
rect 12921 14172 12985 14176
rect 12921 14116 12925 14172
rect 12925 14116 12981 14172
rect 12981 14116 12985 14172
rect 12921 14112 12985 14116
rect 18546 14172 18610 14176
rect 18546 14116 18550 14172
rect 18550 14116 18606 14172
rect 18606 14116 18610 14172
rect 18546 14112 18610 14116
rect 18626 14172 18690 14176
rect 18626 14116 18630 14172
rect 18630 14116 18686 14172
rect 18686 14116 18690 14172
rect 18626 14112 18690 14116
rect 18706 14172 18770 14176
rect 18706 14116 18710 14172
rect 18710 14116 18766 14172
rect 18766 14116 18770 14172
rect 18706 14112 18770 14116
rect 18786 14172 18850 14176
rect 18786 14116 18790 14172
rect 18790 14116 18846 14172
rect 18846 14116 18850 14172
rect 18786 14112 18850 14116
rect 24411 14172 24475 14176
rect 24411 14116 24415 14172
rect 24415 14116 24471 14172
rect 24471 14116 24475 14172
rect 24411 14112 24475 14116
rect 24491 14172 24555 14176
rect 24491 14116 24495 14172
rect 24495 14116 24551 14172
rect 24551 14116 24555 14172
rect 24491 14112 24555 14116
rect 24571 14172 24635 14176
rect 24571 14116 24575 14172
rect 24575 14116 24631 14172
rect 24631 14116 24635 14172
rect 24571 14112 24635 14116
rect 24651 14172 24715 14176
rect 24651 14116 24655 14172
rect 24655 14116 24711 14172
rect 24711 14116 24715 14172
rect 24651 14112 24715 14116
rect 21220 13772 21284 13836
rect 3884 13628 3948 13632
rect 3884 13572 3888 13628
rect 3888 13572 3944 13628
rect 3944 13572 3948 13628
rect 3884 13568 3948 13572
rect 3964 13628 4028 13632
rect 3964 13572 3968 13628
rect 3968 13572 4024 13628
rect 4024 13572 4028 13628
rect 3964 13568 4028 13572
rect 4044 13628 4108 13632
rect 4044 13572 4048 13628
rect 4048 13572 4104 13628
rect 4104 13572 4108 13628
rect 4044 13568 4108 13572
rect 4124 13628 4188 13632
rect 4124 13572 4128 13628
rect 4128 13572 4184 13628
rect 4184 13572 4188 13628
rect 4124 13568 4188 13572
rect 9749 13628 9813 13632
rect 9749 13572 9753 13628
rect 9753 13572 9809 13628
rect 9809 13572 9813 13628
rect 9749 13568 9813 13572
rect 9829 13628 9893 13632
rect 9829 13572 9833 13628
rect 9833 13572 9889 13628
rect 9889 13572 9893 13628
rect 9829 13568 9893 13572
rect 9909 13628 9973 13632
rect 9909 13572 9913 13628
rect 9913 13572 9969 13628
rect 9969 13572 9973 13628
rect 9909 13568 9973 13572
rect 9989 13628 10053 13632
rect 9989 13572 9993 13628
rect 9993 13572 10049 13628
rect 10049 13572 10053 13628
rect 9989 13568 10053 13572
rect 15614 13628 15678 13632
rect 15614 13572 15618 13628
rect 15618 13572 15674 13628
rect 15674 13572 15678 13628
rect 15614 13568 15678 13572
rect 15694 13628 15758 13632
rect 15694 13572 15698 13628
rect 15698 13572 15754 13628
rect 15754 13572 15758 13628
rect 15694 13568 15758 13572
rect 15774 13628 15838 13632
rect 15774 13572 15778 13628
rect 15778 13572 15834 13628
rect 15834 13572 15838 13628
rect 15774 13568 15838 13572
rect 15854 13628 15918 13632
rect 15854 13572 15858 13628
rect 15858 13572 15914 13628
rect 15914 13572 15918 13628
rect 15854 13568 15918 13572
rect 21479 13628 21543 13632
rect 21479 13572 21483 13628
rect 21483 13572 21539 13628
rect 21539 13572 21543 13628
rect 21479 13568 21543 13572
rect 21559 13628 21623 13632
rect 21559 13572 21563 13628
rect 21563 13572 21619 13628
rect 21619 13572 21623 13628
rect 21559 13568 21623 13572
rect 21639 13628 21703 13632
rect 21639 13572 21643 13628
rect 21643 13572 21699 13628
rect 21699 13572 21703 13628
rect 21639 13568 21703 13572
rect 21719 13628 21783 13632
rect 21719 13572 21723 13628
rect 21723 13572 21779 13628
rect 21779 13572 21783 13628
rect 21719 13568 21783 13572
rect 8524 13092 8588 13156
rect 6816 13084 6880 13088
rect 6816 13028 6820 13084
rect 6820 13028 6876 13084
rect 6876 13028 6880 13084
rect 6816 13024 6880 13028
rect 6896 13084 6960 13088
rect 6896 13028 6900 13084
rect 6900 13028 6956 13084
rect 6956 13028 6960 13084
rect 6896 13024 6960 13028
rect 6976 13084 7040 13088
rect 6976 13028 6980 13084
rect 6980 13028 7036 13084
rect 7036 13028 7040 13084
rect 6976 13024 7040 13028
rect 7056 13084 7120 13088
rect 7056 13028 7060 13084
rect 7060 13028 7116 13084
rect 7116 13028 7120 13084
rect 7056 13024 7120 13028
rect 12681 13084 12745 13088
rect 12681 13028 12685 13084
rect 12685 13028 12741 13084
rect 12741 13028 12745 13084
rect 12681 13024 12745 13028
rect 12761 13084 12825 13088
rect 12761 13028 12765 13084
rect 12765 13028 12821 13084
rect 12821 13028 12825 13084
rect 12761 13024 12825 13028
rect 12841 13084 12905 13088
rect 12841 13028 12845 13084
rect 12845 13028 12901 13084
rect 12901 13028 12905 13084
rect 12841 13024 12905 13028
rect 12921 13084 12985 13088
rect 12921 13028 12925 13084
rect 12925 13028 12981 13084
rect 12981 13028 12985 13084
rect 12921 13024 12985 13028
rect 18546 13084 18610 13088
rect 18546 13028 18550 13084
rect 18550 13028 18606 13084
rect 18606 13028 18610 13084
rect 18546 13024 18610 13028
rect 18626 13084 18690 13088
rect 18626 13028 18630 13084
rect 18630 13028 18686 13084
rect 18686 13028 18690 13084
rect 18626 13024 18690 13028
rect 18706 13084 18770 13088
rect 18706 13028 18710 13084
rect 18710 13028 18766 13084
rect 18766 13028 18770 13084
rect 18706 13024 18770 13028
rect 18786 13084 18850 13088
rect 18786 13028 18790 13084
rect 18790 13028 18846 13084
rect 18846 13028 18850 13084
rect 18786 13024 18850 13028
rect 24411 13084 24475 13088
rect 24411 13028 24415 13084
rect 24415 13028 24471 13084
rect 24471 13028 24475 13084
rect 24411 13024 24475 13028
rect 24491 13084 24555 13088
rect 24491 13028 24495 13084
rect 24495 13028 24551 13084
rect 24551 13028 24555 13084
rect 24491 13024 24555 13028
rect 24571 13084 24635 13088
rect 24571 13028 24575 13084
rect 24575 13028 24631 13084
rect 24631 13028 24635 13084
rect 24571 13024 24635 13028
rect 24651 13084 24715 13088
rect 24651 13028 24655 13084
rect 24655 13028 24711 13084
rect 24711 13028 24715 13084
rect 24651 13024 24715 13028
rect 21036 12820 21100 12884
rect 12388 12684 12452 12748
rect 13124 12684 13188 12748
rect 4476 12608 4540 12612
rect 4476 12552 4490 12608
rect 4490 12552 4540 12608
rect 4476 12548 4540 12552
rect 3884 12540 3948 12544
rect 3884 12484 3888 12540
rect 3888 12484 3944 12540
rect 3944 12484 3948 12540
rect 3884 12480 3948 12484
rect 3964 12540 4028 12544
rect 3964 12484 3968 12540
rect 3968 12484 4024 12540
rect 4024 12484 4028 12540
rect 3964 12480 4028 12484
rect 4044 12540 4108 12544
rect 4044 12484 4048 12540
rect 4048 12484 4104 12540
rect 4104 12484 4108 12540
rect 4044 12480 4108 12484
rect 4124 12540 4188 12544
rect 4124 12484 4128 12540
rect 4128 12484 4184 12540
rect 4184 12484 4188 12540
rect 4124 12480 4188 12484
rect 9749 12540 9813 12544
rect 9749 12484 9753 12540
rect 9753 12484 9809 12540
rect 9809 12484 9813 12540
rect 9749 12480 9813 12484
rect 9829 12540 9893 12544
rect 9829 12484 9833 12540
rect 9833 12484 9889 12540
rect 9889 12484 9893 12540
rect 9829 12480 9893 12484
rect 9909 12540 9973 12544
rect 9909 12484 9913 12540
rect 9913 12484 9969 12540
rect 9969 12484 9973 12540
rect 9909 12480 9973 12484
rect 9989 12540 10053 12544
rect 9989 12484 9993 12540
rect 9993 12484 10049 12540
rect 10049 12484 10053 12540
rect 9989 12480 10053 12484
rect 15614 12540 15678 12544
rect 15614 12484 15618 12540
rect 15618 12484 15674 12540
rect 15674 12484 15678 12540
rect 15614 12480 15678 12484
rect 15694 12540 15758 12544
rect 15694 12484 15698 12540
rect 15698 12484 15754 12540
rect 15754 12484 15758 12540
rect 15694 12480 15758 12484
rect 15774 12540 15838 12544
rect 15774 12484 15778 12540
rect 15778 12484 15834 12540
rect 15834 12484 15838 12540
rect 15774 12480 15838 12484
rect 15854 12540 15918 12544
rect 15854 12484 15858 12540
rect 15858 12484 15914 12540
rect 15914 12484 15918 12540
rect 15854 12480 15918 12484
rect 21479 12540 21543 12544
rect 21479 12484 21483 12540
rect 21483 12484 21539 12540
rect 21539 12484 21543 12540
rect 21479 12480 21543 12484
rect 21559 12540 21623 12544
rect 21559 12484 21563 12540
rect 21563 12484 21619 12540
rect 21619 12484 21623 12540
rect 21559 12480 21623 12484
rect 21639 12540 21703 12544
rect 21639 12484 21643 12540
rect 21643 12484 21699 12540
rect 21699 12484 21703 12540
rect 21639 12480 21703 12484
rect 21719 12540 21783 12544
rect 21719 12484 21723 12540
rect 21723 12484 21779 12540
rect 21779 12484 21783 12540
rect 21719 12480 21783 12484
rect 19564 12412 19628 12476
rect 1532 12200 1596 12204
rect 1532 12144 1546 12200
rect 1546 12144 1596 12200
rect 1532 12140 1596 12144
rect 2084 12140 2148 12204
rect 7420 12140 7484 12204
rect 12388 12140 12452 12204
rect 13124 12140 13188 12204
rect 13860 12276 13924 12340
rect 19564 12004 19628 12068
rect 6816 11996 6880 12000
rect 6816 11940 6820 11996
rect 6820 11940 6876 11996
rect 6876 11940 6880 11996
rect 6816 11936 6880 11940
rect 6896 11996 6960 12000
rect 6896 11940 6900 11996
rect 6900 11940 6956 11996
rect 6956 11940 6960 11996
rect 6896 11936 6960 11940
rect 6976 11996 7040 12000
rect 6976 11940 6980 11996
rect 6980 11940 7036 11996
rect 7036 11940 7040 11996
rect 6976 11936 7040 11940
rect 7056 11996 7120 12000
rect 7056 11940 7060 11996
rect 7060 11940 7116 11996
rect 7116 11940 7120 11996
rect 7056 11936 7120 11940
rect 12681 11996 12745 12000
rect 12681 11940 12685 11996
rect 12685 11940 12741 11996
rect 12741 11940 12745 11996
rect 12681 11936 12745 11940
rect 12761 11996 12825 12000
rect 12761 11940 12765 11996
rect 12765 11940 12821 11996
rect 12821 11940 12825 11996
rect 12761 11936 12825 11940
rect 12841 11996 12905 12000
rect 12841 11940 12845 11996
rect 12845 11940 12901 11996
rect 12901 11940 12905 11996
rect 12841 11936 12905 11940
rect 12921 11996 12985 12000
rect 12921 11940 12925 11996
rect 12925 11940 12981 11996
rect 12981 11940 12985 11996
rect 12921 11936 12985 11940
rect 18546 11996 18610 12000
rect 18546 11940 18550 11996
rect 18550 11940 18606 11996
rect 18606 11940 18610 11996
rect 18546 11936 18610 11940
rect 18626 11996 18690 12000
rect 18626 11940 18630 11996
rect 18630 11940 18686 11996
rect 18686 11940 18690 11996
rect 18626 11936 18690 11940
rect 18706 11996 18770 12000
rect 18706 11940 18710 11996
rect 18710 11940 18766 11996
rect 18766 11940 18770 11996
rect 18706 11936 18770 11940
rect 18786 11996 18850 12000
rect 18786 11940 18790 11996
rect 18790 11940 18846 11996
rect 18846 11940 18850 11996
rect 18786 11936 18850 11940
rect 24411 11996 24475 12000
rect 24411 11940 24415 11996
rect 24415 11940 24471 11996
rect 24471 11940 24475 11996
rect 24411 11936 24475 11940
rect 24491 11996 24555 12000
rect 24491 11940 24495 11996
rect 24495 11940 24551 11996
rect 24551 11940 24555 11996
rect 24491 11936 24555 11940
rect 24571 11996 24635 12000
rect 24571 11940 24575 11996
rect 24575 11940 24631 11996
rect 24631 11940 24635 11996
rect 24571 11936 24635 11940
rect 24651 11996 24715 12000
rect 24651 11940 24655 11996
rect 24655 11940 24711 11996
rect 24711 11940 24715 11996
rect 24651 11936 24715 11940
rect 4476 11868 4540 11932
rect 13860 11596 13924 11660
rect 10732 11460 10796 11524
rect 3884 11452 3948 11456
rect 3884 11396 3888 11452
rect 3888 11396 3944 11452
rect 3944 11396 3948 11452
rect 3884 11392 3948 11396
rect 3964 11452 4028 11456
rect 3964 11396 3968 11452
rect 3968 11396 4024 11452
rect 4024 11396 4028 11452
rect 3964 11392 4028 11396
rect 4044 11452 4108 11456
rect 4044 11396 4048 11452
rect 4048 11396 4104 11452
rect 4104 11396 4108 11452
rect 4044 11392 4108 11396
rect 4124 11452 4188 11456
rect 4124 11396 4128 11452
rect 4128 11396 4184 11452
rect 4184 11396 4188 11452
rect 4124 11392 4188 11396
rect 9749 11452 9813 11456
rect 9749 11396 9753 11452
rect 9753 11396 9809 11452
rect 9809 11396 9813 11452
rect 9749 11392 9813 11396
rect 9829 11452 9893 11456
rect 9829 11396 9833 11452
rect 9833 11396 9889 11452
rect 9889 11396 9893 11452
rect 9829 11392 9893 11396
rect 9909 11452 9973 11456
rect 9909 11396 9913 11452
rect 9913 11396 9969 11452
rect 9969 11396 9973 11452
rect 9909 11392 9973 11396
rect 9989 11452 10053 11456
rect 9989 11396 9993 11452
rect 9993 11396 10049 11452
rect 10049 11396 10053 11452
rect 9989 11392 10053 11396
rect 7788 11384 7852 11388
rect 7788 11328 7838 11384
rect 7838 11328 7852 11384
rect 7788 11324 7852 11328
rect 15614 11452 15678 11456
rect 15614 11396 15618 11452
rect 15618 11396 15674 11452
rect 15674 11396 15678 11452
rect 15614 11392 15678 11396
rect 15694 11452 15758 11456
rect 15694 11396 15698 11452
rect 15698 11396 15754 11452
rect 15754 11396 15758 11452
rect 15694 11392 15758 11396
rect 15774 11452 15838 11456
rect 15774 11396 15778 11452
rect 15778 11396 15834 11452
rect 15834 11396 15838 11452
rect 15774 11392 15838 11396
rect 15854 11452 15918 11456
rect 15854 11396 15858 11452
rect 15858 11396 15914 11452
rect 15914 11396 15918 11452
rect 15854 11392 15918 11396
rect 21479 11452 21543 11456
rect 21479 11396 21483 11452
rect 21483 11396 21539 11452
rect 21539 11396 21543 11452
rect 21479 11392 21543 11396
rect 21559 11452 21623 11456
rect 21559 11396 21563 11452
rect 21563 11396 21619 11452
rect 21619 11396 21623 11452
rect 21559 11392 21623 11396
rect 21639 11452 21703 11456
rect 21639 11396 21643 11452
rect 21643 11396 21699 11452
rect 21699 11396 21703 11452
rect 21639 11392 21703 11396
rect 21719 11452 21783 11456
rect 21719 11396 21723 11452
rect 21723 11396 21779 11452
rect 21779 11396 21783 11452
rect 21719 11392 21783 11396
rect 5396 11052 5460 11116
rect 7420 11052 7484 11116
rect 10364 11052 10428 11116
rect 11836 11052 11900 11116
rect 14412 11052 14476 11116
rect 4292 10916 4356 10980
rect 6816 10908 6880 10912
rect 6816 10852 6820 10908
rect 6820 10852 6876 10908
rect 6876 10852 6880 10908
rect 6816 10848 6880 10852
rect 6896 10908 6960 10912
rect 6896 10852 6900 10908
rect 6900 10852 6956 10908
rect 6956 10852 6960 10908
rect 6896 10848 6960 10852
rect 6976 10908 7040 10912
rect 6976 10852 6980 10908
rect 6980 10852 7036 10908
rect 7036 10852 7040 10908
rect 6976 10848 7040 10852
rect 7056 10908 7120 10912
rect 7056 10852 7060 10908
rect 7060 10852 7116 10908
rect 7116 10852 7120 10908
rect 7056 10848 7120 10852
rect 12681 10908 12745 10912
rect 12681 10852 12685 10908
rect 12685 10852 12741 10908
rect 12741 10852 12745 10908
rect 12681 10848 12745 10852
rect 12761 10908 12825 10912
rect 12761 10852 12765 10908
rect 12765 10852 12821 10908
rect 12821 10852 12825 10908
rect 12761 10848 12825 10852
rect 12841 10908 12905 10912
rect 12841 10852 12845 10908
rect 12845 10852 12901 10908
rect 12901 10852 12905 10908
rect 12841 10848 12905 10852
rect 12921 10908 12985 10912
rect 12921 10852 12925 10908
rect 12925 10852 12981 10908
rect 12981 10852 12985 10908
rect 12921 10848 12985 10852
rect 18546 10908 18610 10912
rect 18546 10852 18550 10908
rect 18550 10852 18606 10908
rect 18606 10852 18610 10908
rect 18546 10848 18610 10852
rect 18626 10908 18690 10912
rect 18626 10852 18630 10908
rect 18630 10852 18686 10908
rect 18686 10852 18690 10908
rect 18626 10848 18690 10852
rect 18706 10908 18770 10912
rect 18706 10852 18710 10908
rect 18710 10852 18766 10908
rect 18766 10852 18770 10908
rect 18706 10848 18770 10852
rect 18786 10908 18850 10912
rect 18786 10852 18790 10908
rect 18790 10852 18846 10908
rect 18846 10852 18850 10908
rect 18786 10848 18850 10852
rect 24411 10908 24475 10912
rect 24411 10852 24415 10908
rect 24415 10852 24471 10908
rect 24471 10852 24475 10908
rect 24411 10848 24475 10852
rect 24491 10908 24555 10912
rect 24491 10852 24495 10908
rect 24495 10852 24551 10908
rect 24551 10852 24555 10908
rect 24491 10848 24555 10852
rect 24571 10908 24635 10912
rect 24571 10852 24575 10908
rect 24575 10852 24631 10908
rect 24631 10852 24635 10908
rect 24571 10848 24635 10852
rect 24651 10908 24715 10912
rect 24651 10852 24655 10908
rect 24655 10852 24711 10908
rect 24711 10852 24715 10908
rect 24651 10848 24715 10852
rect 3004 10508 3068 10572
rect 3884 10364 3948 10368
rect 3884 10308 3888 10364
rect 3888 10308 3944 10364
rect 3944 10308 3948 10364
rect 3884 10304 3948 10308
rect 3964 10364 4028 10368
rect 3964 10308 3968 10364
rect 3968 10308 4024 10364
rect 4024 10308 4028 10364
rect 3964 10304 4028 10308
rect 4044 10364 4108 10368
rect 4044 10308 4048 10364
rect 4048 10308 4104 10364
rect 4104 10308 4108 10364
rect 4044 10304 4108 10308
rect 4124 10364 4188 10368
rect 4124 10308 4128 10364
rect 4128 10308 4184 10364
rect 4184 10308 4188 10364
rect 4124 10304 4188 10308
rect 9749 10364 9813 10368
rect 9749 10308 9753 10364
rect 9753 10308 9809 10364
rect 9809 10308 9813 10364
rect 9749 10304 9813 10308
rect 9829 10364 9893 10368
rect 9829 10308 9833 10364
rect 9833 10308 9889 10364
rect 9889 10308 9893 10364
rect 9829 10304 9893 10308
rect 9909 10364 9973 10368
rect 9909 10308 9913 10364
rect 9913 10308 9969 10364
rect 9969 10308 9973 10364
rect 9909 10304 9973 10308
rect 9989 10364 10053 10368
rect 9989 10308 9993 10364
rect 9993 10308 10049 10364
rect 10049 10308 10053 10364
rect 9989 10304 10053 10308
rect 15614 10364 15678 10368
rect 15614 10308 15618 10364
rect 15618 10308 15674 10364
rect 15674 10308 15678 10364
rect 15614 10304 15678 10308
rect 15694 10364 15758 10368
rect 15694 10308 15698 10364
rect 15698 10308 15754 10364
rect 15754 10308 15758 10364
rect 15694 10304 15758 10308
rect 15774 10364 15838 10368
rect 15774 10308 15778 10364
rect 15778 10308 15834 10364
rect 15834 10308 15838 10364
rect 15774 10304 15838 10308
rect 15854 10364 15918 10368
rect 15854 10308 15858 10364
rect 15858 10308 15914 10364
rect 15914 10308 15918 10364
rect 15854 10304 15918 10308
rect 21479 10364 21543 10368
rect 21479 10308 21483 10364
rect 21483 10308 21539 10364
rect 21539 10308 21543 10364
rect 21479 10304 21543 10308
rect 21559 10364 21623 10368
rect 21559 10308 21563 10364
rect 21563 10308 21619 10364
rect 21619 10308 21623 10364
rect 21559 10304 21623 10308
rect 21639 10364 21703 10368
rect 21639 10308 21643 10364
rect 21643 10308 21699 10364
rect 21699 10308 21703 10364
rect 21639 10304 21703 10308
rect 21719 10364 21783 10368
rect 21719 10308 21723 10364
rect 21723 10308 21779 10364
rect 21779 10308 21783 10364
rect 21719 10304 21783 10308
rect 22692 10100 22756 10164
rect 5028 9828 5092 9892
rect 6816 9820 6880 9824
rect 6816 9764 6820 9820
rect 6820 9764 6876 9820
rect 6876 9764 6880 9820
rect 6816 9760 6880 9764
rect 6896 9820 6960 9824
rect 6896 9764 6900 9820
rect 6900 9764 6956 9820
rect 6956 9764 6960 9820
rect 6896 9760 6960 9764
rect 6976 9820 7040 9824
rect 6976 9764 6980 9820
rect 6980 9764 7036 9820
rect 7036 9764 7040 9820
rect 6976 9760 7040 9764
rect 7056 9820 7120 9824
rect 7056 9764 7060 9820
rect 7060 9764 7116 9820
rect 7116 9764 7120 9820
rect 7056 9760 7120 9764
rect 12681 9820 12745 9824
rect 12681 9764 12685 9820
rect 12685 9764 12741 9820
rect 12741 9764 12745 9820
rect 12681 9760 12745 9764
rect 12761 9820 12825 9824
rect 12761 9764 12765 9820
rect 12765 9764 12821 9820
rect 12821 9764 12825 9820
rect 12761 9760 12825 9764
rect 12841 9820 12905 9824
rect 12841 9764 12845 9820
rect 12845 9764 12901 9820
rect 12901 9764 12905 9820
rect 12841 9760 12905 9764
rect 12921 9820 12985 9824
rect 12921 9764 12925 9820
rect 12925 9764 12981 9820
rect 12981 9764 12985 9820
rect 12921 9760 12985 9764
rect 18546 9820 18610 9824
rect 18546 9764 18550 9820
rect 18550 9764 18606 9820
rect 18606 9764 18610 9820
rect 18546 9760 18610 9764
rect 18626 9820 18690 9824
rect 18626 9764 18630 9820
rect 18630 9764 18686 9820
rect 18686 9764 18690 9820
rect 18626 9760 18690 9764
rect 18706 9820 18770 9824
rect 18706 9764 18710 9820
rect 18710 9764 18766 9820
rect 18766 9764 18770 9820
rect 18706 9760 18770 9764
rect 18786 9820 18850 9824
rect 18786 9764 18790 9820
rect 18790 9764 18846 9820
rect 18846 9764 18850 9820
rect 18786 9760 18850 9764
rect 24411 9820 24475 9824
rect 24411 9764 24415 9820
rect 24415 9764 24471 9820
rect 24471 9764 24475 9820
rect 24411 9760 24475 9764
rect 24491 9820 24555 9824
rect 24491 9764 24495 9820
rect 24495 9764 24551 9820
rect 24551 9764 24555 9820
rect 24491 9760 24555 9764
rect 24571 9820 24635 9824
rect 24571 9764 24575 9820
rect 24575 9764 24631 9820
rect 24631 9764 24635 9820
rect 24571 9760 24635 9764
rect 24651 9820 24715 9824
rect 24651 9764 24655 9820
rect 24655 9764 24711 9820
rect 24711 9764 24715 9820
rect 24651 9760 24715 9764
rect 8156 9692 8220 9756
rect 9260 9692 9324 9756
rect 4292 9616 4356 9620
rect 4292 9560 4342 9616
rect 4342 9560 4356 9616
rect 4292 9556 4356 9560
rect 3884 9276 3948 9280
rect 3884 9220 3888 9276
rect 3888 9220 3944 9276
rect 3944 9220 3948 9276
rect 3884 9216 3948 9220
rect 3964 9276 4028 9280
rect 3964 9220 3968 9276
rect 3968 9220 4024 9276
rect 4024 9220 4028 9276
rect 3964 9216 4028 9220
rect 4044 9276 4108 9280
rect 4044 9220 4048 9276
rect 4048 9220 4104 9276
rect 4104 9220 4108 9276
rect 4044 9216 4108 9220
rect 4124 9276 4188 9280
rect 4124 9220 4128 9276
rect 4128 9220 4184 9276
rect 4184 9220 4188 9276
rect 4124 9216 4188 9220
rect 9749 9276 9813 9280
rect 9749 9220 9753 9276
rect 9753 9220 9809 9276
rect 9809 9220 9813 9276
rect 9749 9216 9813 9220
rect 9829 9276 9893 9280
rect 9829 9220 9833 9276
rect 9833 9220 9889 9276
rect 9889 9220 9893 9276
rect 9829 9216 9893 9220
rect 9909 9276 9973 9280
rect 9909 9220 9913 9276
rect 9913 9220 9969 9276
rect 9969 9220 9973 9276
rect 9909 9216 9973 9220
rect 9989 9276 10053 9280
rect 9989 9220 9993 9276
rect 9993 9220 10049 9276
rect 10049 9220 10053 9276
rect 9989 9216 10053 9220
rect 15614 9276 15678 9280
rect 15614 9220 15618 9276
rect 15618 9220 15674 9276
rect 15674 9220 15678 9276
rect 15614 9216 15678 9220
rect 15694 9276 15758 9280
rect 15694 9220 15698 9276
rect 15698 9220 15754 9276
rect 15754 9220 15758 9276
rect 15694 9216 15758 9220
rect 15774 9276 15838 9280
rect 15774 9220 15778 9276
rect 15778 9220 15834 9276
rect 15834 9220 15838 9276
rect 15774 9216 15838 9220
rect 15854 9276 15918 9280
rect 15854 9220 15858 9276
rect 15858 9220 15914 9276
rect 15914 9220 15918 9276
rect 15854 9216 15918 9220
rect 21479 9276 21543 9280
rect 21479 9220 21483 9276
rect 21483 9220 21539 9276
rect 21539 9220 21543 9276
rect 21479 9216 21543 9220
rect 21559 9276 21623 9280
rect 21559 9220 21563 9276
rect 21563 9220 21619 9276
rect 21619 9220 21623 9276
rect 21559 9216 21623 9220
rect 21639 9276 21703 9280
rect 21639 9220 21643 9276
rect 21643 9220 21699 9276
rect 21699 9220 21703 9276
rect 21639 9216 21703 9220
rect 21719 9276 21783 9280
rect 21719 9220 21723 9276
rect 21723 9220 21779 9276
rect 21779 9220 21783 9276
rect 21719 9216 21783 9220
rect 4292 9012 4356 9076
rect 8708 8876 8772 8940
rect 6816 8732 6880 8736
rect 6816 8676 6820 8732
rect 6820 8676 6876 8732
rect 6876 8676 6880 8732
rect 6816 8672 6880 8676
rect 6896 8732 6960 8736
rect 6896 8676 6900 8732
rect 6900 8676 6956 8732
rect 6956 8676 6960 8732
rect 6896 8672 6960 8676
rect 6976 8732 7040 8736
rect 6976 8676 6980 8732
rect 6980 8676 7036 8732
rect 7036 8676 7040 8732
rect 6976 8672 7040 8676
rect 7056 8732 7120 8736
rect 7056 8676 7060 8732
rect 7060 8676 7116 8732
rect 7116 8676 7120 8732
rect 7056 8672 7120 8676
rect 12681 8732 12745 8736
rect 12681 8676 12685 8732
rect 12685 8676 12741 8732
rect 12741 8676 12745 8732
rect 12681 8672 12745 8676
rect 12761 8732 12825 8736
rect 12761 8676 12765 8732
rect 12765 8676 12821 8732
rect 12821 8676 12825 8732
rect 12761 8672 12825 8676
rect 12841 8732 12905 8736
rect 12841 8676 12845 8732
rect 12845 8676 12901 8732
rect 12901 8676 12905 8732
rect 12841 8672 12905 8676
rect 12921 8732 12985 8736
rect 12921 8676 12925 8732
rect 12925 8676 12981 8732
rect 12981 8676 12985 8732
rect 12921 8672 12985 8676
rect 18546 8732 18610 8736
rect 18546 8676 18550 8732
rect 18550 8676 18606 8732
rect 18606 8676 18610 8732
rect 18546 8672 18610 8676
rect 18626 8732 18690 8736
rect 18626 8676 18630 8732
rect 18630 8676 18686 8732
rect 18686 8676 18690 8732
rect 18626 8672 18690 8676
rect 18706 8732 18770 8736
rect 18706 8676 18710 8732
rect 18710 8676 18766 8732
rect 18766 8676 18770 8732
rect 18706 8672 18770 8676
rect 18786 8732 18850 8736
rect 18786 8676 18790 8732
rect 18790 8676 18846 8732
rect 18846 8676 18850 8732
rect 18786 8672 18850 8676
rect 24411 8732 24475 8736
rect 24411 8676 24415 8732
rect 24415 8676 24471 8732
rect 24471 8676 24475 8732
rect 24411 8672 24475 8676
rect 24491 8732 24555 8736
rect 24491 8676 24495 8732
rect 24495 8676 24551 8732
rect 24551 8676 24555 8732
rect 24491 8672 24555 8676
rect 24571 8732 24635 8736
rect 24571 8676 24575 8732
rect 24575 8676 24631 8732
rect 24631 8676 24635 8732
rect 24571 8672 24635 8676
rect 24651 8732 24715 8736
rect 24651 8676 24655 8732
rect 24655 8676 24711 8732
rect 24711 8676 24715 8732
rect 24651 8672 24715 8676
rect 2820 8468 2884 8532
rect 19748 8468 19812 8532
rect 3188 8332 3252 8396
rect 3740 8332 3804 8396
rect 17908 8332 17972 8396
rect 19564 8392 19628 8396
rect 19564 8336 19578 8392
rect 19578 8336 19628 8392
rect 19564 8332 19628 8336
rect 19932 8332 19996 8396
rect 20852 8332 20916 8396
rect 3884 8188 3948 8192
rect 3884 8132 3888 8188
rect 3888 8132 3944 8188
rect 3944 8132 3948 8188
rect 3884 8128 3948 8132
rect 3964 8188 4028 8192
rect 3964 8132 3968 8188
rect 3968 8132 4024 8188
rect 4024 8132 4028 8188
rect 3964 8128 4028 8132
rect 4044 8188 4108 8192
rect 4044 8132 4048 8188
rect 4048 8132 4104 8188
rect 4104 8132 4108 8188
rect 4044 8128 4108 8132
rect 4124 8188 4188 8192
rect 4124 8132 4128 8188
rect 4128 8132 4184 8188
rect 4184 8132 4188 8188
rect 4124 8128 4188 8132
rect 9749 8188 9813 8192
rect 9749 8132 9753 8188
rect 9753 8132 9809 8188
rect 9809 8132 9813 8188
rect 9749 8128 9813 8132
rect 9829 8188 9893 8192
rect 9829 8132 9833 8188
rect 9833 8132 9889 8188
rect 9889 8132 9893 8188
rect 9829 8128 9893 8132
rect 9909 8188 9973 8192
rect 9909 8132 9913 8188
rect 9913 8132 9969 8188
rect 9969 8132 9973 8188
rect 9909 8128 9973 8132
rect 9989 8188 10053 8192
rect 9989 8132 9993 8188
rect 9993 8132 10049 8188
rect 10049 8132 10053 8188
rect 9989 8128 10053 8132
rect 15614 8188 15678 8192
rect 15614 8132 15618 8188
rect 15618 8132 15674 8188
rect 15674 8132 15678 8188
rect 15614 8128 15678 8132
rect 15694 8188 15758 8192
rect 15694 8132 15698 8188
rect 15698 8132 15754 8188
rect 15754 8132 15758 8188
rect 15694 8128 15758 8132
rect 15774 8188 15838 8192
rect 15774 8132 15778 8188
rect 15778 8132 15834 8188
rect 15834 8132 15838 8188
rect 15774 8128 15838 8132
rect 15854 8188 15918 8192
rect 15854 8132 15858 8188
rect 15858 8132 15914 8188
rect 15914 8132 15918 8188
rect 15854 8128 15918 8132
rect 21479 8188 21543 8192
rect 21479 8132 21483 8188
rect 21483 8132 21539 8188
rect 21539 8132 21543 8188
rect 21479 8128 21543 8132
rect 21559 8188 21623 8192
rect 21559 8132 21563 8188
rect 21563 8132 21619 8188
rect 21619 8132 21623 8188
rect 21559 8128 21623 8132
rect 21639 8188 21703 8192
rect 21639 8132 21643 8188
rect 21643 8132 21699 8188
rect 21699 8132 21703 8188
rect 21639 8128 21703 8132
rect 21719 8188 21783 8192
rect 21719 8132 21723 8188
rect 21723 8132 21779 8188
rect 21779 8132 21783 8188
rect 21719 8128 21783 8132
rect 3372 7788 3436 7852
rect 6816 7644 6880 7648
rect 6816 7588 6820 7644
rect 6820 7588 6876 7644
rect 6876 7588 6880 7644
rect 6816 7584 6880 7588
rect 6896 7644 6960 7648
rect 6896 7588 6900 7644
rect 6900 7588 6956 7644
rect 6956 7588 6960 7644
rect 6896 7584 6960 7588
rect 6976 7644 7040 7648
rect 6976 7588 6980 7644
rect 6980 7588 7036 7644
rect 7036 7588 7040 7644
rect 6976 7584 7040 7588
rect 7056 7644 7120 7648
rect 7056 7588 7060 7644
rect 7060 7588 7116 7644
rect 7116 7588 7120 7644
rect 7056 7584 7120 7588
rect 12681 7644 12745 7648
rect 12681 7588 12685 7644
rect 12685 7588 12741 7644
rect 12741 7588 12745 7644
rect 12681 7584 12745 7588
rect 12761 7644 12825 7648
rect 12761 7588 12765 7644
rect 12765 7588 12821 7644
rect 12821 7588 12825 7644
rect 12761 7584 12825 7588
rect 12841 7644 12905 7648
rect 12841 7588 12845 7644
rect 12845 7588 12901 7644
rect 12901 7588 12905 7644
rect 12841 7584 12905 7588
rect 12921 7644 12985 7648
rect 12921 7588 12925 7644
rect 12925 7588 12981 7644
rect 12981 7588 12985 7644
rect 12921 7584 12985 7588
rect 18546 7644 18610 7648
rect 18546 7588 18550 7644
rect 18550 7588 18606 7644
rect 18606 7588 18610 7644
rect 18546 7584 18610 7588
rect 18626 7644 18690 7648
rect 18626 7588 18630 7644
rect 18630 7588 18686 7644
rect 18686 7588 18690 7644
rect 18626 7584 18690 7588
rect 18706 7644 18770 7648
rect 18706 7588 18710 7644
rect 18710 7588 18766 7644
rect 18766 7588 18770 7644
rect 18706 7584 18770 7588
rect 18786 7644 18850 7648
rect 18786 7588 18790 7644
rect 18790 7588 18846 7644
rect 18846 7588 18850 7644
rect 18786 7584 18850 7588
rect 24411 7644 24475 7648
rect 24411 7588 24415 7644
rect 24415 7588 24471 7644
rect 24471 7588 24475 7644
rect 24411 7584 24475 7588
rect 24491 7644 24555 7648
rect 24491 7588 24495 7644
rect 24495 7588 24551 7644
rect 24551 7588 24555 7644
rect 24491 7584 24555 7588
rect 24571 7644 24635 7648
rect 24571 7588 24575 7644
rect 24575 7588 24631 7644
rect 24631 7588 24635 7644
rect 24571 7584 24635 7588
rect 24651 7644 24715 7648
rect 24651 7588 24655 7644
rect 24655 7588 24711 7644
rect 24711 7588 24715 7644
rect 24651 7584 24715 7588
rect 3884 7100 3948 7104
rect 3884 7044 3888 7100
rect 3888 7044 3944 7100
rect 3944 7044 3948 7100
rect 3884 7040 3948 7044
rect 3964 7100 4028 7104
rect 3964 7044 3968 7100
rect 3968 7044 4024 7100
rect 4024 7044 4028 7100
rect 3964 7040 4028 7044
rect 4044 7100 4108 7104
rect 4044 7044 4048 7100
rect 4048 7044 4104 7100
rect 4104 7044 4108 7100
rect 4044 7040 4108 7044
rect 4124 7100 4188 7104
rect 4124 7044 4128 7100
rect 4128 7044 4184 7100
rect 4184 7044 4188 7100
rect 4124 7040 4188 7044
rect 9749 7100 9813 7104
rect 9749 7044 9753 7100
rect 9753 7044 9809 7100
rect 9809 7044 9813 7100
rect 9749 7040 9813 7044
rect 9829 7100 9893 7104
rect 9829 7044 9833 7100
rect 9833 7044 9889 7100
rect 9889 7044 9893 7100
rect 9829 7040 9893 7044
rect 9909 7100 9973 7104
rect 9909 7044 9913 7100
rect 9913 7044 9969 7100
rect 9969 7044 9973 7100
rect 9909 7040 9973 7044
rect 9989 7100 10053 7104
rect 9989 7044 9993 7100
rect 9993 7044 10049 7100
rect 10049 7044 10053 7100
rect 9989 7040 10053 7044
rect 15614 7100 15678 7104
rect 15614 7044 15618 7100
rect 15618 7044 15674 7100
rect 15674 7044 15678 7100
rect 15614 7040 15678 7044
rect 15694 7100 15758 7104
rect 15694 7044 15698 7100
rect 15698 7044 15754 7100
rect 15754 7044 15758 7100
rect 15694 7040 15758 7044
rect 15774 7100 15838 7104
rect 15774 7044 15778 7100
rect 15778 7044 15834 7100
rect 15834 7044 15838 7100
rect 15774 7040 15838 7044
rect 15854 7100 15918 7104
rect 15854 7044 15858 7100
rect 15858 7044 15914 7100
rect 15914 7044 15918 7100
rect 15854 7040 15918 7044
rect 21479 7100 21543 7104
rect 21479 7044 21483 7100
rect 21483 7044 21539 7100
rect 21539 7044 21543 7100
rect 21479 7040 21543 7044
rect 21559 7100 21623 7104
rect 21559 7044 21563 7100
rect 21563 7044 21619 7100
rect 21619 7044 21623 7100
rect 21559 7040 21623 7044
rect 21639 7100 21703 7104
rect 21639 7044 21643 7100
rect 21643 7044 21699 7100
rect 21699 7044 21703 7100
rect 21639 7040 21703 7044
rect 21719 7100 21783 7104
rect 21719 7044 21723 7100
rect 21723 7044 21779 7100
rect 21779 7044 21783 7100
rect 21719 7040 21783 7044
rect 6816 6556 6880 6560
rect 6816 6500 6820 6556
rect 6820 6500 6876 6556
rect 6876 6500 6880 6556
rect 6816 6496 6880 6500
rect 6896 6556 6960 6560
rect 6896 6500 6900 6556
rect 6900 6500 6956 6556
rect 6956 6500 6960 6556
rect 6896 6496 6960 6500
rect 6976 6556 7040 6560
rect 6976 6500 6980 6556
rect 6980 6500 7036 6556
rect 7036 6500 7040 6556
rect 6976 6496 7040 6500
rect 7056 6556 7120 6560
rect 7056 6500 7060 6556
rect 7060 6500 7116 6556
rect 7116 6500 7120 6556
rect 7056 6496 7120 6500
rect 12681 6556 12745 6560
rect 12681 6500 12685 6556
rect 12685 6500 12741 6556
rect 12741 6500 12745 6556
rect 12681 6496 12745 6500
rect 12761 6556 12825 6560
rect 12761 6500 12765 6556
rect 12765 6500 12821 6556
rect 12821 6500 12825 6556
rect 12761 6496 12825 6500
rect 12841 6556 12905 6560
rect 12841 6500 12845 6556
rect 12845 6500 12901 6556
rect 12901 6500 12905 6556
rect 12841 6496 12905 6500
rect 12921 6556 12985 6560
rect 12921 6500 12925 6556
rect 12925 6500 12981 6556
rect 12981 6500 12985 6556
rect 12921 6496 12985 6500
rect 18546 6556 18610 6560
rect 18546 6500 18550 6556
rect 18550 6500 18606 6556
rect 18606 6500 18610 6556
rect 18546 6496 18610 6500
rect 18626 6556 18690 6560
rect 18626 6500 18630 6556
rect 18630 6500 18686 6556
rect 18686 6500 18690 6556
rect 18626 6496 18690 6500
rect 18706 6556 18770 6560
rect 18706 6500 18710 6556
rect 18710 6500 18766 6556
rect 18766 6500 18770 6556
rect 18706 6496 18770 6500
rect 18786 6556 18850 6560
rect 18786 6500 18790 6556
rect 18790 6500 18846 6556
rect 18846 6500 18850 6556
rect 18786 6496 18850 6500
rect 2268 6428 2332 6492
rect 24411 6556 24475 6560
rect 24411 6500 24415 6556
rect 24415 6500 24471 6556
rect 24471 6500 24475 6556
rect 24411 6496 24475 6500
rect 24491 6556 24555 6560
rect 24491 6500 24495 6556
rect 24495 6500 24551 6556
rect 24551 6500 24555 6556
rect 24491 6496 24555 6500
rect 24571 6556 24635 6560
rect 24571 6500 24575 6556
rect 24575 6500 24631 6556
rect 24631 6500 24635 6556
rect 24571 6496 24635 6500
rect 24651 6556 24715 6560
rect 24651 6500 24655 6556
rect 24655 6500 24711 6556
rect 24711 6500 24715 6556
rect 24651 6496 24715 6500
rect 3884 6012 3948 6016
rect 3884 5956 3888 6012
rect 3888 5956 3944 6012
rect 3944 5956 3948 6012
rect 3884 5952 3948 5956
rect 3964 6012 4028 6016
rect 3964 5956 3968 6012
rect 3968 5956 4024 6012
rect 4024 5956 4028 6012
rect 3964 5952 4028 5956
rect 4044 6012 4108 6016
rect 4044 5956 4048 6012
rect 4048 5956 4104 6012
rect 4104 5956 4108 6012
rect 4044 5952 4108 5956
rect 4124 6012 4188 6016
rect 4124 5956 4128 6012
rect 4128 5956 4184 6012
rect 4184 5956 4188 6012
rect 4124 5952 4188 5956
rect 9749 6012 9813 6016
rect 9749 5956 9753 6012
rect 9753 5956 9809 6012
rect 9809 5956 9813 6012
rect 9749 5952 9813 5956
rect 9829 6012 9893 6016
rect 9829 5956 9833 6012
rect 9833 5956 9889 6012
rect 9889 5956 9893 6012
rect 9829 5952 9893 5956
rect 9909 6012 9973 6016
rect 9909 5956 9913 6012
rect 9913 5956 9969 6012
rect 9969 5956 9973 6012
rect 9909 5952 9973 5956
rect 9989 6012 10053 6016
rect 9989 5956 9993 6012
rect 9993 5956 10049 6012
rect 10049 5956 10053 6012
rect 9989 5952 10053 5956
rect 15614 6012 15678 6016
rect 15614 5956 15618 6012
rect 15618 5956 15674 6012
rect 15674 5956 15678 6012
rect 15614 5952 15678 5956
rect 15694 6012 15758 6016
rect 15694 5956 15698 6012
rect 15698 5956 15754 6012
rect 15754 5956 15758 6012
rect 15694 5952 15758 5956
rect 15774 6012 15838 6016
rect 15774 5956 15778 6012
rect 15778 5956 15834 6012
rect 15834 5956 15838 6012
rect 15774 5952 15838 5956
rect 15854 6012 15918 6016
rect 15854 5956 15858 6012
rect 15858 5956 15914 6012
rect 15914 5956 15918 6012
rect 15854 5952 15918 5956
rect 21479 6012 21543 6016
rect 21479 5956 21483 6012
rect 21483 5956 21539 6012
rect 21539 5956 21543 6012
rect 21479 5952 21543 5956
rect 21559 6012 21623 6016
rect 21559 5956 21563 6012
rect 21563 5956 21619 6012
rect 21619 5956 21623 6012
rect 21559 5952 21623 5956
rect 21639 6012 21703 6016
rect 21639 5956 21643 6012
rect 21643 5956 21699 6012
rect 21699 5956 21703 6012
rect 21639 5952 21703 5956
rect 21719 6012 21783 6016
rect 21719 5956 21723 6012
rect 21723 5956 21779 6012
rect 21779 5956 21783 6012
rect 21719 5952 21783 5956
rect 3740 5612 3804 5676
rect 1900 5476 1964 5540
rect 11652 5536 11716 5540
rect 11652 5480 11666 5536
rect 11666 5480 11716 5536
rect 11652 5476 11716 5480
rect 18276 5476 18340 5540
rect 6816 5468 6880 5472
rect 6816 5412 6820 5468
rect 6820 5412 6876 5468
rect 6876 5412 6880 5468
rect 6816 5408 6880 5412
rect 6896 5468 6960 5472
rect 6896 5412 6900 5468
rect 6900 5412 6956 5468
rect 6956 5412 6960 5468
rect 6896 5408 6960 5412
rect 6976 5468 7040 5472
rect 6976 5412 6980 5468
rect 6980 5412 7036 5468
rect 7036 5412 7040 5468
rect 6976 5408 7040 5412
rect 7056 5468 7120 5472
rect 7056 5412 7060 5468
rect 7060 5412 7116 5468
rect 7116 5412 7120 5468
rect 7056 5408 7120 5412
rect 12681 5468 12745 5472
rect 12681 5412 12685 5468
rect 12685 5412 12741 5468
rect 12741 5412 12745 5468
rect 12681 5408 12745 5412
rect 12761 5468 12825 5472
rect 12761 5412 12765 5468
rect 12765 5412 12821 5468
rect 12821 5412 12825 5468
rect 12761 5408 12825 5412
rect 12841 5468 12905 5472
rect 12841 5412 12845 5468
rect 12845 5412 12901 5468
rect 12901 5412 12905 5468
rect 12841 5408 12905 5412
rect 12921 5468 12985 5472
rect 12921 5412 12925 5468
rect 12925 5412 12981 5468
rect 12981 5412 12985 5468
rect 12921 5408 12985 5412
rect 18546 5468 18610 5472
rect 18546 5412 18550 5468
rect 18550 5412 18606 5468
rect 18606 5412 18610 5468
rect 18546 5408 18610 5412
rect 18626 5468 18690 5472
rect 18626 5412 18630 5468
rect 18630 5412 18686 5468
rect 18686 5412 18690 5468
rect 18626 5408 18690 5412
rect 18706 5468 18770 5472
rect 18706 5412 18710 5468
rect 18710 5412 18766 5468
rect 18766 5412 18770 5468
rect 18706 5408 18770 5412
rect 18786 5468 18850 5472
rect 18786 5412 18790 5468
rect 18790 5412 18846 5468
rect 18846 5412 18850 5468
rect 18786 5408 18850 5412
rect 22324 5340 22388 5404
rect 16620 5068 16684 5132
rect 3884 4924 3948 4928
rect 3884 4868 3888 4924
rect 3888 4868 3944 4924
rect 3944 4868 3948 4924
rect 3884 4864 3948 4868
rect 3964 4924 4028 4928
rect 3964 4868 3968 4924
rect 3968 4868 4024 4924
rect 4024 4868 4028 4924
rect 3964 4864 4028 4868
rect 4044 4924 4108 4928
rect 4044 4868 4048 4924
rect 4048 4868 4104 4924
rect 4104 4868 4108 4924
rect 4044 4864 4108 4868
rect 4124 4924 4188 4928
rect 4124 4868 4128 4924
rect 4128 4868 4184 4924
rect 4184 4868 4188 4924
rect 4124 4864 4188 4868
rect 9749 4924 9813 4928
rect 9749 4868 9753 4924
rect 9753 4868 9809 4924
rect 9809 4868 9813 4924
rect 9749 4864 9813 4868
rect 9829 4924 9893 4928
rect 9829 4868 9833 4924
rect 9833 4868 9889 4924
rect 9889 4868 9893 4924
rect 9829 4864 9893 4868
rect 9909 4924 9973 4928
rect 9909 4868 9913 4924
rect 9913 4868 9969 4924
rect 9969 4868 9973 4924
rect 9909 4864 9973 4868
rect 9989 4924 10053 4928
rect 9989 4868 9993 4924
rect 9993 4868 10049 4924
rect 10049 4868 10053 4924
rect 9989 4864 10053 4868
rect 15614 4924 15678 4928
rect 15614 4868 15618 4924
rect 15618 4868 15674 4924
rect 15674 4868 15678 4924
rect 15614 4864 15678 4868
rect 15694 4924 15758 4928
rect 15694 4868 15698 4924
rect 15698 4868 15754 4924
rect 15754 4868 15758 4924
rect 15694 4864 15758 4868
rect 15774 4924 15838 4928
rect 15774 4868 15778 4924
rect 15778 4868 15834 4924
rect 15834 4868 15838 4924
rect 15774 4864 15838 4868
rect 15854 4924 15918 4928
rect 15854 4868 15858 4924
rect 15858 4868 15914 4924
rect 15914 4868 15918 4924
rect 15854 4864 15918 4868
rect 21479 4924 21543 4928
rect 21479 4868 21483 4924
rect 21483 4868 21539 4924
rect 21539 4868 21543 4924
rect 21479 4864 21543 4868
rect 21559 4924 21623 4928
rect 21559 4868 21563 4924
rect 21563 4868 21619 4924
rect 21619 4868 21623 4924
rect 21559 4864 21623 4868
rect 21639 4924 21703 4928
rect 21639 4868 21643 4924
rect 21643 4868 21699 4924
rect 21699 4868 21703 4924
rect 21639 4864 21703 4868
rect 21719 4924 21783 4928
rect 21719 4868 21723 4924
rect 21723 4868 21779 4924
rect 21779 4868 21783 4924
rect 21719 4864 21783 4868
rect 1716 4720 1780 4724
rect 1716 4664 1730 4720
rect 1730 4664 1780 4720
rect 1716 4660 1780 4664
rect 21956 4660 22020 4724
rect 24411 5468 24475 5472
rect 24411 5412 24415 5468
rect 24415 5412 24471 5468
rect 24471 5412 24475 5468
rect 24411 5408 24475 5412
rect 24491 5468 24555 5472
rect 24491 5412 24495 5468
rect 24495 5412 24551 5468
rect 24551 5412 24555 5468
rect 24491 5408 24555 5412
rect 24571 5468 24635 5472
rect 24571 5412 24575 5468
rect 24575 5412 24631 5468
rect 24631 5412 24635 5468
rect 24571 5408 24635 5412
rect 24651 5468 24715 5472
rect 24651 5412 24655 5468
rect 24655 5412 24711 5468
rect 24711 5412 24715 5468
rect 24651 5408 24715 5412
rect 6816 4380 6880 4384
rect 6816 4324 6820 4380
rect 6820 4324 6876 4380
rect 6876 4324 6880 4380
rect 6816 4320 6880 4324
rect 6896 4380 6960 4384
rect 6896 4324 6900 4380
rect 6900 4324 6956 4380
rect 6956 4324 6960 4380
rect 6896 4320 6960 4324
rect 6976 4380 7040 4384
rect 6976 4324 6980 4380
rect 6980 4324 7036 4380
rect 7036 4324 7040 4380
rect 6976 4320 7040 4324
rect 7056 4380 7120 4384
rect 7056 4324 7060 4380
rect 7060 4324 7116 4380
rect 7116 4324 7120 4380
rect 7056 4320 7120 4324
rect 12681 4380 12745 4384
rect 12681 4324 12685 4380
rect 12685 4324 12741 4380
rect 12741 4324 12745 4380
rect 12681 4320 12745 4324
rect 12761 4380 12825 4384
rect 12761 4324 12765 4380
rect 12765 4324 12821 4380
rect 12821 4324 12825 4380
rect 12761 4320 12825 4324
rect 12841 4380 12905 4384
rect 12841 4324 12845 4380
rect 12845 4324 12901 4380
rect 12901 4324 12905 4380
rect 12841 4320 12905 4324
rect 12921 4380 12985 4384
rect 12921 4324 12925 4380
rect 12925 4324 12981 4380
rect 12981 4324 12985 4380
rect 12921 4320 12985 4324
rect 18546 4380 18610 4384
rect 18546 4324 18550 4380
rect 18550 4324 18606 4380
rect 18606 4324 18610 4380
rect 18546 4320 18610 4324
rect 18626 4380 18690 4384
rect 18626 4324 18630 4380
rect 18630 4324 18686 4380
rect 18686 4324 18690 4380
rect 18626 4320 18690 4324
rect 18706 4380 18770 4384
rect 18706 4324 18710 4380
rect 18710 4324 18766 4380
rect 18766 4324 18770 4380
rect 18706 4320 18770 4324
rect 18786 4380 18850 4384
rect 18786 4324 18790 4380
rect 18790 4324 18846 4380
rect 18846 4324 18850 4380
rect 18786 4320 18850 4324
rect 24411 4380 24475 4384
rect 24411 4324 24415 4380
rect 24415 4324 24471 4380
rect 24471 4324 24475 4380
rect 24411 4320 24475 4324
rect 24491 4380 24555 4384
rect 24491 4324 24495 4380
rect 24495 4324 24551 4380
rect 24551 4324 24555 4380
rect 24491 4320 24555 4324
rect 24571 4380 24635 4384
rect 24571 4324 24575 4380
rect 24575 4324 24631 4380
rect 24631 4324 24635 4380
rect 24571 4320 24635 4324
rect 24651 4380 24715 4384
rect 24651 4324 24655 4380
rect 24655 4324 24711 4380
rect 24711 4324 24715 4380
rect 24651 4320 24715 4324
rect 2820 3980 2884 4044
rect 3740 4116 3804 4180
rect 10916 4040 10980 4044
rect 10916 3984 10930 4040
rect 10930 3984 10980 4040
rect 10916 3980 10980 3984
rect 20116 3980 20180 4044
rect 2084 3844 2148 3908
rect 3884 3836 3948 3840
rect 3884 3780 3888 3836
rect 3888 3780 3944 3836
rect 3944 3780 3948 3836
rect 3884 3776 3948 3780
rect 3964 3836 4028 3840
rect 3964 3780 3968 3836
rect 3968 3780 4024 3836
rect 4024 3780 4028 3836
rect 3964 3776 4028 3780
rect 4044 3836 4108 3840
rect 4044 3780 4048 3836
rect 4048 3780 4104 3836
rect 4104 3780 4108 3836
rect 4044 3776 4108 3780
rect 4124 3836 4188 3840
rect 4124 3780 4128 3836
rect 4128 3780 4184 3836
rect 4184 3780 4188 3836
rect 4124 3776 4188 3780
rect 9749 3836 9813 3840
rect 9749 3780 9753 3836
rect 9753 3780 9809 3836
rect 9809 3780 9813 3836
rect 9749 3776 9813 3780
rect 9829 3836 9893 3840
rect 9829 3780 9833 3836
rect 9833 3780 9889 3836
rect 9889 3780 9893 3836
rect 9829 3776 9893 3780
rect 9909 3836 9973 3840
rect 9909 3780 9913 3836
rect 9913 3780 9969 3836
rect 9969 3780 9973 3836
rect 9909 3776 9973 3780
rect 9989 3836 10053 3840
rect 9989 3780 9993 3836
rect 9993 3780 10049 3836
rect 10049 3780 10053 3836
rect 9989 3776 10053 3780
rect 15614 3836 15678 3840
rect 15614 3780 15618 3836
rect 15618 3780 15674 3836
rect 15674 3780 15678 3836
rect 15614 3776 15678 3780
rect 15694 3836 15758 3840
rect 15694 3780 15698 3836
rect 15698 3780 15754 3836
rect 15754 3780 15758 3836
rect 15694 3776 15758 3780
rect 15774 3836 15838 3840
rect 15774 3780 15778 3836
rect 15778 3780 15834 3836
rect 15834 3780 15838 3836
rect 15774 3776 15838 3780
rect 15854 3836 15918 3840
rect 15854 3780 15858 3836
rect 15858 3780 15914 3836
rect 15914 3780 15918 3836
rect 15854 3776 15918 3780
rect 21479 3836 21543 3840
rect 21479 3780 21483 3836
rect 21483 3780 21539 3836
rect 21539 3780 21543 3836
rect 21479 3776 21543 3780
rect 21559 3836 21623 3840
rect 21559 3780 21563 3836
rect 21563 3780 21619 3836
rect 21619 3780 21623 3836
rect 21559 3776 21623 3780
rect 21639 3836 21703 3840
rect 21639 3780 21643 3836
rect 21643 3780 21699 3836
rect 21699 3780 21703 3836
rect 21639 3776 21703 3780
rect 21719 3836 21783 3840
rect 21719 3780 21723 3836
rect 21723 3780 21779 3836
rect 21779 3780 21783 3836
rect 21719 3776 21783 3780
rect 20852 3300 20916 3364
rect 6816 3292 6880 3296
rect 6816 3236 6820 3292
rect 6820 3236 6876 3292
rect 6876 3236 6880 3292
rect 6816 3232 6880 3236
rect 6896 3292 6960 3296
rect 6896 3236 6900 3292
rect 6900 3236 6956 3292
rect 6956 3236 6960 3292
rect 6896 3232 6960 3236
rect 6976 3292 7040 3296
rect 6976 3236 6980 3292
rect 6980 3236 7036 3292
rect 7036 3236 7040 3292
rect 6976 3232 7040 3236
rect 7056 3292 7120 3296
rect 7056 3236 7060 3292
rect 7060 3236 7116 3292
rect 7116 3236 7120 3292
rect 7056 3232 7120 3236
rect 12681 3292 12745 3296
rect 12681 3236 12685 3292
rect 12685 3236 12741 3292
rect 12741 3236 12745 3292
rect 12681 3232 12745 3236
rect 12761 3292 12825 3296
rect 12761 3236 12765 3292
rect 12765 3236 12821 3292
rect 12821 3236 12825 3292
rect 12761 3232 12825 3236
rect 12841 3292 12905 3296
rect 12841 3236 12845 3292
rect 12845 3236 12901 3292
rect 12901 3236 12905 3292
rect 12841 3232 12905 3236
rect 12921 3292 12985 3296
rect 12921 3236 12925 3292
rect 12925 3236 12981 3292
rect 12981 3236 12985 3292
rect 12921 3232 12985 3236
rect 18546 3292 18610 3296
rect 18546 3236 18550 3292
rect 18550 3236 18606 3292
rect 18606 3236 18610 3292
rect 18546 3232 18610 3236
rect 18626 3292 18690 3296
rect 18626 3236 18630 3292
rect 18630 3236 18686 3292
rect 18686 3236 18690 3292
rect 18626 3232 18690 3236
rect 18706 3292 18770 3296
rect 18706 3236 18710 3292
rect 18710 3236 18766 3292
rect 18766 3236 18770 3292
rect 18706 3232 18770 3236
rect 18786 3292 18850 3296
rect 18786 3236 18790 3292
rect 18790 3236 18846 3292
rect 18846 3236 18850 3292
rect 18786 3232 18850 3236
rect 24411 3292 24475 3296
rect 24411 3236 24415 3292
rect 24415 3236 24471 3292
rect 24471 3236 24475 3292
rect 24411 3232 24475 3236
rect 24491 3292 24555 3296
rect 24491 3236 24495 3292
rect 24495 3236 24551 3292
rect 24551 3236 24555 3292
rect 24491 3232 24555 3236
rect 24571 3292 24635 3296
rect 24571 3236 24575 3292
rect 24575 3236 24631 3292
rect 24631 3236 24635 3292
rect 24571 3232 24635 3236
rect 24651 3292 24715 3296
rect 24651 3236 24655 3292
rect 24655 3236 24711 3292
rect 24711 3236 24715 3292
rect 24651 3232 24715 3236
rect 12388 3028 12452 3092
rect 13124 3028 13188 3092
rect 3884 2748 3948 2752
rect 3884 2692 3888 2748
rect 3888 2692 3944 2748
rect 3944 2692 3948 2748
rect 3884 2688 3948 2692
rect 3964 2748 4028 2752
rect 3964 2692 3968 2748
rect 3968 2692 4024 2748
rect 4024 2692 4028 2748
rect 3964 2688 4028 2692
rect 4044 2748 4108 2752
rect 4044 2692 4048 2748
rect 4048 2692 4104 2748
rect 4104 2692 4108 2748
rect 4044 2688 4108 2692
rect 4124 2748 4188 2752
rect 4124 2692 4128 2748
rect 4128 2692 4184 2748
rect 4184 2692 4188 2748
rect 4124 2688 4188 2692
rect 5396 2680 5460 2684
rect 5396 2624 5410 2680
rect 5410 2624 5460 2680
rect 5396 2620 5460 2624
rect 9749 2748 9813 2752
rect 9749 2692 9753 2748
rect 9753 2692 9809 2748
rect 9809 2692 9813 2748
rect 9749 2688 9813 2692
rect 9829 2748 9893 2752
rect 9829 2692 9833 2748
rect 9833 2692 9889 2748
rect 9889 2692 9893 2748
rect 9829 2688 9893 2692
rect 9909 2748 9973 2752
rect 9909 2692 9913 2748
rect 9913 2692 9969 2748
rect 9969 2692 9973 2748
rect 9909 2688 9973 2692
rect 9989 2748 10053 2752
rect 9989 2692 9993 2748
rect 9993 2692 10049 2748
rect 10049 2692 10053 2748
rect 9989 2688 10053 2692
rect 15614 2748 15678 2752
rect 15614 2692 15618 2748
rect 15618 2692 15674 2748
rect 15674 2692 15678 2748
rect 15614 2688 15678 2692
rect 15694 2748 15758 2752
rect 15694 2692 15698 2748
rect 15698 2692 15754 2748
rect 15754 2692 15758 2748
rect 15694 2688 15758 2692
rect 15774 2748 15838 2752
rect 15774 2692 15778 2748
rect 15778 2692 15834 2748
rect 15834 2692 15838 2748
rect 15774 2688 15838 2692
rect 15854 2748 15918 2752
rect 15854 2692 15858 2748
rect 15858 2692 15914 2748
rect 15914 2692 15918 2748
rect 15854 2688 15918 2692
rect 21479 2748 21543 2752
rect 21479 2692 21483 2748
rect 21483 2692 21539 2748
rect 21539 2692 21543 2748
rect 21479 2688 21543 2692
rect 21559 2748 21623 2752
rect 21559 2692 21563 2748
rect 21563 2692 21619 2748
rect 21619 2692 21623 2748
rect 21559 2688 21623 2692
rect 21639 2748 21703 2752
rect 21639 2692 21643 2748
rect 21643 2692 21699 2748
rect 21699 2692 21703 2748
rect 21639 2688 21703 2692
rect 21719 2748 21783 2752
rect 21719 2692 21723 2748
rect 21723 2692 21779 2748
rect 21779 2692 21783 2748
rect 21719 2688 21783 2692
rect 612 2484 676 2548
rect 13308 2620 13372 2684
rect 16988 2620 17052 2684
rect 17172 2680 17236 2684
rect 17172 2624 17186 2680
rect 17186 2624 17236 2680
rect 17172 2620 17236 2624
rect 19564 2680 19628 2684
rect 19564 2624 19614 2680
rect 19614 2624 19628 2680
rect 19564 2620 19628 2624
rect 22140 2680 22204 2684
rect 22140 2624 22190 2680
rect 22190 2624 22204 2680
rect 22140 2620 22204 2624
rect 10364 2484 10428 2548
rect 15332 2484 15396 2548
rect 7420 2212 7484 2276
rect 6816 2204 6880 2208
rect 6816 2148 6820 2204
rect 6820 2148 6876 2204
rect 6876 2148 6880 2204
rect 6816 2144 6880 2148
rect 6896 2204 6960 2208
rect 6896 2148 6900 2204
rect 6900 2148 6956 2204
rect 6956 2148 6960 2204
rect 6896 2144 6960 2148
rect 6976 2204 7040 2208
rect 6976 2148 6980 2204
rect 6980 2148 7036 2204
rect 7036 2148 7040 2204
rect 6976 2144 7040 2148
rect 7056 2204 7120 2208
rect 7056 2148 7060 2204
rect 7060 2148 7116 2204
rect 7116 2148 7120 2204
rect 7056 2144 7120 2148
rect 12020 2348 12084 2412
rect 8156 2272 8220 2276
rect 8156 2216 8170 2272
rect 8170 2216 8220 2272
rect 8156 2212 8220 2216
rect 8892 2272 8956 2276
rect 8892 2216 8906 2272
rect 8906 2216 8956 2272
rect 8892 2212 8956 2216
rect 21220 2348 21284 2412
rect 12681 2204 12745 2208
rect 12681 2148 12685 2204
rect 12685 2148 12741 2204
rect 12741 2148 12745 2204
rect 12681 2144 12745 2148
rect 12761 2204 12825 2208
rect 12761 2148 12765 2204
rect 12765 2148 12821 2204
rect 12821 2148 12825 2204
rect 12761 2144 12825 2148
rect 12841 2204 12905 2208
rect 12841 2148 12845 2204
rect 12845 2148 12901 2204
rect 12901 2148 12905 2204
rect 12841 2144 12905 2148
rect 12921 2204 12985 2208
rect 12921 2148 12925 2204
rect 12925 2148 12981 2204
rect 12981 2148 12985 2204
rect 12921 2144 12985 2148
rect 18546 2204 18610 2208
rect 18546 2148 18550 2204
rect 18550 2148 18606 2204
rect 18606 2148 18610 2204
rect 18546 2144 18610 2148
rect 18626 2204 18690 2208
rect 18626 2148 18630 2204
rect 18630 2148 18686 2204
rect 18686 2148 18690 2204
rect 18626 2144 18690 2148
rect 18706 2204 18770 2208
rect 18706 2148 18710 2204
rect 18710 2148 18766 2204
rect 18766 2148 18770 2204
rect 18706 2144 18770 2148
rect 18786 2204 18850 2208
rect 18786 2148 18790 2204
rect 18790 2148 18846 2204
rect 18846 2148 18850 2204
rect 18786 2144 18850 2148
rect 24411 2204 24475 2208
rect 24411 2148 24415 2204
rect 24415 2148 24471 2204
rect 24471 2148 24475 2204
rect 24411 2144 24475 2148
rect 24491 2204 24555 2208
rect 24491 2148 24495 2204
rect 24495 2148 24551 2204
rect 24551 2148 24555 2204
rect 24491 2144 24555 2148
rect 24571 2204 24635 2208
rect 24571 2148 24575 2204
rect 24575 2148 24631 2204
rect 24631 2148 24635 2204
rect 24571 2144 24635 2148
rect 24651 2204 24715 2208
rect 24651 2148 24655 2204
rect 24655 2148 24711 2204
rect 24711 2148 24715 2204
rect 24651 2144 24715 2148
rect 14412 2136 14476 2140
rect 14412 2080 14462 2136
rect 14462 2080 14476 2136
rect 14412 2076 14476 2080
rect 980 1940 1044 2004
rect 22508 1940 22572 2004
rect 1164 1804 1228 1868
rect 3884 1660 3948 1664
rect 3884 1604 3888 1660
rect 3888 1604 3944 1660
rect 3944 1604 3948 1660
rect 3884 1600 3948 1604
rect 3964 1660 4028 1664
rect 3964 1604 3968 1660
rect 3968 1604 4024 1660
rect 4024 1604 4028 1660
rect 3964 1600 4028 1604
rect 4044 1660 4108 1664
rect 4044 1604 4048 1660
rect 4048 1604 4104 1660
rect 4104 1604 4108 1660
rect 4044 1600 4108 1604
rect 4124 1660 4188 1664
rect 4124 1604 4128 1660
rect 4128 1604 4184 1660
rect 4184 1604 4188 1660
rect 4124 1600 4188 1604
rect 9749 1660 9813 1664
rect 9749 1604 9753 1660
rect 9753 1604 9809 1660
rect 9809 1604 9813 1660
rect 9749 1600 9813 1604
rect 9829 1660 9893 1664
rect 9829 1604 9833 1660
rect 9833 1604 9889 1660
rect 9889 1604 9893 1660
rect 9829 1600 9893 1604
rect 9909 1660 9973 1664
rect 9909 1604 9913 1660
rect 9913 1604 9969 1660
rect 9969 1604 9973 1660
rect 9909 1600 9973 1604
rect 9989 1660 10053 1664
rect 9989 1604 9993 1660
rect 9993 1604 10049 1660
rect 10049 1604 10053 1660
rect 9989 1600 10053 1604
rect 15614 1660 15678 1664
rect 15614 1604 15618 1660
rect 15618 1604 15674 1660
rect 15674 1604 15678 1660
rect 15614 1600 15678 1604
rect 15694 1660 15758 1664
rect 15694 1604 15698 1660
rect 15698 1604 15754 1660
rect 15754 1604 15758 1660
rect 15694 1600 15758 1604
rect 15774 1660 15838 1664
rect 15774 1604 15778 1660
rect 15778 1604 15834 1660
rect 15834 1604 15838 1660
rect 15774 1600 15838 1604
rect 15854 1660 15918 1664
rect 15854 1604 15858 1660
rect 15858 1604 15914 1660
rect 15914 1604 15918 1660
rect 15854 1600 15918 1604
rect 21479 1660 21543 1664
rect 21479 1604 21483 1660
rect 21483 1604 21539 1660
rect 21539 1604 21543 1660
rect 21479 1600 21543 1604
rect 21559 1660 21623 1664
rect 21559 1604 21563 1660
rect 21563 1604 21619 1660
rect 21619 1604 21623 1660
rect 21559 1600 21623 1604
rect 21639 1660 21703 1664
rect 21639 1604 21643 1660
rect 21643 1604 21699 1660
rect 21699 1604 21703 1660
rect 21639 1600 21703 1604
rect 21719 1660 21783 1664
rect 21719 1604 21723 1660
rect 21723 1604 21779 1660
rect 21779 1604 21783 1660
rect 21719 1600 21783 1604
rect 3740 1456 3804 1460
rect 3740 1400 3790 1456
rect 3790 1400 3804 1456
rect 3740 1396 3804 1400
rect 4476 1320 4540 1324
rect 4476 1264 4490 1320
rect 4490 1264 4540 1320
rect 4476 1260 4540 1264
rect 8708 1260 8772 1324
rect 11100 1320 11164 1324
rect 11100 1264 11114 1320
rect 11114 1264 11164 1320
rect 11100 1260 11164 1264
rect 12388 1260 12452 1324
rect 13492 1320 13556 1324
rect 13492 1264 13506 1320
rect 13506 1264 13556 1320
rect 13492 1260 13556 1264
rect 14228 1260 14292 1324
rect 14596 1320 14660 1324
rect 14596 1264 14610 1320
rect 14610 1264 14660 1320
rect 14596 1260 14660 1264
rect 15148 1320 15212 1324
rect 15148 1264 15198 1320
rect 15198 1264 15212 1320
rect 15148 1260 15212 1264
rect 6132 1124 6196 1188
rect 8340 1124 8404 1188
rect 6816 1116 6880 1120
rect 6816 1060 6820 1116
rect 6820 1060 6876 1116
rect 6876 1060 6880 1116
rect 6816 1056 6880 1060
rect 6896 1116 6960 1120
rect 6896 1060 6900 1116
rect 6900 1060 6956 1116
rect 6956 1060 6960 1116
rect 6896 1056 6960 1060
rect 6976 1116 7040 1120
rect 6976 1060 6980 1116
rect 6980 1060 7036 1116
rect 7036 1060 7040 1116
rect 6976 1056 7040 1060
rect 7056 1116 7120 1120
rect 7056 1060 7060 1116
rect 7060 1060 7116 1116
rect 7116 1060 7120 1116
rect 7056 1056 7120 1060
rect 12681 1116 12745 1120
rect 12681 1060 12685 1116
rect 12685 1060 12741 1116
rect 12741 1060 12745 1116
rect 12681 1056 12745 1060
rect 12761 1116 12825 1120
rect 12761 1060 12765 1116
rect 12765 1060 12821 1116
rect 12821 1060 12825 1116
rect 12761 1056 12825 1060
rect 12841 1116 12905 1120
rect 12841 1060 12845 1116
rect 12845 1060 12901 1116
rect 12901 1060 12905 1116
rect 12841 1056 12905 1060
rect 12921 1116 12985 1120
rect 12921 1060 12925 1116
rect 12925 1060 12981 1116
rect 12981 1060 12985 1116
rect 12921 1056 12985 1060
rect 18546 1116 18610 1120
rect 18546 1060 18550 1116
rect 18550 1060 18606 1116
rect 18606 1060 18610 1116
rect 18546 1056 18610 1060
rect 18626 1116 18690 1120
rect 18626 1060 18630 1116
rect 18630 1060 18686 1116
rect 18686 1060 18690 1116
rect 18626 1056 18690 1060
rect 18706 1116 18770 1120
rect 18706 1060 18710 1116
rect 18710 1060 18766 1116
rect 18766 1060 18770 1116
rect 18706 1056 18770 1060
rect 18786 1116 18850 1120
rect 18786 1060 18790 1116
rect 18790 1060 18846 1116
rect 18846 1060 18850 1116
rect 18786 1056 18850 1060
rect 24411 1116 24475 1120
rect 24411 1060 24415 1116
rect 24415 1060 24471 1116
rect 24471 1060 24475 1116
rect 24411 1056 24475 1060
rect 24491 1116 24555 1120
rect 24491 1060 24495 1116
rect 24495 1060 24551 1116
rect 24551 1060 24555 1116
rect 24491 1056 24555 1060
rect 24571 1116 24635 1120
rect 24571 1060 24575 1116
rect 24575 1060 24631 1116
rect 24631 1060 24635 1116
rect 24571 1056 24635 1060
rect 24651 1116 24715 1120
rect 24651 1060 24655 1116
rect 24655 1060 24711 1116
rect 24711 1060 24715 1116
rect 24651 1056 24715 1060
rect 19380 852 19444 916
rect 10548 716 10612 780
rect 796 444 860 508
<< metal4 >>
rect 3876 43008 4196 43568
rect 3876 42944 3884 43008
rect 3948 42944 3964 43008
rect 4028 42944 4044 43008
rect 4108 42944 4124 43008
rect 4188 42944 4196 43008
rect 979 42804 1045 42805
rect 979 42740 980 42804
rect 1044 42740 1045 42804
rect 979 42739 1045 42740
rect 611 40084 677 40085
rect 611 40020 612 40084
rect 676 40020 677 40084
rect 611 40019 677 40020
rect 614 2549 674 40019
rect 795 38860 861 38861
rect 795 38796 796 38860
rect 860 38796 861 38860
rect 795 38795 861 38796
rect 611 2548 677 2549
rect 611 2484 612 2548
rect 676 2484 677 2548
rect 611 2483 677 2484
rect 798 509 858 38795
rect 982 2005 1042 42739
rect 3876 41920 4196 42944
rect 6808 43552 7128 43568
rect 6808 43488 6816 43552
rect 6880 43488 6896 43552
rect 6960 43488 6976 43552
rect 7040 43488 7056 43552
rect 7120 43488 7128 43552
rect 4843 42532 4909 42533
rect 4843 42468 4844 42532
rect 4908 42468 4909 42532
rect 4843 42467 4909 42468
rect 3876 41856 3884 41920
rect 3948 41856 3964 41920
rect 4028 41856 4044 41920
rect 4108 41856 4124 41920
rect 4188 41856 4196 41920
rect 3739 41580 3805 41581
rect 3739 41516 3740 41580
rect 3804 41516 3805 41580
rect 3739 41515 3805 41516
rect 1531 41444 1597 41445
rect 1531 41380 1532 41444
rect 1596 41380 1597 41444
rect 1531 41379 1597 41380
rect 2451 41444 2517 41445
rect 2451 41380 2452 41444
rect 2516 41380 2517 41444
rect 2451 41379 2517 41380
rect 1163 39676 1229 39677
rect 1163 39612 1164 39676
rect 1228 39612 1229 39676
rect 1163 39611 1229 39612
rect 979 2004 1045 2005
rect 979 1940 980 2004
rect 1044 1940 1045 2004
rect 979 1939 1045 1940
rect 1166 1869 1226 39611
rect 1534 30157 1594 41379
rect 2454 38317 2514 41379
rect 2635 40356 2701 40357
rect 2635 40292 2636 40356
rect 2700 40292 2701 40356
rect 2635 40291 2701 40292
rect 2451 38316 2517 38317
rect 2451 38252 2452 38316
rect 2516 38252 2517 38316
rect 2451 38251 2517 38252
rect 2083 32876 2149 32877
rect 2083 32812 2084 32876
rect 2148 32812 2149 32876
rect 2083 32811 2149 32812
rect 1531 30156 1597 30157
rect 1531 30092 1532 30156
rect 1596 30092 1597 30156
rect 1531 30091 1597 30092
rect 1715 29476 1781 29477
rect 1715 29412 1716 29476
rect 1780 29412 1781 29476
rect 1715 29411 1781 29412
rect 1718 20093 1778 29411
rect 1899 21860 1965 21861
rect 1899 21796 1900 21860
rect 1964 21796 1965 21860
rect 1899 21795 1965 21796
rect 1715 20092 1781 20093
rect 1715 20028 1716 20092
rect 1780 20028 1781 20092
rect 1715 20027 1781 20028
rect 1531 19412 1597 19413
rect 1531 19348 1532 19412
rect 1596 19348 1597 19412
rect 1531 19347 1597 19348
rect 1534 12205 1594 19347
rect 1715 17372 1781 17373
rect 1715 17308 1716 17372
rect 1780 17370 1781 17372
rect 1902 17370 1962 21795
rect 2086 20637 2146 32811
rect 2451 32332 2517 32333
rect 2451 32268 2452 32332
rect 2516 32268 2517 32332
rect 2451 32267 2517 32268
rect 2267 26076 2333 26077
rect 2267 26012 2268 26076
rect 2332 26012 2333 26076
rect 2267 26011 2333 26012
rect 2083 20636 2149 20637
rect 2083 20572 2084 20636
rect 2148 20572 2149 20636
rect 2083 20571 2149 20572
rect 2270 19549 2330 26011
rect 2454 23493 2514 32267
rect 2638 31517 2698 40291
rect 3742 39269 3802 41515
rect 3876 40832 4196 41856
rect 3876 40768 3884 40832
rect 3948 40768 3964 40832
rect 4028 40768 4044 40832
rect 4108 40768 4124 40832
rect 4188 40768 4196 40832
rect 3876 39744 4196 40768
rect 4846 40085 4906 42467
rect 6808 42464 7128 43488
rect 6808 42400 6816 42464
rect 6880 42400 6896 42464
rect 6960 42400 6976 42464
rect 7040 42400 7056 42464
rect 7120 42400 7128 42464
rect 5579 42124 5645 42125
rect 5579 42060 5580 42124
rect 5644 42060 5645 42124
rect 5579 42059 5645 42060
rect 4843 40084 4909 40085
rect 4843 40020 4844 40084
rect 4908 40020 4909 40084
rect 4843 40019 4909 40020
rect 3876 39680 3884 39744
rect 3948 39680 3964 39744
rect 4028 39680 4044 39744
rect 4108 39680 4124 39744
rect 4188 39680 4196 39744
rect 3739 39268 3805 39269
rect 3739 39204 3740 39268
rect 3804 39204 3805 39268
rect 3739 39203 3805 39204
rect 3739 38996 3805 38997
rect 3739 38932 3740 38996
rect 3804 38932 3805 38996
rect 3739 38931 3805 38932
rect 3555 38452 3621 38453
rect 3555 38388 3556 38452
rect 3620 38388 3621 38452
rect 3555 38387 3621 38388
rect 3371 38180 3437 38181
rect 3371 38116 3372 38180
rect 3436 38116 3437 38180
rect 3371 38115 3437 38116
rect 3374 33557 3434 38115
rect 3558 36277 3618 38387
rect 3742 36821 3802 38931
rect 3876 38656 4196 39680
rect 5211 39268 5277 39269
rect 5211 39204 5212 39268
rect 5276 39204 5277 39268
rect 5211 39203 5277 39204
rect 3876 38592 3884 38656
rect 3948 38592 3964 38656
rect 4028 38592 4044 38656
rect 4108 38592 4124 38656
rect 4188 38592 4196 38656
rect 3876 37568 4196 38592
rect 4291 38180 4357 38181
rect 4291 38116 4292 38180
rect 4356 38116 4357 38180
rect 4291 38115 4357 38116
rect 3876 37504 3884 37568
rect 3948 37504 3964 37568
rect 4028 37504 4044 37568
rect 4108 37504 4124 37568
rect 4188 37504 4196 37568
rect 3739 36820 3805 36821
rect 3739 36756 3740 36820
rect 3804 36756 3805 36820
rect 3739 36755 3805 36756
rect 3555 36276 3621 36277
rect 3555 36212 3556 36276
rect 3620 36212 3621 36276
rect 3555 36211 3621 36212
rect 3555 36140 3621 36141
rect 3555 36076 3556 36140
rect 3620 36076 3621 36140
rect 3555 36075 3621 36076
rect 3371 33556 3437 33557
rect 3371 33492 3372 33556
rect 3436 33492 3437 33556
rect 3371 33491 3437 33492
rect 2819 31788 2885 31789
rect 2819 31724 2820 31788
rect 2884 31724 2885 31788
rect 2819 31723 2885 31724
rect 2635 31516 2701 31517
rect 2635 31452 2636 31516
rect 2700 31452 2701 31516
rect 2635 31451 2701 31452
rect 2635 31380 2701 31381
rect 2635 31316 2636 31380
rect 2700 31316 2701 31380
rect 2635 31315 2701 31316
rect 2638 24989 2698 31315
rect 2822 25669 2882 31723
rect 2819 25668 2885 25669
rect 2819 25604 2820 25668
rect 2884 25604 2885 25668
rect 2819 25603 2885 25604
rect 2635 24988 2701 24989
rect 2635 24924 2636 24988
rect 2700 24924 2701 24988
rect 2635 24923 2701 24924
rect 2819 24580 2885 24581
rect 2819 24516 2820 24580
rect 2884 24516 2885 24580
rect 2819 24515 2885 24516
rect 2451 23492 2517 23493
rect 2451 23428 2452 23492
rect 2516 23428 2517 23492
rect 2451 23427 2517 23428
rect 2267 19548 2333 19549
rect 2267 19484 2268 19548
rect 2332 19484 2333 19548
rect 2267 19483 2333 19484
rect 1780 17310 1962 17370
rect 1780 17308 1781 17310
rect 1715 17307 1781 17308
rect 1531 12204 1597 12205
rect 1531 12140 1532 12204
rect 1596 12140 1597 12204
rect 1531 12139 1597 12140
rect 1718 4725 1778 17307
rect 1899 15740 1965 15741
rect 1899 15676 1900 15740
rect 1964 15676 1965 15740
rect 1899 15675 1965 15676
rect 1902 5541 1962 15675
rect 2270 14925 2330 19483
rect 2635 18732 2701 18733
rect 2635 18668 2636 18732
rect 2700 18668 2701 18732
rect 2635 18667 2701 18668
rect 2638 15333 2698 18667
rect 2635 15332 2701 15333
rect 2635 15268 2636 15332
rect 2700 15268 2701 15332
rect 2635 15267 2701 15268
rect 2267 14924 2333 14925
rect 2267 14860 2268 14924
rect 2332 14860 2333 14924
rect 2267 14859 2333 14860
rect 2083 12204 2149 12205
rect 2083 12140 2084 12204
rect 2148 12140 2149 12204
rect 2083 12139 2149 12140
rect 1899 5540 1965 5541
rect 1899 5476 1900 5540
rect 1964 5476 1965 5540
rect 1899 5475 1965 5476
rect 1715 4724 1781 4725
rect 1715 4660 1716 4724
rect 1780 4660 1781 4724
rect 1715 4659 1781 4660
rect 2086 3909 2146 12139
rect 2270 6493 2330 14859
rect 2822 8533 2882 24515
rect 3558 23357 3618 36075
rect 3742 33149 3802 36755
rect 3876 36480 4196 37504
rect 3876 36416 3884 36480
rect 3948 36416 3964 36480
rect 4028 36416 4044 36480
rect 4108 36416 4124 36480
rect 4188 36416 4196 36480
rect 3876 35392 4196 36416
rect 3876 35328 3884 35392
rect 3948 35328 3964 35392
rect 4028 35328 4044 35392
rect 4108 35328 4124 35392
rect 4188 35328 4196 35392
rect 3876 34304 4196 35328
rect 3876 34240 3884 34304
rect 3948 34240 3964 34304
rect 4028 34240 4044 34304
rect 4108 34240 4124 34304
rect 4188 34240 4196 34304
rect 3876 33216 4196 34240
rect 3876 33152 3884 33216
rect 3948 33152 3964 33216
rect 4028 33152 4044 33216
rect 4108 33152 4124 33216
rect 4188 33152 4196 33216
rect 3739 33148 3805 33149
rect 3739 33084 3740 33148
rect 3804 33084 3805 33148
rect 3739 33083 3805 33084
rect 3876 32128 4196 33152
rect 4294 33149 4354 38115
rect 4659 37092 4725 37093
rect 4659 37028 4660 37092
rect 4724 37028 4725 37092
rect 4659 37027 4725 37028
rect 4475 36548 4541 36549
rect 4475 36484 4476 36548
rect 4540 36484 4541 36548
rect 4475 36483 4541 36484
rect 4478 33965 4538 36483
rect 4475 33964 4541 33965
rect 4475 33900 4476 33964
rect 4540 33900 4541 33964
rect 4475 33899 4541 33900
rect 4291 33148 4357 33149
rect 4291 33084 4292 33148
rect 4356 33084 4357 33148
rect 4291 33083 4357 33084
rect 3876 32064 3884 32128
rect 3948 32064 3964 32128
rect 4028 32064 4044 32128
rect 4108 32064 4124 32128
rect 4188 32064 4196 32128
rect 3876 31040 4196 32064
rect 3876 30976 3884 31040
rect 3948 30976 3964 31040
rect 4028 30976 4044 31040
rect 4108 30976 4124 31040
rect 4188 30976 4196 31040
rect 3876 29952 4196 30976
rect 3876 29888 3884 29952
rect 3948 29888 3964 29952
rect 4028 29888 4044 29952
rect 4108 29888 4124 29952
rect 4188 29888 4196 29952
rect 3876 28864 4196 29888
rect 3876 28800 3884 28864
rect 3948 28800 3964 28864
rect 4028 28800 4044 28864
rect 4108 28800 4124 28864
rect 4188 28800 4196 28864
rect 3876 27776 4196 28800
rect 3876 27712 3884 27776
rect 3948 27712 3964 27776
rect 4028 27712 4044 27776
rect 4108 27712 4124 27776
rect 4188 27712 4196 27776
rect 3739 27028 3805 27029
rect 3739 26964 3740 27028
rect 3804 26964 3805 27028
rect 3739 26963 3805 26964
rect 3555 23356 3621 23357
rect 3555 23292 3556 23356
rect 3620 23292 3621 23356
rect 3555 23291 3621 23292
rect 3187 20908 3253 20909
rect 3187 20844 3188 20908
rect 3252 20844 3253 20908
rect 3187 20843 3253 20844
rect 3003 17508 3069 17509
rect 3003 17444 3004 17508
rect 3068 17444 3069 17508
rect 3003 17443 3069 17444
rect 3006 10573 3066 17443
rect 3003 10572 3069 10573
rect 3003 10508 3004 10572
rect 3068 10508 3069 10572
rect 3003 10507 3069 10508
rect 2819 8532 2885 8533
rect 2819 8468 2820 8532
rect 2884 8468 2885 8532
rect 2819 8467 2885 8468
rect 2267 6492 2333 6493
rect 2267 6428 2268 6492
rect 2332 6428 2333 6492
rect 2267 6427 2333 6428
rect 2822 4045 2882 8467
rect 3190 8397 3250 20843
rect 3742 19957 3802 26963
rect 3876 26688 4196 27712
rect 4294 27573 4354 33083
rect 4291 27572 4357 27573
rect 4291 27508 4292 27572
rect 4356 27508 4357 27572
rect 4291 27507 4357 27508
rect 4662 27301 4722 37027
rect 5214 35733 5274 39203
rect 5395 37500 5461 37501
rect 5395 37436 5396 37500
rect 5460 37436 5461 37500
rect 5395 37435 5461 37436
rect 5211 35732 5277 35733
rect 5211 35668 5212 35732
rect 5276 35668 5277 35732
rect 5211 35667 5277 35668
rect 5398 35050 5458 37435
rect 5214 34990 5458 35050
rect 5214 34237 5274 34990
rect 5211 34236 5277 34237
rect 5211 34172 5212 34236
rect 5276 34172 5277 34236
rect 5211 34171 5277 34172
rect 5214 30293 5274 34171
rect 5582 31789 5642 42059
rect 6131 41444 6197 41445
rect 6131 41380 6132 41444
rect 6196 41380 6197 41444
rect 6131 41379 6197 41380
rect 5947 35732 6013 35733
rect 5947 35668 5948 35732
rect 6012 35668 6013 35732
rect 5947 35667 6013 35668
rect 5950 32197 6010 35667
rect 6134 34509 6194 41379
rect 6808 41376 7128 42400
rect 9741 43008 10061 43568
rect 12673 43552 12993 43568
rect 12673 43488 12681 43552
rect 12745 43488 12761 43552
rect 12825 43488 12841 43552
rect 12905 43488 12921 43552
rect 12985 43488 12993 43552
rect 11651 43076 11717 43077
rect 11651 43012 11652 43076
rect 11716 43012 11717 43076
rect 11651 43011 11717 43012
rect 9741 42944 9749 43008
rect 9813 42944 9829 43008
rect 9893 42944 9909 43008
rect 9973 42944 9989 43008
rect 10053 42944 10061 43008
rect 8891 41988 8957 41989
rect 8891 41924 8892 41988
rect 8956 41924 8957 41988
rect 8891 41923 8957 41924
rect 6808 41312 6816 41376
rect 6880 41312 6896 41376
rect 6960 41312 6976 41376
rect 7040 41312 7056 41376
rect 7120 41312 7128 41376
rect 6808 40288 7128 41312
rect 6808 40224 6816 40288
rect 6880 40224 6896 40288
rect 6960 40224 6976 40288
rect 7040 40224 7056 40288
rect 7120 40224 7128 40288
rect 6808 39200 7128 40224
rect 6808 39136 6816 39200
rect 6880 39136 6896 39200
rect 6960 39136 6976 39200
rect 7040 39136 7056 39200
rect 7120 39136 7128 39200
rect 6315 39132 6381 39133
rect 6315 39068 6316 39132
rect 6380 39068 6381 39132
rect 6315 39067 6381 39068
rect 6131 34508 6197 34509
rect 6131 34444 6132 34508
rect 6196 34444 6197 34508
rect 6131 34443 6197 34444
rect 6131 33148 6197 33149
rect 6131 33084 6132 33148
rect 6196 33084 6197 33148
rect 6131 33083 6197 33084
rect 5947 32196 6013 32197
rect 5947 32132 5948 32196
rect 6012 32132 6013 32196
rect 5947 32131 6013 32132
rect 5579 31788 5645 31789
rect 5579 31724 5580 31788
rect 5644 31724 5645 31788
rect 5579 31723 5645 31724
rect 5579 31516 5645 31517
rect 5579 31452 5580 31516
rect 5644 31452 5645 31516
rect 5579 31451 5645 31452
rect 5211 30292 5277 30293
rect 5211 30228 5212 30292
rect 5276 30228 5277 30292
rect 5211 30227 5277 30228
rect 5027 29884 5093 29885
rect 5027 29820 5028 29884
rect 5092 29820 5093 29884
rect 5027 29819 5093 29820
rect 4659 27300 4725 27301
rect 4659 27236 4660 27300
rect 4724 27236 4725 27300
rect 4659 27235 4725 27236
rect 4475 27164 4541 27165
rect 4475 27100 4476 27164
rect 4540 27100 4541 27164
rect 4475 27099 4541 27100
rect 3876 26624 3884 26688
rect 3948 26624 3964 26688
rect 4028 26624 4044 26688
rect 4108 26624 4124 26688
rect 4188 26624 4196 26688
rect 3876 25600 4196 26624
rect 3876 25536 3884 25600
rect 3948 25536 3964 25600
rect 4028 25536 4044 25600
rect 4108 25536 4124 25600
rect 4188 25536 4196 25600
rect 3876 24512 4196 25536
rect 3876 24448 3884 24512
rect 3948 24448 3964 24512
rect 4028 24448 4044 24512
rect 4108 24448 4124 24512
rect 4188 24448 4196 24512
rect 3876 23424 4196 24448
rect 3876 23360 3884 23424
rect 3948 23360 3964 23424
rect 4028 23360 4044 23424
rect 4108 23360 4124 23424
rect 4188 23360 4196 23424
rect 3876 22336 4196 23360
rect 3876 22272 3884 22336
rect 3948 22272 3964 22336
rect 4028 22272 4044 22336
rect 4108 22272 4124 22336
rect 4188 22272 4196 22336
rect 3876 21248 4196 22272
rect 4478 21997 4538 27099
rect 4662 26893 4722 27235
rect 4659 26892 4725 26893
rect 4659 26828 4660 26892
rect 4724 26828 4725 26892
rect 4659 26827 4725 26828
rect 5030 24173 5090 29819
rect 5214 26213 5274 30227
rect 5582 29069 5642 31451
rect 5579 29068 5645 29069
rect 5579 29004 5580 29068
rect 5644 29004 5645 29068
rect 5579 29003 5645 29004
rect 5763 27708 5829 27709
rect 5763 27644 5764 27708
rect 5828 27644 5829 27708
rect 5763 27643 5829 27644
rect 5766 26621 5826 27643
rect 5763 26620 5829 26621
rect 5763 26556 5764 26620
rect 5828 26556 5829 26620
rect 5763 26555 5829 26556
rect 5211 26212 5277 26213
rect 5211 26148 5212 26212
rect 5276 26148 5277 26212
rect 5211 26147 5277 26148
rect 5211 26076 5277 26077
rect 5211 26012 5212 26076
rect 5276 26012 5277 26076
rect 5211 26011 5277 26012
rect 5027 24172 5093 24173
rect 5027 24108 5028 24172
rect 5092 24108 5093 24172
rect 5027 24107 5093 24108
rect 5027 23492 5093 23493
rect 5027 23428 5028 23492
rect 5092 23428 5093 23492
rect 5027 23427 5093 23428
rect 4475 21996 4541 21997
rect 4475 21932 4476 21996
rect 4540 21932 4541 21996
rect 4475 21931 4541 21932
rect 3876 21184 3884 21248
rect 3948 21184 3964 21248
rect 4028 21184 4044 21248
rect 4108 21184 4124 21248
rect 4188 21184 4196 21248
rect 3876 20160 4196 21184
rect 3876 20096 3884 20160
rect 3948 20096 3964 20160
rect 4028 20096 4044 20160
rect 4108 20096 4124 20160
rect 4188 20096 4196 20160
rect 3739 19956 3805 19957
rect 3739 19892 3740 19956
rect 3804 19892 3805 19956
rect 3739 19891 3805 19892
rect 3371 19684 3437 19685
rect 3371 19620 3372 19684
rect 3436 19620 3437 19684
rect 3371 19619 3437 19620
rect 3187 8396 3253 8397
rect 3187 8332 3188 8396
rect 3252 8332 3253 8396
rect 3187 8331 3253 8332
rect 3374 7853 3434 19619
rect 3876 19072 4196 20096
rect 4291 19140 4357 19141
rect 4291 19076 4292 19140
rect 4356 19076 4357 19140
rect 4291 19075 4357 19076
rect 3876 19008 3884 19072
rect 3948 19008 3964 19072
rect 4028 19008 4044 19072
rect 4108 19008 4124 19072
rect 4188 19008 4196 19072
rect 3876 17984 4196 19008
rect 3876 17920 3884 17984
rect 3948 17920 3964 17984
rect 4028 17920 4044 17984
rect 4108 17920 4124 17984
rect 4188 17920 4196 17984
rect 3876 16896 4196 17920
rect 3876 16832 3884 16896
rect 3948 16832 3964 16896
rect 4028 16832 4044 16896
rect 4108 16832 4124 16896
rect 4188 16832 4196 16896
rect 3876 15808 4196 16832
rect 3876 15744 3884 15808
rect 3948 15744 3964 15808
rect 4028 15744 4044 15808
rect 4108 15744 4124 15808
rect 4188 15744 4196 15808
rect 3876 14720 4196 15744
rect 3876 14656 3884 14720
rect 3948 14656 3964 14720
rect 4028 14656 4044 14720
rect 4108 14656 4124 14720
rect 4188 14656 4196 14720
rect 3876 13632 4196 14656
rect 3876 13568 3884 13632
rect 3948 13568 3964 13632
rect 4028 13568 4044 13632
rect 4108 13568 4124 13632
rect 4188 13568 4196 13632
rect 3876 12544 4196 13568
rect 3876 12480 3884 12544
rect 3948 12480 3964 12544
rect 4028 12480 4044 12544
rect 4108 12480 4124 12544
rect 4188 12480 4196 12544
rect 3876 11456 4196 12480
rect 3876 11392 3884 11456
rect 3948 11392 3964 11456
rect 4028 11392 4044 11456
rect 4108 11392 4124 11456
rect 4188 11392 4196 11456
rect 3876 10368 4196 11392
rect 4294 10981 4354 19075
rect 4478 12613 4538 21931
rect 4475 12612 4541 12613
rect 4475 12548 4476 12612
rect 4540 12548 4541 12612
rect 4475 12547 4541 12548
rect 4475 11932 4541 11933
rect 4475 11868 4476 11932
rect 4540 11868 4541 11932
rect 4475 11867 4541 11868
rect 4291 10980 4357 10981
rect 4291 10916 4292 10980
rect 4356 10916 4357 10980
rect 4291 10915 4357 10916
rect 3876 10304 3884 10368
rect 3948 10304 3964 10368
rect 4028 10304 4044 10368
rect 4108 10304 4124 10368
rect 4188 10304 4196 10368
rect 3876 9280 4196 10304
rect 4291 9620 4357 9621
rect 4291 9556 4292 9620
rect 4356 9556 4357 9620
rect 4291 9555 4357 9556
rect 3876 9216 3884 9280
rect 3948 9216 3964 9280
rect 4028 9216 4044 9280
rect 4108 9216 4124 9280
rect 4188 9216 4196 9280
rect 3739 8396 3805 8397
rect 3739 8332 3740 8396
rect 3804 8332 3805 8396
rect 3739 8331 3805 8332
rect 3371 7852 3437 7853
rect 3371 7788 3372 7852
rect 3436 7788 3437 7852
rect 3371 7787 3437 7788
rect 3742 5677 3802 8331
rect 3876 8192 4196 9216
rect 4294 9077 4354 9555
rect 4291 9076 4357 9077
rect 4291 9012 4292 9076
rect 4356 9012 4357 9076
rect 4291 9011 4357 9012
rect 3876 8128 3884 8192
rect 3948 8128 3964 8192
rect 4028 8128 4044 8192
rect 4108 8128 4124 8192
rect 4188 8128 4196 8192
rect 3876 7104 4196 8128
rect 3876 7040 3884 7104
rect 3948 7040 3964 7104
rect 4028 7040 4044 7104
rect 4108 7040 4124 7104
rect 4188 7040 4196 7104
rect 3876 6016 4196 7040
rect 3876 5952 3884 6016
rect 3948 5952 3964 6016
rect 4028 5952 4044 6016
rect 4108 5952 4124 6016
rect 4188 5952 4196 6016
rect 3739 5676 3805 5677
rect 3739 5612 3740 5676
rect 3804 5612 3805 5676
rect 3739 5611 3805 5612
rect 3876 4928 4196 5952
rect 3876 4864 3884 4928
rect 3948 4864 3964 4928
rect 4028 4864 4044 4928
rect 4108 4864 4124 4928
rect 4188 4864 4196 4928
rect 3739 4180 3805 4181
rect 3739 4116 3740 4180
rect 3804 4116 3805 4180
rect 3739 4115 3805 4116
rect 2819 4044 2885 4045
rect 2819 3980 2820 4044
rect 2884 3980 2885 4044
rect 2819 3979 2885 3980
rect 2083 3908 2149 3909
rect 2083 3844 2084 3908
rect 2148 3844 2149 3908
rect 2083 3843 2149 3844
rect 1163 1868 1229 1869
rect 1163 1804 1164 1868
rect 1228 1804 1229 1868
rect 1163 1803 1229 1804
rect 3742 1461 3802 4115
rect 3876 3840 4196 4864
rect 3876 3776 3884 3840
rect 3948 3776 3964 3840
rect 4028 3776 4044 3840
rect 4108 3776 4124 3840
rect 4188 3776 4196 3840
rect 3876 2752 4196 3776
rect 3876 2688 3884 2752
rect 3948 2688 3964 2752
rect 4028 2688 4044 2752
rect 4108 2688 4124 2752
rect 4188 2688 4196 2752
rect 3876 1664 4196 2688
rect 3876 1600 3884 1664
rect 3948 1600 3964 1664
rect 4028 1600 4044 1664
rect 4108 1600 4124 1664
rect 4188 1600 4196 1664
rect 3739 1460 3805 1461
rect 3739 1396 3740 1460
rect 3804 1396 3805 1460
rect 3739 1395 3805 1396
rect 3876 1040 4196 1600
rect 4478 1325 4538 11867
rect 5030 9893 5090 23427
rect 5214 15877 5274 26011
rect 5950 25669 6010 32131
rect 6134 27709 6194 33083
rect 6318 28525 6378 39067
rect 6808 38112 7128 39136
rect 6808 38048 6816 38112
rect 6880 38048 6896 38112
rect 6960 38048 6976 38112
rect 7040 38048 7056 38112
rect 7120 38048 7128 38112
rect 6808 37024 7128 38048
rect 6808 36960 6816 37024
rect 6880 36960 6896 37024
rect 6960 36960 6976 37024
rect 7040 36960 7056 37024
rect 7120 36960 7128 37024
rect 6808 35936 7128 36960
rect 6808 35872 6816 35936
rect 6880 35872 6896 35936
rect 6960 35872 6976 35936
rect 7040 35872 7056 35936
rect 7120 35872 7128 35936
rect 6808 34848 7128 35872
rect 6808 34784 6816 34848
rect 6880 34784 6896 34848
rect 6960 34784 6976 34848
rect 7040 34784 7056 34848
rect 7120 34784 7128 34848
rect 6808 33760 7128 34784
rect 7971 34508 8037 34509
rect 7971 34444 7972 34508
rect 8036 34444 8037 34508
rect 7971 34443 8037 34444
rect 7603 34100 7669 34101
rect 7603 34036 7604 34100
rect 7668 34036 7669 34100
rect 7603 34035 7669 34036
rect 6808 33696 6816 33760
rect 6880 33696 6896 33760
rect 6960 33696 6976 33760
rect 7040 33696 7056 33760
rect 7120 33696 7128 33760
rect 6499 33556 6565 33557
rect 6499 33492 6500 33556
rect 6564 33492 6565 33556
rect 6499 33491 6565 33492
rect 6502 29069 6562 33491
rect 6808 32672 7128 33696
rect 6808 32608 6816 32672
rect 6880 32608 6896 32672
rect 6960 32608 6976 32672
rect 7040 32608 7056 32672
rect 7120 32608 7128 32672
rect 6808 31584 7128 32608
rect 7606 31653 7666 34035
rect 7787 32468 7853 32469
rect 7787 32404 7788 32468
rect 7852 32404 7853 32468
rect 7787 32403 7853 32404
rect 7603 31652 7669 31653
rect 7603 31588 7604 31652
rect 7668 31588 7669 31652
rect 7603 31587 7669 31588
rect 6808 31520 6816 31584
rect 6880 31520 6896 31584
rect 6960 31520 6976 31584
rect 7040 31520 7056 31584
rect 7120 31520 7128 31584
rect 6808 30496 7128 31520
rect 6808 30432 6816 30496
rect 6880 30432 6896 30496
rect 6960 30432 6976 30496
rect 7040 30432 7056 30496
rect 7120 30432 7128 30496
rect 6808 29408 7128 30432
rect 6808 29344 6816 29408
rect 6880 29344 6896 29408
rect 6960 29344 6976 29408
rect 7040 29344 7056 29408
rect 7120 29344 7128 29408
rect 6499 29068 6565 29069
rect 6499 29004 6500 29068
rect 6564 29004 6565 29068
rect 6499 29003 6565 29004
rect 6315 28524 6381 28525
rect 6315 28460 6316 28524
rect 6380 28460 6381 28524
rect 6315 28459 6381 28460
rect 6131 27708 6197 27709
rect 6131 27644 6132 27708
rect 6196 27644 6197 27708
rect 6131 27643 6197 27644
rect 6318 27570 6378 28459
rect 6134 27510 6378 27570
rect 6134 26893 6194 27510
rect 6131 26892 6197 26893
rect 6131 26828 6132 26892
rect 6196 26828 6197 26892
rect 6131 26827 6197 26828
rect 6315 26892 6381 26893
rect 6315 26828 6316 26892
rect 6380 26828 6381 26892
rect 6315 26827 6381 26828
rect 5947 25668 6013 25669
rect 5947 25604 5948 25668
rect 6012 25604 6013 25668
rect 5947 25603 6013 25604
rect 5395 25396 5461 25397
rect 5395 25332 5396 25396
rect 5460 25332 5461 25396
rect 5395 25331 5461 25332
rect 5398 20637 5458 25331
rect 5763 24988 5829 24989
rect 5763 24924 5764 24988
rect 5828 24924 5829 24988
rect 5763 24923 5829 24924
rect 5395 20636 5461 20637
rect 5395 20572 5396 20636
rect 5460 20572 5461 20636
rect 5395 20571 5461 20572
rect 5395 19956 5461 19957
rect 5395 19892 5396 19956
rect 5460 19892 5461 19956
rect 5395 19891 5461 19892
rect 5398 16149 5458 19891
rect 5579 19684 5645 19685
rect 5579 19620 5580 19684
rect 5644 19620 5645 19684
rect 5579 19619 5645 19620
rect 5395 16148 5461 16149
rect 5395 16084 5396 16148
rect 5460 16084 5461 16148
rect 5395 16083 5461 16084
rect 5211 15876 5277 15877
rect 5211 15812 5212 15876
rect 5276 15812 5277 15876
rect 5211 15811 5277 15812
rect 5582 14925 5642 19619
rect 5766 17917 5826 24923
rect 6318 18053 6378 26827
rect 6315 18052 6381 18053
rect 6315 17988 6316 18052
rect 6380 17988 6381 18052
rect 6315 17987 6381 17988
rect 5763 17916 5829 17917
rect 5763 17852 5764 17916
rect 5828 17852 5829 17916
rect 5763 17851 5829 17852
rect 6502 17237 6562 29003
rect 6808 28320 7128 29344
rect 6808 28256 6816 28320
rect 6880 28256 6896 28320
rect 6960 28256 6976 28320
rect 7040 28256 7056 28320
rect 7120 28256 7128 28320
rect 6808 27232 7128 28256
rect 7603 27300 7669 27301
rect 7603 27236 7604 27300
rect 7668 27236 7669 27300
rect 7603 27235 7669 27236
rect 6808 27168 6816 27232
rect 6880 27168 6896 27232
rect 6960 27168 6976 27232
rect 7040 27168 7056 27232
rect 7120 27168 7128 27232
rect 6808 26144 7128 27168
rect 7419 27164 7485 27165
rect 7419 27100 7420 27164
rect 7484 27100 7485 27164
rect 7419 27099 7485 27100
rect 6808 26080 6816 26144
rect 6880 26080 6896 26144
rect 6960 26080 6976 26144
rect 7040 26080 7056 26144
rect 7120 26080 7128 26144
rect 6808 25056 7128 26080
rect 6808 24992 6816 25056
rect 6880 24992 6896 25056
rect 6960 24992 6976 25056
rect 7040 24992 7056 25056
rect 7120 24992 7128 25056
rect 6808 23968 7128 24992
rect 6808 23904 6816 23968
rect 6880 23904 6896 23968
rect 6960 23904 6976 23968
rect 7040 23904 7056 23968
rect 7120 23904 7128 23968
rect 6808 22880 7128 23904
rect 6808 22816 6816 22880
rect 6880 22816 6896 22880
rect 6960 22816 6976 22880
rect 7040 22816 7056 22880
rect 7120 22816 7128 22880
rect 6808 21792 7128 22816
rect 6808 21728 6816 21792
rect 6880 21728 6896 21792
rect 6960 21728 6976 21792
rect 7040 21728 7056 21792
rect 7120 21728 7128 21792
rect 6808 20704 7128 21728
rect 6808 20640 6816 20704
rect 6880 20640 6896 20704
rect 6960 20640 6976 20704
rect 7040 20640 7056 20704
rect 7120 20640 7128 20704
rect 6808 19616 7128 20640
rect 6808 19552 6816 19616
rect 6880 19552 6896 19616
rect 6960 19552 6976 19616
rect 7040 19552 7056 19616
rect 7120 19552 7128 19616
rect 6808 18528 7128 19552
rect 6808 18464 6816 18528
rect 6880 18464 6896 18528
rect 6960 18464 6976 18528
rect 7040 18464 7056 18528
rect 7120 18464 7128 18528
rect 6808 17440 7128 18464
rect 6808 17376 6816 17440
rect 6880 17376 6896 17440
rect 6960 17376 6976 17440
rect 7040 17376 7056 17440
rect 7120 17376 7128 17440
rect 6499 17236 6565 17237
rect 6499 17172 6500 17236
rect 6564 17172 6565 17236
rect 6499 17171 6565 17172
rect 6808 16352 7128 17376
rect 6808 16288 6816 16352
rect 6880 16288 6896 16352
rect 6960 16288 6976 16352
rect 7040 16288 7056 16352
rect 7120 16288 7128 16352
rect 6808 15264 7128 16288
rect 6808 15200 6816 15264
rect 6880 15200 6896 15264
rect 6960 15200 6976 15264
rect 7040 15200 7056 15264
rect 7120 15200 7128 15264
rect 5579 14924 5645 14925
rect 5579 14860 5580 14924
rect 5644 14860 5645 14924
rect 5579 14859 5645 14860
rect 6131 14380 6197 14381
rect 6131 14316 6132 14380
rect 6196 14316 6197 14380
rect 6131 14315 6197 14316
rect 5395 11116 5461 11117
rect 5395 11052 5396 11116
rect 5460 11052 5461 11116
rect 5395 11051 5461 11052
rect 5027 9892 5093 9893
rect 5027 9828 5028 9892
rect 5092 9828 5093 9892
rect 5027 9827 5093 9828
rect 5398 2685 5458 11051
rect 5395 2684 5461 2685
rect 5395 2620 5396 2684
rect 5460 2620 5461 2684
rect 5395 2619 5461 2620
rect 4475 1324 4541 1325
rect 4475 1260 4476 1324
rect 4540 1260 4541 1324
rect 4475 1259 4541 1260
rect 6134 1189 6194 14315
rect 6808 14176 7128 15200
rect 6808 14112 6816 14176
rect 6880 14112 6896 14176
rect 6960 14112 6976 14176
rect 7040 14112 7056 14176
rect 7120 14112 7128 14176
rect 6808 13088 7128 14112
rect 6808 13024 6816 13088
rect 6880 13024 6896 13088
rect 6960 13024 6976 13088
rect 7040 13024 7056 13088
rect 7120 13024 7128 13088
rect 6808 12000 7128 13024
rect 7422 12205 7482 27099
rect 7606 21861 7666 27235
rect 7603 21860 7669 21861
rect 7603 21796 7604 21860
rect 7668 21796 7669 21860
rect 7603 21795 7669 21796
rect 7419 12204 7485 12205
rect 7419 12140 7420 12204
rect 7484 12140 7485 12204
rect 7419 12139 7485 12140
rect 6808 11936 6816 12000
rect 6880 11936 6896 12000
rect 6960 11936 6976 12000
rect 7040 11936 7056 12000
rect 7120 11936 7128 12000
rect 6808 10912 7128 11936
rect 7790 11389 7850 32403
rect 7974 30021 8034 34443
rect 8155 32332 8221 32333
rect 8155 32268 8156 32332
rect 8220 32268 8221 32332
rect 8155 32267 8221 32268
rect 7971 30020 8037 30021
rect 7971 29956 7972 30020
rect 8036 29956 8037 30020
rect 7971 29955 8037 29956
rect 7974 26213 8034 29955
rect 7971 26212 8037 26213
rect 7971 26148 7972 26212
rect 8036 26148 8037 26212
rect 7971 26147 8037 26148
rect 8158 22110 8218 32267
rect 8707 29884 8773 29885
rect 8707 29820 8708 29884
rect 8772 29820 8773 29884
rect 8707 29819 8773 29820
rect 8710 28525 8770 29819
rect 8707 28524 8773 28525
rect 8707 28460 8708 28524
rect 8772 28460 8773 28524
rect 8707 28459 8773 28460
rect 8158 22050 8586 22110
rect 8526 21589 8586 22050
rect 8523 21588 8589 21589
rect 8523 21524 8524 21588
rect 8588 21524 8589 21588
rect 8523 21523 8589 21524
rect 8339 15196 8405 15197
rect 8339 15132 8340 15196
rect 8404 15132 8405 15196
rect 8339 15131 8405 15132
rect 7787 11388 7853 11389
rect 7787 11324 7788 11388
rect 7852 11324 7853 11388
rect 7787 11323 7853 11324
rect 7419 11116 7485 11117
rect 7419 11052 7420 11116
rect 7484 11052 7485 11116
rect 7419 11051 7485 11052
rect 6808 10848 6816 10912
rect 6880 10848 6896 10912
rect 6960 10848 6976 10912
rect 7040 10848 7056 10912
rect 7120 10848 7128 10912
rect 6808 9824 7128 10848
rect 6808 9760 6816 9824
rect 6880 9760 6896 9824
rect 6960 9760 6976 9824
rect 7040 9760 7056 9824
rect 7120 9760 7128 9824
rect 6808 8736 7128 9760
rect 6808 8672 6816 8736
rect 6880 8672 6896 8736
rect 6960 8672 6976 8736
rect 7040 8672 7056 8736
rect 7120 8672 7128 8736
rect 6808 7648 7128 8672
rect 6808 7584 6816 7648
rect 6880 7584 6896 7648
rect 6960 7584 6976 7648
rect 7040 7584 7056 7648
rect 7120 7584 7128 7648
rect 6808 6560 7128 7584
rect 6808 6496 6816 6560
rect 6880 6496 6896 6560
rect 6960 6496 6976 6560
rect 7040 6496 7056 6560
rect 7120 6496 7128 6560
rect 6808 5472 7128 6496
rect 6808 5408 6816 5472
rect 6880 5408 6896 5472
rect 6960 5408 6976 5472
rect 7040 5408 7056 5472
rect 7120 5408 7128 5472
rect 6808 4384 7128 5408
rect 6808 4320 6816 4384
rect 6880 4320 6896 4384
rect 6960 4320 6976 4384
rect 7040 4320 7056 4384
rect 7120 4320 7128 4384
rect 6808 3296 7128 4320
rect 6808 3232 6816 3296
rect 6880 3232 6896 3296
rect 6960 3232 6976 3296
rect 7040 3232 7056 3296
rect 7120 3232 7128 3296
rect 6808 2208 7128 3232
rect 7422 2277 7482 11051
rect 8155 9756 8221 9757
rect 8155 9692 8156 9756
rect 8220 9692 8221 9756
rect 8155 9691 8221 9692
rect 8158 2277 8218 9691
rect 7419 2276 7485 2277
rect 7419 2212 7420 2276
rect 7484 2212 7485 2276
rect 7419 2211 7485 2212
rect 8155 2276 8221 2277
rect 8155 2212 8156 2276
rect 8220 2212 8221 2276
rect 8155 2211 8221 2212
rect 6808 2144 6816 2208
rect 6880 2144 6896 2208
rect 6960 2144 6976 2208
rect 7040 2144 7056 2208
rect 7120 2144 7128 2208
rect 6131 1188 6197 1189
rect 6131 1124 6132 1188
rect 6196 1124 6197 1188
rect 6131 1123 6197 1124
rect 6808 1120 7128 2144
rect 8342 1189 8402 15131
rect 8526 13157 8586 21523
rect 8707 21044 8773 21045
rect 8707 20980 8708 21044
rect 8772 20980 8773 21044
rect 8707 20979 8773 20980
rect 8710 18461 8770 20979
rect 8707 18460 8773 18461
rect 8707 18396 8708 18460
rect 8772 18396 8773 18460
rect 8707 18395 8773 18396
rect 8523 13156 8589 13157
rect 8523 13092 8524 13156
rect 8588 13092 8589 13156
rect 8523 13091 8589 13092
rect 8707 8940 8773 8941
rect 8707 8876 8708 8940
rect 8772 8876 8773 8940
rect 8707 8875 8773 8876
rect 8710 1325 8770 8875
rect 8894 2277 8954 41923
rect 9741 41920 10061 42944
rect 10363 42124 10429 42125
rect 10363 42060 10364 42124
rect 10428 42060 10429 42124
rect 10363 42059 10429 42060
rect 9741 41856 9749 41920
rect 9813 41856 9829 41920
rect 9893 41856 9909 41920
rect 9973 41856 9989 41920
rect 10053 41856 10061 41920
rect 9075 41852 9141 41853
rect 9075 41788 9076 41852
rect 9140 41788 9141 41852
rect 9075 41787 9141 41788
rect 9078 16557 9138 41787
rect 9259 41580 9325 41581
rect 9259 41516 9260 41580
rect 9324 41516 9325 41580
rect 9259 41515 9325 41516
rect 9443 41580 9509 41581
rect 9443 41516 9444 41580
rect 9508 41516 9509 41580
rect 9443 41515 9509 41516
rect 9075 16556 9141 16557
rect 9075 16492 9076 16556
rect 9140 16492 9141 16556
rect 9075 16491 9141 16492
rect 9262 9757 9322 41515
rect 9446 20773 9506 41515
rect 9741 40832 10061 41856
rect 9741 40768 9749 40832
rect 9813 40768 9829 40832
rect 9893 40768 9909 40832
rect 9973 40768 9989 40832
rect 10053 40768 10061 40832
rect 9741 39744 10061 40768
rect 9741 39680 9749 39744
rect 9813 39680 9829 39744
rect 9893 39680 9909 39744
rect 9973 39680 9989 39744
rect 10053 39680 10061 39744
rect 9741 38656 10061 39680
rect 9741 38592 9749 38656
rect 9813 38592 9829 38656
rect 9893 38592 9909 38656
rect 9973 38592 9989 38656
rect 10053 38592 10061 38656
rect 9741 37568 10061 38592
rect 9741 37504 9749 37568
rect 9813 37504 9829 37568
rect 9893 37504 9909 37568
rect 9973 37504 9989 37568
rect 10053 37504 10061 37568
rect 9741 36480 10061 37504
rect 9741 36416 9749 36480
rect 9813 36416 9829 36480
rect 9893 36416 9909 36480
rect 9973 36416 9989 36480
rect 10053 36416 10061 36480
rect 9741 35392 10061 36416
rect 10179 36140 10245 36141
rect 10179 36076 10180 36140
rect 10244 36076 10245 36140
rect 10179 36075 10245 36076
rect 9741 35328 9749 35392
rect 9813 35328 9829 35392
rect 9893 35328 9909 35392
rect 9973 35328 9989 35392
rect 10053 35328 10061 35392
rect 9741 34304 10061 35328
rect 9741 34240 9749 34304
rect 9813 34240 9829 34304
rect 9893 34240 9909 34304
rect 9973 34240 9989 34304
rect 10053 34240 10061 34304
rect 9741 33216 10061 34240
rect 9741 33152 9749 33216
rect 9813 33152 9829 33216
rect 9893 33152 9909 33216
rect 9973 33152 9989 33216
rect 10053 33152 10061 33216
rect 9741 32128 10061 33152
rect 10182 32605 10242 36075
rect 10179 32604 10245 32605
rect 10179 32540 10180 32604
rect 10244 32540 10245 32604
rect 10179 32539 10245 32540
rect 9741 32064 9749 32128
rect 9813 32064 9829 32128
rect 9893 32064 9909 32128
rect 9973 32064 9989 32128
rect 10053 32064 10061 32128
rect 9741 31040 10061 32064
rect 10182 31245 10242 32539
rect 10179 31244 10245 31245
rect 10179 31180 10180 31244
rect 10244 31180 10245 31244
rect 10179 31179 10245 31180
rect 9741 30976 9749 31040
rect 9813 30976 9829 31040
rect 9893 30976 9909 31040
rect 9973 30976 9989 31040
rect 10053 30976 10061 31040
rect 9741 29952 10061 30976
rect 10179 30428 10245 30429
rect 10179 30364 10180 30428
rect 10244 30364 10245 30428
rect 10179 30363 10245 30364
rect 9741 29888 9749 29952
rect 9813 29888 9829 29952
rect 9893 29888 9909 29952
rect 9973 29888 9989 29952
rect 10053 29888 10061 29952
rect 9741 28864 10061 29888
rect 9741 28800 9749 28864
rect 9813 28800 9829 28864
rect 9893 28800 9909 28864
rect 9973 28800 9989 28864
rect 10053 28800 10061 28864
rect 9741 27776 10061 28800
rect 9741 27712 9749 27776
rect 9813 27712 9829 27776
rect 9893 27712 9909 27776
rect 9973 27712 9989 27776
rect 10053 27712 10061 27776
rect 9741 26688 10061 27712
rect 10182 27029 10242 30363
rect 10179 27028 10245 27029
rect 10179 26964 10180 27028
rect 10244 26964 10245 27028
rect 10179 26963 10245 26964
rect 10366 26893 10426 42059
rect 10915 41444 10981 41445
rect 10915 41380 10916 41444
rect 10980 41380 10981 41444
rect 10915 41379 10981 41380
rect 10547 27572 10613 27573
rect 10547 27508 10548 27572
rect 10612 27508 10613 27572
rect 10547 27507 10613 27508
rect 10363 26892 10429 26893
rect 10363 26828 10364 26892
rect 10428 26828 10429 26892
rect 10363 26827 10429 26828
rect 9741 26624 9749 26688
rect 9813 26624 9829 26688
rect 9893 26624 9909 26688
rect 9973 26624 9989 26688
rect 10053 26624 10061 26688
rect 9741 25600 10061 26624
rect 10550 26618 10610 27507
rect 10731 26892 10797 26893
rect 10731 26828 10732 26892
rect 10796 26828 10797 26892
rect 10731 26827 10797 26828
rect 10366 26558 10610 26618
rect 10179 26348 10245 26349
rect 10179 26284 10180 26348
rect 10244 26284 10245 26348
rect 10179 26283 10245 26284
rect 9741 25536 9749 25600
rect 9813 25536 9829 25600
rect 9893 25536 9909 25600
rect 9973 25536 9989 25600
rect 10053 25536 10061 25600
rect 9741 24512 10061 25536
rect 9741 24448 9749 24512
rect 9813 24448 9829 24512
rect 9893 24448 9909 24512
rect 9973 24448 9989 24512
rect 10053 24448 10061 24512
rect 9741 23424 10061 24448
rect 9741 23360 9749 23424
rect 9813 23360 9829 23424
rect 9893 23360 9909 23424
rect 9973 23360 9989 23424
rect 10053 23360 10061 23424
rect 9741 22336 10061 23360
rect 9741 22272 9749 22336
rect 9813 22272 9829 22336
rect 9893 22272 9909 22336
rect 9973 22272 9989 22336
rect 10053 22272 10061 22336
rect 9741 21248 10061 22272
rect 9741 21184 9749 21248
rect 9813 21184 9829 21248
rect 9893 21184 9909 21248
rect 9973 21184 9989 21248
rect 10053 21184 10061 21248
rect 9443 20772 9509 20773
rect 9443 20708 9444 20772
rect 9508 20708 9509 20772
rect 9443 20707 9509 20708
rect 9741 20160 10061 21184
rect 10182 20229 10242 26283
rect 10179 20228 10245 20229
rect 10179 20164 10180 20228
rect 10244 20164 10245 20228
rect 10179 20163 10245 20164
rect 9741 20096 9749 20160
rect 9813 20096 9829 20160
rect 9893 20096 9909 20160
rect 9973 20096 9989 20160
rect 10053 20096 10061 20160
rect 9741 19072 10061 20096
rect 10366 19957 10426 26558
rect 10547 22268 10613 22269
rect 10547 22204 10548 22268
rect 10612 22204 10613 22268
rect 10547 22203 10613 22204
rect 10363 19956 10429 19957
rect 10363 19892 10364 19956
rect 10428 19892 10429 19956
rect 10363 19891 10429 19892
rect 9741 19008 9749 19072
rect 9813 19008 9829 19072
rect 9893 19008 9909 19072
rect 9973 19008 9989 19072
rect 10053 19008 10061 19072
rect 9741 17984 10061 19008
rect 9741 17920 9749 17984
rect 9813 17920 9829 17984
rect 9893 17920 9909 17984
rect 9973 17920 9989 17984
rect 10053 17920 10061 17984
rect 9741 16896 10061 17920
rect 9741 16832 9749 16896
rect 9813 16832 9829 16896
rect 9893 16832 9909 16896
rect 9973 16832 9989 16896
rect 10053 16832 10061 16896
rect 9741 15808 10061 16832
rect 9741 15744 9749 15808
rect 9813 15744 9829 15808
rect 9893 15744 9909 15808
rect 9973 15744 9989 15808
rect 10053 15744 10061 15808
rect 9741 14720 10061 15744
rect 9741 14656 9749 14720
rect 9813 14656 9829 14720
rect 9893 14656 9909 14720
rect 9973 14656 9989 14720
rect 10053 14656 10061 14720
rect 9741 13632 10061 14656
rect 9741 13568 9749 13632
rect 9813 13568 9829 13632
rect 9893 13568 9909 13632
rect 9973 13568 9989 13632
rect 10053 13568 10061 13632
rect 9741 12544 10061 13568
rect 9741 12480 9749 12544
rect 9813 12480 9829 12544
rect 9893 12480 9909 12544
rect 9973 12480 9989 12544
rect 10053 12480 10061 12544
rect 9741 11456 10061 12480
rect 9741 11392 9749 11456
rect 9813 11392 9829 11456
rect 9893 11392 9909 11456
rect 9973 11392 9989 11456
rect 10053 11392 10061 11456
rect 9741 10368 10061 11392
rect 10363 11116 10429 11117
rect 10363 11052 10364 11116
rect 10428 11052 10429 11116
rect 10363 11051 10429 11052
rect 9741 10304 9749 10368
rect 9813 10304 9829 10368
rect 9893 10304 9909 10368
rect 9973 10304 9989 10368
rect 10053 10304 10061 10368
rect 9259 9756 9325 9757
rect 9259 9692 9260 9756
rect 9324 9692 9325 9756
rect 9259 9691 9325 9692
rect 9741 9280 10061 10304
rect 9741 9216 9749 9280
rect 9813 9216 9829 9280
rect 9893 9216 9909 9280
rect 9973 9216 9989 9280
rect 10053 9216 10061 9280
rect 9741 8192 10061 9216
rect 9741 8128 9749 8192
rect 9813 8128 9829 8192
rect 9893 8128 9909 8192
rect 9973 8128 9989 8192
rect 10053 8128 10061 8192
rect 9741 7104 10061 8128
rect 9741 7040 9749 7104
rect 9813 7040 9829 7104
rect 9893 7040 9909 7104
rect 9973 7040 9989 7104
rect 10053 7040 10061 7104
rect 9741 6016 10061 7040
rect 9741 5952 9749 6016
rect 9813 5952 9829 6016
rect 9893 5952 9909 6016
rect 9973 5952 9989 6016
rect 10053 5952 10061 6016
rect 9741 4928 10061 5952
rect 9741 4864 9749 4928
rect 9813 4864 9829 4928
rect 9893 4864 9909 4928
rect 9973 4864 9989 4928
rect 10053 4864 10061 4928
rect 9741 3840 10061 4864
rect 9741 3776 9749 3840
rect 9813 3776 9829 3840
rect 9893 3776 9909 3840
rect 9973 3776 9989 3840
rect 10053 3776 10061 3840
rect 9741 2752 10061 3776
rect 9741 2688 9749 2752
rect 9813 2688 9829 2752
rect 9893 2688 9909 2752
rect 9973 2688 9989 2752
rect 10053 2688 10061 2752
rect 8891 2276 8957 2277
rect 8891 2212 8892 2276
rect 8956 2212 8957 2276
rect 8891 2211 8957 2212
rect 9741 1664 10061 2688
rect 10366 2549 10426 11051
rect 10363 2548 10429 2549
rect 10363 2484 10364 2548
rect 10428 2484 10429 2548
rect 10363 2483 10429 2484
rect 9741 1600 9749 1664
rect 9813 1600 9829 1664
rect 9893 1600 9909 1664
rect 9973 1600 9989 1664
rect 10053 1600 10061 1664
rect 8707 1324 8773 1325
rect 8707 1260 8708 1324
rect 8772 1260 8773 1324
rect 8707 1259 8773 1260
rect 8339 1188 8405 1189
rect 8339 1124 8340 1188
rect 8404 1124 8405 1188
rect 8339 1123 8405 1124
rect 6808 1056 6816 1120
rect 6880 1056 6896 1120
rect 6960 1056 6976 1120
rect 7040 1056 7056 1120
rect 7120 1056 7128 1120
rect 6808 1040 7128 1056
rect 9741 1040 10061 1600
rect 10550 781 10610 22203
rect 10734 11525 10794 26827
rect 10918 23085 10978 41379
rect 11467 38724 11533 38725
rect 11467 38660 11468 38724
rect 11532 38660 11533 38724
rect 11467 38659 11533 38660
rect 11099 32332 11165 32333
rect 11099 32268 11100 32332
rect 11164 32268 11165 32332
rect 11099 32267 11165 32268
rect 10915 23084 10981 23085
rect 10915 23020 10916 23084
rect 10980 23020 10981 23084
rect 10915 23019 10981 23020
rect 10915 16556 10981 16557
rect 10915 16492 10916 16556
rect 10980 16492 10981 16556
rect 10915 16491 10981 16492
rect 10731 11524 10797 11525
rect 10731 11460 10732 11524
rect 10796 11460 10797 11524
rect 10731 11459 10797 11460
rect 10918 4045 10978 16491
rect 10915 4044 10981 4045
rect 10915 3980 10916 4044
rect 10980 3980 10981 4044
rect 10915 3979 10981 3980
rect 11102 1325 11162 32267
rect 11470 30429 11530 38659
rect 11467 30428 11533 30429
rect 11467 30364 11468 30428
rect 11532 30364 11533 30428
rect 11467 30363 11533 30364
rect 11283 26620 11349 26621
rect 11283 26556 11284 26620
rect 11348 26556 11349 26620
rect 11283 26555 11349 26556
rect 11286 23629 11346 26555
rect 11283 23628 11349 23629
rect 11283 23564 11284 23628
rect 11348 23564 11349 23628
rect 11283 23563 11349 23564
rect 11286 21045 11346 23563
rect 11283 21044 11349 21045
rect 11283 20980 11284 21044
rect 11348 20980 11349 21044
rect 11283 20979 11349 20980
rect 11654 5541 11714 43011
rect 11835 42940 11901 42941
rect 11835 42876 11836 42940
rect 11900 42876 11901 42940
rect 11835 42875 11901 42876
rect 11838 11117 11898 42875
rect 12673 42464 12993 43488
rect 15606 43008 15926 43568
rect 15606 42944 15614 43008
rect 15678 42944 15694 43008
rect 15758 42944 15774 43008
rect 15838 42944 15854 43008
rect 15918 42944 15926 43008
rect 14963 42940 15029 42941
rect 14963 42876 14964 42940
rect 15028 42876 15029 42940
rect 14963 42875 15029 42876
rect 15331 42940 15397 42941
rect 15331 42876 15332 42940
rect 15396 42876 15397 42940
rect 15331 42875 15397 42876
rect 12673 42400 12681 42464
rect 12745 42400 12761 42464
rect 12825 42400 12841 42464
rect 12905 42400 12921 42464
rect 12985 42400 12993 42464
rect 12673 41376 12993 42400
rect 12673 41312 12681 41376
rect 12745 41312 12761 41376
rect 12825 41312 12841 41376
rect 12905 41312 12921 41376
rect 12985 41312 12993 41376
rect 12673 40288 12993 41312
rect 12673 40224 12681 40288
rect 12745 40224 12761 40288
rect 12825 40224 12841 40288
rect 12905 40224 12921 40288
rect 12985 40224 12993 40288
rect 12673 39200 12993 40224
rect 13307 39948 13373 39949
rect 13307 39884 13308 39948
rect 13372 39884 13373 39948
rect 13307 39883 13373 39884
rect 12673 39136 12681 39200
rect 12745 39136 12761 39200
rect 12825 39136 12841 39200
rect 12905 39136 12921 39200
rect 12985 39136 12993 39200
rect 12673 38112 12993 39136
rect 12673 38048 12681 38112
rect 12745 38048 12761 38112
rect 12825 38048 12841 38112
rect 12905 38048 12921 38112
rect 12985 38048 12993 38112
rect 12673 37024 12993 38048
rect 12673 36960 12681 37024
rect 12745 36960 12761 37024
rect 12825 36960 12841 37024
rect 12905 36960 12921 37024
rect 12985 36960 12993 37024
rect 12673 35936 12993 36960
rect 12673 35872 12681 35936
rect 12745 35872 12761 35936
rect 12825 35872 12841 35936
rect 12905 35872 12921 35936
rect 12985 35872 12993 35936
rect 12673 34848 12993 35872
rect 12673 34784 12681 34848
rect 12745 34784 12761 34848
rect 12825 34784 12841 34848
rect 12905 34784 12921 34848
rect 12985 34784 12993 34848
rect 12673 33760 12993 34784
rect 12673 33696 12681 33760
rect 12745 33696 12761 33760
rect 12825 33696 12841 33760
rect 12905 33696 12921 33760
rect 12985 33696 12993 33760
rect 12673 32672 12993 33696
rect 12673 32608 12681 32672
rect 12745 32608 12761 32672
rect 12825 32608 12841 32672
rect 12905 32608 12921 32672
rect 12985 32608 12993 32672
rect 12673 31584 12993 32608
rect 12673 31520 12681 31584
rect 12745 31520 12761 31584
rect 12825 31520 12841 31584
rect 12905 31520 12921 31584
rect 12985 31520 12993 31584
rect 12673 30496 12993 31520
rect 12673 30432 12681 30496
rect 12745 30432 12761 30496
rect 12825 30432 12841 30496
rect 12905 30432 12921 30496
rect 12985 30432 12993 30496
rect 12019 30428 12085 30429
rect 12019 30364 12020 30428
rect 12084 30364 12085 30428
rect 12019 30363 12085 30364
rect 11835 11116 11901 11117
rect 11835 11052 11836 11116
rect 11900 11052 11901 11116
rect 11835 11051 11901 11052
rect 11651 5540 11717 5541
rect 11651 5476 11652 5540
rect 11716 5476 11717 5540
rect 11651 5475 11717 5476
rect 12022 2413 12082 30363
rect 12673 29408 12993 30432
rect 12673 29344 12681 29408
rect 12745 29344 12761 29408
rect 12825 29344 12841 29408
rect 12905 29344 12921 29408
rect 12985 29344 12993 29408
rect 12673 28320 12993 29344
rect 13123 29068 13189 29069
rect 13123 29004 13124 29068
rect 13188 29004 13189 29068
rect 13123 29003 13189 29004
rect 12673 28256 12681 28320
rect 12745 28256 12761 28320
rect 12825 28256 12841 28320
rect 12905 28256 12921 28320
rect 12985 28256 12993 28320
rect 12673 27232 12993 28256
rect 12673 27168 12681 27232
rect 12745 27168 12761 27232
rect 12825 27168 12841 27232
rect 12905 27168 12921 27232
rect 12985 27168 12993 27232
rect 12673 26144 12993 27168
rect 12673 26080 12681 26144
rect 12745 26080 12761 26144
rect 12825 26080 12841 26144
rect 12905 26080 12921 26144
rect 12985 26080 12993 26144
rect 12673 25056 12993 26080
rect 12673 24992 12681 25056
rect 12745 24992 12761 25056
rect 12825 24992 12841 25056
rect 12905 24992 12921 25056
rect 12985 24992 12993 25056
rect 12673 23968 12993 24992
rect 12673 23904 12681 23968
rect 12745 23904 12761 23968
rect 12825 23904 12841 23968
rect 12905 23904 12921 23968
rect 12985 23904 12993 23968
rect 12673 22880 12993 23904
rect 12673 22816 12681 22880
rect 12745 22816 12761 22880
rect 12825 22816 12841 22880
rect 12905 22816 12921 22880
rect 12985 22816 12993 22880
rect 12387 22132 12453 22133
rect 12387 22068 12388 22132
rect 12452 22068 12453 22132
rect 12387 22067 12453 22068
rect 12390 21997 12450 22067
rect 12387 21996 12453 21997
rect 12387 21932 12388 21996
rect 12452 21932 12453 21996
rect 12387 21931 12453 21932
rect 12673 21792 12993 22816
rect 13126 22133 13186 29003
rect 13310 22269 13370 39883
rect 13675 37364 13741 37365
rect 13675 37300 13676 37364
rect 13740 37300 13741 37364
rect 13675 37299 13741 37300
rect 13307 22268 13373 22269
rect 13307 22204 13308 22268
rect 13372 22204 13373 22268
rect 13307 22203 13373 22204
rect 13123 22132 13189 22133
rect 13123 22068 13124 22132
rect 13188 22068 13189 22132
rect 13123 22067 13189 22068
rect 13491 22132 13557 22133
rect 13491 22068 13492 22132
rect 13556 22068 13557 22132
rect 13491 22067 13557 22068
rect 13123 21996 13189 21997
rect 13123 21932 13124 21996
rect 13188 21932 13189 21996
rect 13123 21931 13189 21932
rect 12673 21728 12681 21792
rect 12745 21728 12761 21792
rect 12825 21728 12841 21792
rect 12905 21728 12921 21792
rect 12985 21728 12993 21792
rect 12673 20704 12993 21728
rect 12673 20640 12681 20704
rect 12745 20640 12761 20704
rect 12825 20640 12841 20704
rect 12905 20640 12921 20704
rect 12985 20640 12993 20704
rect 12673 19616 12993 20640
rect 12673 19552 12681 19616
rect 12745 19552 12761 19616
rect 12825 19552 12841 19616
rect 12905 19552 12921 19616
rect 12985 19552 12993 19616
rect 12673 18528 12993 19552
rect 12673 18464 12681 18528
rect 12745 18464 12761 18528
rect 12825 18464 12841 18528
rect 12905 18464 12921 18528
rect 12985 18464 12993 18528
rect 12673 17440 12993 18464
rect 12673 17376 12681 17440
rect 12745 17376 12761 17440
rect 12825 17376 12841 17440
rect 12905 17376 12921 17440
rect 12985 17376 12993 17440
rect 12673 16352 12993 17376
rect 12673 16288 12681 16352
rect 12745 16288 12761 16352
rect 12825 16288 12841 16352
rect 12905 16288 12921 16352
rect 12985 16288 12993 16352
rect 12673 15264 12993 16288
rect 12673 15200 12681 15264
rect 12745 15200 12761 15264
rect 12825 15200 12841 15264
rect 12905 15200 12921 15264
rect 12985 15200 12993 15264
rect 12673 14176 12993 15200
rect 12673 14112 12681 14176
rect 12745 14112 12761 14176
rect 12825 14112 12841 14176
rect 12905 14112 12921 14176
rect 12985 14112 12993 14176
rect 12673 13088 12993 14112
rect 12673 13024 12681 13088
rect 12745 13024 12761 13088
rect 12825 13024 12841 13088
rect 12905 13024 12921 13088
rect 12985 13024 12993 13088
rect 12387 12748 12453 12749
rect 12387 12684 12388 12748
rect 12452 12684 12453 12748
rect 12387 12683 12453 12684
rect 12390 12205 12450 12683
rect 12387 12204 12453 12205
rect 12387 12140 12388 12204
rect 12452 12140 12453 12204
rect 12387 12139 12453 12140
rect 12673 12000 12993 13024
rect 13126 12749 13186 21931
rect 13307 20772 13373 20773
rect 13307 20708 13308 20772
rect 13372 20708 13373 20772
rect 13307 20707 13373 20708
rect 13123 12748 13189 12749
rect 13123 12684 13124 12748
rect 13188 12684 13189 12748
rect 13123 12683 13189 12684
rect 13123 12204 13189 12205
rect 13123 12140 13124 12204
rect 13188 12140 13189 12204
rect 13123 12139 13189 12140
rect 12673 11936 12681 12000
rect 12745 11936 12761 12000
rect 12825 11936 12841 12000
rect 12905 11936 12921 12000
rect 12985 11936 12993 12000
rect 12673 10912 12993 11936
rect 12673 10848 12681 10912
rect 12745 10848 12761 10912
rect 12825 10848 12841 10912
rect 12905 10848 12921 10912
rect 12985 10848 12993 10912
rect 12673 9824 12993 10848
rect 12673 9760 12681 9824
rect 12745 9760 12761 9824
rect 12825 9760 12841 9824
rect 12905 9760 12921 9824
rect 12985 9760 12993 9824
rect 12673 8736 12993 9760
rect 12673 8672 12681 8736
rect 12745 8672 12761 8736
rect 12825 8672 12841 8736
rect 12905 8672 12921 8736
rect 12985 8672 12993 8736
rect 12673 7648 12993 8672
rect 12673 7584 12681 7648
rect 12745 7584 12761 7648
rect 12825 7584 12841 7648
rect 12905 7584 12921 7648
rect 12985 7584 12993 7648
rect 12673 6560 12993 7584
rect 12673 6496 12681 6560
rect 12745 6496 12761 6560
rect 12825 6496 12841 6560
rect 12905 6496 12921 6560
rect 12985 6496 12993 6560
rect 12673 5472 12993 6496
rect 12673 5408 12681 5472
rect 12745 5408 12761 5472
rect 12825 5408 12841 5472
rect 12905 5408 12921 5472
rect 12985 5408 12993 5472
rect 12673 4384 12993 5408
rect 12673 4320 12681 4384
rect 12745 4320 12761 4384
rect 12825 4320 12841 4384
rect 12905 4320 12921 4384
rect 12985 4320 12993 4384
rect 12673 3296 12993 4320
rect 12673 3232 12681 3296
rect 12745 3232 12761 3296
rect 12825 3232 12841 3296
rect 12905 3232 12921 3296
rect 12985 3232 12993 3296
rect 12387 3092 12453 3093
rect 12387 3028 12388 3092
rect 12452 3028 12453 3092
rect 12387 3027 12453 3028
rect 12019 2412 12085 2413
rect 12019 2348 12020 2412
rect 12084 2348 12085 2412
rect 12019 2347 12085 2348
rect 12390 1325 12450 3027
rect 12673 2208 12993 3232
rect 13126 3093 13186 12139
rect 13123 3092 13189 3093
rect 13123 3028 13124 3092
rect 13188 3028 13189 3092
rect 13123 3027 13189 3028
rect 13310 2685 13370 20707
rect 13307 2684 13373 2685
rect 13307 2620 13308 2684
rect 13372 2620 13373 2684
rect 13307 2619 13373 2620
rect 12673 2144 12681 2208
rect 12745 2144 12761 2208
rect 12825 2144 12841 2208
rect 12905 2144 12921 2208
rect 12985 2144 12993 2208
rect 11099 1324 11165 1325
rect 11099 1260 11100 1324
rect 11164 1260 11165 1324
rect 11099 1259 11165 1260
rect 12387 1324 12453 1325
rect 12387 1260 12388 1324
rect 12452 1260 12453 1324
rect 12387 1259 12453 1260
rect 12673 1120 12993 2144
rect 13494 1325 13554 22067
rect 13678 20773 13738 37299
rect 14043 28524 14109 28525
rect 14043 28460 14044 28524
rect 14108 28460 14109 28524
rect 14043 28459 14109 28460
rect 14046 26621 14106 28459
rect 14043 26620 14109 26621
rect 14043 26556 14044 26620
rect 14108 26556 14109 26620
rect 14043 26555 14109 26556
rect 14779 26620 14845 26621
rect 14779 26556 14780 26620
rect 14844 26556 14845 26620
rect 14779 26555 14845 26556
rect 14227 23492 14293 23493
rect 14227 23428 14228 23492
rect 14292 23428 14293 23492
rect 14227 23427 14293 23428
rect 13675 20772 13741 20773
rect 13675 20708 13676 20772
rect 13740 20708 13741 20772
rect 13675 20707 13741 20708
rect 13859 17780 13925 17781
rect 13859 17716 13860 17780
rect 13924 17716 13925 17780
rect 13859 17715 13925 17716
rect 13862 12341 13922 17715
rect 13859 12340 13925 12341
rect 13859 12276 13860 12340
rect 13924 12276 13925 12340
rect 13859 12275 13925 12276
rect 13862 11661 13922 12275
rect 13859 11660 13925 11661
rect 13859 11596 13860 11660
rect 13924 11596 13925 11660
rect 13859 11595 13925 11596
rect 14230 1325 14290 23427
rect 14411 22676 14477 22677
rect 14411 22612 14412 22676
rect 14476 22612 14477 22676
rect 14411 22611 14477 22612
rect 14414 20637 14474 22611
rect 14595 20772 14661 20773
rect 14595 20708 14596 20772
rect 14660 20708 14661 20772
rect 14595 20707 14661 20708
rect 14411 20636 14477 20637
rect 14411 20572 14412 20636
rect 14476 20572 14477 20636
rect 14411 20571 14477 20572
rect 14411 11116 14477 11117
rect 14411 11052 14412 11116
rect 14476 11052 14477 11116
rect 14411 11051 14477 11052
rect 14414 2141 14474 11051
rect 14411 2140 14477 2141
rect 14411 2076 14412 2140
rect 14476 2076 14477 2140
rect 14411 2075 14477 2076
rect 14598 1325 14658 20707
rect 14782 15469 14842 26555
rect 14966 20501 15026 42875
rect 15147 31924 15213 31925
rect 15147 31860 15148 31924
rect 15212 31860 15213 31924
rect 15147 31859 15213 31860
rect 15150 28117 15210 31859
rect 15147 28116 15213 28117
rect 15147 28052 15148 28116
rect 15212 28052 15213 28116
rect 15147 28051 15213 28052
rect 14963 20500 15029 20501
rect 14963 20436 14964 20500
rect 15028 20436 15029 20500
rect 14963 20435 15029 20436
rect 14963 20228 15029 20229
rect 14963 20164 14964 20228
rect 15028 20164 15029 20228
rect 14963 20163 15029 20164
rect 14966 16149 15026 20163
rect 15147 19412 15213 19413
rect 15147 19348 15148 19412
rect 15212 19348 15213 19412
rect 15147 19347 15213 19348
rect 14963 16148 15029 16149
rect 14963 16084 14964 16148
rect 15028 16084 15029 16148
rect 14963 16083 15029 16084
rect 14779 15468 14845 15469
rect 14779 15404 14780 15468
rect 14844 15404 14845 15468
rect 14779 15403 14845 15404
rect 15150 1325 15210 19347
rect 15334 2549 15394 42875
rect 15606 41920 15926 42944
rect 18538 43552 18858 43568
rect 18538 43488 18546 43552
rect 18610 43488 18626 43552
rect 18690 43488 18706 43552
rect 18770 43488 18786 43552
rect 18850 43488 18858 43552
rect 17723 42940 17789 42941
rect 17723 42876 17724 42940
rect 17788 42876 17789 42940
rect 17723 42875 17789 42876
rect 16619 42668 16685 42669
rect 16619 42604 16620 42668
rect 16684 42604 16685 42668
rect 16619 42603 16685 42604
rect 15606 41856 15614 41920
rect 15678 41856 15694 41920
rect 15758 41856 15774 41920
rect 15838 41856 15854 41920
rect 15918 41856 15926 41920
rect 15606 40832 15926 41856
rect 15606 40768 15614 40832
rect 15678 40768 15694 40832
rect 15758 40768 15774 40832
rect 15838 40768 15854 40832
rect 15918 40768 15926 40832
rect 15606 39744 15926 40768
rect 15606 39680 15614 39744
rect 15678 39680 15694 39744
rect 15758 39680 15774 39744
rect 15838 39680 15854 39744
rect 15918 39680 15926 39744
rect 15606 38656 15926 39680
rect 15606 38592 15614 38656
rect 15678 38592 15694 38656
rect 15758 38592 15774 38656
rect 15838 38592 15854 38656
rect 15918 38592 15926 38656
rect 15606 37568 15926 38592
rect 15606 37504 15614 37568
rect 15678 37504 15694 37568
rect 15758 37504 15774 37568
rect 15838 37504 15854 37568
rect 15918 37504 15926 37568
rect 15606 36480 15926 37504
rect 15606 36416 15614 36480
rect 15678 36416 15694 36480
rect 15758 36416 15774 36480
rect 15838 36416 15854 36480
rect 15918 36416 15926 36480
rect 15606 35392 15926 36416
rect 15606 35328 15614 35392
rect 15678 35328 15694 35392
rect 15758 35328 15774 35392
rect 15838 35328 15854 35392
rect 15918 35328 15926 35392
rect 15606 34304 15926 35328
rect 15606 34240 15614 34304
rect 15678 34240 15694 34304
rect 15758 34240 15774 34304
rect 15838 34240 15854 34304
rect 15918 34240 15926 34304
rect 15606 33216 15926 34240
rect 15606 33152 15614 33216
rect 15678 33152 15694 33216
rect 15758 33152 15774 33216
rect 15838 33152 15854 33216
rect 15918 33152 15926 33216
rect 15606 32128 15926 33152
rect 15606 32064 15614 32128
rect 15678 32064 15694 32128
rect 15758 32064 15774 32128
rect 15838 32064 15854 32128
rect 15918 32064 15926 32128
rect 15606 31040 15926 32064
rect 15606 30976 15614 31040
rect 15678 30976 15694 31040
rect 15758 30976 15774 31040
rect 15838 30976 15854 31040
rect 15918 30976 15926 31040
rect 15606 29952 15926 30976
rect 15606 29888 15614 29952
rect 15678 29888 15694 29952
rect 15758 29888 15774 29952
rect 15838 29888 15854 29952
rect 15918 29888 15926 29952
rect 15606 28864 15926 29888
rect 16435 29612 16501 29613
rect 16435 29548 16436 29612
rect 16500 29548 16501 29612
rect 16435 29547 16501 29548
rect 15606 28800 15614 28864
rect 15678 28800 15694 28864
rect 15758 28800 15774 28864
rect 15838 28800 15854 28864
rect 15918 28800 15926 28864
rect 15606 27776 15926 28800
rect 16251 28116 16317 28117
rect 16251 28052 16252 28116
rect 16316 28052 16317 28116
rect 16251 28051 16317 28052
rect 15606 27712 15614 27776
rect 15678 27712 15694 27776
rect 15758 27712 15774 27776
rect 15838 27712 15854 27776
rect 15918 27712 15926 27776
rect 15606 26688 15926 27712
rect 15606 26624 15614 26688
rect 15678 26624 15694 26688
rect 15758 26624 15774 26688
rect 15838 26624 15854 26688
rect 15918 26624 15926 26688
rect 15606 25600 15926 26624
rect 15606 25536 15614 25600
rect 15678 25536 15694 25600
rect 15758 25536 15774 25600
rect 15838 25536 15854 25600
rect 15918 25536 15926 25600
rect 15606 24512 15926 25536
rect 15606 24448 15614 24512
rect 15678 24448 15694 24512
rect 15758 24448 15774 24512
rect 15838 24448 15854 24512
rect 15918 24448 15926 24512
rect 15606 23424 15926 24448
rect 15606 23360 15614 23424
rect 15678 23360 15694 23424
rect 15758 23360 15774 23424
rect 15838 23360 15854 23424
rect 15918 23360 15926 23424
rect 15606 22336 15926 23360
rect 15606 22272 15614 22336
rect 15678 22272 15694 22336
rect 15758 22272 15774 22336
rect 15838 22272 15854 22336
rect 15918 22272 15926 22336
rect 15606 21248 15926 22272
rect 15606 21184 15614 21248
rect 15678 21184 15694 21248
rect 15758 21184 15774 21248
rect 15838 21184 15854 21248
rect 15918 21184 15926 21248
rect 15606 20160 15926 21184
rect 15606 20096 15614 20160
rect 15678 20096 15694 20160
rect 15758 20096 15774 20160
rect 15838 20096 15854 20160
rect 15918 20096 15926 20160
rect 15606 19072 15926 20096
rect 15606 19008 15614 19072
rect 15678 19008 15694 19072
rect 15758 19008 15774 19072
rect 15838 19008 15854 19072
rect 15918 19008 15926 19072
rect 15606 17984 15926 19008
rect 15606 17920 15614 17984
rect 15678 17920 15694 17984
rect 15758 17920 15774 17984
rect 15838 17920 15854 17984
rect 15918 17920 15926 17984
rect 15606 16896 15926 17920
rect 16254 17781 16314 28051
rect 16438 19413 16498 29547
rect 16435 19412 16501 19413
rect 16435 19348 16436 19412
rect 16500 19348 16501 19412
rect 16435 19347 16501 19348
rect 16251 17780 16317 17781
rect 16251 17716 16252 17780
rect 16316 17716 16317 17780
rect 16251 17715 16317 17716
rect 15606 16832 15614 16896
rect 15678 16832 15694 16896
rect 15758 16832 15774 16896
rect 15838 16832 15854 16896
rect 15918 16832 15926 16896
rect 15606 15808 15926 16832
rect 15606 15744 15614 15808
rect 15678 15744 15694 15808
rect 15758 15744 15774 15808
rect 15838 15744 15854 15808
rect 15918 15744 15926 15808
rect 15606 14720 15926 15744
rect 15606 14656 15614 14720
rect 15678 14656 15694 14720
rect 15758 14656 15774 14720
rect 15838 14656 15854 14720
rect 15918 14656 15926 14720
rect 15606 13632 15926 14656
rect 15606 13568 15614 13632
rect 15678 13568 15694 13632
rect 15758 13568 15774 13632
rect 15838 13568 15854 13632
rect 15918 13568 15926 13632
rect 15606 12544 15926 13568
rect 15606 12480 15614 12544
rect 15678 12480 15694 12544
rect 15758 12480 15774 12544
rect 15838 12480 15854 12544
rect 15918 12480 15926 12544
rect 15606 11456 15926 12480
rect 15606 11392 15614 11456
rect 15678 11392 15694 11456
rect 15758 11392 15774 11456
rect 15838 11392 15854 11456
rect 15918 11392 15926 11456
rect 15606 10368 15926 11392
rect 15606 10304 15614 10368
rect 15678 10304 15694 10368
rect 15758 10304 15774 10368
rect 15838 10304 15854 10368
rect 15918 10304 15926 10368
rect 15606 9280 15926 10304
rect 15606 9216 15614 9280
rect 15678 9216 15694 9280
rect 15758 9216 15774 9280
rect 15838 9216 15854 9280
rect 15918 9216 15926 9280
rect 15606 8192 15926 9216
rect 15606 8128 15614 8192
rect 15678 8128 15694 8192
rect 15758 8128 15774 8192
rect 15838 8128 15854 8192
rect 15918 8128 15926 8192
rect 15606 7104 15926 8128
rect 15606 7040 15614 7104
rect 15678 7040 15694 7104
rect 15758 7040 15774 7104
rect 15838 7040 15854 7104
rect 15918 7040 15926 7104
rect 15606 6016 15926 7040
rect 15606 5952 15614 6016
rect 15678 5952 15694 6016
rect 15758 5952 15774 6016
rect 15838 5952 15854 6016
rect 15918 5952 15926 6016
rect 15606 4928 15926 5952
rect 16622 5133 16682 42603
rect 16987 42124 17053 42125
rect 16987 42060 16988 42124
rect 17052 42060 17053 42124
rect 16987 42059 17053 42060
rect 16619 5132 16685 5133
rect 16619 5068 16620 5132
rect 16684 5068 16685 5132
rect 16619 5067 16685 5068
rect 15606 4864 15614 4928
rect 15678 4864 15694 4928
rect 15758 4864 15774 4928
rect 15838 4864 15854 4928
rect 15918 4864 15926 4928
rect 15606 3840 15926 4864
rect 15606 3776 15614 3840
rect 15678 3776 15694 3840
rect 15758 3776 15774 3840
rect 15838 3776 15854 3840
rect 15918 3776 15926 3840
rect 15606 2752 15926 3776
rect 15606 2688 15614 2752
rect 15678 2688 15694 2752
rect 15758 2688 15774 2752
rect 15838 2688 15854 2752
rect 15918 2688 15926 2752
rect 15331 2548 15397 2549
rect 15331 2484 15332 2548
rect 15396 2484 15397 2548
rect 15331 2483 15397 2484
rect 15606 1664 15926 2688
rect 16990 2685 17050 42059
rect 17171 41988 17237 41989
rect 17171 41924 17172 41988
rect 17236 41924 17237 41988
rect 17171 41923 17237 41924
rect 17174 2685 17234 41923
rect 17726 15197 17786 42875
rect 18538 42464 18858 43488
rect 18538 42400 18546 42464
rect 18610 42400 18626 42464
rect 18690 42400 18706 42464
rect 18770 42400 18786 42464
rect 18850 42400 18858 42464
rect 18275 41988 18341 41989
rect 18275 41924 18276 41988
rect 18340 41924 18341 41988
rect 18275 41923 18341 41924
rect 17907 35052 17973 35053
rect 17907 34988 17908 35052
rect 17972 34988 17973 35052
rect 17907 34987 17973 34988
rect 17723 15196 17789 15197
rect 17723 15132 17724 15196
rect 17788 15132 17789 15196
rect 17723 15131 17789 15132
rect 17910 8397 17970 34987
rect 18091 29204 18157 29205
rect 18091 29140 18092 29204
rect 18156 29140 18157 29204
rect 18091 29139 18157 29140
rect 18094 19413 18154 29139
rect 18091 19412 18157 19413
rect 18091 19348 18092 19412
rect 18156 19348 18157 19412
rect 18091 19347 18157 19348
rect 17907 8396 17973 8397
rect 17907 8332 17908 8396
rect 17972 8332 17973 8396
rect 17907 8331 17973 8332
rect 18278 5541 18338 41923
rect 18538 41376 18858 42400
rect 21471 43008 21791 43568
rect 24403 43552 24723 43568
rect 24403 43488 24411 43552
rect 24475 43488 24491 43552
rect 24555 43488 24571 43552
rect 24635 43488 24651 43552
rect 24715 43488 24723 43552
rect 21955 43212 22021 43213
rect 21955 43148 21956 43212
rect 22020 43148 22021 43212
rect 21955 43147 22021 43148
rect 21471 42944 21479 43008
rect 21543 42944 21559 43008
rect 21623 42944 21639 43008
rect 21703 42944 21719 43008
rect 21783 42944 21791 43008
rect 19563 41988 19629 41989
rect 19563 41924 19564 41988
rect 19628 41924 19629 41988
rect 19563 41923 19629 41924
rect 19931 41988 19997 41989
rect 19931 41924 19932 41988
rect 19996 41924 19997 41988
rect 19931 41923 19997 41924
rect 18538 41312 18546 41376
rect 18610 41312 18626 41376
rect 18690 41312 18706 41376
rect 18770 41312 18786 41376
rect 18850 41312 18858 41376
rect 18538 40288 18858 41312
rect 18538 40224 18546 40288
rect 18610 40224 18626 40288
rect 18690 40224 18706 40288
rect 18770 40224 18786 40288
rect 18850 40224 18858 40288
rect 18538 39200 18858 40224
rect 19379 39540 19445 39541
rect 19379 39476 19380 39540
rect 19444 39476 19445 39540
rect 19379 39475 19445 39476
rect 18538 39136 18546 39200
rect 18610 39136 18626 39200
rect 18690 39136 18706 39200
rect 18770 39136 18786 39200
rect 18850 39136 18858 39200
rect 18538 38112 18858 39136
rect 18538 38048 18546 38112
rect 18610 38048 18626 38112
rect 18690 38048 18706 38112
rect 18770 38048 18786 38112
rect 18850 38048 18858 38112
rect 18538 37024 18858 38048
rect 18538 36960 18546 37024
rect 18610 36960 18626 37024
rect 18690 36960 18706 37024
rect 18770 36960 18786 37024
rect 18850 36960 18858 37024
rect 18538 35936 18858 36960
rect 18538 35872 18546 35936
rect 18610 35872 18626 35936
rect 18690 35872 18706 35936
rect 18770 35872 18786 35936
rect 18850 35872 18858 35936
rect 18538 34848 18858 35872
rect 18538 34784 18546 34848
rect 18610 34784 18626 34848
rect 18690 34784 18706 34848
rect 18770 34784 18786 34848
rect 18850 34784 18858 34848
rect 18538 33760 18858 34784
rect 18538 33696 18546 33760
rect 18610 33696 18626 33760
rect 18690 33696 18706 33760
rect 18770 33696 18786 33760
rect 18850 33696 18858 33760
rect 18538 32672 18858 33696
rect 18538 32608 18546 32672
rect 18610 32608 18626 32672
rect 18690 32608 18706 32672
rect 18770 32608 18786 32672
rect 18850 32608 18858 32672
rect 18538 31584 18858 32608
rect 18538 31520 18546 31584
rect 18610 31520 18626 31584
rect 18690 31520 18706 31584
rect 18770 31520 18786 31584
rect 18850 31520 18858 31584
rect 18538 30496 18858 31520
rect 18538 30432 18546 30496
rect 18610 30432 18626 30496
rect 18690 30432 18706 30496
rect 18770 30432 18786 30496
rect 18850 30432 18858 30496
rect 18538 29408 18858 30432
rect 18538 29344 18546 29408
rect 18610 29344 18626 29408
rect 18690 29344 18706 29408
rect 18770 29344 18786 29408
rect 18850 29344 18858 29408
rect 18538 28320 18858 29344
rect 18538 28256 18546 28320
rect 18610 28256 18626 28320
rect 18690 28256 18706 28320
rect 18770 28256 18786 28320
rect 18850 28256 18858 28320
rect 18538 27232 18858 28256
rect 18538 27168 18546 27232
rect 18610 27168 18626 27232
rect 18690 27168 18706 27232
rect 18770 27168 18786 27232
rect 18850 27168 18858 27232
rect 18538 26144 18858 27168
rect 18538 26080 18546 26144
rect 18610 26080 18626 26144
rect 18690 26080 18706 26144
rect 18770 26080 18786 26144
rect 18850 26080 18858 26144
rect 18538 25056 18858 26080
rect 18538 24992 18546 25056
rect 18610 24992 18626 25056
rect 18690 24992 18706 25056
rect 18770 24992 18786 25056
rect 18850 24992 18858 25056
rect 18538 23968 18858 24992
rect 18538 23904 18546 23968
rect 18610 23904 18626 23968
rect 18690 23904 18706 23968
rect 18770 23904 18786 23968
rect 18850 23904 18858 23968
rect 18538 22880 18858 23904
rect 18538 22816 18546 22880
rect 18610 22816 18626 22880
rect 18690 22816 18706 22880
rect 18770 22816 18786 22880
rect 18850 22816 18858 22880
rect 18538 21792 18858 22816
rect 18538 21728 18546 21792
rect 18610 21728 18626 21792
rect 18690 21728 18706 21792
rect 18770 21728 18786 21792
rect 18850 21728 18858 21792
rect 18538 20704 18858 21728
rect 18538 20640 18546 20704
rect 18610 20640 18626 20704
rect 18690 20640 18706 20704
rect 18770 20640 18786 20704
rect 18850 20640 18858 20704
rect 18538 19616 18858 20640
rect 18538 19552 18546 19616
rect 18610 19552 18626 19616
rect 18690 19552 18706 19616
rect 18770 19552 18786 19616
rect 18850 19552 18858 19616
rect 18538 18528 18858 19552
rect 18538 18464 18546 18528
rect 18610 18464 18626 18528
rect 18690 18464 18706 18528
rect 18770 18464 18786 18528
rect 18850 18464 18858 18528
rect 18538 17440 18858 18464
rect 18538 17376 18546 17440
rect 18610 17376 18626 17440
rect 18690 17376 18706 17440
rect 18770 17376 18786 17440
rect 18850 17376 18858 17440
rect 18538 16352 18858 17376
rect 18538 16288 18546 16352
rect 18610 16288 18626 16352
rect 18690 16288 18706 16352
rect 18770 16288 18786 16352
rect 18850 16288 18858 16352
rect 18538 15264 18858 16288
rect 18538 15200 18546 15264
rect 18610 15200 18626 15264
rect 18690 15200 18706 15264
rect 18770 15200 18786 15264
rect 18850 15200 18858 15264
rect 18538 14176 18858 15200
rect 18538 14112 18546 14176
rect 18610 14112 18626 14176
rect 18690 14112 18706 14176
rect 18770 14112 18786 14176
rect 18850 14112 18858 14176
rect 18538 13088 18858 14112
rect 18538 13024 18546 13088
rect 18610 13024 18626 13088
rect 18690 13024 18706 13088
rect 18770 13024 18786 13088
rect 18850 13024 18858 13088
rect 18538 12000 18858 13024
rect 18538 11936 18546 12000
rect 18610 11936 18626 12000
rect 18690 11936 18706 12000
rect 18770 11936 18786 12000
rect 18850 11936 18858 12000
rect 18538 10912 18858 11936
rect 18538 10848 18546 10912
rect 18610 10848 18626 10912
rect 18690 10848 18706 10912
rect 18770 10848 18786 10912
rect 18850 10848 18858 10912
rect 18538 9824 18858 10848
rect 18538 9760 18546 9824
rect 18610 9760 18626 9824
rect 18690 9760 18706 9824
rect 18770 9760 18786 9824
rect 18850 9760 18858 9824
rect 18538 8736 18858 9760
rect 18538 8672 18546 8736
rect 18610 8672 18626 8736
rect 18690 8672 18706 8736
rect 18770 8672 18786 8736
rect 18850 8672 18858 8736
rect 18538 7648 18858 8672
rect 18538 7584 18546 7648
rect 18610 7584 18626 7648
rect 18690 7584 18706 7648
rect 18770 7584 18786 7648
rect 18850 7584 18858 7648
rect 18538 6560 18858 7584
rect 18538 6496 18546 6560
rect 18610 6496 18626 6560
rect 18690 6496 18706 6560
rect 18770 6496 18786 6560
rect 18850 6496 18858 6560
rect 18275 5540 18341 5541
rect 18275 5476 18276 5540
rect 18340 5476 18341 5540
rect 18275 5475 18341 5476
rect 18538 5472 18858 6496
rect 18538 5408 18546 5472
rect 18610 5408 18626 5472
rect 18690 5408 18706 5472
rect 18770 5408 18786 5472
rect 18850 5408 18858 5472
rect 18538 4384 18858 5408
rect 18538 4320 18546 4384
rect 18610 4320 18626 4384
rect 18690 4320 18706 4384
rect 18770 4320 18786 4384
rect 18850 4320 18858 4384
rect 18538 3296 18858 4320
rect 18538 3232 18546 3296
rect 18610 3232 18626 3296
rect 18690 3232 18706 3296
rect 18770 3232 18786 3296
rect 18850 3232 18858 3296
rect 16987 2684 17053 2685
rect 16987 2620 16988 2684
rect 17052 2620 17053 2684
rect 16987 2619 17053 2620
rect 17171 2684 17237 2685
rect 17171 2620 17172 2684
rect 17236 2620 17237 2684
rect 17171 2619 17237 2620
rect 15606 1600 15614 1664
rect 15678 1600 15694 1664
rect 15758 1600 15774 1664
rect 15838 1600 15854 1664
rect 15918 1600 15926 1664
rect 13491 1324 13557 1325
rect 13491 1260 13492 1324
rect 13556 1260 13557 1324
rect 13491 1259 13557 1260
rect 14227 1324 14293 1325
rect 14227 1260 14228 1324
rect 14292 1260 14293 1324
rect 14227 1259 14293 1260
rect 14595 1324 14661 1325
rect 14595 1260 14596 1324
rect 14660 1260 14661 1324
rect 14595 1259 14661 1260
rect 15147 1324 15213 1325
rect 15147 1260 15148 1324
rect 15212 1260 15213 1324
rect 15147 1259 15213 1260
rect 12673 1056 12681 1120
rect 12745 1056 12761 1120
rect 12825 1056 12841 1120
rect 12905 1056 12921 1120
rect 12985 1056 12993 1120
rect 12673 1040 12993 1056
rect 15606 1040 15926 1600
rect 18538 2208 18858 3232
rect 18538 2144 18546 2208
rect 18610 2144 18626 2208
rect 18690 2144 18706 2208
rect 18770 2144 18786 2208
rect 18850 2144 18858 2208
rect 18538 1120 18858 2144
rect 18538 1056 18546 1120
rect 18610 1056 18626 1120
rect 18690 1056 18706 1120
rect 18770 1056 18786 1120
rect 18850 1056 18858 1120
rect 18538 1040 18858 1056
rect 19382 917 19442 39475
rect 19566 31770 19626 41923
rect 19566 31710 19810 31770
rect 19563 12476 19629 12477
rect 19563 12412 19564 12476
rect 19628 12412 19629 12476
rect 19563 12411 19629 12412
rect 19566 12069 19626 12411
rect 19563 12068 19629 12069
rect 19563 12004 19564 12068
rect 19628 12004 19629 12068
rect 19563 12003 19629 12004
rect 19750 8533 19810 31710
rect 19747 8532 19813 8533
rect 19747 8468 19748 8532
rect 19812 8468 19813 8532
rect 19747 8467 19813 8468
rect 19934 8397 19994 41923
rect 21471 41920 21791 42944
rect 21471 41856 21479 41920
rect 21543 41856 21559 41920
rect 21623 41856 21639 41920
rect 21703 41856 21719 41920
rect 21783 41856 21791 41920
rect 21219 41580 21285 41581
rect 21219 41516 21220 41580
rect 21284 41516 21285 41580
rect 21219 41515 21285 41516
rect 21035 39404 21101 39405
rect 21035 39340 21036 39404
rect 21100 39340 21101 39404
rect 21035 39339 21101 39340
rect 20851 29068 20917 29069
rect 20851 29004 20852 29068
rect 20916 29004 20917 29068
rect 20851 29003 20917 29004
rect 20115 25940 20181 25941
rect 20115 25876 20116 25940
rect 20180 25876 20181 25940
rect 20115 25875 20181 25876
rect 19563 8396 19629 8397
rect 19563 8332 19564 8396
rect 19628 8332 19629 8396
rect 19563 8331 19629 8332
rect 19931 8396 19997 8397
rect 19931 8332 19932 8396
rect 19996 8332 19997 8396
rect 19931 8331 19997 8332
rect 19566 2685 19626 8331
rect 20118 4045 20178 25875
rect 20854 16557 20914 29003
rect 20851 16556 20917 16557
rect 20851 16492 20852 16556
rect 20916 16492 20917 16556
rect 20851 16491 20917 16492
rect 21038 12885 21098 39339
rect 21222 21997 21282 41515
rect 21471 40832 21791 41856
rect 21471 40768 21479 40832
rect 21543 40768 21559 40832
rect 21623 40768 21639 40832
rect 21703 40768 21719 40832
rect 21783 40768 21791 40832
rect 21471 39744 21791 40768
rect 21958 39813 22018 43147
rect 22139 42668 22205 42669
rect 22139 42604 22140 42668
rect 22204 42604 22205 42668
rect 22139 42603 22205 42604
rect 21955 39812 22021 39813
rect 21955 39748 21956 39812
rect 22020 39748 22021 39812
rect 21955 39747 22021 39748
rect 21471 39680 21479 39744
rect 21543 39680 21559 39744
rect 21623 39680 21639 39744
rect 21703 39680 21719 39744
rect 21783 39680 21791 39744
rect 21471 38656 21791 39680
rect 21471 38592 21479 38656
rect 21543 38592 21559 38656
rect 21623 38592 21639 38656
rect 21703 38592 21719 38656
rect 21783 38592 21791 38656
rect 21471 37568 21791 38592
rect 21471 37504 21479 37568
rect 21543 37504 21559 37568
rect 21623 37504 21639 37568
rect 21703 37504 21719 37568
rect 21783 37504 21791 37568
rect 21471 36480 21791 37504
rect 21471 36416 21479 36480
rect 21543 36416 21559 36480
rect 21623 36416 21639 36480
rect 21703 36416 21719 36480
rect 21783 36416 21791 36480
rect 21471 35392 21791 36416
rect 21471 35328 21479 35392
rect 21543 35328 21559 35392
rect 21623 35328 21639 35392
rect 21703 35328 21719 35392
rect 21783 35328 21791 35392
rect 21471 34304 21791 35328
rect 21471 34240 21479 34304
rect 21543 34240 21559 34304
rect 21623 34240 21639 34304
rect 21703 34240 21719 34304
rect 21783 34240 21791 34304
rect 21471 33216 21791 34240
rect 21471 33152 21479 33216
rect 21543 33152 21559 33216
rect 21623 33152 21639 33216
rect 21703 33152 21719 33216
rect 21783 33152 21791 33216
rect 21471 32128 21791 33152
rect 21471 32064 21479 32128
rect 21543 32064 21559 32128
rect 21623 32064 21639 32128
rect 21703 32064 21719 32128
rect 21783 32064 21791 32128
rect 21471 31040 21791 32064
rect 21471 30976 21479 31040
rect 21543 30976 21559 31040
rect 21623 30976 21639 31040
rect 21703 30976 21719 31040
rect 21783 30976 21791 31040
rect 21471 29952 21791 30976
rect 21471 29888 21479 29952
rect 21543 29888 21559 29952
rect 21623 29888 21639 29952
rect 21703 29888 21719 29952
rect 21783 29888 21791 29952
rect 21471 28864 21791 29888
rect 21471 28800 21479 28864
rect 21543 28800 21559 28864
rect 21623 28800 21639 28864
rect 21703 28800 21719 28864
rect 21783 28800 21791 28864
rect 21471 27776 21791 28800
rect 21471 27712 21479 27776
rect 21543 27712 21559 27776
rect 21623 27712 21639 27776
rect 21703 27712 21719 27776
rect 21783 27712 21791 27776
rect 21471 26688 21791 27712
rect 21471 26624 21479 26688
rect 21543 26624 21559 26688
rect 21623 26624 21639 26688
rect 21703 26624 21719 26688
rect 21783 26624 21791 26688
rect 21471 25600 21791 26624
rect 21471 25536 21479 25600
rect 21543 25536 21559 25600
rect 21623 25536 21639 25600
rect 21703 25536 21719 25600
rect 21783 25536 21791 25600
rect 21471 24512 21791 25536
rect 21471 24448 21479 24512
rect 21543 24448 21559 24512
rect 21623 24448 21639 24512
rect 21703 24448 21719 24512
rect 21783 24448 21791 24512
rect 21471 23424 21791 24448
rect 21955 24172 22021 24173
rect 21955 24108 21956 24172
rect 22020 24108 22021 24172
rect 21955 24107 22021 24108
rect 21471 23360 21479 23424
rect 21543 23360 21559 23424
rect 21623 23360 21639 23424
rect 21703 23360 21719 23424
rect 21783 23360 21791 23424
rect 21471 22336 21791 23360
rect 21471 22272 21479 22336
rect 21543 22272 21559 22336
rect 21623 22272 21639 22336
rect 21703 22272 21719 22336
rect 21783 22272 21791 22336
rect 21219 21996 21285 21997
rect 21219 21932 21220 21996
rect 21284 21932 21285 21996
rect 21219 21931 21285 21932
rect 21471 21248 21791 22272
rect 21471 21184 21479 21248
rect 21543 21184 21559 21248
rect 21623 21184 21639 21248
rect 21703 21184 21719 21248
rect 21783 21184 21791 21248
rect 21471 20160 21791 21184
rect 21471 20096 21479 20160
rect 21543 20096 21559 20160
rect 21623 20096 21639 20160
rect 21703 20096 21719 20160
rect 21783 20096 21791 20160
rect 21471 19072 21791 20096
rect 21471 19008 21479 19072
rect 21543 19008 21559 19072
rect 21623 19008 21639 19072
rect 21703 19008 21719 19072
rect 21783 19008 21791 19072
rect 21471 17984 21791 19008
rect 21471 17920 21479 17984
rect 21543 17920 21559 17984
rect 21623 17920 21639 17984
rect 21703 17920 21719 17984
rect 21783 17920 21791 17984
rect 21471 16896 21791 17920
rect 21471 16832 21479 16896
rect 21543 16832 21559 16896
rect 21623 16832 21639 16896
rect 21703 16832 21719 16896
rect 21783 16832 21791 16896
rect 21471 15808 21791 16832
rect 21471 15744 21479 15808
rect 21543 15744 21559 15808
rect 21623 15744 21639 15808
rect 21703 15744 21719 15808
rect 21783 15744 21791 15808
rect 21471 14720 21791 15744
rect 21471 14656 21479 14720
rect 21543 14656 21559 14720
rect 21623 14656 21639 14720
rect 21703 14656 21719 14720
rect 21783 14656 21791 14720
rect 21219 13836 21285 13837
rect 21219 13772 21220 13836
rect 21284 13772 21285 13836
rect 21219 13771 21285 13772
rect 21035 12884 21101 12885
rect 21035 12820 21036 12884
rect 21100 12820 21101 12884
rect 21035 12819 21101 12820
rect 20851 8396 20917 8397
rect 20851 8332 20852 8396
rect 20916 8332 20917 8396
rect 20851 8331 20917 8332
rect 20115 4044 20181 4045
rect 20115 3980 20116 4044
rect 20180 3980 20181 4044
rect 20115 3979 20181 3980
rect 20854 3365 20914 8331
rect 20851 3364 20917 3365
rect 20851 3300 20852 3364
rect 20916 3300 20917 3364
rect 20851 3299 20917 3300
rect 19563 2684 19629 2685
rect 19563 2620 19564 2684
rect 19628 2620 19629 2684
rect 19563 2619 19629 2620
rect 21222 2413 21282 13771
rect 21471 13632 21791 14656
rect 21471 13568 21479 13632
rect 21543 13568 21559 13632
rect 21623 13568 21639 13632
rect 21703 13568 21719 13632
rect 21783 13568 21791 13632
rect 21471 12544 21791 13568
rect 21471 12480 21479 12544
rect 21543 12480 21559 12544
rect 21623 12480 21639 12544
rect 21703 12480 21719 12544
rect 21783 12480 21791 12544
rect 21471 11456 21791 12480
rect 21471 11392 21479 11456
rect 21543 11392 21559 11456
rect 21623 11392 21639 11456
rect 21703 11392 21719 11456
rect 21783 11392 21791 11456
rect 21471 10368 21791 11392
rect 21471 10304 21479 10368
rect 21543 10304 21559 10368
rect 21623 10304 21639 10368
rect 21703 10304 21719 10368
rect 21783 10304 21791 10368
rect 21471 9280 21791 10304
rect 21471 9216 21479 9280
rect 21543 9216 21559 9280
rect 21623 9216 21639 9280
rect 21703 9216 21719 9280
rect 21783 9216 21791 9280
rect 21471 8192 21791 9216
rect 21471 8128 21479 8192
rect 21543 8128 21559 8192
rect 21623 8128 21639 8192
rect 21703 8128 21719 8192
rect 21783 8128 21791 8192
rect 21471 7104 21791 8128
rect 21471 7040 21479 7104
rect 21543 7040 21559 7104
rect 21623 7040 21639 7104
rect 21703 7040 21719 7104
rect 21783 7040 21791 7104
rect 21471 6016 21791 7040
rect 21471 5952 21479 6016
rect 21543 5952 21559 6016
rect 21623 5952 21639 6016
rect 21703 5952 21719 6016
rect 21783 5952 21791 6016
rect 21471 4928 21791 5952
rect 21471 4864 21479 4928
rect 21543 4864 21559 4928
rect 21623 4864 21639 4928
rect 21703 4864 21719 4928
rect 21783 4864 21791 4928
rect 21471 3840 21791 4864
rect 21958 4725 22018 24107
rect 21955 4724 22021 4725
rect 21955 4660 21956 4724
rect 22020 4660 22021 4724
rect 21955 4659 22021 4660
rect 21471 3776 21479 3840
rect 21543 3776 21559 3840
rect 21623 3776 21639 3840
rect 21703 3776 21719 3840
rect 21783 3776 21791 3840
rect 21471 2752 21791 3776
rect 21471 2688 21479 2752
rect 21543 2688 21559 2752
rect 21623 2688 21639 2752
rect 21703 2688 21719 2752
rect 21783 2688 21791 2752
rect 21219 2412 21285 2413
rect 21219 2348 21220 2412
rect 21284 2348 21285 2412
rect 21219 2347 21285 2348
rect 21471 1664 21791 2688
rect 22142 2685 22202 42603
rect 24403 42464 24723 43488
rect 24403 42400 24411 42464
rect 24475 42400 24491 42464
rect 24555 42400 24571 42464
rect 24635 42400 24651 42464
rect 24715 42400 24723 42464
rect 24403 41376 24723 42400
rect 24403 41312 24411 41376
rect 24475 41312 24491 41376
rect 24555 41312 24571 41376
rect 24635 41312 24651 41376
rect 24715 41312 24723 41376
rect 24403 40288 24723 41312
rect 24403 40224 24411 40288
rect 24475 40224 24491 40288
rect 24555 40224 24571 40288
rect 24635 40224 24651 40288
rect 24715 40224 24723 40288
rect 24403 39200 24723 40224
rect 24403 39136 24411 39200
rect 24475 39136 24491 39200
rect 24555 39136 24571 39200
rect 24635 39136 24651 39200
rect 24715 39136 24723 39200
rect 24403 38112 24723 39136
rect 24403 38048 24411 38112
rect 24475 38048 24491 38112
rect 24555 38048 24571 38112
rect 24635 38048 24651 38112
rect 24715 38048 24723 38112
rect 24403 37024 24723 38048
rect 24403 36960 24411 37024
rect 24475 36960 24491 37024
rect 24555 36960 24571 37024
rect 24635 36960 24651 37024
rect 24715 36960 24723 37024
rect 24403 35936 24723 36960
rect 24403 35872 24411 35936
rect 24475 35872 24491 35936
rect 24555 35872 24571 35936
rect 24635 35872 24651 35936
rect 24715 35872 24723 35936
rect 22507 35596 22573 35597
rect 22507 35532 22508 35596
rect 22572 35532 22573 35596
rect 22507 35531 22573 35532
rect 22323 34644 22389 34645
rect 22323 34580 22324 34644
rect 22388 34580 22389 34644
rect 22323 34579 22389 34580
rect 22326 5405 22386 34579
rect 22323 5404 22389 5405
rect 22323 5340 22324 5404
rect 22388 5340 22389 5404
rect 22323 5339 22389 5340
rect 22139 2684 22205 2685
rect 22139 2620 22140 2684
rect 22204 2620 22205 2684
rect 22139 2619 22205 2620
rect 22510 2005 22570 35531
rect 24403 34848 24723 35872
rect 24403 34784 24411 34848
rect 24475 34784 24491 34848
rect 24555 34784 24571 34848
rect 24635 34784 24651 34848
rect 24715 34784 24723 34848
rect 24403 33760 24723 34784
rect 24403 33696 24411 33760
rect 24475 33696 24491 33760
rect 24555 33696 24571 33760
rect 24635 33696 24651 33760
rect 24715 33696 24723 33760
rect 24403 32672 24723 33696
rect 24403 32608 24411 32672
rect 24475 32608 24491 32672
rect 24555 32608 24571 32672
rect 24635 32608 24651 32672
rect 24715 32608 24723 32672
rect 24403 31584 24723 32608
rect 24403 31520 24411 31584
rect 24475 31520 24491 31584
rect 24555 31520 24571 31584
rect 24635 31520 24651 31584
rect 24715 31520 24723 31584
rect 24403 30496 24723 31520
rect 24403 30432 24411 30496
rect 24475 30432 24491 30496
rect 24555 30432 24571 30496
rect 24635 30432 24651 30496
rect 24715 30432 24723 30496
rect 24403 29408 24723 30432
rect 24403 29344 24411 29408
rect 24475 29344 24491 29408
rect 24555 29344 24571 29408
rect 24635 29344 24651 29408
rect 24715 29344 24723 29408
rect 24403 28320 24723 29344
rect 24403 28256 24411 28320
rect 24475 28256 24491 28320
rect 24555 28256 24571 28320
rect 24635 28256 24651 28320
rect 24715 28256 24723 28320
rect 22691 27980 22757 27981
rect 22691 27916 22692 27980
rect 22756 27916 22757 27980
rect 22691 27915 22757 27916
rect 22694 10165 22754 27915
rect 24403 27232 24723 28256
rect 24403 27168 24411 27232
rect 24475 27168 24491 27232
rect 24555 27168 24571 27232
rect 24635 27168 24651 27232
rect 24715 27168 24723 27232
rect 24403 26144 24723 27168
rect 24403 26080 24411 26144
rect 24475 26080 24491 26144
rect 24555 26080 24571 26144
rect 24635 26080 24651 26144
rect 24715 26080 24723 26144
rect 24403 25056 24723 26080
rect 24403 24992 24411 25056
rect 24475 24992 24491 25056
rect 24555 24992 24571 25056
rect 24635 24992 24651 25056
rect 24715 24992 24723 25056
rect 24403 23968 24723 24992
rect 24403 23904 24411 23968
rect 24475 23904 24491 23968
rect 24555 23904 24571 23968
rect 24635 23904 24651 23968
rect 24715 23904 24723 23968
rect 24403 22880 24723 23904
rect 24403 22816 24411 22880
rect 24475 22816 24491 22880
rect 24555 22816 24571 22880
rect 24635 22816 24651 22880
rect 24715 22816 24723 22880
rect 24403 21792 24723 22816
rect 24403 21728 24411 21792
rect 24475 21728 24491 21792
rect 24555 21728 24571 21792
rect 24635 21728 24651 21792
rect 24715 21728 24723 21792
rect 24403 20704 24723 21728
rect 24403 20640 24411 20704
rect 24475 20640 24491 20704
rect 24555 20640 24571 20704
rect 24635 20640 24651 20704
rect 24715 20640 24723 20704
rect 24403 19616 24723 20640
rect 24403 19552 24411 19616
rect 24475 19552 24491 19616
rect 24555 19552 24571 19616
rect 24635 19552 24651 19616
rect 24715 19552 24723 19616
rect 24403 18528 24723 19552
rect 24403 18464 24411 18528
rect 24475 18464 24491 18528
rect 24555 18464 24571 18528
rect 24635 18464 24651 18528
rect 24715 18464 24723 18528
rect 24403 17440 24723 18464
rect 24403 17376 24411 17440
rect 24475 17376 24491 17440
rect 24555 17376 24571 17440
rect 24635 17376 24651 17440
rect 24715 17376 24723 17440
rect 24403 16352 24723 17376
rect 24403 16288 24411 16352
rect 24475 16288 24491 16352
rect 24555 16288 24571 16352
rect 24635 16288 24651 16352
rect 24715 16288 24723 16352
rect 24403 15264 24723 16288
rect 24403 15200 24411 15264
rect 24475 15200 24491 15264
rect 24555 15200 24571 15264
rect 24635 15200 24651 15264
rect 24715 15200 24723 15264
rect 24403 14176 24723 15200
rect 24403 14112 24411 14176
rect 24475 14112 24491 14176
rect 24555 14112 24571 14176
rect 24635 14112 24651 14176
rect 24715 14112 24723 14176
rect 24403 13088 24723 14112
rect 24403 13024 24411 13088
rect 24475 13024 24491 13088
rect 24555 13024 24571 13088
rect 24635 13024 24651 13088
rect 24715 13024 24723 13088
rect 24403 12000 24723 13024
rect 24403 11936 24411 12000
rect 24475 11936 24491 12000
rect 24555 11936 24571 12000
rect 24635 11936 24651 12000
rect 24715 11936 24723 12000
rect 24403 10912 24723 11936
rect 24403 10848 24411 10912
rect 24475 10848 24491 10912
rect 24555 10848 24571 10912
rect 24635 10848 24651 10912
rect 24715 10848 24723 10912
rect 22691 10164 22757 10165
rect 22691 10100 22692 10164
rect 22756 10100 22757 10164
rect 22691 10099 22757 10100
rect 24403 9824 24723 10848
rect 24403 9760 24411 9824
rect 24475 9760 24491 9824
rect 24555 9760 24571 9824
rect 24635 9760 24651 9824
rect 24715 9760 24723 9824
rect 24403 8736 24723 9760
rect 24403 8672 24411 8736
rect 24475 8672 24491 8736
rect 24555 8672 24571 8736
rect 24635 8672 24651 8736
rect 24715 8672 24723 8736
rect 24403 7648 24723 8672
rect 24403 7584 24411 7648
rect 24475 7584 24491 7648
rect 24555 7584 24571 7648
rect 24635 7584 24651 7648
rect 24715 7584 24723 7648
rect 24403 6560 24723 7584
rect 24403 6496 24411 6560
rect 24475 6496 24491 6560
rect 24555 6496 24571 6560
rect 24635 6496 24651 6560
rect 24715 6496 24723 6560
rect 24403 5472 24723 6496
rect 24403 5408 24411 5472
rect 24475 5408 24491 5472
rect 24555 5408 24571 5472
rect 24635 5408 24651 5472
rect 24715 5408 24723 5472
rect 24403 4384 24723 5408
rect 24403 4320 24411 4384
rect 24475 4320 24491 4384
rect 24555 4320 24571 4384
rect 24635 4320 24651 4384
rect 24715 4320 24723 4384
rect 24403 3296 24723 4320
rect 24403 3232 24411 3296
rect 24475 3232 24491 3296
rect 24555 3232 24571 3296
rect 24635 3232 24651 3296
rect 24715 3232 24723 3296
rect 24403 2208 24723 3232
rect 24403 2144 24411 2208
rect 24475 2144 24491 2208
rect 24555 2144 24571 2208
rect 24635 2144 24651 2208
rect 24715 2144 24723 2208
rect 22507 2004 22573 2005
rect 22507 1940 22508 2004
rect 22572 1940 22573 2004
rect 22507 1939 22573 1940
rect 21471 1600 21479 1664
rect 21543 1600 21559 1664
rect 21623 1600 21639 1664
rect 21703 1600 21719 1664
rect 21783 1600 21791 1664
rect 21471 1040 21791 1600
rect 24403 1120 24723 2144
rect 24403 1056 24411 1120
rect 24475 1056 24491 1120
rect 24555 1056 24571 1120
rect 24635 1056 24651 1120
rect 24715 1056 24723 1120
rect 24403 1040 24723 1056
rect 19379 916 19445 917
rect 19379 852 19380 916
rect 19444 852 19445 916
rect 19379 851 19445 852
rect 10547 780 10613 781
rect 10547 716 10548 780
rect 10612 716 10613 780
rect 10547 715 10613 716
rect 795 508 861 509
rect 795 444 796 508
rect 860 444 861 508
rect 795 443 861 444
use sky130_fd_sc_hd__diode_2  ANTENNA_1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 6532 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1688980957
transform 1 0 9568 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1688980957
transform 1 0 3956 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1688980957
transform 1 0 3588 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1688980957
transform 1 0 16376 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp 1688980957
transform 1 0 12052 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp 1688980957
transform 1 0 22724 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_8
timestamp 1688980957
transform 1 0 23184 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_9
timestamp 1688980957
transform 1 0 9200 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_10
timestamp 1688980957
transform 1 0 11592 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_11
timestamp 1688980957
transform 1 0 5888 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_12
timestamp 1688980957
transform 1 0 5520 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_13
timestamp 1688980957
transform 1 0 8096 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_14
timestamp 1688980957
transform 1 0 10028 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_15
timestamp 1688980957
transform 1 0 9108 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_16
timestamp 1688980957
transform 1 0 14444 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_17
timestamp 1688980957
transform 1 0 2484 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_18
timestamp 1688980957
transform 1 0 15640 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_19
timestamp 1688980957
transform 1 0 9016 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_20
timestamp 1688980957
transform 1 0 23092 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_21
timestamp 1688980957
transform 1 0 23276 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_22
timestamp 1688980957
transform 1 0 4048 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_23
timestamp 1688980957
transform 1 0 2208 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_24
timestamp 1688980957
transform 1 0 4416 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_25
timestamp 1688980957
transform 1 0 1564 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_26
timestamp 1688980957
transform 1 0 23644 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_0__0_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 23092 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_1__0_
timestamp 1688980957
transform 1 0 23184 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_2__0_
timestamp 1688980957
transform 1 0 23184 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_3__0_
timestamp 1688980957
transform 1 0 23460 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_4__0_
timestamp 1688980957
transform 1 0 23460 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_5__0_
timestamp 1688980957
transform 1 0 23184 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_6__0_
timestamp 1688980957
transform 1 0 23276 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_7__0_
timestamp 1688980957
transform 1 0 22724 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_8__0_
timestamp 1688980957
transform 1 0 23276 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_9__0_
timestamp 1688980957
transform 1 0 22724 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_10__0_
timestamp 1688980957
transform 1 0 22540 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_11__0_
timestamp 1688980957
transform 1 0 23092 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_12__0_
timestamp 1688980957
transform 1 0 22908 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_13__0_
timestamp 1688980957
transform 1 0 23184 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_14__0_
timestamp 1688980957
transform 1 0 22632 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_15__0_
timestamp 1688980957
transform 1 0 22816 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_16__0_
timestamp 1688980957
transform 1 0 21804 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_17__0_
timestamp 1688980957
transform 1 0 22632 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_18__0_
timestamp 1688980957
transform 1 0 20424 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_19__0_
timestamp 1688980957
transform 1 0 20976 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_20__0_
timestamp 1688980957
transform 1 0 20148 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_21__0_
timestamp 1688980957
transform 1 0 23368 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_22__0_
timestamp 1688980957
transform 1 0 21896 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_23__0_
timestamp 1688980957
transform 1 0 19688 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_24__0_
timestamp 1688980957
transform 1 0 18584 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_25__0_
timestamp 1688980957
transform 1 0 21804 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_26__0_
timestamp 1688980957
transform 1 0 22264 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_27__0_
timestamp 1688980957
transform 1 0 20332 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_28__0_
timestamp 1688980957
transform 1 0 18400 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_29__0_
timestamp 1688980957
transform 1 0 23368 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_30__0_
timestamp 1688980957
transform 1 0 21068 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_31__0_
timestamp 1688980957
transform 1 0 20516 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_0__0_
timestamp 1688980957
transform 1 0 23644 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_1__0_
timestamp 1688980957
transform 1 0 23644 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_2__0_
timestamp 1688980957
transform 1 0 22908 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_3__0_
timestamp 1688980957
transform 1 0 22632 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_4__0_
timestamp 1688980957
transform 1 0 23644 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_5__0_
timestamp 1688980957
transform 1 0 23644 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_6__0_
timestamp 1688980957
transform 1 0 23000 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_7__0_
timestamp 1688980957
transform 1 0 23644 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_8__0_
timestamp 1688980957
transform 1 0 23368 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_9__0_
timestamp 1688980957
transform 1 0 23460 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_10__0_
timestamp 1688980957
transform 1 0 23184 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_11__0_
timestamp 1688980957
transform 1 0 23644 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_12__0_
timestamp 1688980957
transform 1 0 23552 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_13__0_
timestamp 1688980957
transform 1 0 23644 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_14__0_
timestamp 1688980957
transform 1 0 23368 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_15__0_
timestamp 1688980957
transform 1 0 23368 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_16__0_
timestamp 1688980957
transform 1 0 22356 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_17__0_
timestamp 1688980957
transform 1 0 23092 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_18__0_
timestamp 1688980957
transform 1 0 21252 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_19__0_
timestamp 1688980957
transform 1 0 21712 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_20__0_
timestamp 1688980957
transform 1 0 20792 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_21__0_
timestamp 1688980957
transform 1 0 23644 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_22__0_
timestamp 1688980957
transform 1 0 22632 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_23__0_
timestamp 1688980957
transform 1 0 20332 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_24__0_
timestamp 1688980957
transform 1 0 19320 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_25__0_
timestamp 1688980957
transform 1 0 22356 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_26__0_
timestamp 1688980957
transform 1 0 21988 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_27__0_
timestamp 1688980957
transform 1 0 23184 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_28__0_
timestamp 1688980957
transform 1 0 19044 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_29__0_
timestamp 1688980957
transform 1 0 23092 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_30__0_
timestamp 1688980957
transform 1 0 21712 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_31__0_
timestamp 1688980957
transform 1 0 21160 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1380 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_43
timestamp 1688980957
transform 1 0 5060 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_91
timestamp 1688980957
transform 1 0 9476 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_107
timestamp 1688980957
transform 1 0 10948 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_138 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 13800 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_151
timestamp 1688980957
transform 1 0 14996 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_9
timestamp 1688980957
transform 1 0 1932 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_17
timestamp 1688980957
transform 1 0 2668 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_85
timestamp 1688980957
transform 1 0 8924 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_89
timestamp 1688980957
transform 1 0 9292 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_140 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 13984 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_144
timestamp 1688980957
transform 1 0 14352 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_147
timestamp 1688980957
transform 1 0 14628 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_153
timestamp 1688980957
transform 1 0 15180 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_167
timestamp 1688980957
transform 1 0 16468 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_213
timestamp 1688980957
transform 1 0 20700 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_241
timestamp 1688980957
transform 1 0 23276 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_247
timestamp 1688980957
transform 1 0 23828 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_3
timestamp 1688980957
transform 1 0 1380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_11
timestamp 1688980957
transform 1 0 2116 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_75
timestamp 1688980957
transform 1 0 8004 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 1688980957
transform 1 0 8740 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_112
timestamp 1688980957
transform 1 0 11408 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_116
timestamp 1688980957
transform 1 0 11776 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_139
timestamp 1688980957
transform 1 0 13892 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_141 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_153
timestamp 1688980957
transform 1 0 15180 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_157
timestamp 1688980957
transform 1 0 15548 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_175
timestamp 1688980957
transform 1 0 17204 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_232
timestamp 1688980957
transform 1 0 22448 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_3
timestamp 1688980957
transform 1 0 1380 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_17
timestamp 1688980957
transform 1 0 2668 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_39
timestamp 1688980957
transform 1 0 4692 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_100
timestamp 1688980957
transform 1 0 10304 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_104
timestamp 1688980957
transform 1 0 10672 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_111
timestamp 1688980957
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_113
timestamp 1688980957
transform 1 0 11500 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_129
timestamp 1688980957
transform 1 0 12972 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_141
timestamp 1688980957
transform 1 0 14076 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_153
timestamp 1688980957
transform 1 0 15180 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_165
timestamp 1688980957
transform 1 0 16284 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_169
timestamp 1688980957
transform 1 0 16652 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_251
timestamp 1688980957
transform 1 0 24196 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_77
timestamp 1688980957
transform 1 0 8188 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_103 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 10580 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_121
timestamp 1688980957
transform 1 0 12236 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_139
timestamp 1688980957
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_141
timestamp 1688980957
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_153
timestamp 1688980957
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_165 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 16284 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_173
timestamp 1688980957
transform 1 0 17020 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_195
timestamp 1688980957
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_235
timestamp 1688980957
transform 1 0 22724 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_250
timestamp 1688980957
transform 1 0 24104 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_57
timestamp 1688980957
transform 1 0 6348 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_86
timestamp 1688980957
transform 1 0 9016 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_94
timestamp 1688980957
transform 1 0 9752 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_99
timestamp 1688980957
transform 1 0 10212 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_107
timestamp 1688980957
transform 1 0 10948 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_111
timestamp 1688980957
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_128
timestamp 1688980957
transform 1 0 12880 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_145
timestamp 1688980957
transform 1 0 14444 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_157
timestamp 1688980957
transform 1 0 15548 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_165
timestamp 1688980957
transform 1 0 16284 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_169
timestamp 1688980957
transform 1 0 16652 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_177
timestamp 1688980957
transform 1 0 17388 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_187
timestamp 1688980957
transform 1 0 18308 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_204
timestamp 1688980957
transform 1 0 19872 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_212
timestamp 1688980957
transform 1 0 20608 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_219
timestamp 1688980957
transform 1 0 21252 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_247
timestamp 1688980957
transform 1 0 23828 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1688980957
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_51
timestamp 1688980957
transform 1 0 5796 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_82
timestamp 1688980957
transform 1 0 8648 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_85
timestamp 1688980957
transform 1 0 8924 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_102 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 10488 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_108
timestamp 1688980957
transform 1 0 11040 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_127
timestamp 1688980957
transform 1 0 12788 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_139
timestamp 1688980957
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_141
timestamp 1688980957
transform 1 0 14076 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_147
timestamp 1688980957
transform 1 0 14628 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_163
timestamp 1688980957
transform 1 0 16100 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_197
timestamp 1688980957
transform 1 0 19228 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_48
timestamp 1688980957
transform 1 0 5520 0 -1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_57
timestamp 1688980957
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_69
timestamp 1688980957
transform 1 0 7452 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_110
timestamp 1688980957
transform 1 0 11224 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_113
timestamp 1688980957
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_125
timestamp 1688980957
transform 1 0 12604 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_163
timestamp 1688980957
transform 1 0 16100 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_167
timestamp 1688980957
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_169
timestamp 1688980957
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_181
timestamp 1688980957
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_193
timestamp 1688980957
transform 1 0 18860 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_214
timestamp 1688980957
transform 1 0 20792 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_250
timestamp 1688980957
transform 1 0 24104 0 -1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_3
timestamp 1688980957
transform 1 0 1380 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_29
timestamp 1688980957
transform 1 0 3772 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_33
timestamp 1688980957
transform 1 0 4140 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_72
timestamp 1688980957
transform 1 0 7728 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_85
timestamp 1688980957
transform 1 0 8924 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_93
timestamp 1688980957
transform 1 0 9660 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_111
timestamp 1688980957
transform 1 0 11316 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_123
timestamp 1688980957
transform 1 0 12420 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_135
timestamp 1688980957
transform 1 0 13524 0 1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_139
timestamp 1688980957
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_141
timestamp 1688980957
transform 1 0 14076 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_166
timestamp 1688980957
transform 1 0 16376 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_178
timestamp 1688980957
transform 1 0 17480 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_210
timestamp 1688980957
transform 1 0 20424 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_39
timestamp 1688980957
transform 1 0 4692 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_57
timestamp 1688980957
transform 1 0 6348 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_90
timestamp 1688980957
transform 1 0 9384 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_102
timestamp 1688980957
transform 1 0 10488 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_110
timestamp 1688980957
transform 1 0 11224 0 -1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_113
timestamp 1688980957
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_125
timestamp 1688980957
transform 1 0 12604 0 -1 6528
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_146
timestamp 1688980957
transform 1 0 14536 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_158
timestamp 1688980957
transform 1 0 15640 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_166
timestamp 1688980957
transform 1 0 16376 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_212
timestamp 1688980957
transform 1 0 20608 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_9
timestamp 1688980957
transform 1 0 1932 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_29
timestamp 1688980957
transform 1 0 3772 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_33
timestamp 1688980957
transform 1 0 4140 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_70
timestamp 1688980957
transform 1 0 7544 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_82
timestamp 1688980957
transform 1 0 8648 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_85
timestamp 1688980957
transform 1 0 8924 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_93
timestamp 1688980957
transform 1 0 9660 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_141
timestamp 1688980957
transform 1 0 14076 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_157
timestamp 1688980957
transform 1 0 15548 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_165
timestamp 1688980957
transform 1 0 16284 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_191
timestamp 1688980957
transform 1 0 18676 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_195
timestamp 1688980957
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_200
timestamp 1688980957
transform 1 0 19504 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_208
timestamp 1688980957
transform 1 0 20240 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_231
timestamp 1688980957
transform 1 0 22356 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_236
timestamp 1688980957
transform 1 0 22816 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_250
timestamp 1688980957
transform 1 0 24104 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_3
timestamp 1688980957
transform 1 0 1380 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_19
timestamp 1688980957
transform 1 0 2852 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_55
timestamp 1688980957
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_57
timestamp 1688980957
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_69
timestamp 1688980957
transform 1 0 7452 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_111
timestamp 1688980957
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_131
timestamp 1688980957
transform 1 0 13156 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_143
timestamp 1688980957
transform 1 0 14260 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_166
timestamp 1688980957
transform 1 0 16376 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_169
timestamp 1688980957
transform 1 0 16652 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_186
timestamp 1688980957
transform 1 0 18216 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_198
timestamp 1688980957
transform 1 0 19320 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_202
timestamp 1688980957
transform 1 0 19688 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_218
timestamp 1688980957
transform 1 0 21160 0 -1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_225
timestamp 1688980957
transform 1 0 21804 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_237
timestamp 1688980957
transform 1 0 22908 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_242
timestamp 1688980957
transform 1 0 23368 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_3
timestamp 1688980957
transform 1 0 1380 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_56
timestamp 1688980957
transform 1 0 6256 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_64
timestamp 1688980957
transform 1 0 6992 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_82
timestamp 1688980957
transform 1 0 8648 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_85
timestamp 1688980957
transform 1 0 8924 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_102
timestamp 1688980957
transform 1 0 10488 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_106
timestamp 1688980957
transform 1 0 10856 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_141
timestamp 1688980957
transform 1 0 14076 0 1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_164
timestamp 1688980957
transform 1 0 16192 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_176
timestamp 1688980957
transform 1 0 17296 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_188
timestamp 1688980957
transform 1 0 18400 0 1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_197
timestamp 1688980957
transform 1 0 19228 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_209
timestamp 1688980957
transform 1 0 20332 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_248
timestamp 1688980957
transform 1 0 23920 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_3
timestamp 1688980957
transform 1 0 1380 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_25
timestamp 1688980957
transform 1 0 3404 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_29
timestamp 1688980957
transform 1 0 3772 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_51
timestamp 1688980957
transform 1 0 5796 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_55
timestamp 1688980957
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_72
timestamp 1688980957
transform 1 0 7728 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_90
timestamp 1688980957
transform 1 0 9384 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_102
timestamp 1688980957
transform 1 0 10488 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_110
timestamp 1688980957
transform 1 0 11224 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_113
timestamp 1688980957
transform 1 0 11500 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_125
timestamp 1688980957
transform 1 0 12604 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_137
timestamp 1688980957
transform 1 0 13708 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_149
timestamp 1688980957
transform 1 0 14812 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_196
timestamp 1688980957
transform 1 0 19136 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_206
timestamp 1688980957
transform 1 0 20056 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_210
timestamp 1688980957
transform 1 0 20424 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_217
timestamp 1688980957
transform 1 0 21068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_223
timestamp 1688980957
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_225
timestamp 1688980957
transform 1 0 21804 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_3
timestamp 1688980957
transform 1 0 1380 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_7
timestamp 1688980957
transform 1 0 1748 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_23
timestamp 1688980957
transform 1 0 3220 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_27
timestamp 1688980957
transform 1 0 3588 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_29
timestamp 1688980957
transform 1 0 3772 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_85
timestamp 1688980957
transform 1 0 8924 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_91
timestamp 1688980957
transform 1 0 9476 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_107
timestamp 1688980957
transform 1 0 10948 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_111
timestamp 1688980957
transform 1 0 11316 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_127
timestamp 1688980957
transform 1 0 12788 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_139
timestamp 1688980957
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_14_141
timestamp 1688980957
transform 1 0 14076 0 1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_14_153
timestamp 1688980957
transform 1 0 15180 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_157
timestamp 1688980957
transform 1 0 15548 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_195
timestamp 1688980957
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_3
timestamp 1688980957
transform 1 0 1380 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_11
timestamp 1688980957
transform 1 0 2116 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_57
timestamp 1688980957
transform 1 0 6348 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_65
timestamp 1688980957
transform 1 0 7084 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_82
timestamp 1688980957
transform 1 0 8648 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_88
timestamp 1688980957
transform 1 0 9200 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_107
timestamp 1688980957
transform 1 0 10948 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_111
timestamp 1688980957
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_113
timestamp 1688980957
transform 1 0 11500 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_121
timestamp 1688980957
transform 1 0 12236 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_137
timestamp 1688980957
transform 1 0 13708 0 -1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_15_156
timestamp 1688980957
transform 1 0 15456 0 -1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_169
timestamp 1688980957
transform 1 0 16652 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_188
timestamp 1688980957
transform 1 0 18400 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_228
timestamp 1688980957
transform 1 0 22080 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_251
timestamp 1688980957
transform 1 0 24196 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_24
timestamp 1688980957
transform 1 0 3312 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_53
timestamp 1688980957
transform 1 0 5980 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_61
timestamp 1688980957
transform 1 0 6716 0 1 9792
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_100
timestamp 1688980957
transform 1 0 10304 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_112
timestamp 1688980957
transform 1 0 11408 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_136
timestamp 1688980957
transform 1 0 13616 0 1 9792
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_16_162
timestamp 1688980957
transform 1 0 16008 0 1 9792
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_174
timestamp 1688980957
transform 1 0 17112 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_195
timestamp 1688980957
transform 1 0 19044 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_197
timestamp 1688980957
transform 1 0 19228 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_206
timestamp 1688980957
transform 1 0 20056 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_212
timestamp 1688980957
transform 1 0 20608 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_220
timestamp 1688980957
transform 1 0 21344 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_228
timestamp 1688980957
transform 1 0 22080 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_54
timestamp 1688980957
transform 1 0 6072 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_57
timestamp 1688980957
transform 1 0 6348 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_69
timestamp 1688980957
transform 1 0 7452 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_81
timestamp 1688980957
transform 1 0 8556 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_93
timestamp 1688980957
transform 1 0 9660 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_128
timestamp 1688980957
transform 1 0 12880 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_149
timestamp 1688980957
transform 1 0 14812 0 -1 10880
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_184
timestamp 1688980957
transform 1 0 18032 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_196
timestamp 1688980957
transform 1 0 19136 0 -1 10880
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_208
timestamp 1688980957
transform 1 0 20240 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_17_220
timestamp 1688980957
transform 1 0 21344 0 -1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_17_231
timestamp 1688980957
transform 1 0 22356 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_3
timestamp 1688980957
transform 1 0 1380 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_21
timestamp 1688980957
transform 1 0 3036 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_41
timestamp 1688980957
transform 1 0 4876 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_64
timestamp 1688980957
transform 1 0 6992 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_68
timestamp 1688980957
transform 1 0 7360 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_100
timestamp 1688980957
transform 1 0 10304 0 1 10880
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_122
timestamp 1688980957
transform 1 0 12328 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_134
timestamp 1688980957
transform 1 0 13432 0 1 10880
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_18_141
timestamp 1688980957
transform 1 0 14076 0 1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_153
timestamp 1688980957
transform 1 0 15180 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_157
timestamp 1688980957
transform 1 0 15548 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_179
timestamp 1688980957
transform 1 0 17572 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_186
timestamp 1688980957
transform 1 0 18216 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_194
timestamp 1688980957
transform 1 0 18952 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_18_197
timestamp 1688980957
transform 1 0 19228 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_234
timestamp 1688980957
transform 1 0 22632 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_250
timestamp 1688980957
transform 1 0 24104 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_3
timestamp 1688980957
transform 1 0 1380 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_25
timestamp 1688980957
transform 1 0 3404 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_48
timestamp 1688980957
transform 1 0 5520 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_72
timestamp 1688980957
transform 1 0 7728 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_94
timestamp 1688980957
transform 1 0 9752 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_19_106
timestamp 1688980957
transform 1 0 10856 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_113
timestamp 1688980957
transform 1 0 11500 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_121
timestamp 1688980957
transform 1 0 12236 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_138
timestamp 1688980957
transform 1 0 13800 0 -1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_19_154
timestamp 1688980957
transform 1 0 15272 0 -1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_166
timestamp 1688980957
transform 1 0 16376 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_169
timestamp 1688980957
transform 1 0 16652 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_173
timestamp 1688980957
transform 1 0 17020 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_215
timestamp 1688980957
transform 1 0 20884 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_223
timestamp 1688980957
transform 1 0 21620 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_228
timestamp 1688980957
transform 1 0 22080 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_232
timestamp 1688980957
transform 1 0 22448 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_251
timestamp 1688980957
transform 1 0 24196 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_9
timestamp 1688980957
transform 1 0 1932 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_29
timestamp 1688980957
transform 1 0 3772 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_43
timestamp 1688980957
transform 1 0 5060 0 1 11968
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_62
timestamp 1688980957
transform 1 0 6808 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_74
timestamp 1688980957
transform 1 0 7912 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_82
timestamp 1688980957
transform 1 0 8648 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_20_85
timestamp 1688980957
transform 1 0 8924 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_91
timestamp 1688980957
transform 1 0 9476 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_107
timestamp 1688980957
transform 1 0 10948 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_141
timestamp 1688980957
transform 1 0 14076 0 1 11968
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_20_160
timestamp 1688980957
transform 1 0 15824 0 1 11968
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_172
timestamp 1688980957
transform 1 0 16928 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_180
timestamp 1688980957
transform 1 0 17664 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_191
timestamp 1688980957
transform 1 0 18676 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_215
timestamp 1688980957
transform 1 0 20884 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_232
timestamp 1688980957
transform 1 0 22448 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_250
timestamp 1688980957
transform 1 0 24104 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_3
timestamp 1688980957
transform 1 0 1380 0 -1 13056
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_44
timestamp 1688980957
transform 1 0 5152 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_57
timestamp 1688980957
transform 1 0 6348 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_61
timestamp 1688980957
transform 1 0 6716 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_77
timestamp 1688980957
transform 1 0 8188 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_107
timestamp 1688980957
transform 1 0 10948 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_111
timestamp 1688980957
transform 1 0 11316 0 -1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_21_128
timestamp 1688980957
transform 1 0 12880 0 -1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_140
timestamp 1688980957
transform 1 0 13984 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_161
timestamp 1688980957
transform 1 0 15916 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_167
timestamp 1688980957
transform 1 0 16468 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_169
timestamp 1688980957
transform 1 0 16652 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_188
timestamp 1688980957
transform 1 0 18400 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_196
timestamp 1688980957
transform 1 0 19136 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_206
timestamp 1688980957
transform 1 0 20056 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_225
timestamp 1688980957
transform 1 0 21804 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_230
timestamp 1688980957
transform 1 0 22264 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_250
timestamp 1688980957
transform 1 0 24104 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_3
timestamp 1688980957
transform 1 0 1380 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_19
timestamp 1688980957
transform 1 0 2852 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_27
timestamp 1688980957
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_29
timestamp 1688980957
transform 1 0 3772 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_47
timestamp 1688980957
transform 1 0 5428 0 1 13056
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_72
timestamp 1688980957
transform 1 0 7728 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_103
timestamp 1688980957
transform 1 0 10580 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_122
timestamp 1688980957
transform 1 0 12328 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_141
timestamp 1688980957
transform 1 0 14076 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_153
timestamp 1688980957
transform 1 0 15180 0 1 13056
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_177
timestamp 1688980957
transform 1 0 17388 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_189
timestamp 1688980957
transform 1 0 18492 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_195
timestamp 1688980957
transform 1 0 19044 0 1 13056
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_22_197
timestamp 1688980957
transform 1 0 19228 0 1 13056
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_22_209
timestamp 1688980957
transform 1 0 20332 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_213
timestamp 1688980957
transform 1 0 20700 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_22_245
timestamp 1688980957
transform 1 0 23644 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_3
timestamp 1688980957
transform 1 0 1380 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_40
timestamp 1688980957
transform 1 0 4784 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_57
timestamp 1688980957
transform 1 0 6348 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_86
timestamp 1688980957
transform 1 0 9016 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_94
timestamp 1688980957
transform 1 0 9752 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_152
timestamp 1688980957
transform 1 0 15088 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_187
timestamp 1688980957
transform 1 0 18308 0 -1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_193
timestamp 1688980957
transform 1 0 18860 0 -1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_205
timestamp 1688980957
transform 1 0 19964 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_217
timestamp 1688980957
transform 1 0 21068 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_223
timestamp 1688980957
transform 1 0 21620 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_225
timestamp 1688980957
transform 1 0 21804 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_9
timestamp 1688980957
transform 1 0 1932 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_17
timestamp 1688980957
transform 1 0 2668 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_25
timestamp 1688980957
transform 1 0 3404 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_56
timestamp 1688980957
transform 1 0 6256 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_83
timestamp 1688980957
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_100
timestamp 1688980957
transform 1 0 10304 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_112
timestamp 1688980957
transform 1 0 11408 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_118
timestamp 1688980957
transform 1 0 11960 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_24_134
timestamp 1688980957
transform 1 0 13432 0 1 14144
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_156
timestamp 1688980957
transform 1 0 15456 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_168
timestamp 1688980957
transform 1 0 16560 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_195
timestamp 1688980957
transform 1 0 19044 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_222
timestamp 1688980957
transform 1 0 21528 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_239
timestamp 1688980957
transform 1 0 23092 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_250
timestamp 1688980957
transform 1 0 24104 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_18
timestamp 1688980957
transform 1 0 2760 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_32
timestamp 1688980957
transform 1 0 4048 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_53
timestamp 1688980957
transform 1 0 5980 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_57
timestamp 1688980957
transform 1 0 6348 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_101
timestamp 1688980957
transform 1 0 10396 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_109
timestamp 1688980957
transform 1 0 11132 0 -1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_113
timestamp 1688980957
transform 1 0 11500 0 -1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_125
timestamp 1688980957
transform 1 0 12604 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_137
timestamp 1688980957
transform 1 0 13708 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_164
timestamp 1688980957
transform 1 0 16192 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_169
timestamp 1688980957
transform 1 0 16652 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_188
timestamp 1688980957
transform 1 0 18400 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_194
timestamp 1688980957
transform 1 0 18952 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_219
timestamp 1688980957
transform 1 0 21252 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_223
timestamp 1688980957
transform 1 0 21620 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_225
timestamp 1688980957
transform 1 0 21804 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_229
timestamp 1688980957
transform 1 0 22172 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_246
timestamp 1688980957
transform 1 0 23736 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_3
timestamp 1688980957
transform 1 0 1380 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_7
timestamp 1688980957
transform 1 0 1748 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_27
timestamp 1688980957
transform 1 0 3588 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_35
timestamp 1688980957
transform 1 0 4324 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_52
timestamp 1688980957
transform 1 0 5888 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_64
timestamp 1688980957
transform 1 0 6992 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_76
timestamp 1688980957
transform 1 0 8096 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_85
timestamp 1688980957
transform 1 0 8924 0 1 15232
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_94
timestamp 1688980957
transform 1 0 9752 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_106
timestamp 1688980957
transform 1 0 10856 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_118
timestamp 1688980957
transform 1 0 11960 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_124
timestamp 1688980957
transform 1 0 12512 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_141
timestamp 1688980957
transform 1 0 14076 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_145
timestamp 1688980957
transform 1 0 14444 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_161
timestamp 1688980957
transform 1 0 15916 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_173
timestamp 1688980957
transform 1 0 17020 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_177
timestamp 1688980957
transform 1 0 17388 0 1 15232
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_181
timestamp 1688980957
transform 1 0 17756 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_193
timestamp 1688980957
transform 1 0 18860 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_197
timestamp 1688980957
transform 1 0 19228 0 1 15232
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_204
timestamp 1688980957
transform 1 0 19872 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_216
timestamp 1688980957
transform 1 0 20976 0 1 15232
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_228
timestamp 1688980957
transform 1 0 22080 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_26_240
timestamp 1688980957
transform 1 0 23184 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_3
timestamp 1688980957
transform 1 0 1380 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_21
timestamp 1688980957
transform 1 0 3036 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_44
timestamp 1688980957
transform 1 0 5152 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_57
timestamp 1688980957
transform 1 0 6348 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_90
timestamp 1688980957
transform 1 0 9384 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_27_113
timestamp 1688980957
transform 1 0 11500 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_121
timestamp 1688980957
transform 1 0 12236 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_144
timestamp 1688980957
transform 1 0 14352 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_167
timestamp 1688980957
transform 1 0 16468 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_27_169
timestamp 1688980957
transform 1 0 16652 0 -1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_27_180
timestamp 1688980957
transform 1 0 17664 0 -1 16320
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_196
timestamp 1688980957
transform 1 0 19136 0 -1 16320
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_208
timestamp 1688980957
transform 1 0 20240 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_220
timestamp 1688980957
transform 1 0 21344 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_240
timestamp 1688980957
transform 1 0 23184 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_3
timestamp 1688980957
transform 1 0 1380 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_26
timestamp 1688980957
transform 1 0 3496 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_33
timestamp 1688980957
transform 1 0 4140 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_76
timestamp 1688980957
transform 1 0 8096 0 1 16320
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_85
timestamp 1688980957
transform 1 0 8924 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_97
timestamp 1688980957
transform 1 0 10028 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_113
timestamp 1688980957
transform 1 0 11500 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_132
timestamp 1688980957
transform 1 0 13248 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_137
timestamp 1688980957
transform 1 0 13708 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_28_141
timestamp 1688980957
transform 1 0 14076 0 1 16320
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_28_159
timestamp 1688980957
transform 1 0 15732 0 1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_171
timestamp 1688980957
transform 1 0 16836 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_188
timestamp 1688980957
transform 1 0 18400 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_203
timestamp 1688980957
transform 1 0 19780 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_208
timestamp 1688980957
transform 1 0 20240 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_219
timestamp 1688980957
transform 1 0 21252 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_223
timestamp 1688980957
transform 1 0 21620 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_39
timestamp 1688980957
transform 1 0 4692 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_90
timestamp 1688980957
transform 1 0 9384 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_106
timestamp 1688980957
transform 1 0 10856 0 -1 17408
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_128
timestamp 1688980957
transform 1 0 12880 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_140
timestamp 1688980957
transform 1 0 13984 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_146
timestamp 1688980957
transform 1 0 14536 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_184
timestamp 1688980957
transform 1 0 18032 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_192
timestamp 1688980957
transform 1 0 18768 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_228
timestamp 1688980957
transform 1 0 22080 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_239
timestamp 1688980957
transform 1 0 23092 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_250
timestamp 1688980957
transform 1 0 24104 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_29
timestamp 1688980957
transform 1 0 3772 0 1 17408
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_41
timestamp 1688980957
transform 1 0 4876 0 1 17408
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_53
timestamp 1688980957
transform 1 0 5980 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_65
timestamp 1688980957
transform 1 0 7084 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_30_81
timestamp 1688980957
transform 1 0 8556 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_85
timestamp 1688980957
transform 1 0 8924 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_93
timestamp 1688980957
transform 1 0 9660 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_131
timestamp 1688980957
transform 1 0 13156 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_139
timestamp 1688980957
transform 1 0 13892 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_156
timestamp 1688980957
transform 1 0 15456 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_160
timestamp 1688980957
transform 1 0 15824 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_168
timestamp 1688980957
transform 1 0 16560 0 1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_30_184
timestamp 1688980957
transform 1 0 18032 0 1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_197
timestamp 1688980957
transform 1 0 19228 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_201
timestamp 1688980957
transform 1 0 19596 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_209
timestamp 1688980957
transform 1 0 20332 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_226
timestamp 1688980957
transform 1 0 21896 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_243
timestamp 1688980957
transform 1 0 23460 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_48
timestamp 1688980957
transform 1 0 5520 0 -1 18496
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_57
timestamp 1688980957
transform 1 0 6348 0 -1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_69
timestamp 1688980957
transform 1 0 7452 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_81
timestamp 1688980957
transform 1 0 8556 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_89
timestamp 1688980957
transform 1 0 9292 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_105
timestamp 1688980957
transform 1 0 10764 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_111
timestamp 1688980957
transform 1 0 11316 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_113
timestamp 1688980957
transform 1 0 11500 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_154
timestamp 1688980957
transform 1 0 15272 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_166
timestamp 1688980957
transform 1 0 16376 0 -1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_31_190
timestamp 1688980957
transform 1 0 18584 0 -1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_202
timestamp 1688980957
transform 1 0 19688 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_31_210
timestamp 1688980957
transform 1 0 20424 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_216
timestamp 1688980957
transform 1 0 20976 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_225
timestamp 1688980957
transform 1 0 21804 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_233
timestamp 1688980957
transform 1 0 22540 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_27
timestamp 1688980957
transform 1 0 3588 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_44
timestamp 1688980957
transform 1 0 5152 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_67
timestamp 1688980957
transform 1 0 7268 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_79
timestamp 1688980957
transform 1 0 8372 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_83
timestamp 1688980957
transform 1 0 8740 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_103
timestamp 1688980957
transform 1 0 10580 0 1 18496
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_121
timestamp 1688980957
transform 1 0 12236 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_32_133
timestamp 1688980957
transform 1 0 13340 0 1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_139
timestamp 1688980957
transform 1 0 13892 0 1 18496
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_141
timestamp 1688980957
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_153
timestamp 1688980957
transform 1 0 15180 0 1 18496
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_165
timestamp 1688980957
transform 1 0 16284 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32_177
timestamp 1688980957
transform 1 0 17388 0 1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_195
timestamp 1688980957
transform 1 0 19044 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_203
timestamp 1688980957
transform 1 0 19780 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_214
timestamp 1688980957
transform 1 0 20792 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_226
timestamp 1688980957
transform 1 0 21896 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_251
timestamp 1688980957
transform 1 0 24196 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_22
timestamp 1688980957
transform 1 0 3128 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_38
timestamp 1688980957
transform 1 0 4600 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_33_57
timestamp 1688980957
transform 1 0 6348 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_78
timestamp 1688980957
transform 1 0 8280 0 -1 19584
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_100
timestamp 1688980957
transform 1 0 10304 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_113
timestamp 1688980957
transform 1 0 11500 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_121
timestamp 1688980957
transform 1 0 12236 0 -1 19584
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_138
timestamp 1688980957
transform 1 0 13800 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_33_165
timestamp 1688980957
transform 1 0 16284 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_220
timestamp 1688980957
transform 1 0 21344 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_250
timestamp 1688980957
transform 1 0 24104 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_7
timestamp 1688980957
transform 1 0 1748 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_27
timestamp 1688980957
transform 1 0 3588 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_29
timestamp 1688980957
transform 1 0 3772 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_41
timestamp 1688980957
transform 1 0 4876 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_49
timestamp 1688980957
transform 1 0 5612 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_85
timestamp 1688980957
transform 1 0 8924 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_34_122
timestamp 1688980957
transform 1 0 12328 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_141
timestamp 1688980957
transform 1 0 14076 0 1 19584
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_168
timestamp 1688980957
transform 1 0 16560 0 1 19584
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_180
timestamp 1688980957
transform 1 0 17664 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_192
timestamp 1688980957
transform 1 0 18768 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_34_232
timestamp 1688980957
transform 1 0 22448 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_238
timestamp 1688980957
transform 1 0 23000 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_15
timestamp 1688980957
transform 1 0 2484 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_42
timestamp 1688980957
transform 1 0 4968 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_54
timestamp 1688980957
transform 1 0 6072 0 -1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_57
timestamp 1688980957
transform 1 0 6348 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_69
timestamp 1688980957
transform 1 0 7452 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_85
timestamp 1688980957
transform 1 0 8924 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_97
timestamp 1688980957
transform 1 0 10028 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_109
timestamp 1688980957
transform 1 0 11132 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_113
timestamp 1688980957
transform 1 0 11500 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_118
timestamp 1688980957
transform 1 0 11960 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_125
timestamp 1688980957
transform 1 0 12604 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_163
timestamp 1688980957
transform 1 0 16100 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_167
timestamp 1688980957
transform 1 0 16468 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_169
timestamp 1688980957
transform 1 0 16652 0 -1 20672
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_181
timestamp 1688980957
transform 1 0 17756 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_193
timestamp 1688980957
transform 1 0 18860 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_201
timestamp 1688980957
transform 1 0 19596 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_205
timestamp 1688980957
transform 1 0 19964 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_210
timestamp 1688980957
transform 1 0 20424 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_215
timestamp 1688980957
transform 1 0 20884 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_221
timestamp 1688980957
transform 1 0 21436 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_231
timestamp 1688980957
transform 1 0 22356 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_235
timestamp 1688980957
transform 1 0 22724 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_251
timestamp 1688980957
transform 1 0 24196 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_29
timestamp 1688980957
transform 1 0 3772 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_41
timestamp 1688980957
transform 1 0 4876 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_36_79
timestamp 1688980957
transform 1 0 8372 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_83
timestamp 1688980957
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_85
timestamp 1688980957
transform 1 0 8924 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_97
timestamp 1688980957
transform 1 0 10028 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_109
timestamp 1688980957
transform 1 0 11132 0 1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_127
timestamp 1688980957
transform 1 0 12788 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_139
timestamp 1688980957
transform 1 0 13892 0 1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_141
timestamp 1688980957
transform 1 0 14076 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_153
timestamp 1688980957
transform 1 0 15180 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_161
timestamp 1688980957
transform 1 0 15916 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_188
timestamp 1688980957
transform 1 0 18400 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_197
timestamp 1688980957
transform 1 0 19228 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_205
timestamp 1688980957
transform 1 0 19964 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_36_222
timestamp 1688980957
transform 1 0 21528 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_228
timestamp 1688980957
transform 1 0 22080 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_245
timestamp 1688980957
transform 1 0 23644 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_24
timestamp 1688980957
transform 1 0 3312 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_28
timestamp 1688980957
transform 1 0 3680 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_50
timestamp 1688980957
transform 1 0 5704 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_57
timestamp 1688980957
transform 1 0 6348 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_63
timestamp 1688980957
transform 1 0 6900 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_79
timestamp 1688980957
transform 1 0 8372 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_113
timestamp 1688980957
transform 1 0 11500 0 -1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_134
timestamp 1688980957
transform 1 0 13432 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_146
timestamp 1688980957
transform 1 0 14536 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_152
timestamp 1688980957
transform 1 0 15088 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_199
timestamp 1688980957
transform 1 0 19412 0 -1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_205
timestamp 1688980957
transform 1 0 19964 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_217
timestamp 1688980957
transform 1 0 21068 0 -1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_223
timestamp 1688980957
transform 1 0 21620 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_225
timestamp 1688980957
transform 1 0 21804 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_233
timestamp 1688980957
transform 1 0 22540 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37_238
timestamp 1688980957
transform 1 0 23000 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_3
timestamp 1688980957
transform 1 0 1380 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_25
timestamp 1688980957
transform 1 0 3404 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_29
timestamp 1688980957
transform 1 0 3772 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_46
timestamp 1688980957
transform 1 0 5336 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_83
timestamp 1688980957
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_85
timestamp 1688980957
transform 1 0 8924 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_89
timestamp 1688980957
transform 1 0 9292 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_38_93
timestamp 1688980957
transform 1 0 9660 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_115
timestamp 1688980957
transform 1 0 11684 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_134
timestamp 1688980957
transform 1 0 13432 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_38_162
timestamp 1688980957
transform 1 0 16008 0 1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_170
timestamp 1688980957
transform 1 0 16744 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_176
timestamp 1688980957
transform 1 0 17296 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_184
timestamp 1688980957
transform 1 0 18032 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_188
timestamp 1688980957
transform 1 0 18400 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_215
timestamp 1688980957
transform 1 0 20884 0 1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_221
timestamp 1688980957
transform 1 0 21436 0 1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_233
timestamp 1688980957
transform 1 0 22540 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_38_245
timestamp 1688980957
transform 1 0 23644 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_22
timestamp 1688980957
transform 1 0 3128 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_39
timestamp 1688980957
transform 1 0 4692 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_57
timestamp 1688980957
transform 1 0 6348 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_80
timestamp 1688980957
transform 1 0 8464 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_85
timestamp 1688980957
transform 1 0 8924 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_93
timestamp 1688980957
transform 1 0 9660 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_109
timestamp 1688980957
transform 1 0 11132 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_113
timestamp 1688980957
transform 1 0 11500 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_121
timestamp 1688980957
transform 1 0 12236 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_39_159
timestamp 1688980957
transform 1 0 15732 0 -1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_167
timestamp 1688980957
transform 1 0 16468 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_172
timestamp 1688980957
transform 1 0 16928 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_184
timestamp 1688980957
transform 1 0 18032 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_204
timestamp 1688980957
transform 1 0 19872 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_235
timestamp 1688980957
transform 1 0 22724 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_243
timestamp 1688980957
transform 1 0 23460 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_11
timestamp 1688980957
transform 1 0 2116 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_29
timestamp 1688980957
transform 1 0 3772 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_41
timestamp 1688980957
transform 1 0 4876 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_53
timestamp 1688980957
transform 1 0 5980 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_65
timestamp 1688980957
transform 1 0 7084 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_77
timestamp 1688980957
transform 1 0 8188 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_83
timestamp 1688980957
transform 1 0 8740 0 1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_85
timestamp 1688980957
transform 1 0 8924 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_97
timestamp 1688980957
transform 1 0 10028 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_109
timestamp 1688980957
transform 1 0 11132 0 1 22848
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_121
timestamp 1688980957
transform 1 0 12236 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_133
timestamp 1688980957
transform 1 0 13340 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_139
timestamp 1688980957
transform 1 0 13892 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_141
timestamp 1688980957
transform 1 0 14076 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_160
timestamp 1688980957
transform 1 0 15824 0 1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_178
timestamp 1688980957
transform 1 0 17480 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_190
timestamp 1688980957
transform 1 0 18584 0 1 22848
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_40_197
timestamp 1688980957
transform 1 0 19228 0 1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_209
timestamp 1688980957
transform 1 0 20332 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_231
timestamp 1688980957
transform 1 0 22356 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_12
timestamp 1688980957
transform 1 0 2208 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_32
timestamp 1688980957
transform 1 0 4048 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_51
timestamp 1688980957
transform 1 0 5796 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_55
timestamp 1688980957
transform 1 0 6164 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_108
timestamp 1688980957
transform 1 0 11040 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_113
timestamp 1688980957
transform 1 0 11500 0 -1 23936
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_129
timestamp 1688980957
transform 1 0 12972 0 -1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_141
timestamp 1688980957
transform 1 0 14076 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_194
timestamp 1688980957
transform 1 0 18952 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_198
timestamp 1688980957
transform 1 0 19320 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_214
timestamp 1688980957
transform 1 0 20792 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_223
timestamp 1688980957
transform 1 0 21620 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_41_225
timestamp 1688980957
transform 1 0 21804 0 -1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_19
timestamp 1688980957
transform 1 0 2852 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_27
timestamp 1688980957
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_29
timestamp 1688980957
transform 1 0 3772 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_33
timestamp 1688980957
transform 1 0 4140 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_55
timestamp 1688980957
transform 1 0 6164 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_63
timestamp 1688980957
transform 1 0 6900 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_82
timestamp 1688980957
transform 1 0 8648 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_85
timestamp 1688980957
transform 1 0 8924 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_108
timestamp 1688980957
transform 1 0 11040 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_137
timestamp 1688980957
transform 1 0 13708 0 1 23936
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_141
timestamp 1688980957
transform 1 0 14076 0 1 23936
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_42_153
timestamp 1688980957
transform 1 0 15180 0 1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_165
timestamp 1688980957
transform 1 0 16284 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_173
timestamp 1688980957
transform 1 0 17020 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_194
timestamp 1688980957
transform 1 0 18952 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_223
timestamp 1688980957
transform 1 0 21620 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_231
timestamp 1688980957
transform 1 0 22356 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_236
timestamp 1688980957
transform 1 0 22816 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_21
timestamp 1688980957
transform 1 0 3036 0 -1 25024
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_44
timestamp 1688980957
transform 1 0 5152 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_90
timestamp 1688980957
transform 1 0 9384 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_107
timestamp 1688980957
transform 1 0 10948 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_111
timestamp 1688980957
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_113
timestamp 1688980957
transform 1 0 11500 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_157
timestamp 1688980957
transform 1 0 15548 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_165
timestamp 1688980957
transform 1 0 16284 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_169
timestamp 1688980957
transform 1 0 16652 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_173
timestamp 1688980957
transform 1 0 17020 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_202
timestamp 1688980957
transform 1 0 19688 0 -1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_209
timestamp 1688980957
transform 1 0 20332 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_221
timestamp 1688980957
transform 1 0 21436 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_43_225
timestamp 1688980957
transform 1 0 21804 0 -1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_233
timestamp 1688980957
transform 1 0 22540 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_24
timestamp 1688980957
transform 1 0 3312 0 1 25024
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_29
timestamp 1688980957
transform 1 0 3772 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_41
timestamp 1688980957
transform 1 0 4876 0 1 25024
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_64
timestamp 1688980957
transform 1 0 6992 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_76
timestamp 1688980957
transform 1 0 8096 0 1 25024
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_85
timestamp 1688980957
transform 1 0 8924 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_97
timestamp 1688980957
transform 1 0 10028 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_108
timestamp 1688980957
transform 1 0 11040 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_112
timestamp 1688980957
transform 1 0 11408 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_134
timestamp 1688980957
transform 1 0 13432 0 1 25024
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_177
timestamp 1688980957
transform 1 0 17388 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_189
timestamp 1688980957
transform 1 0 18492 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_195
timestamp 1688980957
transform 1 0 19044 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_44_197
timestamp 1688980957
transform 1 0 19228 0 1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_209
timestamp 1688980957
transform 1 0 20332 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_217
timestamp 1688980957
transform 1 0 21068 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_222
timestamp 1688980957
transform 1 0 21528 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_244
timestamp 1688980957
transform 1 0 23552 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_21
timestamp 1688980957
transform 1 0 3036 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_37
timestamp 1688980957
transform 1 0 4508 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_57
timestamp 1688980957
transform 1 0 6348 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_69
timestamp 1688980957
transform 1 0 7452 0 -1 26112
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_81
timestamp 1688980957
transform 1 0 8556 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_111
timestamp 1688980957
transform 1 0 11316 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_45_128
timestamp 1688980957
transform 1 0 12880 0 -1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_136
timestamp 1688980957
transform 1 0 13616 0 -1 26112
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_154
timestamp 1688980957
transform 1 0 15272 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_166
timestamp 1688980957
transform 1 0 16376 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_45_184
timestamp 1688980957
transform 1 0 18032 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_203
timestamp 1688980957
transform 1 0 19780 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_207
timestamp 1688980957
transform 1 0 20148 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_45_232
timestamp 1688980957
transform 1 0 22448 0 -1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_237
timestamp 1688980957
transform 1 0 22908 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_9
timestamp 1688980957
transform 1 0 1932 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_26
timestamp 1688980957
transform 1 0 3496 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_50
timestamp 1688980957
transform 1 0 5704 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_113
timestamp 1688980957
transform 1 0 11500 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_132
timestamp 1688980957
transform 1 0 13248 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_46_141
timestamp 1688980957
transform 1 0 14076 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_145
timestamp 1688980957
transform 1 0 14444 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_161
timestamp 1688980957
transform 1 0 15916 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_46_183
timestamp 1688980957
transform 1 0 17940 0 1 26112
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_191
timestamp 1688980957
transform 1 0 18676 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_195
timestamp 1688980957
transform 1 0 19044 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_197
timestamp 1688980957
transform 1 0 19228 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_202
timestamp 1688980957
transform 1 0 19688 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_207
timestamp 1688980957
transform 1 0 20148 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_227
timestamp 1688980957
transform 1 0 21988 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_239
timestamp 1688980957
transform 1 0 23092 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_245
timestamp 1688980957
transform 1 0 23644 0 1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_42
timestamp 1688980957
transform 1 0 4968 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_54
timestamp 1688980957
transform 1 0 6072 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_57
timestamp 1688980957
transform 1 0 6348 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_61
timestamp 1688980957
transform 1 0 6716 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47_80
timestamp 1688980957
transform 1 0 8464 0 -1 27200
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_98
timestamp 1688980957
transform 1 0 10120 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_110
timestamp 1688980957
transform 1 0 11224 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_113
timestamp 1688980957
transform 1 0 11500 0 -1 27200
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_136
timestamp 1688980957
transform 1 0 13616 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_148
timestamp 1688980957
transform 1 0 14720 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_160
timestamp 1688980957
transform 1 0 15824 0 -1 27200
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_169
timestamp 1688980957
transform 1 0 16652 0 -1 27200
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_181
timestamp 1688980957
transform 1 0 17756 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_193
timestamp 1688980957
transform 1 0 18860 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_212
timestamp 1688980957
transform 1 0 20608 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_216
timestamp 1688980957
transform 1 0 20976 0 -1 27200
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_47_225
timestamp 1688980957
transform 1 0 21804 0 -1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_47_237
timestamp 1688980957
transform 1 0 22908 0 -1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47_242
timestamp 1688980957
transform 1 0 23368 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_3
timestamp 1688980957
transform 1 0 1380 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_26
timestamp 1688980957
transform 1 0 3496 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_32
timestamp 1688980957
transform 1 0 4048 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_48_40
timestamp 1688980957
transform 1 0 4784 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_48_58
timestamp 1688980957
transform 1 0 6440 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_79
timestamp 1688980957
transform 1 0 8372 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_83
timestamp 1688980957
transform 1 0 8740 0 1 27200
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_85
timestamp 1688980957
transform 1 0 8924 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_97
timestamp 1688980957
transform 1 0 10028 0 1 27200
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_120
timestamp 1688980957
transform 1 0 12144 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_132
timestamp 1688980957
transform 1 0 13248 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_171
timestamp 1688980957
transform 1 0 16836 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_194
timestamp 1688980957
transform 1 0 18952 0 1 27200
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_197
timestamp 1688980957
transform 1 0 19228 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_209
timestamp 1688980957
transform 1 0 20332 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_213
timestamp 1688980957
transform 1 0 20700 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_230
timestamp 1688980957
transform 1 0 22264 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_243
timestamp 1688980957
transform 1 0 23460 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_31
timestamp 1688980957
transform 1 0 3956 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_37
timestamp 1688980957
transform 1 0 4508 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_57
timestamp 1688980957
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_69
timestamp 1688980957
transform 1 0 7452 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_49_94
timestamp 1688980957
transform 1 0 9752 0 -1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_100
timestamp 1688980957
transform 1 0 10304 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_49_108
timestamp 1688980957
transform 1 0 11040 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_146
timestamp 1688980957
transform 1 0 14536 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_169
timestamp 1688980957
transform 1 0 16652 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49_177
timestamp 1688980957
transform 1 0 17388 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49_183
timestamp 1688980957
transform 1 0 17940 0 -1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_196
timestamp 1688980957
transform 1 0 19136 0 -1 28288
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_208
timestamp 1688980957
transform 1 0 20240 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_220
timestamp 1688980957
transform 1 0 21344 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_225
timestamp 1688980957
transform 1 0 21804 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_246
timestamp 1688980957
transform 1 0 23736 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_7
timestamp 1688980957
transform 1 0 1748 0 1 28288
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_62
timestamp 1688980957
transform 1 0 6808 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_50_74
timestamp 1688980957
transform 1 0 7912 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_82
timestamp 1688980957
transform 1 0 8648 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_50_85
timestamp 1688980957
transform 1 0 8924 0 1 28288
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_91
timestamp 1688980957
transform 1 0 9476 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_107
timestamp 1688980957
transform 1 0 10948 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_138
timestamp 1688980957
transform 1 0 13800 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_50_144
timestamp 1688980957
transform 1 0 14352 0 1 28288
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_162
timestamp 1688980957
transform 1 0 16008 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_174
timestamp 1688980957
transform 1 0 17112 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_195
timestamp 1688980957
transform 1 0 19044 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_197
timestamp 1688980957
transform 1 0 19228 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_216
timestamp 1688980957
transform 1 0 20976 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_50_231
timestamp 1688980957
transform 1 0 22356 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_237
timestamp 1688980957
transform 1 0 22908 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_241
timestamp 1688980957
transform 1 0 23276 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_246
timestamp 1688980957
transform 1 0 23736 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_17
timestamp 1688980957
transform 1 0 2668 0 -1 29376
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_40
timestamp 1688980957
transform 1 0 4784 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_52
timestamp 1688980957
transform 1 0 5888 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_93
timestamp 1688980957
transform 1 0 9660 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_107
timestamp 1688980957
transform 1 0 10948 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_111
timestamp 1688980957
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_113
timestamp 1688980957
transform 1 0 11500 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_51_125
timestamp 1688980957
transform 1 0 12604 0 -1 29376
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_149
timestamp 1688980957
transform 1 0 14812 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_161
timestamp 1688980957
transform 1 0 15916 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_190
timestamp 1688980957
transform 1 0 18584 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_220
timestamp 1688980957
transform 1 0 21344 0 -1 29376
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_51_225
timestamp 1688980957
transform 1 0 21804 0 -1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_51_237
timestamp 1688980957
transform 1 0 22908 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_7
timestamp 1688980957
transform 1 0 1748 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_26
timestamp 1688980957
transform 1 0 3496 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_39
timestamp 1688980957
transform 1 0 4692 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_52_74
timestamp 1688980957
transform 1 0 7912 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_82
timestamp 1688980957
transform 1 0 8648 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_118
timestamp 1688980957
transform 1 0 11960 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_52_130
timestamp 1688980957
transform 1 0 13064 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_138
timestamp 1688980957
transform 1 0 13800 0 1 29376
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_141
timestamp 1688980957
transform 1 0 14076 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_153
timestamp 1688980957
transform 1 0 15180 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_189
timestamp 1688980957
transform 1 0 18492 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_195
timestamp 1688980957
transform 1 0 19044 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_52_197
timestamp 1688980957
transform 1 0 19228 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_203
timestamp 1688980957
transform 1 0 19780 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_209
timestamp 1688980957
transform 1 0 20332 0 1 29376
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_213
timestamp 1688980957
transform 1 0 20700 0 1 29376
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_52_225
timestamp 1688980957
transform 1 0 21804 0 1 29376
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_52_237
timestamp 1688980957
transform 1 0 22908 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_243
timestamp 1688980957
transform 1 0 23460 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53_3
timestamp 1688980957
transform 1 0 1380 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_55
timestamp 1688980957
transform 1 0 6164 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_53_57
timestamp 1688980957
transform 1 0 6348 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53_65
timestamp 1688980957
transform 1 0 7084 0 -1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_83
timestamp 1688980957
transform 1 0 8740 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_53_95
timestamp 1688980957
transform 1 0 9844 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_113
timestamp 1688980957
transform 1 0 11500 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53_136
timestamp 1688980957
transform 1 0 13616 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_53_157
timestamp 1688980957
transform 1 0 15548 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_53_165
timestamp 1688980957
transform 1 0 16284 0 -1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_169
timestamp 1688980957
transform 1 0 16652 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_181
timestamp 1688980957
transform 1 0 17756 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_193
timestamp 1688980957
transform 1 0 18860 0 -1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_205
timestamp 1688980957
transform 1 0 19964 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_53_217
timestamp 1688980957
transform 1 0 21068 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_223
timestamp 1688980957
transform 1 0 21620 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_228
timestamp 1688980957
transform 1 0 22080 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_53_233
timestamp 1688980957
transform 1 0 22540 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_244
timestamp 1688980957
transform 1 0 23552 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_54_29
timestamp 1688980957
transform 1 0 3772 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_34
timestamp 1688980957
transform 1 0 4232 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_54_54
timestamp 1688980957
transform 1 0 6072 0 1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_72
timestamp 1688980957
transform 1 0 7728 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_85
timestamp 1688980957
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_97
timestamp 1688980957
transform 1 0 10028 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_103
timestamp 1688980957
transform 1 0 10580 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_119
timestamp 1688980957
transform 1 0 12052 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_138
timestamp 1688980957
transform 1 0 13800 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_141
timestamp 1688980957
transform 1 0 14076 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_174
timestamp 1688980957
transform 1 0 17112 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_180
timestamp 1688980957
transform 1 0 17664 0 1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_204
timestamp 1688980957
transform 1 0 19872 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_216
timestamp 1688980957
transform 1 0 20976 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_244
timestamp 1688980957
transform 1 0 23552 0 1 30464
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_57
timestamp 1688980957
transform 1 0 6348 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_55_84
timestamp 1688980957
transform 1 0 8832 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_55_88
timestamp 1688980957
transform 1 0 9200 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_105
timestamp 1688980957
transform 1 0 10764 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_111
timestamp 1688980957
transform 1 0 11316 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_113
timestamp 1688980957
transform 1 0 11500 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_55_118
timestamp 1688980957
transform 1 0 11960 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_126
timestamp 1688980957
transform 1 0 12696 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_55_157
timestamp 1688980957
transform 1 0 15548 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_55_165
timestamp 1688980957
transform 1 0 16284 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_169
timestamp 1688980957
transform 1 0 16652 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_55_191
timestamp 1688980957
transform 1 0 18676 0 -1 31552
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_225
timestamp 1688980957
transform 1 0 21804 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_55_237
timestamp 1688980957
transform 1 0 22908 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_241
timestamp 1688980957
transform 1 0 23276 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_9
timestamp 1688980957
transform 1 0 1932 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_44
timestamp 1688980957
transform 1 0 5152 0 1 31552
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_103
timestamp 1688980957
transform 1 0 10580 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_115
timestamp 1688980957
transform 1 0 11684 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_121
timestamp 1688980957
transform 1 0 12236 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_56_137
timestamp 1688980957
transform 1 0 13708 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_56_141
timestamp 1688980957
transform 1 0 14076 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_149
timestamp 1688980957
transform 1 0 14812 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_56_183
timestamp 1688980957
transform 1 0 17940 0 1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_56_190
timestamp 1688980957
transform 1 0 18584 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_195
timestamp 1688980957
transform 1 0 19044 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_197
timestamp 1688980957
transform 1 0 19228 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_56_201
timestamp 1688980957
transform 1 0 19596 0 1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_56_220
timestamp 1688980957
transform 1 0 21344 0 1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_56_232
timestamp 1688980957
transform 1 0 22448 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_56_238
timestamp 1688980957
transform 1 0 23000 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_57_33
timestamp 1688980957
transform 1 0 4140 0 -1 32640
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_57
timestamp 1688980957
transform 1 0 6348 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_69
timestamp 1688980957
transform 1 0 7452 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_91
timestamp 1688980957
transform 1 0 9476 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_57_103
timestamp 1688980957
transform 1 0 10580 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_111
timestamp 1688980957
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_113
timestamp 1688980957
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_125
timestamp 1688980957
transform 1 0 12604 0 -1 32640
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_152
timestamp 1688980957
transform 1 0 15088 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57_164
timestamp 1688980957
transform 1 0 16192 0 -1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_169
timestamp 1688980957
transform 1 0 16652 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_181
timestamp 1688980957
transform 1 0 17756 0 -1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_209
timestamp 1688980957
transform 1 0 20332 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_57_221
timestamp 1688980957
transform 1 0 21436 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_57_225
timestamp 1688980957
transform 1 0 21804 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57_236
timestamp 1688980957
transform 1 0 22816 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57_243
timestamp 1688980957
transform 1 0 23460 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58_3
timestamp 1688980957
transform 1 0 1380 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_58_23
timestamp 1688980957
transform 1 0 3220 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_27
timestamp 1688980957
transform 1 0 3588 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_40
timestamp 1688980957
transform 1 0 4784 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_52
timestamp 1688980957
transform 1 0 5888 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_64
timestamp 1688980957
transform 1 0 6992 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_58_80
timestamp 1688980957
transform 1 0 8464 0 1 32640
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_85
timestamp 1688980957
transform 1 0 8924 0 1 32640
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_97
timestamp 1688980957
transform 1 0 10028 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_58_109
timestamp 1688980957
transform 1 0 11132 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_117
timestamp 1688980957
transform 1 0 11868 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58_122
timestamp 1688980957
transform 1 0 12328 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_139
timestamp 1688980957
transform 1 0 13892 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_177
timestamp 1688980957
transform 1 0 17388 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_189
timestamp 1688980957
transform 1 0 18492 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_195
timestamp 1688980957
transform 1 0 19044 0 1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_58_197
timestamp 1688980957
transform 1 0 19228 0 1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_58_209
timestamp 1688980957
transform 1 0 20332 0 1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_58_242
timestamp 1688980957
transform 1 0 23368 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_24
timestamp 1688980957
transform 1 0 3312 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_30
timestamp 1688980957
transform 1 0 3864 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_49
timestamp 1688980957
transform 1 0 5612 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_55
timestamp 1688980957
transform 1 0 6164 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_57
timestamp 1688980957
transform 1 0 6348 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_59_69
timestamp 1688980957
transform 1 0 7452 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_86
timestamp 1688980957
transform 1 0 9016 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_92
timestamp 1688980957
transform 1 0 9568 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_96
timestamp 1688980957
transform 1 0 9936 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_131
timestamp 1688980957
transform 1 0 13156 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_169
timestamp 1688980957
transform 1 0 16652 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_181
timestamp 1688980957
transform 1 0 17756 0 -1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_193
timestamp 1688980957
transform 1 0 18860 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_59_205
timestamp 1688980957
transform 1 0 19964 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_59_234
timestamp 1688980957
transform 1 0 22632 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_243
timestamp 1688980957
transform 1 0 23460 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_247
timestamp 1688980957
transform 1 0 23828 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_27
timestamp 1688980957
transform 1 0 3588 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_29
timestamp 1688980957
transform 1 0 3772 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_60_48
timestamp 1688980957
transform 1 0 5520 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_56
timestamp 1688980957
transform 1 0 6256 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_75
timestamp 1688980957
transform 1 0 8004 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_85
timestamp 1688980957
transform 1 0 8924 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_60_107
timestamp 1688980957
transform 1 0 10948 0 1 33728
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_125
timestamp 1688980957
transform 1 0 12604 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_60_137
timestamp 1688980957
transform 1 0 13708 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_60_141
timestamp 1688980957
transform 1 0 14076 0 1 33728
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_164
timestamp 1688980957
transform 1 0 16192 0 1 33728
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_176
timestamp 1688980957
transform 1 0 17296 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_60_188
timestamp 1688980957
transform 1 0 18400 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_60_197
timestamp 1688980957
transform 1 0 19228 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_60_214
timestamp 1688980957
transform 1 0 20792 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_220
timestamp 1688980957
transform 1 0 21344 0 1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_224
timestamp 1688980957
transform 1 0 21712 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_60_236
timestamp 1688980957
transform 1 0 22816 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_244
timestamp 1688980957
transform 1 0 23552 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_61_3
timestamp 1688980957
transform 1 0 1380 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_61_37
timestamp 1688980957
transform 1 0 4508 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_61_54
timestamp 1688980957
transform 1 0 6072 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_61_57
timestamp 1688980957
transform 1 0 6348 0 -1 34816
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_75
timestamp 1688980957
transform 1 0 8004 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_61_87
timestamp 1688980957
transform 1 0 9108 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_91
timestamp 1688980957
transform 1 0 9476 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_96
timestamp 1688980957
transform 1 0 9936 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_61_108
timestamp 1688980957
transform 1 0 11040 0 -1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_113
timestamp 1688980957
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_125
timestamp 1688980957
transform 1 0 12604 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_137
timestamp 1688980957
transform 1 0 13708 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_149
timestamp 1688980957
transform 1 0 14812 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_161
timestamp 1688980957
transform 1 0 15916 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_167
timestamp 1688980957
transform 1 0 16468 0 -1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_169
timestamp 1688980957
transform 1 0 16652 0 -1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_181
timestamp 1688980957
transform 1 0 17756 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_61_219
timestamp 1688980957
transform 1 0 21252 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_223
timestamp 1688980957
transform 1 0 21620 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_61_228
timestamp 1688980957
transform 1 0 22080 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_61_237
timestamp 1688980957
transform 1 0 22908 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_241
timestamp 1688980957
transform 1 0 23276 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_245
timestamp 1688980957
transform 1 0 23644 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_62_3
timestamp 1688980957
transform 1 0 1380 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_27
timestamp 1688980957
transform 1 0 3588 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_62_41
timestamp 1688980957
transform 1 0 4876 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_62_76
timestamp 1688980957
transform 1 0 8096 0 1 34816
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_85
timestamp 1688980957
transform 1 0 8924 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_97
timestamp 1688980957
transform 1 0 10028 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_124
timestamp 1688980957
transform 1 0 12512 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_62_136
timestamp 1688980957
transform 1 0 13616 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_141
timestamp 1688980957
transform 1 0 14076 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_147
timestamp 1688980957
transform 1 0 14628 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_154
timestamp 1688980957
transform 1 0 15272 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_166
timestamp 1688980957
transform 1 0 16376 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_178
timestamp 1688980957
transform 1 0 17480 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_62_190
timestamp 1688980957
transform 1 0 18584 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_197
timestamp 1688980957
transform 1 0 19228 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_62_201
timestamp 1688980957
transform 1 0 19596 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_208
timestamp 1688980957
transform 1 0 20240 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_212
timestamp 1688980957
transform 1 0 20608 0 1 34816
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_224
timestamp 1688980957
transform 1 0 21712 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_62_239
timestamp 1688980957
transform 1 0 23092 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_62_243
timestamp 1688980957
transform 1 0 23460 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_18
timestamp 1688980957
transform 1 0 2760 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_63_37
timestamp 1688980957
transform 1 0 4508 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_63_57
timestamp 1688980957
transform 1 0 6348 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_63_65
timestamp 1688980957
transform 1 0 7084 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_63_101
timestamp 1688980957
transform 1 0 10396 0 -1 35904
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_156
timestamp 1688980957
transform 1 0 15456 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_169
timestamp 1688980957
transform 1 0 16652 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_181
timestamp 1688980957
transform 1 0 17756 0 -1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_193
timestamp 1688980957
transform 1 0 18860 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_63_205
timestamp 1688980957
transform 1 0 19964 0 -1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_212
timestamp 1688980957
transform 1 0 20608 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_63_228
timestamp 1688980957
transform 1 0 22080 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_63_237
timestamp 1688980957
transform 1 0 22908 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_64_9
timestamp 1688980957
transform 1 0 1932 0 1 35904
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_53
timestamp 1688980957
transform 1 0 5980 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_64_65
timestamp 1688980957
transform 1 0 7084 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_85
timestamp 1688980957
transform 1 0 8924 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_116
timestamp 1688980957
transform 1 0 11776 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_128
timestamp 1688980957
transform 1 0 12880 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_64_141
timestamp 1688980957
transform 1 0 14076 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_145
timestamp 1688980957
transform 1 0 14444 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_149
timestamp 1688980957
transform 1 0 14812 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_161
timestamp 1688980957
transform 1 0 15916 0 1 35904
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_173
timestamp 1688980957
transform 1 0 17020 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_64_185
timestamp 1688980957
transform 1 0 18124 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_193
timestamp 1688980957
transform 1 0 18860 0 1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_197
timestamp 1688980957
transform 1 0 19228 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_209
timestamp 1688980957
transform 1 0 20332 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_64_213
timestamp 1688980957
transform 1 0 20700 0 1 35904
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_222
timestamp 1688980957
transform 1 0 21528 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_64_234
timestamp 1688980957
transform 1 0 22632 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_238
timestamp 1688980957
transform 1 0 23000 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_245
timestamp 1688980957
transform 1 0 23644 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_65_39
timestamp 1688980957
transform 1 0 4692 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_65_57
timestamp 1688980957
transform 1 0 6348 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_65_65
timestamp 1688980957
transform 1 0 7084 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_65_85
timestamp 1688980957
transform 1 0 8924 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_65_93
timestamp 1688980957
transform 1 0 9660 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_111
timestamp 1688980957
transform 1 0 11316 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_113
timestamp 1688980957
transform 1 0 11500 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_125
timestamp 1688980957
transform 1 0 12604 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_137
timestamp 1688980957
transform 1 0 13708 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_149
timestamp 1688980957
transform 1 0 14812 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_65_161
timestamp 1688980957
transform 1 0 15916 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_167
timestamp 1688980957
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_169
timestamp 1688980957
transform 1 0 16652 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_181
timestamp 1688980957
transform 1 0 17756 0 -1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_193
timestamp 1688980957
transform 1 0 18860 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_65_205
timestamp 1688980957
transform 1 0 19964 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_65_210
timestamp 1688980957
transform 1 0 20424 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_65_219
timestamp 1688980957
transform 1 0 21252 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_223
timestamp 1688980957
transform 1 0 21620 0 -1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_225
timestamp 1688980957
transform 1 0 21804 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_65_237
timestamp 1688980957
transform 1 0 22908 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_65_246
timestamp 1688980957
transform 1 0 23736 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_66_24
timestamp 1688980957
transform 1 0 3312 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_66_35
timestamp 1688980957
transform 1 0 4324 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_39
timestamp 1688980957
transform 1 0 4692 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_66_58
timestamp 1688980957
transform 1 0 6440 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_62
timestamp 1688980957
transform 1 0 6808 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66_78
timestamp 1688980957
transform 1 0 8280 0 1 36992
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_85
timestamp 1688980957
transform 1 0 8924 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_66_97
timestamp 1688980957
transform 1 0 10028 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_101
timestamp 1688980957
transform 1 0 10396 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_120
timestamp 1688980957
transform 1 0 12144 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_66_132
timestamp 1688980957
transform 1 0 13248 0 1 36992
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_141
timestamp 1688980957
transform 1 0 14076 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_153
timestamp 1688980957
transform 1 0 15180 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_165
timestamp 1688980957
transform 1 0 16284 0 1 36992
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_177
timestamp 1688980957
transform 1 0 17388 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66_189
timestamp 1688980957
transform 1 0 18492 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_195
timestamp 1688980957
transform 1 0 19044 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_197
timestamp 1688980957
transform 1 0 19228 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_66_209
timestamp 1688980957
transform 1 0 20332 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_213
timestamp 1688980957
transform 1 0 20700 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66_217
timestamp 1688980957
transform 1 0 21068 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_223
timestamp 1688980957
transform 1 0 21620 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_227
timestamp 1688980957
transform 1 0 21988 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_66_239
timestamp 1688980957
transform 1 0 23092 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_3
timestamp 1688980957
transform 1 0 1380 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_19
timestamp 1688980957
transform 1 0 2852 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_50
timestamp 1688980957
transform 1 0 5704 0 -1 38080
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_57
timestamp 1688980957
transform 1 0 6348 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_67_69
timestamp 1688980957
transform 1 0 7452 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_67_77
timestamp 1688980957
transform 1 0 8188 0 -1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_94
timestamp 1688980957
transform 1 0 9752 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_106
timestamp 1688980957
transform 1 0 10856 0 -1 38080
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_128
timestamp 1688980957
transform 1 0 12880 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_140
timestamp 1688980957
transform 1 0 13984 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_152
timestamp 1688980957
transform 1 0 15088 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_67_164
timestamp 1688980957
transform 1 0 16192 0 -1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_169
timestamp 1688980957
transform 1 0 16652 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_181
timestamp 1688980957
transform 1 0 17756 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_193
timestamp 1688980957
transform 1 0 18860 0 -1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_205
timestamp 1688980957
transform 1 0 19964 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_217
timestamp 1688980957
transform 1 0 21068 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_223
timestamp 1688980957
transform 1 0 21620 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_225
timestamp 1688980957
transform 1 0 21804 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_229
timestamp 1688980957
transform 1 0 22172 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_241
timestamp 1688980957
transform 1 0 23276 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_68_26
timestamp 1688980957
transform 1 0 3496 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_68_50
timestamp 1688980957
transform 1 0 5704 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_68_79
timestamp 1688980957
transform 1 0 8372 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_83
timestamp 1688980957
transform 1 0 8740 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_103
timestamp 1688980957
transform 1 0 10580 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_115
timestamp 1688980957
transform 1 0 11684 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_127
timestamp 1688980957
transform 1 0 12788 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_139
timestamp 1688980957
transform 1 0 13892 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_141
timestamp 1688980957
transform 1 0 14076 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_153
timestamp 1688980957
transform 1 0 15180 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_165
timestamp 1688980957
transform 1 0 16284 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_177
timestamp 1688980957
transform 1 0 17388 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_189
timestamp 1688980957
transform 1 0 18492 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_68_193
timestamp 1688980957
transform 1 0 18860 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_68_197
timestamp 1688980957
transform 1 0 19228 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_201
timestamp 1688980957
transform 1 0 19596 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_205
timestamp 1688980957
transform 1 0 19964 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_217
timestamp 1688980957
transform 1 0 21068 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_68_229
timestamp 1688980957
transform 1 0 22172 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_233
timestamp 1688980957
transform 1 0 22540 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_68_237
timestamp 1688980957
transform 1 0 22908 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_68_245
timestamp 1688980957
transform 1 0 23644 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_69_57
timestamp 1688980957
transform 1 0 6348 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_82
timestamp 1688980957
transform 1 0 8648 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_69_86
timestamp 1688980957
transform 1 0 9016 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_69_90
timestamp 1688980957
transform 1 0 9384 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_69_110
timestamp 1688980957
transform 1 0 11224 0 -1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_117
timestamp 1688980957
transform 1 0 11868 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_129
timestamp 1688980957
transform 1 0 12972 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_141
timestamp 1688980957
transform 1 0 14076 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_153
timestamp 1688980957
transform 1 0 15180 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_69_165
timestamp 1688980957
transform 1 0 16284 0 -1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_169
timestamp 1688980957
transform 1 0 16652 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_181
timestamp 1688980957
transform 1 0 17756 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_193
timestamp 1688980957
transform 1 0 18860 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_69_205
timestamp 1688980957
transform 1 0 19964 0 -1 39168
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_212
timestamp 1688980957
transform 1 0 20608 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_69_228
timestamp 1688980957
transform 1 0 22080 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_236
timestamp 1688980957
transform 1 0 22816 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_69_243
timestamp 1688980957
transform 1 0 23460 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_3
timestamp 1688980957
transform 1 0 1380 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_70_56
timestamp 1688980957
transform 1 0 6256 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_70_77
timestamp 1688980957
transform 1 0 8188 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_83
timestamp 1688980957
transform 1 0 8740 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_110
timestamp 1688980957
transform 1 0 11224 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_122
timestamp 1688980957
transform 1 0 12328 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_70_134
timestamp 1688980957
transform 1 0 13432 0 1 39168
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_141
timestamp 1688980957
transform 1 0 14076 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_153
timestamp 1688980957
transform 1 0 15180 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_165
timestamp 1688980957
transform 1 0 16284 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_177
timestamp 1688980957
transform 1 0 17388 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_70_189
timestamp 1688980957
transform 1 0 18492 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_195
timestamp 1688980957
transform 1 0 19044 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_197
timestamp 1688980957
transform 1 0 19228 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_201
timestamp 1688980957
transform 1 0 19596 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_213
timestamp 1688980957
transform 1 0 20700 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_70_225
timestamp 1688980957
transform 1 0 21804 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_70_234
timestamp 1688980957
transform 1 0 22632 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_71_3
timestamp 1688980957
transform 1 0 1380 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_71_46
timestamp 1688980957
transform 1 0 5336 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_71_50
timestamp 1688980957
transform 1 0 5704 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_71_54
timestamp 1688980957
transform 1 0 6072 0 -1 40256
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_72
timestamp 1688980957
transform 1 0 7728 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_84
timestamp 1688980957
transform 1 0 8832 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_96
timestamp 1688980957
transform 1 0 9936 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_71_108
timestamp 1688980957
transform 1 0 11040 0 -1 40256
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_113
timestamp 1688980957
transform 1 0 11500 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_125
timestamp 1688980957
transform 1 0 12604 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_137
timestamp 1688980957
transform 1 0 13708 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_149
timestamp 1688980957
transform 1 0 14812 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_71_161
timestamp 1688980957
transform 1 0 15916 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_167
timestamp 1688980957
transform 1 0 16468 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_169
timestamp 1688980957
transform 1 0 16652 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_181
timestamp 1688980957
transform 1 0 17756 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_193
timestamp 1688980957
transform 1 0 18860 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_205
timestamp 1688980957
transform 1 0 19964 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_71_217
timestamp 1688980957
transform 1 0 21068 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_71_225
timestamp 1688980957
transform 1 0 21804 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_71_233
timestamp 1688980957
transform 1 0 22540 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_3
timestamp 1688980957
transform 1 0 1380 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_72_56
timestamp 1688980957
transform 1 0 6256 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_72_61
timestamp 1688980957
transform 1 0 6716 0 1 40256
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_69
timestamp 1688980957
transform 1 0 7452 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_72_81
timestamp 1688980957
transform 1 0 8556 0 1 40256
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_85
timestamp 1688980957
transform 1 0 8924 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_97
timestamp 1688980957
transform 1 0 10028 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_109
timestamp 1688980957
transform 1 0 11132 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_121
timestamp 1688980957
transform 1 0 12236 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_72_133
timestamp 1688980957
transform 1 0 13340 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_139
timestamp 1688980957
transform 1 0 13892 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_141
timestamp 1688980957
transform 1 0 14076 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_153
timestamp 1688980957
transform 1 0 15180 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_165
timestamp 1688980957
transform 1 0 16284 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_72_177
timestamp 1688980957
transform 1 0 17388 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_72_185
timestamp 1688980957
transform 1 0 18124 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_72_191
timestamp 1688980957
transform 1 0 18676 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_195
timestamp 1688980957
transform 1 0 19044 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_197
timestamp 1688980957
transform 1 0 19228 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_72_209
timestamp 1688980957
transform 1 0 20332 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_72_232
timestamp 1688980957
transform 1 0 22448 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_72_237
timestamp 1688980957
transform 1 0 22908 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_73_63
timestamp 1688980957
transform 1 0 6900 0 -1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_86
timestamp 1688980957
transform 1 0 9016 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_98
timestamp 1688980957
transform 1 0 10120 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_73_110
timestamp 1688980957
transform 1 0 11224 0 -1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_113
timestamp 1688980957
transform 1 0 11500 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_125
timestamp 1688980957
transform 1 0 12604 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_137
timestamp 1688980957
transform 1 0 13708 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_149
timestamp 1688980957
transform 1 0 14812 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_73_161
timestamp 1688980957
transform 1 0 15916 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_167
timestamp 1688980957
transform 1 0 16468 0 -1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_169
timestamp 1688980957
transform 1 0 16652 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_181
timestamp 1688980957
transform 1 0 17756 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_73_193
timestamp 1688980957
transform 1 0 18860 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_73_198
timestamp 1688980957
transform 1 0 19320 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_73_206
timestamp 1688980957
transform 1 0 20056 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_73_225
timestamp 1688980957
transform 1 0 21804 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_233
timestamp 1688980957
transform 1 0 22540 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_73_250
timestamp 1688980957
transform 1 0 24104 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_29
timestamp 1688980957
transform 1 0 3772 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_74_34
timestamp 1688980957
transform 1 0 4232 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_74_38
timestamp 1688980957
transform 1 0 4600 0 1 41344
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_91
timestamp 1688980957
transform 1 0 9476 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_103
timestamp 1688980957
transform 1 0 10580 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_115
timestamp 1688980957
transform 1 0 11684 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_127
timestamp 1688980957
transform 1 0 12788 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_139
timestamp 1688980957
transform 1 0 13892 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_141
timestamp 1688980957
transform 1 0 14076 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_153
timestamp 1688980957
transform 1 0 15180 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_165
timestamp 1688980957
transform 1 0 16284 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_177
timestamp 1688980957
transform 1 0 17388 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_74_189
timestamp 1688980957
transform 1 0 18492 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_195
timestamp 1688980957
transform 1 0 19044 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_74_207
timestamp 1688980957
transform 1 0 20148 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_227
timestamp 1688980957
transform 1 0 21988 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_75_48
timestamp 1688980957
transform 1 0 5520 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_57
timestamp 1688980957
transform 1 0 6348 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_83
timestamp 1688980957
transform 1 0 8740 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_75_90
timestamp 1688980957
transform 1 0 9384 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_75_94
timestamp 1688980957
transform 1 0 9752 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_75_102
timestamp 1688980957
transform 1 0 10488 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_75_110
timestamp 1688980957
transform 1 0 11224 0 -1 42432
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_113
timestamp 1688980957
transform 1 0 11500 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_125
timestamp 1688980957
transform 1 0 12604 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_137
timestamp 1688980957
transform 1 0 13708 0 -1 42432
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_149
timestamp 1688980957
transform 1 0 14812 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_75_161
timestamp 1688980957
transform 1 0 15916 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_167
timestamp 1688980957
transform 1 0 16468 0 -1 42432
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_169
timestamp 1688980957
transform 1 0 16652 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_75_181
timestamp 1688980957
transform 1 0 17756 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_225
timestamp 1688980957
transform 1 0 21804 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_75_250
timestamp 1688980957
transform 1 0 24104 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_3
timestamp 1688980957
transform 1 0 1380 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_76_10
timestamp 1688980957
transform 1 0 2024 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_76_14
timestamp 1688980957
transform 1 0 2392 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_76_62
timestamp 1688980957
transform 1 0 6808 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_76_70
timestamp 1688980957
transform 1 0 7544 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_76_107
timestamp 1688980957
transform 1 0 10948 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_76_119
timestamp 1688980957
transform 1 0 12052 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_76_128
timestamp 1688980957
transform 1 0 12880 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_136
timestamp 1688980957
transform 1 0 13616 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_76_141
timestamp 1688980957
transform 1 0 14076 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_76_146
timestamp 1688980957
transform 1 0 14536 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_76_155
timestamp 1688980957
transform 1 0 15364 0 1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_163
timestamp 1688980957
transform 1 0 16100 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_247
timestamp 1688980957
transform 1 0 23828 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_77_7
timestamp 1688980957
transform 1 0 1748 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_15
timestamp 1688980957
transform 1 0 2484 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_61
timestamp 1688980957
transform 1 0 6716 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_77_74
timestamp 1688980957
transform 1 0 7912 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_77_78
timestamp 1688980957
transform 1 0 8280 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_111
timestamp 1688980957
transform 1 0 11316 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_77_117
timestamp 1688980957
transform 1 0 11868 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_126
timestamp 1688980957
transform 1 0 12696 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_77_138
timestamp 1688980957
transform 1 0 13800 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_144
timestamp 1688980957
transform 1 0 14352 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_167
timestamp 1688980957
transform 1 0 16468 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_206
timestamp 1688980957
transform 1 0 20056 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_217
timestamp 1688980957
transform 1 0 21068 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_77_250
timestamp 1688980957
transform 1 0 24104 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  input1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4508 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input2 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2760 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input3
timestamp 1688980957
transform 1 0 3772 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input4
timestamp 1688980957
transform 1 0 2760 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input5 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2760 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input6
timestamp 1688980957
transform 1 0 1380 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input7
timestamp 1688980957
transform 1 0 1748 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input8
timestamp 1688980957
transform 1 0 1932 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input9
timestamp 1688980957
transform 1 0 2760 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input10
timestamp 1688980957
transform 1 0 1748 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input11
timestamp 1688980957
transform 1 0 1380 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input12
timestamp 1688980957
transform 1 0 1656 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input13
timestamp 1688980957
transform 1 0 1380 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input14
timestamp 1688980957
transform 1 0 2116 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input15
timestamp 1688980957
transform 1 0 3312 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input16
timestamp 1688980957
transform 1 0 1380 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input17
timestamp 1688980957
transform 1 0 1380 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input18
timestamp 1688980957
transform 1 0 1748 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input19
timestamp 1688980957
transform 1 0 1380 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input20
timestamp 1688980957
transform 1 0 3036 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input21
timestamp 1688980957
transform 1 0 3312 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input22
timestamp 1688980957
transform 1 0 3864 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input23
timestamp 1688980957
transform 1 0 2024 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input24
timestamp 1688980957
transform 1 0 1380 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input25 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1380 0 -1 29376
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input26
timestamp 1688980957
transform 1 0 2760 0 1 30464
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input27
timestamp 1688980957
transform 1 0 2300 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input28
timestamp 1688980957
transform 1 0 3772 0 1 29376
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input29
timestamp 1688980957
transform 1 0 3220 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input30
timestamp 1688980957
transform 1 0 1380 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input31
timestamp 1688980957
transform 1 0 3588 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input32
timestamp 1688980957
transform 1 0 2944 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input33
timestamp 1688980957
transform 1 0 1380 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input34
timestamp 1688980957
transform 1 0 3036 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input35
timestamp 1688980957
transform 1 0 3312 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input36
timestamp 1688980957
transform 1 0 2944 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input37
timestamp 1688980957
transform 1 0 3220 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input38
timestamp 1688980957
transform 1 0 3772 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input39
timestamp 1688980957
transform 1 0 3680 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input40
timestamp 1688980957
transform 1 0 1380 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input41
timestamp 1688980957
transform 1 0 2576 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input42
timestamp 1688980957
transform 1 0 1380 0 1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input43
timestamp 1688980957
transform 1 0 2300 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input44
timestamp 1688980957
transform 1 0 1380 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input45
timestamp 1688980957
transform 1 0 1656 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input46
timestamp 1688980957
transform 1 0 2760 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input47
timestamp 1688980957
transform 1 0 3036 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input48
timestamp 1688980957
transform 1 0 2760 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  input49 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1380 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input50
timestamp 1688980957
transform 1 0 3036 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input51
timestamp 1688980957
transform 1 0 1380 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input52
timestamp 1688980957
transform 1 0 3772 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input53
timestamp 1688980957
transform 1 0 4324 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input54
timestamp 1688980957
transform 1 0 2760 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input55
timestamp 1688980957
transform 1 0 3312 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input56
timestamp 1688980957
transform 1 0 3864 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input57
timestamp 1688980957
transform 1 0 3772 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input58
timestamp 1688980957
transform 1 0 5428 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input59
timestamp 1688980957
transform 1 0 2392 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input60
timestamp 1688980957
transform 1 0 2392 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input61
timestamp 1688980957
transform 1 0 1380 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input62
timestamp 1688980957
transform 1 0 2944 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input63
timestamp 1688980957
transform 1 0 3772 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input64
timestamp 1688980957
transform 1 0 3772 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input65
timestamp 1688980957
transform 1 0 4324 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input66
timestamp 1688980957
transform 1 0 5152 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_8  input67 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1380 0 1 38080
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  input68
timestamp 1688980957
transform 1 0 2760 0 -1 39168
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_4  input69
timestamp 1688980957
transform 1 0 10396 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input70
timestamp 1688980957
transform 1 0 1748 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input71
timestamp 1688980957
transform 1 0 5336 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_8  input72
timestamp 1688980957
transform 1 0 1380 0 -1 41344
box -38 -48 1050 592
use sky130_fd_sc_hd__clkbuf_8  input73
timestamp 1688980957
transform 1 0 2944 0 -1 40256
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_4  input74
timestamp 1688980957
transform 1 0 3312 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_8  input75
timestamp 1688980957
transform 1 0 1380 0 -1 31552
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_4  input76
timestamp 1688980957
transform 1 0 1380 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_8  input77
timestamp 1688980957
transform 1 0 3772 0 1 32640
box -38 -48 1050 592
use sky130_fd_sc_hd__buf_4  input78
timestamp 1688980957
transform 1 0 1932 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input79
timestamp 1688980957
transform 1 0 2760 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input80
timestamp 1688980957
transform 1 0 2484 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__buf_8  input81 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 20332 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  input82
timestamp 1688980957
transform 1 0 18768 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input83
timestamp 1688980957
transform 1 0 23460 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input84
timestamp 1688980957
transform 1 0 21344 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input85
timestamp 1688980957
transform 1 0 23920 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input86
timestamp 1688980957
transform 1 0 23644 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input87
timestamp 1688980957
transform 1 0 23644 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input88
timestamp 1688980957
transform 1 0 20792 0 -1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input89
timestamp 1688980957
transform 1 0 21896 0 1 4352
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input90
timestamp 1688980957
transform 1 0 21804 0 -1 3264
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input91
timestamp 1688980957
transform 1 0 23920 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_16  input92 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 20608 0 1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_8  input93
timestamp 1688980957
transform 1 0 19504 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  input94
timestamp 1688980957
transform 1 0 23000 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_16  input95
timestamp 1688980957
transform 1 0 21804 0 1 1088
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_8  input96
timestamp 1688980957
transform 1 0 22540 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  input97
timestamp 1688980957
transform 1 0 20608 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  input98
timestamp 1688980957
transform 1 0 19504 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  input99
timestamp 1688980957
transform 1 0 18032 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  input100
timestamp 1688980957
transform 1 0 22816 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  input101
timestamp 1688980957
transform 1 0 6348 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input102
timestamp 1688980957
transform 1 0 1472 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input103
timestamp 1688980957
transform 1 0 1380 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input104 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2116 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  input105
timestamp 1688980957
transform 1 0 5520 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input106
timestamp 1688980957
transform 1 0 2576 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input107
timestamp 1688980957
transform 1 0 4140 0 1 1088
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input108
timestamp 1688980957
transform 1 0 2944 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input109
timestamp 1688980957
transform 1 0 5980 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input110
timestamp 1688980957
transform 1 0 7268 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input111
timestamp 1688980957
transform 1 0 5152 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input112
timestamp 1688980957
transform 1 0 5612 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input113
timestamp 1688980957
transform 1 0 2760 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input114
timestamp 1688980957
transform 1 0 1380 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input115
timestamp 1688980957
transform 1 0 1840 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input116
timestamp 1688980957
transform 1 0 2300 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input117
timestamp 1688980957
transform 1 0 3404 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input118
timestamp 1688980957
transform 1 0 2760 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input119
timestamp 1688980957
transform 1 0 2208 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input120
timestamp 1688980957
transform 1 0 5244 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input121
timestamp 1688980957
transform 1 0 6348 0 1 1088
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_1  input122
timestamp 1688980957
transform 1 0 8464 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input123
timestamp 1688980957
transform 1 0 9476 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input124
timestamp 1688980957
transform 1 0 8924 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input125
timestamp 1688980957
transform 1 0 9200 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input126
timestamp 1688980957
transform 1 0 8556 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input127
timestamp 1688980957
transform 1 0 13708 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input128
timestamp 1688980957
transform 1 0 3312 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input129
timestamp 1688980957
transform 1 0 5520 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input130
timestamp 1688980957
transform 1 0 7268 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input131
timestamp 1688980957
transform 1 0 7636 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input132
timestamp 1688980957
transform 1 0 6992 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input133
timestamp 1688980957
transform 1 0 6716 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input134
timestamp 1688980957
transform 1 0 7268 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input135
timestamp 1688980957
transform 1 0 7912 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input136
timestamp 1688980957
transform 1 0 8188 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input137
timestamp 1688980957
transform 1 0 24012 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input138
timestamp 1688980957
transform 1 0 24012 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input139
timestamp 1688980957
transform 1 0 24012 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input140
timestamp 1688980957
transform 1 0 23368 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input141
timestamp 1688980957
transform 1 0 24012 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input142
timestamp 1688980957
transform 1 0 23368 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input143
timestamp 1688980957
transform 1 0 23736 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input144
timestamp 1688980957
transform 1 0 23460 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input145
timestamp 1688980957
transform 1 0 21160 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input146
timestamp 1688980957
transform 1 0 22540 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input147
timestamp 1688980957
transform 1 0 20884 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input148
timestamp 1688980957
transform 1 0 22540 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input149
timestamp 1688980957
transform 1 0 22264 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input150
timestamp 1688980957
transform 1 0 17756 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input151
timestamp 1688980957
transform 1 0 21804 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input152
timestamp 1688980957
transform 1 0 20424 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input153
timestamp 1688980957
transform 1 0 9844 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input154
timestamp 1688980957
transform 1 0 10212 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input155
timestamp 1688980957
transform 1 0 10580 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input156
timestamp 1688980957
transform 1 0 10948 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input157
timestamp 1688980957
transform 1 0 11500 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input158
timestamp 1688980957
transform 1 0 11500 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input159
timestamp 1688980957
transform 1 0 11776 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input160
timestamp 1688980957
transform 1 0 12052 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input161
timestamp 1688980957
transform 1 0 12328 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input162
timestamp 1688980957
transform 1 0 12604 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input163
timestamp 1688980957
transform 1 0 12788 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input164
timestamp 1688980957
transform 1 0 13064 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input165
timestamp 1688980957
transform 1 0 13432 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input166
timestamp 1688980957
transform 1 0 13708 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input167
timestamp 1688980957
transform 1 0 14076 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input168
timestamp 1688980957
transform 1 0 14260 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input169
timestamp 1688980957
transform 1 0 14444 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input170
timestamp 1688980957
transform 1 0 14812 0 -1 43520
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input171
timestamp 1688980957
transform 1 0 15088 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input172
timestamp 1688980957
transform 1 0 15732 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input173
timestamp 1688980957
transform 1 0 16100 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input174
timestamp 1688980957
transform 1 0 19504 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input175
timestamp 1688980957
transform 1 0 19780 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input176
timestamp 1688980957
transform 1 0 20792 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input177
timestamp 1688980957
transform 1 0 19964 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input178
timestamp 1688980957
transform 1 0 20516 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input179
timestamp 1688980957
transform 1 0 21436 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input180
timestamp 1688980957
transform 1 0 16652 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input181
timestamp 1688980957
transform 1 0 17020 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input182
timestamp 1688980957
transform 1 0 17388 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input183
timestamp 1688980957
transform 1 0 17756 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input184
timestamp 1688980957
transform 1 0 18032 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input185
timestamp 1688980957
transform 1 0 18308 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input186
timestamp 1688980957
transform 1 0 18584 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input187
timestamp 1688980957
transform 1 0 18860 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input188
timestamp 1688980957
transform 1 0 19228 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  inst_clk_buf
timestamp 1688980957
transform 1 0 18676 0 -1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_1  Inst_Config_accessConfig_access__0_
timestamp 1688980957
transform 1 0 23644 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_Config_accessConfig_access__1_
timestamp 1688980957
transform 1 0 22540 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_Config_accessConfig_access__2_
timestamp 1688980957
transform 1 0 22264 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_Config_accessConfig_access__3_
timestamp 1688980957
transform 1 0 24012 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_A0_OutPass4_frame_config_mux__0_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 16928 0 1 16320
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_A0_OutPass4_frame_config_mux__1_
timestamp 1688980957
transform 1 0 20424 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_A0_OutPass4_frame_config_mux__2_
timestamp 1688980957
transform 1 0 21988 0 1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_A0_OutPass4_frame_config_mux__3_
timestamp 1688980957
transform 1 0 21804 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_A0_OutPass4_frame_config_mux_cus_mux21_inst0__2_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 18860 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_A0_OutPass4_frame_config_mux_cus_mux21_inst0__3_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 19504 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_A0_OutPass4_frame_config_mux_cus_mux21_inst0__4_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 18492 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_A0_OutPass4_frame_config_mux_cus_mux21_inst0_break_comb_loop_inst0__0_
timestamp 1688980957
transform 1 0 17388 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_A0_OutPass4_frame_config_mux_cus_mux21_inst0_break_comb_loop_inst1__0_
timestamp 1688980957
transform 1 0 19228 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_A0_OutPass4_frame_config_mux_cus_mux21_inst1__2_
timestamp 1688980957
transform 1 0 22080 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_A0_OutPass4_frame_config_mux_cus_mux21_inst1__3_
timestamp 1688980957
transform 1 0 22356 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_A0_OutPass4_frame_config_mux_cus_mux21_inst1__4_
timestamp 1688980957
transform 1 0 21712 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_A0_OutPass4_frame_config_mux_cus_mux21_inst1_break_comb_loop_inst0__0_
timestamp 1688980957
transform 1 0 20700 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_A0_OutPass4_frame_config_mux_cus_mux21_inst1_break_comb_loop_inst1__0_
timestamp 1688980957
transform 1 0 21804 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_A0_OutPass4_frame_config_mux_cus_mux21_inst2__2_
timestamp 1688980957
transform 1 0 22264 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_A0_OutPass4_frame_config_mux_cus_mux21_inst2__3_
timestamp 1688980957
transform 1 0 24012 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_A0_OutPass4_frame_config_mux_cus_mux21_inst2__4_
timestamp 1688980957
transform 1 0 23736 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_A0_OutPass4_frame_config_mux_cus_mux21_inst2_break_comb_loop_inst0__0_
timestamp 1688980957
transform 1 0 22540 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_A0_OutPass4_frame_config_mux_cus_mux21_inst2_break_comb_loop_inst1__0_
timestamp 1688980957
transform 1 0 22816 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_A0_OutPass4_frame_config_mux_cus_mux21_inst3__2_
timestamp 1688980957
transform 1 0 22908 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_A0_OutPass4_frame_config_mux_cus_mux21_inst3__3_
timestamp 1688980957
transform 1 0 22632 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_A0_OutPass4_frame_config_mux_cus_mux21_inst3__4_
timestamp 1688980957
transform 1 0 23828 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_A0_OutPass4_frame_config_mux_cus_mux21_inst3_break_comb_loop_inst0__0_
timestamp 1688980957
transform 1 0 22172 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_A0_OutPass4_frame_config_mux_cus_mux21_inst3_break_comb_loop_inst1__0_
timestamp 1688980957
transform 1 0 23276 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_A1_OutPass4_frame_config_mux__0_
timestamp 1688980957
transform 1 0 16928 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_A1_OutPass4_frame_config_mux__1_
timestamp 1688980957
transform 1 0 22264 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_A1_OutPass4_frame_config_mux__2_
timestamp 1688980957
transform 1 0 19136 0 -1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_A1_OutPass4_frame_config_mux__3_
timestamp 1688980957
transform 1 0 18860 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_A1_OutPass4_frame_config_mux_cus_mux21_inst0__2_
timestamp 1688980957
transform 1 0 18032 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_A1_OutPass4_frame_config_mux_cus_mux21_inst0__3_
timestamp 1688980957
transform 1 0 18676 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_A1_OutPass4_frame_config_mux_cus_mux21_inst0__4_
timestamp 1688980957
transform 1 0 19228 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_A1_OutPass4_frame_config_mux_cus_mux21_inst0_break_comb_loop_inst0__0_
timestamp 1688980957
transform 1 0 17480 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_A1_OutPass4_frame_config_mux_cus_mux21_inst0_break_comb_loop_inst1__0_
timestamp 1688980957
transform 1 0 18584 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_A1_OutPass4_frame_config_mux_cus_mux21_inst1__2_
timestamp 1688980957
transform 1 0 22632 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_A1_OutPass4_frame_config_mux_cus_mux21_inst1__3_
timestamp 1688980957
transform 1 0 22264 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_A1_OutPass4_frame_config_mux_cus_mux21_inst1__4_
timestamp 1688980957
transform 1 0 23736 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_A1_OutPass4_frame_config_mux_cus_mux21_inst1_break_comb_loop_inst0__0_
timestamp 1688980957
transform 1 0 22816 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_A1_OutPass4_frame_config_mux_cus_mux21_inst1_break_comb_loop_inst1__0_
timestamp 1688980957
transform 1 0 22540 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_A1_OutPass4_frame_config_mux_cus_mux21_inst2__2_
timestamp 1688980957
transform 1 0 20976 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_A1_OutPass4_frame_config_mux_cus_mux21_inst2__3_
timestamp 1688980957
transform 1 0 21252 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_A1_OutPass4_frame_config_mux_cus_mux21_inst2__4_
timestamp 1688980957
transform 1 0 20608 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_A1_OutPass4_frame_config_mux_cus_mux21_inst2_break_comb_loop_inst0__0_
timestamp 1688980957
transform 1 0 19596 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_A1_OutPass4_frame_config_mux_cus_mux21_inst2_break_comb_loop_inst1__0_
timestamp 1688980957
transform 1 0 20976 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_A1_OutPass4_frame_config_mux_cus_mux21_inst3__2_
timestamp 1688980957
transform 1 0 19964 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_A1_OutPass4_frame_config_mux_cus_mux21_inst3__3_
timestamp 1688980957
transform 1 0 20976 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_A1_OutPass4_frame_config_mux_cus_mux21_inst3__4_
timestamp 1688980957
transform 1 0 20332 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_A1_OutPass4_frame_config_mux_cus_mux21_inst3_break_comb_loop_inst0__0_
timestamp 1688980957
transform 1 0 19320 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_A1_OutPass4_frame_config_mux_cus_mux21_inst3_break_comb_loop_inst1__0_
timestamp 1688980957
transform 1 0 20700 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_C_OutPass4_frame_config_mux__0_
timestamp 1688980957
transform 1 0 20792 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_C_OutPass4_frame_config_mux__1_
timestamp 1688980957
transform 1 0 18860 0 -1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_C_OutPass4_frame_config_mux__2_
timestamp 1688980957
transform 1 0 18860 0 -1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_C_OutPass4_frame_config_mux__3_
timestamp 1688980957
transform 1 0 19228 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_C_OutPass4_frame_config_mux_cus_mux21_inst0__2_
timestamp 1688980957
transform 1 0 21988 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_C_OutPass4_frame_config_mux_cus_mux21_inst0__3_
timestamp 1688980957
transform 1 0 22080 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_C_OutPass4_frame_config_mux_cus_mux21_inst0__4_
timestamp 1688980957
transform 1 0 22448 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_C_OutPass4_frame_config_mux_cus_mux21_inst0_break_comb_loop_inst0__0_
timestamp 1688980957
transform 1 0 21344 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_C_OutPass4_frame_config_mux_cus_mux21_inst0_break_comb_loop_inst1__0_
timestamp 1688980957
transform 1 0 22356 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_C_OutPass4_frame_config_mux_cus_mux21_inst1__2_
timestamp 1688980957
transform 1 0 19872 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_C_OutPass4_frame_config_mux_cus_mux21_inst1__3_
timestamp 1688980957
transform 1 0 20792 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  Inst_FAB2RAM_C_OutPass4_frame_config_mux_cus_mux21_inst1__4_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 20148 0 1 31552
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_C_OutPass4_frame_config_mux_cus_mux21_inst1_break_comb_loop_inst0__0_
timestamp 1688980957
transform 1 0 19320 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_C_OutPass4_frame_config_mux_cus_mux21_inst1_break_comb_loop_inst1__0_
timestamp 1688980957
transform 1 0 21068 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_C_OutPass4_frame_config_mux_cus_mux21_inst2__2_
timestamp 1688980957
transform 1 0 19964 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_C_OutPass4_frame_config_mux_cus_mux21_inst2__3_
timestamp 1688980957
transform 1 0 20976 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  Inst_FAB2RAM_C_OutPass4_frame_config_mux_cus_mux21_inst2__4_
timestamp 1688980957
transform 1 0 20332 0 -1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_C_OutPass4_frame_config_mux_cus_mux21_inst2_break_comb_loop_inst0__0_
timestamp 1688980957
transform 1 0 19320 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_C_OutPass4_frame_config_mux_cus_mux21_inst2_break_comb_loop_inst1__0_
timestamp 1688980957
transform 1 0 20332 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_C_OutPass4_frame_config_mux_cus_mux21_inst3__2_
timestamp 1688980957
transform 1 0 19688 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_C_OutPass4_frame_config_mux_cus_mux21_inst3__3_
timestamp 1688980957
transform 1 0 20516 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_C_OutPass4_frame_config_mux_cus_mux21_inst3__4_
timestamp 1688980957
transform 1 0 20148 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_C_OutPass4_frame_config_mux_cus_mux21_inst3_break_comb_loop_inst0__0_
timestamp 1688980957
transform 1 0 18860 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_C_OutPass4_frame_config_mux_cus_mux21_inst3_break_comb_loop_inst1__0_
timestamp 1688980957
transform 1 0 20148 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_D0_OutPass4_frame_config_mux__0_
timestamp 1688980957
transform 1 0 22080 0 1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_D0_OutPass4_frame_config_mux__1_
timestamp 1688980957
transform 1 0 20240 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_D0_OutPass4_frame_config_mux__2_
timestamp 1688980957
transform 1 0 20792 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_D0_OutPass4_frame_config_mux__3_
timestamp 1688980957
transform 1 0 17296 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_D0_OutPass4_frame_config_mux_cus_mux21_inst0__2_
timestamp 1688980957
transform 1 0 24012 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_D0_OutPass4_frame_config_mux_cus_mux21_inst0__3_
timestamp 1688980957
transform 1 0 23276 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_D0_OutPass4_frame_config_mux_cus_mux21_inst0__4_
timestamp 1688980957
transform 1 0 23644 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D0_OutPass4_frame_config_mux_cus_mux21_inst0_break_comb_loop_inst0__0_
timestamp 1688980957
transform 1 0 22632 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D0_OutPass4_frame_config_mux_cus_mux21_inst0_break_comb_loop_inst1__0_
timestamp 1688980957
transform 1 0 24012 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_D0_OutPass4_frame_config_mux_cus_mux21_inst1__2_
timestamp 1688980957
transform 1 0 21804 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_D0_OutPass4_frame_config_mux_cus_mux21_inst1__3_
timestamp 1688980957
transform 1 0 22724 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_D0_OutPass4_frame_config_mux_cus_mux21_inst1__4_
timestamp 1688980957
transform 1 0 22172 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D0_OutPass4_frame_config_mux_cus_mux21_inst1_break_comb_loop_inst0__0_
timestamp 1688980957
transform 1 0 21068 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D0_OutPass4_frame_config_mux_cus_mux21_inst1_break_comb_loop_inst1__0_
timestamp 1688980957
transform 1 0 23000 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_D0_OutPass4_frame_config_mux_cus_mux21_inst2__2_
timestamp 1688980957
transform 1 0 22080 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_D0_OutPass4_frame_config_mux_cus_mux21_inst2__3_
timestamp 1688980957
transform 1 0 22632 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_D0_OutPass4_frame_config_mux_cus_mux21_inst2__4_
timestamp 1688980957
transform 1 0 23368 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D0_OutPass4_frame_config_mux_cus_mux21_inst2_break_comb_loop_inst0__0_
timestamp 1688980957
transform 1 0 21436 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D0_OutPass4_frame_config_mux_cus_mux21_inst2_break_comb_loop_inst1__0_
timestamp 1688980957
transform 1 0 22356 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_D0_OutPass4_frame_config_mux_cus_mux21_inst3__2_
timestamp 1688980957
transform 1 0 18216 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_D0_OutPass4_frame_config_mux_cus_mux21_inst3__3_
timestamp 1688980957
transform 1 0 18860 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_D0_OutPass4_frame_config_mux_cus_mux21_inst3__4_
timestamp 1688980957
transform 1 0 18492 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D0_OutPass4_frame_config_mux_cus_mux21_inst3_break_comb_loop_inst0__0_
timestamp 1688980957
transform 1 0 17664 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D0_OutPass4_frame_config_mux_cus_mux21_inst3_break_comb_loop_inst1__0_
timestamp 1688980957
transform 1 0 18768 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_D1_OutPass4_frame_config_mux__0_
timestamp 1688980957
transform 1 0 20240 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_D1_OutPass4_frame_config_mux__1_
timestamp 1688980957
transform 1 0 21988 0 -1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_D1_OutPass4_frame_config_mux__2_
timestamp 1688980957
transform 1 0 20240 0 1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_D1_OutPass4_frame_config_mux__3_
timestamp 1688980957
transform 1 0 18308 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_D1_OutPass4_frame_config_mux_cus_mux21_inst0__2_
timestamp 1688980957
transform 1 0 21344 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_D1_OutPass4_frame_config_mux_cus_mux21_inst0__3_
timestamp 1688980957
transform 1 0 22448 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_D1_OutPass4_frame_config_mux_cus_mux21_inst0__4_
timestamp 1688980957
transform 1 0 21804 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D1_OutPass4_frame_config_mux_cus_mux21_inst0_break_comb_loop_inst0__0_
timestamp 1688980957
transform 1 0 20700 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D1_OutPass4_frame_config_mux_cus_mux21_inst0_break_comb_loop_inst1__0_
timestamp 1688980957
transform 1 0 22172 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_D1_OutPass4_frame_config_mux_cus_mux21_inst1__2_
timestamp 1688980957
transform 1 0 23184 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_D1_OutPass4_frame_config_mux_cus_mux21_inst1__3_
timestamp 1688980957
transform 1 0 22908 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_D1_OutPass4_frame_config_mux_cus_mux21_inst1__4_
timestamp 1688980957
transform 1 0 23920 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D1_OutPass4_frame_config_mux_cus_mux21_inst1_break_comb_loop_inst0__0_
timestamp 1688980957
transform 1 0 22540 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D1_OutPass4_frame_config_mux_cus_mux21_inst1_break_comb_loop_inst1__0_
timestamp 1688980957
transform 1 0 23460 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_D1_OutPass4_frame_config_mux_cus_mux21_inst2__2_
timestamp 1688980957
transform 1 0 21252 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_D1_OutPass4_frame_config_mux_cus_mux21_inst2__3_
timestamp 1688980957
transform 1 0 22172 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_D1_OutPass4_frame_config_mux_cus_mux21_inst2__4_
timestamp 1688980957
transform 1 0 21804 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D1_OutPass4_frame_config_mux_cus_mux21_inst2_break_comb_loop_inst0__0_
timestamp 1688980957
transform 1 0 20700 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D1_OutPass4_frame_config_mux_cus_mux21_inst2_break_comb_loop_inst1__0_
timestamp 1688980957
transform 1 0 21712 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_D1_OutPass4_frame_config_mux_cus_mux21_inst3__2_
timestamp 1688980957
transform 1 0 19412 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_D1_OutPass4_frame_config_mux_cus_mux21_inst3__3_
timestamp 1688980957
transform 1 0 20332 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_D1_OutPass4_frame_config_mux_cus_mux21_inst3__4_
timestamp 1688980957
transform 1 0 19780 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D1_OutPass4_frame_config_mux_cus_mux21_inst3_break_comb_loop_inst0__0_
timestamp 1688980957
transform 1 0 18768 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D1_OutPass4_frame_config_mux_cus_mux21_inst3_break_comb_loop_inst1__0_
timestamp 1688980957
transform 1 0 19872 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_D2_OutPass4_frame_config_mux__0_
timestamp 1688980957
transform 1 0 17112 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_D2_OutPass4_frame_config_mux__1_
timestamp 1688980957
transform 1 0 20240 0 -1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_D2_OutPass4_frame_config_mux__2_
timestamp 1688980957
transform 1 0 18952 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_D2_OutPass4_frame_config_mux__3_
timestamp 1688980957
transform 1 0 17204 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_D2_OutPass4_frame_config_mux_cus_mux21_inst0__2_
timestamp 1688980957
transform 1 0 18584 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_D2_OutPass4_frame_config_mux_cus_mux21_inst0__3_
timestamp 1688980957
transform 1 0 19136 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_D2_OutPass4_frame_config_mux_cus_mux21_inst0__4_
timestamp 1688980957
transform 1 0 18584 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D2_OutPass4_frame_config_mux_cus_mux21_inst0_break_comb_loop_inst0__0_
timestamp 1688980957
transform 1 0 17296 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D2_OutPass4_frame_config_mux_cus_mux21_inst0_break_comb_loop_inst1__0_
timestamp 1688980957
transform 1 0 18860 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_D2_OutPass4_frame_config_mux_cus_mux21_inst1__2_
timestamp 1688980957
transform 1 0 22080 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_D2_OutPass4_frame_config_mux_cus_mux21_inst1__3_
timestamp 1688980957
transform 1 0 22816 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_D2_OutPass4_frame_config_mux_cus_mux21_inst1__4_
timestamp 1688980957
transform 1 0 22448 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D2_OutPass4_frame_config_mux_cus_mux21_inst1_break_comb_loop_inst0__0_
timestamp 1688980957
transform 1 0 21804 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D2_OutPass4_frame_config_mux_cus_mux21_inst1_break_comb_loop_inst1__0_
timestamp 1688980957
transform 1 0 22356 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_D2_OutPass4_frame_config_mux_cus_mux21_inst2__2_
timestamp 1688980957
transform 1 0 20792 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_D2_OutPass4_frame_config_mux_cus_mux21_inst2__3_
timestamp 1688980957
transform 1 0 21068 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_D2_OutPass4_frame_config_mux_cus_mux21_inst2__4_
timestamp 1688980957
transform 1 0 20424 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D2_OutPass4_frame_config_mux_cus_mux21_inst2_break_comb_loop_inst0__0_
timestamp 1688980957
transform 1 0 19504 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D2_OutPass4_frame_config_mux_cus_mux21_inst2_break_comb_loop_inst1__0_
timestamp 1688980957
transform 1 0 20424 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_D2_OutPass4_frame_config_mux_cus_mux21_inst3__2_
timestamp 1688980957
transform 1 0 18308 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_D2_OutPass4_frame_config_mux_cus_mux21_inst3__3_
timestamp 1688980957
transform 1 0 19596 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_D2_OutPass4_frame_config_mux_cus_mux21_inst3__4_
timestamp 1688980957
transform 1 0 19228 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D2_OutPass4_frame_config_mux_cus_mux21_inst3_break_comb_loop_inst0__0_
timestamp 1688980957
transform 1 0 17664 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D2_OutPass4_frame_config_mux_cus_mux21_inst3_break_comb_loop_inst1__0_
timestamp 1688980957
transform 1 0 18768 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_D3_OutPass4_frame_config_mux__0_
timestamp 1688980957
transform 1 0 19228 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_D3_OutPass4_frame_config_mux__1_
timestamp 1688980957
transform 1 0 22172 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_D3_OutPass4_frame_config_mux__2_
timestamp 1688980957
transform 1 0 20056 0 1 20672
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_D3_OutPass4_frame_config_mux__3_
timestamp 1688980957
transform 1 0 18124 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_D3_OutPass4_frame_config_mux_cus_mux21_inst0__2_
timestamp 1688980957
transform 1 0 20056 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_D3_OutPass4_frame_config_mux_cus_mux21_inst0__3_
timestamp 1688980957
transform 1 0 21068 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_D3_OutPass4_frame_config_mux_cus_mux21_inst0__4_
timestamp 1688980957
transform 1 0 20700 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D3_OutPass4_frame_config_mux_cus_mux21_inst0_break_comb_loop_inst0__0_
timestamp 1688980957
transform 1 0 19412 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D3_OutPass4_frame_config_mux_cus_mux21_inst0_break_comb_loop_inst1__0_
timestamp 1688980957
transform 1 0 21344 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_D3_OutPass4_frame_config_mux_cus_mux21_inst1__2_
timestamp 1688980957
transform 1 0 23368 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_D3_OutPass4_frame_config_mux_cus_mux21_inst1__3_
timestamp 1688980957
transform 1 0 23092 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_D3_OutPass4_frame_config_mux_cus_mux21_inst1__4_
timestamp 1688980957
transform 1 0 23920 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D3_OutPass4_frame_config_mux_cus_mux21_inst1_break_comb_loop_inst0__0_
timestamp 1688980957
transform 1 0 22724 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D3_OutPass4_frame_config_mux_cus_mux21_inst1_break_comb_loop_inst1__0_
timestamp 1688980957
transform 1 0 23644 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_D3_OutPass4_frame_config_mux_cus_mux21_inst2__2_
timestamp 1688980957
transform 1 0 21160 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_D3_OutPass4_frame_config_mux_cus_mux21_inst2__3_
timestamp 1688980957
transform 1 0 22080 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_D3_OutPass4_frame_config_mux_cus_mux21_inst2__4_
timestamp 1688980957
transform 1 0 22080 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D3_OutPass4_frame_config_mux_cus_mux21_inst2_break_comb_loop_inst0__0_
timestamp 1688980957
transform 1 0 20608 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D3_OutPass4_frame_config_mux_cus_mux21_inst2_break_comb_loop_inst1__0_
timestamp 1688980957
transform 1 0 21804 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_D3_OutPass4_frame_config_mux_cus_mux21_inst3__2_
timestamp 1688980957
transform 1 0 18860 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_D3_OutPass4_frame_config_mux_cus_mux21_inst3__3_
timestamp 1688980957
transform 1 0 20608 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_D3_OutPass4_frame_config_mux_cus_mux21_inst3__4_
timestamp 1688980957
transform 1 0 19596 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D3_OutPass4_frame_config_mux_cus_mux21_inst3_break_comb_loop_inst0__0_
timestamp 1688980957
transform 1 0 18584 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D3_OutPass4_frame_config_mux_cus_mux21_inst3_break_comb_loop_inst1__0_
timestamp 1688980957
transform 1 0 19596 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  Inst_RAM2FAB_D0_InPass4_frame_config_mux__0_
timestamp 1688980957
transform 1 0 16928 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_RAM2FAB_D0_InPass4_frame_config_mux__1_
timestamp 1688980957
transform 1 0 17572 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_RAM2FAB_D0_InPass4_frame_config_mux__2_
timestamp 1688980957
transform 1 0 22264 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_RAM2FAB_D0_InPass4_frame_config_mux__3_
timestamp 1688980957
transform 1 0 19228 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  Inst_RAM2FAB_D0_InPass4_frame_config_mux_cus_mux21_inst0__2_
timestamp 1688980957
transform 1 0 16376 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM2FAB_D0_InPass4_frame_config_mux_cus_mux21_inst0__3_
timestamp 1688980957
transform 1 0 18032 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_4  Inst_RAM2FAB_D0_InPass4_frame_config_mux_cus_mux21_inst0__4_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 17020 0 -1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D0_InPass4_frame_config_mux_cus_mux21_inst0_break_comb_loop_inst0__0_
timestamp 1688980957
transform 1 0 16652 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D0_InPass4_frame_config_mux_cus_mux21_inst0_break_comb_loop_inst1__0_
timestamp 1688980957
transform 1 0 18400 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_RAM2FAB_D0_InPass4_frame_config_mux_cus_mux21_inst1__2_
timestamp 1688980957
transform 1 0 18032 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM2FAB_D0_InPass4_frame_config_mux_cus_mux21_inst1__3_
timestamp 1688980957
transform 1 0 18308 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_4  Inst_RAM2FAB_D0_InPass4_frame_config_mux_cus_mux21_inst1__4_
timestamp 1688980957
transform 1 0 17848 0 1 9792
box -38 -48 1234 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D0_InPass4_frame_config_mux_cus_mux21_inst1_break_comb_loop_inst0__0_
timestamp 1688980957
transform 1 0 18584 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D0_InPass4_frame_config_mux_cus_mux21_inst1_break_comb_loop_inst1__0_
timestamp 1688980957
transform 1 0 18860 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_RAM2FAB_D0_InPass4_frame_config_mux_cus_mux21_inst2__2_
timestamp 1688980957
transform 1 0 21988 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM2FAB_D0_InPass4_frame_config_mux_cus_mux21_inst2__3_
timestamp 1688980957
transform 1 0 23092 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_4  Inst_RAM2FAB_D0_InPass4_frame_config_mux_cus_mux21_inst2__4_
timestamp 1688980957
transform 1 0 22172 0 1 8704
box -38 -48 1234 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D0_InPass4_frame_config_mux_cus_mux21_inst2_break_comb_loop_inst0__0_
timestamp 1688980957
transform 1 0 22816 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D0_InPass4_frame_config_mux_cus_mux21_inst2_break_comb_loop_inst1__0_
timestamp 1688980957
transform 1 0 23736 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_RAM2FAB_D0_InPass4_frame_config_mux_cus_mux21_inst3__2_
timestamp 1688980957
transform 1 0 19504 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM2FAB_D0_InPass4_frame_config_mux_cus_mux21_inst3__3_
timestamp 1688980957
transform 1 0 19780 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_4  Inst_RAM2FAB_D0_InPass4_frame_config_mux_cus_mux21_inst3__4_
timestamp 1688980957
transform 1 0 19964 0 -1 9792
box -38 -48 1234 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D0_InPass4_frame_config_mux_cus_mux21_inst3_break_comb_loop_inst0__0_
timestamp 1688980957
transform 1 0 19780 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D0_InPass4_frame_config_mux_cus_mux21_inst3_break_comb_loop_inst1__0_
timestamp 1688980957
transform 1 0 20148 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  Inst_RAM2FAB_D1_InPass4_frame_config_mux__0_
timestamp 1688980957
transform 1 0 17388 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_RAM2FAB_D1_InPass4_frame_config_mux__1_
timestamp 1688980957
transform 1 0 21160 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_RAM2FAB_D1_InPass4_frame_config_mux__2_
timestamp 1688980957
transform 1 0 20792 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_RAM2FAB_D1_InPass4_frame_config_mux__3_
timestamp 1688980957
transform 1 0 18584 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  Inst_RAM2FAB_D1_InPass4_frame_config_mux_cus_mux21_inst0__2_
timestamp 1688980957
transform 1 0 17940 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM2FAB_D1_InPass4_frame_config_mux_cus_mux21_inst0__3_
timestamp 1688980957
transform 1 0 18400 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  Inst_RAM2FAB_D1_InPass4_frame_config_mux_cus_mux21_inst0__4_
timestamp 1688980957
transform 1 0 17756 0 1 11968
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D1_InPass4_frame_config_mux_cus_mux21_inst0_break_comb_loop_inst0__0_
timestamp 1688980957
transform 1 0 17112 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D1_InPass4_frame_config_mux_cus_mux21_inst0_break_comb_loop_inst1__0_
timestamp 1688980957
transform 1 0 18860 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_RAM2FAB_D1_InPass4_frame_config_mux_cus_mux21_inst1__2_
timestamp 1688980957
transform 1 0 21804 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM2FAB_D1_InPass4_frame_config_mux_cus_mux21_inst1__3_
timestamp 1688980957
transform 1 0 21804 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_4  Inst_RAM2FAB_D1_InPass4_frame_config_mux_cus_mux21_inst1__4_
timestamp 1688980957
transform 1 0 21252 0 1 11968
box -38 -48 1234 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D1_InPass4_frame_config_mux_cus_mux21_inst1_break_comb_loop_inst0__0_
timestamp 1688980957
transform 1 0 22080 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D1_InPass4_frame_config_mux_cus_mux21_inst1_break_comb_loop_inst1__0_
timestamp 1688980957
transform 1 0 22172 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_RAM2FAB_D1_InPass4_frame_config_mux_cus_mux21_inst2__2_
timestamp 1688980957
transform 1 0 20884 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM2FAB_D1_InPass4_frame_config_mux_cus_mux21_inst2__3_
timestamp 1688980957
transform 1 0 21804 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_4  Inst_RAM2FAB_D1_InPass4_frame_config_mux_cus_mux21_inst2__4_
timestamp 1688980957
transform 1 0 20608 0 1 6528
box -38 -48 1234 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D1_InPass4_frame_config_mux_cus_mux21_inst2_break_comb_loop_inst0__0_
timestamp 1688980957
transform 1 0 20332 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D1_InPass4_frame_config_mux_cus_mux21_inst2_break_comb_loop_inst1__0_
timestamp 1688980957
transform 1 0 22080 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_RAM2FAB_D1_InPass4_frame_config_mux_cus_mux21_inst3__2_
timestamp 1688980957
transform 1 0 19228 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM2FAB_D1_InPass4_frame_config_mux_cus_mux21_inst3__3_
timestamp 1688980957
transform 1 0 20056 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_4  Inst_RAM2FAB_D1_InPass4_frame_config_mux_cus_mux21_inst3__4_
timestamp 1688980957
transform 1 0 19228 0 1 5440
box -38 -48 1234 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D1_InPass4_frame_config_mux_cus_mux21_inst3_break_comb_loop_inst0__0_
timestamp 1688980957
transform 1 0 18308 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D1_InPass4_frame_config_mux_cus_mux21_inst3_break_comb_loop_inst1__0_
timestamp 1688980957
transform 1 0 20332 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  Inst_RAM2FAB_D2_InPass4_frame_config_mux__0_
timestamp 1688980957
transform 1 0 19228 0 -1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_RAM2FAB_D2_InPass4_frame_config_mux__1_
timestamp 1688980957
transform 1 0 20424 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_RAM2FAB_D2_InPass4_frame_config_mux__2_
timestamp 1688980957
transform 1 0 19136 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_RAM2FAB_D2_InPass4_frame_config_mux__3_
timestamp 1688980957
transform 1 0 20700 0 1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  Inst_RAM2FAB_D2_InPass4_frame_config_mux_cus_mux21_inst0__2_
timestamp 1688980957
transform 1 0 19228 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM2FAB_D2_InPass4_frame_config_mux_cus_mux21_inst0__3_
timestamp 1688980957
transform 1 0 16744 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  Inst_RAM2FAB_D2_InPass4_frame_config_mux_cus_mux21_inst0__4_
timestamp 1688980957
transform 1 0 19228 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D2_InPass4_frame_config_mux_cus_mux21_inst0_break_comb_loop_inst0__0_
timestamp 1688980957
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D2_InPass4_frame_config_mux_cus_mux21_inst0_break_comb_loop_inst1__0_
timestamp 1688980957
transform 1 0 19872 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_RAM2FAB_D2_InPass4_frame_config_mux_cus_mux21_inst1__2_
timestamp 1688980957
transform 1 0 20148 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM2FAB_D2_InPass4_frame_config_mux_cus_mux21_inst1__3_
timestamp 1688980957
transform 1 0 21436 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_4  Inst_RAM2FAB_D2_InPass4_frame_config_mux_cus_mux21_inst1__4_
timestamp 1688980957
transform 1 0 21804 0 -1 5440
box -38 -48 1234 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D2_InPass4_frame_config_mux_cus_mux21_inst1_break_comb_loop_inst0__0_
timestamp 1688980957
transform 1 0 19136 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D2_InPass4_frame_config_mux_cus_mux21_inst1_break_comb_loop_inst1__0_
timestamp 1688980957
transform 1 0 19320 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_RAM2FAB_D2_InPass4_frame_config_mux_cus_mux21_inst2__2_
timestamp 1688980957
transform 1 0 18860 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM2FAB_D2_InPass4_frame_config_mux_cus_mux21_inst2__3_
timestamp 1688980957
transform 1 0 20608 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  Inst_RAM2FAB_D2_InPass4_frame_config_mux_cus_mux21_inst2__4_
timestamp 1688980957
transform 1 0 19412 0 -1 13056
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D2_InPass4_frame_config_mux_cus_mux21_inst2_break_comb_loop_inst0__0_
timestamp 1688980957
transform 1 0 19504 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D2_InPass4_frame_config_mux_cus_mux21_inst2_break_comb_loop_inst1__0_
timestamp 1688980957
transform 1 0 20608 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_RAM2FAB_D2_InPass4_frame_config_mux_cus_mux21_inst3__2_
timestamp 1688980957
transform 1 0 21160 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM2FAB_D2_InPass4_frame_config_mux_cus_mux21_inst3__3_
timestamp 1688980957
transform 1 0 21436 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  Inst_RAM2FAB_D2_InPass4_frame_config_mux_cus_mux21_inst3__4_
timestamp 1688980957
transform 1 0 20700 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D2_InPass4_frame_config_mux_cus_mux21_inst3_break_comb_loop_inst0__0_
timestamp 1688980957
transform 1 0 20792 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D2_InPass4_frame_config_mux_cus_mux21_inst3_break_comb_loop_inst1__0_
timestamp 1688980957
transform 1 0 21804 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  Inst_RAM2FAB_D3_InPass4_frame_config_mux__0_
timestamp 1688980957
transform 1 0 17296 0 1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_RAM2FAB_D3_InPass4_frame_config_mux__1_
timestamp 1688980957
transform 1 0 22816 0 1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_RAM2FAB_D3_InPass4_frame_config_mux__2_
timestamp 1688980957
transform 1 0 22724 0 -1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_RAM2FAB_D3_InPass4_frame_config_mux__3_
timestamp 1688980957
transform 1 0 21804 0 -1 2176
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  Inst_RAM2FAB_D3_InPass4_frame_config_mux_cus_mux21_inst0__2_
timestamp 1688980957
transform 1 0 17664 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM2FAB_D3_InPass4_frame_config_mux_cus_mux21_inst0__3_
timestamp 1688980957
transform 1 0 17388 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  Inst_RAM2FAB_D3_InPass4_frame_config_mux_cus_mux21_inst0__4_
timestamp 1688980957
transform 1 0 17664 0 -1 4352
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D3_InPass4_frame_config_mux_cus_mux21_inst0_break_comb_loop_inst0__0_
timestamp 1688980957
transform 1 0 17296 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D3_InPass4_frame_config_mux_cus_mux21_inst0_break_comb_loop_inst1__0_
timestamp 1688980957
transform 1 0 20056 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_RAM2FAB_D3_InPass4_frame_config_mux_cus_mux21_inst1__2_
timestamp 1688980957
transform 1 0 23460 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM2FAB_D3_InPass4_frame_config_mux_cus_mux21_inst1__3_
timestamp 1688980957
transform 1 0 23736 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_4  Inst_RAM2FAB_D3_InPass4_frame_config_mux_cus_mux21_inst1__4_
timestamp 1688980957
transform 1 0 22908 0 1 6528
box -38 -48 1234 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D3_InPass4_frame_config_mux_cus_mux21_inst1_break_comb_loop_inst0__0_
timestamp 1688980957
transform 1 0 23092 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D3_InPass4_frame_config_mux_cus_mux21_inst1_break_comb_loop_inst1__0_
timestamp 1688980957
transform 1 0 23644 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_RAM2FAB_D3_InPass4_frame_config_mux_cus_mux21_inst2__2_
timestamp 1688980957
transform 1 0 18860 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM2FAB_D3_InPass4_frame_config_mux_cus_mux21_inst2__3_
timestamp 1688980957
transform 1 0 20516 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_4  Inst_RAM2FAB_D3_InPass4_frame_config_mux_cus_mux21_inst2__4_
timestamp 1688980957
transform 1 0 22908 0 1 3264
box -38 -48 1234 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D3_InPass4_frame_config_mux_cus_mux21_inst2_break_comb_loop_inst0__0_
timestamp 1688980957
transform 1 0 21804 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D3_InPass4_frame_config_mux_cus_mux21_inst2_break_comb_loop_inst1__0_
timestamp 1688980957
transform 1 0 15824 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_RAM2FAB_D3_InPass4_frame_config_mux_cus_mux21_inst3__2_
timestamp 1688980957
transform 1 0 17112 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM2FAB_D3_InPass4_frame_config_mux_cus_mux21_inst3__3_
timestamp 1688980957
transform 1 0 21160 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  Inst_RAM2FAB_D3_InPass4_frame_config_mux_cus_mux21_inst3__4_
timestamp 1688980957
transform 1 0 22080 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__buf_1  Inst_RAM2FAB_D3_InPass4_frame_config_mux_cus_mux21_inst3_break_comb_loop_inst0__0_
timestamp 1688980957
transform 1 0 21436 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D3_InPass4_frame_config_mux_cus_mux21_inst3_break_comb_loop_inst1__0_
timestamp 1688980957
transform 1 0 19596 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame0_bit0 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 9108 0 1 4352
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame0_bit1
timestamp 1688980957
transform 1 0 9936 0 1 5440
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame0_bit2
timestamp 1688980957
transform 1 0 2944 0 -1 41344
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame0_bit3
timestamp 1688980957
transform 1 0 4140 0 -1 42432
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame0_bit4
timestamp 1688980957
transform 1 0 2300 0 1 35904
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame0_bit5
timestamp 1688980957
transform 1 0 3772 0 1 38080
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame0_bit6
timestamp 1688980957
transform 1 0 10948 0 1 7616
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame0_bit7
timestamp 1688980957
transform 1 0 11224 0 1 6528
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame0_bit8
timestamp 1688980957
transform 1 0 9568 0 1 1088
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame0_bit9
timestamp 1688980957
transform 1 0 10028 0 -1 2176
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame0_bit10
timestamp 1688980957
transform 1 0 9200 0 1 38080
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame0_bit11
timestamp 1688980957
transform 1 0 9844 0 1 39168
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame0_bit12
timestamp 1688980957
transform 1 0 3956 0 -1 30464
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame0_bit13
timestamp 1688980957
transform 1 0 4876 0 -1 31552
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame0_bit14
timestamp 1688980957
transform 1 0 10028 0 -1 33728
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame0_bit15
timestamp 1688980957
transform 1 0 11224 0 1 33728
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame0_bit16
timestamp 1688980957
transform 1 0 10856 0 1 3264
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame0_bit17
timestamp 1688980957
transform 1 0 11500 0 -1 4352
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame0_bit18
timestamp 1688980957
transform 1 0 6900 0 -1 19584
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame0_bit19
timestamp 1688980957
transform 1 0 7544 0 -1 20672
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame0_bit20
timestamp 1688980957
transform 1 0 10028 0 -1 30464
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame0_bit21
timestamp 1688980957
transform 1 0 10672 0 1 30464
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame0_bit22
timestamp 1688980957
transform 1 0 11592 0 -1 3264
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame0_bit23
timestamp 1688980957
transform 1 0 12328 0 -1 2176
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame0_bit24
timestamp 1688980957
transform 1 0 8924 0 1 13056
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame0_bit25
timestamp 1688980957
transform 1 0 9568 0 1 11968
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame0_bit26
timestamp 1688980957
transform 1 0 3772 0 -1 43520
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame0_bit27
timestamp 1688980957
transform 1 0 2300 0 1 41344
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame0_bit28
timestamp 1688980957
transform 1 0 2300 0 1 39168
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame0_bit29
timestamp 1688980957
transform 1 0 2944 0 -1 38080
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame0_bit30
timestamp 1688980957
transform 1 0 12420 0 1 28288
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame0_bit31
timestamp 1688980957
transform 1 0 13156 0 -1 28288
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame1_bit0
timestamp 1688980957
transform 1 0 10028 0 -1 14144
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame1_bit1
timestamp 1688980957
transform 1 0 10948 0 1 13056
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame1_bit2
timestamp 1688980957
transform 1 0 6808 0 -1 42432
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame1_bit3
timestamp 1688980957
transform 1 0 7452 0 1 41344
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame1_bit4
timestamp 1688980957
transform 1 0 10396 0 1 35904
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame1_bit5
timestamp 1688980957
transform 1 0 11132 0 1 34816
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame1_bit6
timestamp 1688980957
transform 1 0 15732 0 1 29376
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame1_bit7
timestamp 1688980957
transform 1 0 17112 0 1 29376
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame1_bit8
timestamp 1688980957
transform 1 0 7544 0 -1 3264
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame1_bit9
timestamp 1688980957
transform 1 0 8924 0 -1 3264
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame1_bit10
timestamp 1688980957
transform 1 0 3956 0 -1 40256
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame1_bit11
timestamp 1688980957
transform 1 0 4876 0 -1 39168
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame1_bit12
timestamp 1688980957
transform 1 0 2300 0 1 28288
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame1_bit13
timestamp 1688980957
transform 1 0 3404 0 -1 29376
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame1_bit14
timestamp 1688980957
transform 1 0 12052 0 1 14144
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame1_bit15
timestamp 1688980957
transform 1 0 12604 0 1 13056
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame1_bit16
timestamp 1688980957
transform 1 0 8924 0 1 9792
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame1_bit17
timestamp 1688980957
transform 1 0 9568 0 1 8704
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame1_bit18
timestamp 1688980957
transform 1 0 4324 0 -1 38080
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame1_bit19
timestamp 1688980957
transform 1 0 4876 0 -1 36992
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame1_bit20
timestamp 1688980957
transform 1 0 2300 0 1 31552
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame1_bit21
timestamp 1688980957
transform 1 0 3772 0 1 31552
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame1_bit22
timestamp 1688980957
transform 1 0 11408 0 1 8704
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame1_bit23
timestamp 1688980957
transform 1 0 12328 0 -1 9792
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame1_bit24
timestamp 1688980957
transform 1 0 9108 0 1 7616
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame1_bit25
timestamp 1688980957
transform 1 0 9844 0 1 6528
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame1_bit26
timestamp 1688980957
transform 1 0 4048 0 1 42432
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame1_bit27
timestamp 1688980957
transform 1 0 5428 0 1 42432
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame1_bit28
timestamp 1688980957
transform 1 0 3128 0 -1 34816
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame1_bit29
timestamp 1688980957
transform 1 0 4232 0 -1 33728
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame1_bit30
timestamp 1688980957
transform 1 0 12604 0 1 6528
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame1_bit31
timestamp 1688980957
transform 1 0 13156 0 -1 6528
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame2_bit0
timestamp 1688980957
transform 1 0 11592 0 -1 23936
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame2_bit1
timestamp 1688980957
transform 1 0 12236 0 -1 27200
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame2_bit2
timestamp 1688980957
transform 1 0 6716 0 1 34816
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame2_bit3
timestamp 1688980957
transform 1 0 6624 0 -1 34816
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame2_bit4
timestamp 1688980957
transform 1 0 4876 0 1 29376
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame2_bit5
timestamp 1688980957
transform 1 0 6348 0 -1 29376
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame2_bit6
timestamp 1688980957
transform 1 0 14904 0 1 31552
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame2_bit7
timestamp 1688980957
transform 1 0 16284 0 1 31552
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame2_bit8
timestamp 1688980957
transform 1 0 12236 0 -1 25024
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame2_bit9
timestamp 1688980957
transform 1 0 13892 0 -1 26112
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame2_bit10
timestamp 1688980957
transform 1 0 6348 0 -1 23936
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame2_bit11
timestamp 1688980957
transform 1 0 8004 0 -1 25024
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame2_bit12
timestamp 1688980957
transform 1 0 7452 0 1 26112
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame2_bit13
timestamp 1688980957
transform 1 0 8740 0 -1 27200
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame2_bit14
timestamp 1688980957
transform 1 0 15180 0 -1 23936
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame2_bit15
timestamp 1688980957
transform 1 0 16100 0 1 22848
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame2_bit16
timestamp 1688980957
transform 1 0 14352 0 1 16320
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame2_bit17
timestamp 1688980957
transform 1 0 15088 0 -1 16320
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame2_bit18
timestamp 1688980957
transform 1 0 9844 0 1 17408
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame2_bit19
timestamp 1688980957
transform 1 0 11500 0 -1 17408
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame2_bit20
timestamp 1688980957
transform 1 0 8648 0 -1 19584
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame2_bit21
timestamp 1688980957
transform 1 0 9384 0 -1 18496
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame2_bit22
timestamp 1688980957
transform 1 0 14444 0 -1 20672
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame2_bit23
timestamp 1688980957
transform 1 0 14904 0 -1 19584
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame2_bit24
timestamp 1688980957
transform 1 0 11868 0 1 16320
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame2_bit25
timestamp 1688980957
transform 1 0 12604 0 1 15232
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame2_bit26
timestamp 1688980957
transform 1 0 7084 0 -1 15232
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame2_bit27
timestamp 1688980957
transform 1 0 8924 0 1 14144
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame2_bit28
timestamp 1688980957
transform 1 0 9292 0 1 19584
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame2_bit29
timestamp 1688980957
transform 1 0 10856 0 1 18496
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame2_bit30
timestamp 1688980957
transform 1 0 15180 0 -1 21760
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame2_bit31
timestamp 1688980957
transform 1 0 16652 0 -1 21760
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame3_bit0
timestamp 1688980957
transform 1 0 13892 0 -1 11968
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame3_bit1
timestamp 1688980957
transform 1 0 14536 0 -1 13056
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame3_bit2
timestamp 1688980957
transform 1 0 4876 0 -1 14144
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame3_bit3
timestamp 1688980957
transform 1 0 6348 0 -1 11968
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame3_bit4
timestamp 1688980957
transform 1 0 6348 0 -1 17408
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame3_bit5
timestamp 1688980957
transform 1 0 6624 0 -1 16320
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame3_bit6
timestamp 1688980957
transform 1 0 7452 0 1 10880
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame3_bit7
timestamp 1688980957
transform 1 0 8924 0 1 10880
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame3_bit8
timestamp 1688980957
transform 1 0 14076 0 1 14144
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame3_bit9
timestamp 1688980957
transform 1 0 14536 0 1 15232
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame3_bit10
timestamp 1688980957
transform 1 0 4876 0 -1 19584
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame3_bit11
timestamp 1688980957
transform 1 0 5796 0 1 19584
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame3_bit12
timestamp 1688980957
transform 1 0 4876 0 -1 22848
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame3_bit13
timestamp 1688980957
transform 1 0 6992 0 1 20672
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame3_bit14
timestamp 1688980957
transform 1 0 6808 0 -1 13056
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame3_bit15
timestamp 1688980957
transform 1 0 7360 0 1 14144
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame3_bit16
timestamp 1688980957
transform 1 0 11500 0 -1 26112
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame3_bit17
timestamp 1688980957
transform 1 0 11868 0 1 26112
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame3_bit18
timestamp 1688980957
transform 1 0 4876 0 -1 32640
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame3_bit19
timestamp 1688980957
transform 1 0 6348 0 1 30464
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame3_bit20
timestamp 1688980957
transform 1 0 5428 0 1 28288
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame3_bit21
timestamp 1688980957
transform 1 0 5060 0 1 27200
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame3_bit22
timestamp 1688980957
transform 1 0 14628 0 1 28288
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame3_bit23
timestamp 1688980957
transform 1 0 15456 0 1 27200
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame3_bit24
timestamp 1688980957
transform 1 0 14076 0 1 27200
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame3_bit25
timestamp 1688980957
transform 1 0 14536 0 1 26112
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame3_bit26
timestamp 1688980957
transform 1 0 4876 0 -1 26112
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame3_bit27
timestamp 1688980957
transform 1 0 5612 0 1 25024
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame3_bit28
timestamp 1688980957
transform 1 0 6072 0 1 26112
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame3_bit29
timestamp 1688980957
transform 1 0 6992 0 1 27200
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame3_bit30
timestamp 1688980957
transform 1 0 16008 0 1 25024
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame3_bit31
timestamp 1688980957
transform 1 0 16652 0 -1 26112
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame4_bit0
timestamp 1688980957
transform 1 0 13432 0 -1 10880
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame4_bit1
timestamp 1688980957
transform 1 0 14076 0 -1 9792
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame4_bit2
timestamp 1688980957
transform 1 0 4692 0 -1 10880
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame4_bit3
timestamp 1688980957
transform 1 0 5428 0 1 11968
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame4_bit4
timestamp 1688980957
transform 1 0 1932 0 -1 17408
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame4_bit5
timestamp 1688980957
transform 1 0 3312 0 -1 17408
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame4_bit6
timestamp 1688980957
transform 1 0 7268 0 1 7616
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame4_bit7
timestamp 1688980957
transform 1 0 8004 0 -1 8704
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame4_bit8
timestamp 1688980957
transform 1 0 15180 0 -1 10880
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame4_bit9
timestamp 1688980957
transform 1 0 16652 0 -1 10880
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame4_bit10
timestamp 1688980957
transform 1 0 1932 0 -1 10880
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame4_bit11
timestamp 1688980957
transform 1 0 3312 0 -1 10880
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame4_bit12
timestamp 1688980957
transform 1 0 4508 0 1 15232
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame4_bit13
timestamp 1688980957
transform 1 0 4876 0 -1 17408
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame4_bit14
timestamp 1688980957
transform 1 0 7452 0 1 8704
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame4_bit15
timestamp 1688980957
transform 1 0 7268 0 -1 9792
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame4_bit16
timestamp 1688980957
transform 1 0 15180 0 -1 14144
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame4_bit17
timestamp 1688980957
transform 1 0 16652 0 -1 14144
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame4_bit18
timestamp 1688980957
transform 1 0 3220 0 -1 19584
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame4_bit19
timestamp 1688980957
transform 1 0 3772 0 1 18496
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame4_bit20
timestamp 1688980957
transform 1 0 3312 0 -1 22848
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame4_bit21
timestamp 1688980957
transform 1 0 3956 0 1 21760
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame4_bit22
timestamp 1688980957
transform 1 0 4876 0 -1 3264
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame4_bit23
timestamp 1688980957
transform 1 0 5888 0 1 2176
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame4_bit24
timestamp 1688980957
transform 1 0 10028 0 -1 10880
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame4_bit25
timestamp 1688980957
transform 1 0 11500 0 -1 10880
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame4_bit26
timestamp 1688980957
transform 1 0 4692 0 -1 34816
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame4_bit27
timestamp 1688980957
transform 1 0 4876 0 -1 35904
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame4_bit28
timestamp 1688980957
transform 1 0 3128 0 -1 26112
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame4_bit29
timestamp 1688980957
transform 1 0 3588 0 -1 27200
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame4_bit30
timestamp 1688980957
transform 1 0 11500 0 -1 13056
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame4_bit31
timestamp 1688980957
transform 1 0 12420 0 -1 11968
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame5_bit0
timestamp 1688980957
transform 1 0 14720 0 -1 5440
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame5_bit1
timestamp 1688980957
transform 1 0 14720 0 1 4352
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame5_bit2
timestamp 1688980957
transform 1 0 1380 0 1 9792
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame5_bit3
timestamp 1688980957
transform 1 0 1656 0 1 10880
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame5_bit4
timestamp 1688980957
transform 1 0 1380 0 1 4352
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame5_bit5
timestamp 1688980957
transform 1 0 1380 0 -1 5440
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame5_bit6
timestamp 1688980957
transform 1 0 1748 0 1 3264
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame5_bit7
timestamp 1688980957
transform 1 0 2300 0 1 2176
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame5_bit8
timestamp 1688980957
transform 1 0 4232 0 -1 2176
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame5_bit9
timestamp 1688980957
transform 1 0 4600 0 -1 4352
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame5_bit10
timestamp 1688980957
transform 1 0 1840 0 1 8704
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame5_bit11
timestamp 1688980957
transform 1 0 2300 0 1 7616
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame5_bit12
timestamp 1688980957
transform 1 0 1380 0 1 17408
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame5_bit13
timestamp 1688980957
transform 1 0 1656 0 -1 16320
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame5_bit14
timestamp 1688980957
transform 1 0 4876 0 -1 9792
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame5_bit15
timestamp 1688980957
transform 1 0 6348 0 -1 8704
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame5_bit16
timestamp 1688980957
transform 1 0 14168 0 1 6528
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame5_bit17
timestamp 1688980957
transform 1 0 14812 0 1 7616
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame5_bit18
timestamp 1688980957
transform 1 0 1380 0 -1 15232
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame5_bit19
timestamp 1688980957
transform 1 0 1472 0 1 13056
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame5_bit20
timestamp 1688980957
transform 1 0 1380 0 -1 6528
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame5_bit21
timestamp 1688980957
transform 1 0 1472 0 -1 7616
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame5_bit22
timestamp 1688980957
transform 1 0 3772 0 1 2176
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame5_bit23
timestamp 1688980957
transform 1 0 2852 0 -1 2176
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame5_bit24
timestamp 1688980957
transform 1 0 15180 0 -1 8704
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame5_bit25
timestamp 1688980957
transform 1 0 16652 0 -1 8704
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame5_bit26
timestamp 1688980957
transform 1 0 1380 0 -1 19584
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame5_bit27
timestamp 1688980957
transform 1 0 1656 0 -1 18496
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame5_bit28
timestamp 1688980957
transform 1 0 1380 0 -1 21760
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame5_bit29
timestamp 1688980957
transform 1 0 1380 0 -1 22848
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame5_bit30
timestamp 1688980957
transform 1 0 6624 0 -1 6528
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame5_bit31
timestamp 1688980957
transform 1 0 8004 0 -1 6528
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame6_bit0
timestamp 1688980957
transform 1 0 10764 0 1 27200
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame6_bit1
timestamp 1688980957
transform 1 0 11040 0 1 28288
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame6_bit2
timestamp 1688980957
transform 1 0 11960 0 -1 18496
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame6_bit3
timestamp 1688980957
transform 1 0 14076 0 1 17408
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame6_bit4
timestamp 1688980957
transform 1 0 12420 0 -1 22848
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame6_bit5
timestamp 1688980957
transform 1 0 14444 0 1 22848
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame6_bit6
timestamp 1688980957
transform 1 0 18032 0 -1 21760
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame6_bit7
timestamp 1688980957
transform 1 0 5428 0 1 21760
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame6_bit8
timestamp 1688980957
transform 1 0 6992 0 -1 21760
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame6_bit9
timestamp 1688980957
transform 1 0 8648 0 -1 21760
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame6_bit10
timestamp 1688980957
transform 1 0 7360 0 -1 30464
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame6_bit11
timestamp 1688980957
transform 1 0 8924 0 1 29376
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame6_bit12
timestamp 1688980957
transform 1 0 9568 0 1 28288
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame6_bit13
timestamp 1688980957
transform 1 0 16652 0 -1 17408
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame6_bit14
timestamp 1688980957
transform 1 0 16652 0 1 17408
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame6_bit15
timestamp 1688980957
transform 1 0 18584 0 -1 19584
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame6_bit16
timestamp 1688980957
transform 1 0 5888 0 1 4352
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame6_bit17
timestamp 1688980957
transform 1 0 7268 0 1 4352
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame6_bit18
timestamp 1688980957
transform 1 0 4048 0 1 13056
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame6_bit19
timestamp 1688980957
transform 1 0 4600 0 -1 15232
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame6_bit20
timestamp 1688980957
transform 1 0 3772 0 1 7616
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame6_bit21
timestamp 1688980957
transform 1 0 4140 0 1 8704
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame6_bit22
timestamp 1688980957
transform 1 0 12512 0 1 3264
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame6_bit23
timestamp 1688980957
transform 1 0 13064 0 -1 4352
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame6_bit24
timestamp 1688980957
transform 1 0 4140 0 -1 5440
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame6_bit25
timestamp 1688980957
transform 1 0 4232 0 1 6528
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame6_bit26
timestamp 1688980957
transform 1 0 2300 0 1 6528
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame6_bit27
timestamp 1688980957
transform 1 0 3128 0 -1 7616
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame6_bit28
timestamp 1688980957
transform 1 0 2300 0 1 11968
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame6_bit29
timestamp 1688980957
transform 1 0 3404 0 -1 14144
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame6_bit30
timestamp 1688980957
transform 1 0 4876 0 -1 6528
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame6_bit31
timestamp 1688980957
transform 1 0 6348 0 1 5440
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame7_bit0
timestamp 1688980957
transform 1 0 7728 0 -1 23936
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame7_bit1
timestamp 1688980957
transform 1 0 9568 0 -1 25024
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame7_bit2
timestamp 1688980957
transform 1 0 9660 0 -1 26112
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame7_bit3
timestamp 1688980957
transform 1 0 6348 0 -1 40256
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame7_bit4
timestamp 1688980957
transform 1 0 6808 0 1 39168
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame7_bit5
timestamp 1688980957
transform 1 0 8372 0 -1 38080
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame7_bit6
timestamp 1688980957
transform 1 0 7084 0 1 32640
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame7_bit7
timestamp 1688980957
transform 1 0 7636 0 -1 33728
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame7_bit8
timestamp 1688980957
transform 1 0 9292 0 1 33728
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame7_bit9
timestamp 1688980957
transform 1 0 12512 0 1 32640
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame7_bit10
timestamp 1688980957
transform 1 0 13248 0 -1 33728
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame7_bit11
timestamp 1688980957
transform 1 0 13432 0 -1 35904
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame7_bit12
timestamp 1688980957
transform 1 0 9476 0 -1 17408
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame7_bit13
timestamp 1688980957
transform 1 0 10120 0 1 16320
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame7_bit14
timestamp 1688980957
transform 1 0 6900 0 1 36992
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame7_bit15
timestamp 1688980957
transform 1 0 7360 0 -1 35904
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame7_bit16
timestamp 1688980957
transform 1 0 7452 0 1 35904
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame7_bit17
timestamp 1688980957
transform 1 0 9016 0 1 35904
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame7_bit18
timestamp 1688980957
transform 1 0 12788 0 -1 31552
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame7_bit19
timestamp 1688980957
transform 1 0 14168 0 -1 31552
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame7_bit20
timestamp 1688980957
transform 1 0 11408 0 1 20672
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame7_bit21
timestamp 1688980957
transform 1 0 12052 0 -1 21760
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame7_bit22
timestamp 1688980957
transform 1 0 9936 0 -1 36992
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame7_bit23
timestamp 1688980957
transform 1 0 11500 0 -1 38080
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame7_bit24
timestamp 1688980957
transform 1 0 7452 0 -1 31552
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame7_bit25
timestamp 1688980957
transform 1 0 9384 0 -1 31552
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame7_bit26
timestamp 1688980957
transform 1 0 11868 0 -1 30464
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame7_bit27
timestamp 1688980957
transform 1 0 12328 0 1 31552
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame7_bit28
timestamp 1688980957
transform 1 0 12420 0 -1 19584
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame7_bit29
timestamp 1688980957
transform 1 0 12604 0 1 19584
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame7_bit30
timestamp 1688980957
transform 1 0 7176 0 1 17408
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame7_bit31
timestamp 1688980957
transform 1 0 8004 0 -1 16320
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame8_bit0
timestamp 1688980957
transform 1 0 22264 0 1 13056
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame8_bit1
timestamp 1688980957
transform 1 0 18860 0 -1 31552
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame8_bit2
timestamp 1688980957
transform 1 0 19412 0 1 33728
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame8_bit3
timestamp 1688980957
transform 1 0 19964 0 -1 19584
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame8_bit4
timestamp 1688980957
transform 1 0 22816 0 -1 9792
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame8_bit5
timestamp 1688980957
transform 1 0 22632 0 -1 10880
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame8_bit6
timestamp 1688980957
transform 1 0 22724 0 1 10880
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame8_bit7
timestamp 1688980957
transform 1 0 22816 0 -1 11968
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame8_bit8
timestamp 1688980957
transform 1 0 9752 0 -1 22848
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame8_bit9
timestamp 1688980957
transform 1 0 10028 0 -1 21760
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame8_bit10
timestamp 1688980957
transform 1 0 1380 0 -1 39168
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame8_bit11
timestamp 1688980957
transform 1 0 1564 0 -1 40256
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame8_bit12
timestamp 1688980957
transform 1 0 1380 0 -1 35904
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame8_bit13
timestamp 1688980957
transform 1 0 1748 0 -1 34816
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame8_bit14
timestamp 1688980957
transform 1 0 14812 0 1 33728
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame8_bit15
timestamp 1688980957
transform 1 0 16008 0 1 32640
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame8_bit16
timestamp 1688980957
transform 1 0 2116 0 1 26112
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame8_bit17
timestamp 1688980957
transform 1 0 2300 0 1 22848
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame8_bit18
timestamp 1688980957
transform 1 0 1380 0 -1 36992
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame8_bit19
timestamp 1688980957
transform 1 0 1472 0 -1 38080
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame8_bit20
timestamp 1688980957
transform 1 0 1380 0 -1 33728
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame8_bit21
timestamp 1688980957
transform 1 0 1564 0 1 32640
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame8_bit22
timestamp 1688980957
transform 1 0 1380 0 1 30464
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame8_bit23
timestamp 1688980957
transform 1 0 1840 0 1 29376
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame8_bit24
timestamp 1688980957
transform 1 0 3772 0 -1 25024
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame8_bit25
timestamp 1688980957
transform 1 0 4416 0 -1 23936
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame8_bit26
timestamp 1688980957
transform 1 0 1380 0 -1 26112
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame8_bit27
timestamp 1688980957
transform 1 0 1656 0 -1 25024
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame8_bit28
timestamp 1688980957
transform 1 0 1380 0 -1 27200
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame8_bit29
timestamp 1688980957
transform 1 0 1564 0 1 27200
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame8_bit30
timestamp 1688980957
transform 1 0 1932 0 1 19584
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame8_bit31
timestamp 1688980957
transform 1 0 2668 0 -1 20672
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame9_bit0
timestamp 1688980957
transform 1 0 18492 0 -1 4352
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame9_bit1
timestamp 1688980957
transform 1 0 19412 0 -1 5440
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame9_bit2
timestamp 1688980957
transform 1 0 19228 0 1 11968
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame9_bit3
timestamp 1688980957
transform 1 0 19780 0 1 10880
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame9_bit4
timestamp 1688980957
transform 1 0 17204 0 1 4352
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame9_bit5
timestamp 1688980957
transform 1 0 22080 0 -1 6528
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame9_bit6
timestamp 1688980957
transform 1 0 22080 0 -1 4352
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame9_bit7
timestamp 1688980957
transform 1 0 20700 0 1 3264
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame9_bit8
timestamp 1688980957
transform 1 0 22632 0 -1 25024
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame9_bit9
timestamp 1688980957
transform 1 0 21344 0 1 30464
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame9_bit10
timestamp 1688980957
transform 1 0 21988 0 -1 28288
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame9_bit11
timestamp 1688980957
transform 1 0 17572 0 1 27200
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame9_bit12
timestamp 1688980957
transform 1 0 20976 0 1 22848
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame9_bit13
timestamp 1688980957
transform 1 0 22540 0 1 22848
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame9_bit14
timestamp 1688980957
transform 1 0 20332 0 -1 26112
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame9_bit15
timestamp 1688980957
transform 1 0 18952 0 -1 27200
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame9_bit16
timestamp 1688980957
transform 1 0 17572 0 1 23936
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame9_bit17
timestamp 1688980957
transform 1 0 21068 0 1 32640
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame9_bit18
timestamp 1688980957
transform 1 0 19596 0 1 28288
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame9_bit19
timestamp 1688980957
transform 1 0 17756 0 1 30464
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame9_bit20
timestamp 1688980957
transform 1 0 19412 0 -1 23936
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame9_bit21
timestamp 1688980957
transform 1 0 22816 0 -1 20672
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame9_bit22
timestamp 1688980957
transform 1 0 20700 0 1 19584
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame9_bit23
timestamp 1688980957
transform 1 0 19228 0 1 21760
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame9_bit24
timestamp 1688980957
transform 1 0 17756 0 -1 16320
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame9_bit25
timestamp 1688980957
transform 1 0 21804 0 -1 16320
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame9_bit26
timestamp 1688980957
transform 1 0 22632 0 1 16320
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame9_bit27
timestamp 1688980957
transform 1 0 22448 0 1 18496
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame9_bit28
timestamp 1688980957
transform 1 0 17664 0 1 14144
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame9_bit29
timestamp 1688980957
transform 1 0 22908 0 -1 14144
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame9_bit30
timestamp 1688980957
transform 1 0 19596 0 1 14144
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame9_bit31
timestamp 1688980957
transform 1 0 20332 0 -1 17408
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame10_bit24
timestamp 1688980957
transform 1 0 16652 0 -1 6528
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame10_bit25
timestamp 1688980957
transform 1 0 17020 0 -1 9792
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame10_bit26
timestamp 1688980957
transform 1 0 21436 0 1 7616
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame10_bit27
timestamp 1688980957
transform 1 0 18584 0 -1 9792
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame10_bit28
timestamp 1688980957
transform 1 0 17020 0 -1 13056
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame10_bit29
timestamp 1688980957
transform 1 0 20332 0 -1 13056
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame10_bit30
timestamp 1688980957
transform 1 0 19780 0 -1 7616
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem_Inst_frame10_bit31
timestamp 1688980957
transform 1 0 17756 0 1 5440
box -38 -48 1418 592
use sky130_fd_sc_hd__buf_2  Inst_RAM_IO_switch_matrix__32_
timestamp 1688980957
transform 1 0 3772 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM_IO_switch_matrix__33_
timestamp 1688980957
transform 1 0 4324 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_RAM_IO_switch_matrix__34_
timestamp 1688980957
transform 1 0 2944 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_RAM_IO_switch_matrix__35_
timestamp 1688980957
transform 1 0 3956 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  Inst_RAM_IO_switch_matrix__36_
timestamp 1688980957
transform 1 0 4876 0 1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  Inst_RAM_IO_switch_matrix__37_
timestamp 1688980957
transform 1 0 4048 0 -1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  Inst_RAM_IO_switch_matrix__38_
timestamp 1688980957
transform 1 0 5888 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  Inst_RAM_IO_switch_matrix__39_
timestamp 1688980957
transform 1 0 5152 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM_IO_switch_matrix__40_
timestamp 1688980957
transform 1 0 11500 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  Inst_RAM_IO_switch_matrix__41_
timestamp 1688980957
transform 1 0 11500 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  Inst_RAM_IO_switch_matrix__42_
timestamp 1688980957
transform 1 0 11592 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  Inst_RAM_IO_switch_matrix__43_
timestamp 1688980957
transform 1 0 11960 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM_IO_switch_matrix__44_
timestamp 1688980957
transform 1 0 11500 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_RAM_IO_switch_matrix__45_
timestamp 1688980957
transform 1 0 12328 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  Inst_RAM_IO_switch_matrix__46_
timestamp 1688980957
transform 1 0 13248 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM_IO_switch_matrix__47_
timestamp 1688980957
transform 1 0 13616 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_FAB2RAM_A0_I0_395 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 15548 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_FAB2RAM_A0_I0 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14628 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_FAB2RAM_A0_I1_396
timestamp 1688980957
transform 1 0 11684 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_FAB2RAM_A0_I1
timestamp 1688980957
transform 1 0 11224 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_FAB2RAM_A0_I2_397
timestamp 1688980957
transform 1 0 10028 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_FAB2RAM_A0_I2 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 8924 0 1 18496
box -38 -48 1694 592
use sky130_fd_sc_hd__conb_1  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_FAB2RAM_A0_I3_398
timestamp 1688980957
transform 1 0 15824 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_FAB2RAM_A0_I3
timestamp 1688980957
transform 1 0 14628 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_FAB2RAM_A1_I0_399
timestamp 1688980957
transform 1 0 13432 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_FAB2RAM_A1_I0
timestamp 1688980957
transform 1 0 12420 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_FAB2RAM_A1_I1_400
timestamp 1688980957
transform 1 0 9476 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_FAB2RAM_A1_I1
timestamp 1688980957
transform 1 0 8464 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_FAB2RAM_A1_I2_401
timestamp 1688980957
transform 1 0 11684 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_FAB2RAM_A1_I2
timestamp 1688980957
transform 1 0 10672 0 1 19584
box -38 -48 1694 592
use sky130_fd_sc_hd__conb_1  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_FAB2RAM_A1_I3_402
timestamp 1688980957
transform 1 0 17020 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_FAB2RAM_A1_I3
timestamp 1688980957
transform 1 0 16100 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_FAB2RAM_C_I0_403
timestamp 1688980957
transform 1 0 11684 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_FAB2RAM_C_I0
timestamp 1688980957
transform 1 0 11500 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_FAB2RAM_C_I1
timestamp 1688980957
transform 1 0 7360 0 -1 41344
box -38 -48 1694 592
use sky130_fd_sc_hd__conb_1  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_FAB2RAM_C_I1_404
timestamp 1688980957
transform 1 0 7084 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_FAB2RAM_C_I2
timestamp 1688980957
transform 1 0 11500 0 -1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_FAB2RAM_C_I2_405
timestamp 1688980957
transform 1 0 11132 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_FAB2RAM_C_I3_409
timestamp 1688980957
transform 1 0 16284 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_FAB2RAM_C_I3
timestamp 1688980957
transform 1 0 16652 0 -1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_FAB2RAM_D0_I0
timestamp 1688980957
transform 1 0 11500 0 1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_FAB2RAM_D0_I1
timestamp 1688980957
transform 1 0 5244 0 1 31552
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_FAB2RAM_D0_I2
timestamp 1688980957
transform 1 0 4600 0 -1 28288
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_FAB2RAM_D0_I3
timestamp 1688980957
transform 1 0 14628 0 -1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_FAB2RAM_D1_I0
timestamp 1688980957
transform 1 0 14076 0 1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_FAB2RAM_D1_I1
timestamp 1688980957
transform 1 0 6348 0 -1 25024
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_FAB2RAM_D1_I2
timestamp 1688980957
transform 1 0 6808 0 -1 27200
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_FAB2RAM_D1_I3
timestamp 1688980957
transform 1 0 16008 0 1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_FAB2RAM_D2_I0
timestamp 1688980957
transform 1 0 11776 0 1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_FAB2RAM_D2_I1
timestamp 1688980957
transform 1 0 6348 0 1 33728
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_FAB2RAM_D2_I2
timestamp 1688980957
transform 1 0 6256 0 1 29376
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_FAB2RAM_D2_I3
timestamp 1688980957
transform 1 0 15180 0 1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_FAB2RAM_D3_I0
timestamp 1688980957
transform 1 0 13616 0 -1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_FAB2RAM_D3_I1
timestamp 1688980957
transform 1 0 6992 0 1 23936
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_FAB2RAM_D3_I2
timestamp 1688980957
transform 1 0 8924 0 1 26112
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_FAB2RAM_D3_I3
timestamp 1688980957
transform 1 0 16652 0 -1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_J_NS1_BEG0_406
timestamp 1688980957
transform 1 0 10304 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_J_NS1_BEG0
timestamp 1688980957
transform 1 0 9292 0 -1 13056
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_J_NS1_BEG1
timestamp 1688980957
transform 1 0 2484 0 -1 42432
box -38 -48 1694 592
use sky130_fd_sc_hd__conb_1  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_J_NS1_BEG1_407
timestamp 1688980957
transform 1 0 1472 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_J_NS1_BEG2_408
timestamp 1688980957
transform 1 0 4416 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_J_NS1_BEG2
timestamp 1688980957
transform 1 0 2852 0 -1 35904
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_J_NS1_BEG3
timestamp 1688980957
transform 1 0 12880 0 -1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_J_NS1_BEG3_394
timestamp 1688980957
transform 1 0 14076 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_J_NS2_BEG0
timestamp 1688980957
transform 1 0 9752 0 1 2176
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_J_NS2_BEG1
timestamp 1688980957
transform 1 0 9568 0 -1 39168
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_J_NS2_BEG2
timestamp 1688980957
transform 1 0 4416 0 1 30464
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_J_NS2_BEG3
timestamp 1688980957
transform 1 0 11500 0 -1 33728
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_J_NS2_BEG4
timestamp 1688980957
transform 1 0 11132 0 1 4352
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_J_NS2_BEG5
timestamp 1688980957
transform 1 0 7176 0 1 19584
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_J_NS2_BEG6
timestamp 1688980957
transform 1 0 10304 0 1 29376
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_J_NS2_BEG7
timestamp 1688980957
transform 1 0 11960 0 1 2176
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_J_NS4_BEG0
timestamp 1688980957
transform 1 0 8924 0 1 3264
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_J_NS4_BEG1
timestamp 1688980957
transform 1 0 4600 0 1 39168
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_J_NS4_BEG2
timestamp 1688980957
transform 1 0 3772 0 1 28288
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_J_NS4_BEG3
timestamp 1688980957
transform 1 0 13432 0 -1 14144
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_J_NS4_BEG4
timestamp 1688980957
transform 1 0 9292 0 -1 9792
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_J_NS4_BEG5
timestamp 1688980957
transform 1 0 4784 0 1 36992
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_J_NS4_BEG6
timestamp 1688980957
transform 1 0 3220 0 -1 31552
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_J_NS4_BEG7
timestamp 1688980957
transform 1 0 11960 0 1 9792
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_J_NS4_BEG8
timestamp 1688980957
transform 1 0 9660 0 -1 7616
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_J_NS4_BEG9
timestamp 1688980957
transform 1 0 4876 0 1 41344
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_J_NS4_BEG10
timestamp 1688980957
transform 1 0 3864 0 1 33728
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_J_NS4_BEG11
timestamp 1688980957
transform 1 0 12328 0 1 7616
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_J_NS4_BEG12
timestamp 1688980957
transform 1 0 9568 0 -1 5440
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_J_NS4_BEG13
timestamp 1688980957
transform 1 0 4324 0 -1 41344
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_J_NS4_BEG14
timestamp 1688980957
transform 1 0 3772 0 1 35904
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_J_NS4_BEG15
timestamp 1688980957
transform 1 0 11500 0 -1 7616
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_N1BEG0
timestamp 1688980957
transform 1 0 10028 0 1 21760
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_N1BEG1
timestamp 1688980957
transform 1 0 1472 0 1 40256
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_N1BEG2
timestamp 1688980957
transform 1 0 1656 0 1 34816
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_N1BEG3
timestamp 1688980957
transform 1 0 14628 0 -1 33728
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_N2BEG0
timestamp 1688980957
transform 1 0 2392 0 -1 23936
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_N2BEG1
timestamp 1688980957
transform 1 0 1380 0 1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_N2BEG2
timestamp 1688980957
transform 1 0 1380 0 -1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_N2BEG3
timestamp 1688980957
transform 1 0 1656 0 -1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_N2BEG4
timestamp 1688980957
transform 1 0 4232 0 1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_N2BEG5
timestamp 1688980957
transform 1 0 1380 0 1 25024
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_N2BEG6
timestamp 1688980957
transform 1 0 1380 0 -1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_N2BEG7
timestamp 1688980957
transform 1 0 2024 0 1 20672
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_S1BEG0
timestamp 1688980957
transform 1 0 9476 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_S1BEG1
timestamp 1688980957
transform 1 0 7268 0 -1 36992
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_S1BEG2
timestamp 1688980957
transform 1 0 8740 0 -1 35904
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_S1BEG3
timestamp 1688980957
transform 1 0 13892 0 -1 30464
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_S2BEG0
timestamp 1688980957
transform 1 0 11776 0 1 21760
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_S2BEG1
timestamp 1688980957
transform 1 0 10488 0 1 36992
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_S2BEG2
timestamp 1688980957
transform 1 0 8924 0 1 31552
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_S2BEG3
timestamp 1688980957
transform 1 0 12144 0 1 30464
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_S2BEG4
timestamp 1688980957
transform 1 0 12788 0 -1 20672
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_S2BEG5
timestamp 1688980957
transform 1 0 7728 0 -1 17408
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_S2BEG6
timestamp 1688980957
transform 1 0 11500 0 -1 28288
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_S2BEG7
timestamp 1688980957
transform 1 0 13340 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_W1BEG0
timestamp 1688980957
transform 1 0 7084 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_W1BEG1
timestamp 1688980957
transform 1 0 4324 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_W1BEG2
timestamp 1688980957
transform 1 0 3864 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_W1BEG3
timestamp 1688980957
transform 1 0 12788 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_W2BEG0
timestamp 1688980957
transform 1 0 4416 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_W2BEG1
timestamp 1688980957
transform 1 0 2760 0 -1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_W2BEG2
timestamp 1688980957
transform 1 0 2668 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_W2BEG3
timestamp 1688980957
transform 1 0 5612 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_W2BEG4
timestamp 1688980957
transform 1 0 14444 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_W2BEG5
timestamp 1688980957
transform 1 0 1472 0 -1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_W2BEG6
timestamp 1688980957
transform 1 0 1472 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_W2BEG7
timestamp 1688980957
transform 1 0 2668 0 -1 4352
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_W2BEGb0
timestamp 1688980957
transform 1 0 3772 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_W2BEGb1
timestamp 1688980957
transform 1 0 2392 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_W2BEGb2
timestamp 1688980957
transform 1 0 1564 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_W2BEGb3
timestamp 1688980957
transform 1 0 5520 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_W2BEGb4
timestamp 1688980957
transform 1 0 14444 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_W2BEGb5
timestamp 1688980957
transform 1 0 1472 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_W2BEGb6
timestamp 1688980957
transform 1 0 1472 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_W2BEGb7
timestamp 1688980957
transform 1 0 2760 0 -1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_W6BEG0
timestamp 1688980957
transform 1 0 10396 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_W6BEG1
timestamp 1688980957
transform 1 0 5060 0 1 34816
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_W6BEG2
timestamp 1688980957
transform 1 0 3772 0 1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_W6BEG3
timestamp 1688980957
transform 1 0 12052 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_W6BEG4
timestamp 1688980957
transform 1 0 14168 0 1 11968
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_W6BEG5
timestamp 1688980957
transform 1 0 5796 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_W6BEG6
timestamp 1688980957
transform 1 0 6164 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_W6BEG7
timestamp 1688980957
transform 1 0 7820 0 -1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_W6BEG8
timestamp 1688980957
transform 1 0 14260 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_W6BEG9
timestamp 1688980957
transform 1 0 5336 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_W6BEG10
timestamp 1688980957
transform 1 0 5060 0 1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_W6BEG11
timestamp 1688980957
transform 1 0 7084 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_WW4BEG0
timestamp 1688980957
transform 1 0 15640 0 1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_WW4BEG1
timestamp 1688980957
transform 1 0 1656 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_WW4BEG2
timestamp 1688980957
transform 1 0 1472 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_WW4BEG3
timestamp 1688980957
transform 1 0 7636 0 -1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_WW4BEG4
timestamp 1688980957
transform 1 0 14076 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_WW4BEG5
timestamp 1688980957
transform 1 0 5060 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_WW4BEG6
timestamp 1688980957
transform 1 0 3220 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_WW4BEG7
timestamp 1688980957
transform 1 0 7728 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_WW4BEG8
timestamp 1688980957
transform 1 0 15640 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_WW4BEG9
timestamp 1688980957
transform 1 0 3588 0 -1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_WW4BEG10
timestamp 1688980957
transform 1 0 4232 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_WW4BEG11
timestamp 1688980957
transform 1 0 6900 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_WW4BEG12
timestamp 1688980957
transform 1 0 15456 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_WW4BEG13
timestamp 1688980957
transform 1 0 3588 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_WW4BEG14
timestamp 1688980957
transform 1 0 3772 0 -1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix_inst_cus_mux41_buf_WW4BEG15
timestamp 1688980957
transform 1 0 5704 0 1 3264
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_2  Inst_RAM_IO_switch_matrix_inst_cus_mux81_buf_N4BEG0_cus_mux21_inst__2_
timestamp 1688980957
transform 1 0 10948 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM_IO_switch_matrix_inst_cus_mux81_buf_N4BEG0_cus_mux21_inst__3_
timestamp 1688980957
transform 1 0 11224 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_RAM_IO_switch_matrix_inst_cus_mux81_buf_N4BEG0_cus_mux21_inst__4_
timestamp 1688980957
transform 1 0 10580 0 1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM_IO_switch_matrix_inst_cus_mux81_buf_N4BEG0_cus_mux21_inst_break_comb_loop_inst0__0_
timestamp 1688980957
transform 1 0 10764 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM_IO_switch_matrix_inst_cus_mux81_buf_N4BEG0_cus_mux21_inst_break_comb_loop_inst1__0_
timestamp 1688980957
transform 1 0 11040 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix_inst_cus_mux81_buf_N4BEG0_cus_mux41_buf_inst0
timestamp 1688980957
transform 1 0 9108 0 -1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix_inst_cus_mux81_buf_N4BEG0_cus_mux41_buf_inst1
timestamp 1688980957
transform 1 0 9108 0 1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_2  Inst_RAM_IO_switch_matrix_inst_cus_mux81_buf_N4BEG1_cus_mux21_inst__2_
timestamp 1688980957
transform 1 0 9568 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM_IO_switch_matrix_inst_cus_mux81_buf_N4BEG1_cus_mux21_inst__3_
timestamp 1688980957
transform 1 0 9292 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_RAM_IO_switch_matrix_inst_cus_mux81_buf_N4BEG1_cus_mux21_inst__4_
timestamp 1688980957
transform 1 0 8924 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM_IO_switch_matrix_inst_cus_mux81_buf_N4BEG1_cus_mux21_inst_break_comb_loop_inst0__0_
timestamp 1688980957
transform 1 0 8740 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM_IO_switch_matrix_inst_cus_mux81_buf_N4BEG1_cus_mux21_inst_break_comb_loop_inst1__0_
timestamp 1688980957
transform 1 0 8924 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix_inst_cus_mux81_buf_N4BEG1_cus_mux41_buf_inst0
timestamp 1688980957
transform 1 0 6440 0 1 38080
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix_inst_cus_mux81_buf_N4BEG1_cus_mux41_buf_inst1
timestamp 1688980957
transform 1 0 6716 0 -1 39168
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_2  Inst_RAM_IO_switch_matrix_inst_cus_mux81_buf_N4BEG2_cus_mux21_inst__2_
timestamp 1688980957
transform 1 0 8556 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM_IO_switch_matrix_inst_cus_mux81_buf_N4BEG2_cus_mux21_inst__3_
timestamp 1688980957
transform 1 0 10672 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_RAM_IO_switch_matrix_inst_cus_mux81_buf_N4BEG2_cus_mux21_inst__4_
timestamp 1688980957
transform 1 0 9568 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM_IO_switch_matrix_inst_cus_mux81_buf_N4BEG2_cus_mux21_inst_break_comb_loop_inst0__0_
timestamp 1688980957
transform 1 0 9016 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM_IO_switch_matrix_inst_cus_mux81_buf_N4BEG2_cus_mux21_inst_break_comb_loop_inst1__0_
timestamp 1688980957
transform 1 0 9660 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix_inst_cus_mux81_buf_N4BEG2_cus_mux41_buf_inst0
timestamp 1688980957
transform 1 0 6900 0 1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix_inst_cus_mux81_buf_N4BEG2_cus_mux41_buf_inst1
timestamp 1688980957
transform 1 0 7544 0 -1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_2  Inst_RAM_IO_switch_matrix_inst_cus_mux81_buf_N4BEG3_cus_mux21_inst__2_
timestamp 1688980957
transform 1 0 15180 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM_IO_switch_matrix_inst_cus_mux81_buf_N4BEG3_cus_mux21_inst__3_
timestamp 1688980957
transform 1 0 14536 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_RAM_IO_switch_matrix_inst_cus_mux81_buf_N4BEG3_cus_mux21_inst__4_
timestamp 1688980957
transform 1 0 14812 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM_IO_switch_matrix_inst_cus_mux81_buf_N4BEG3_cus_mux21_inst_break_comb_loop_inst0__0_
timestamp 1688980957
transform 1 0 14720 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM_IO_switch_matrix_inst_cus_mux81_buf_N4BEG3_cus_mux21_inst_break_comb_loop_inst1__0_
timestamp 1688980957
transform 1 0 14996 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix_inst_cus_mux81_buf_N4BEG3_cus_mux41_buf_inst0
timestamp 1688980957
transform 1 0 13156 0 -1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix_inst_cus_mux81_buf_N4BEG3_cus_mux41_buf_inst1
timestamp 1688980957
transform 1 0 14076 0 1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_2  Inst_RAM_IO_switch_matrix_inst_cus_mux81_buf_S4BEG0_cus_mux21_inst__2_
timestamp 1688980957
transform 1 0 17480 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM_IO_switch_matrix_inst_cus_mux81_buf_S4BEG0_cus_mux21_inst__3_
timestamp 1688980957
transform 1 0 18124 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_RAM_IO_switch_matrix_inst_cus_mux81_buf_S4BEG0_cus_mux21_inst__4_
timestamp 1688980957
transform 1 0 18032 0 1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM_IO_switch_matrix_inst_cus_mux81_buf_S4BEG0_cus_mux21_inst_break_comb_loop_inst0__0_
timestamp 1688980957
transform 1 0 16652 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM_IO_switch_matrix_inst_cus_mux81_buf_S4BEG0_cus_mux21_inst_break_comb_loop_inst1__0_
timestamp 1688980957
transform 1 0 17756 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix_inst_cus_mux81_buf_S4BEG0_cus_mux41_buf_inst0
timestamp 1688980957
transform 1 0 13800 0 -1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix_inst_cus_mux81_buf_S4BEG0_cus_mux41_buf_inst1
timestamp 1688980957
transform 1 0 14076 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_2  Inst_RAM_IO_switch_matrix_inst_cus_mux81_buf_S4BEG1_cus_mux21_inst__2_
timestamp 1688980957
transform 1 0 9108 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM_IO_switch_matrix_inst_cus_mux81_buf_S4BEG1_cus_mux21_inst__3_
timestamp 1688980957
transform 1 0 9384 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  Inst_RAM_IO_switch_matrix_inst_cus_mux81_buf_S4BEG1_cus_mux21_inst__4_
timestamp 1688980957
transform 1 0 9384 0 1 20672
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM_IO_switch_matrix_inst_cus_mux81_buf_S4BEG1_cus_mux21_inst_break_comb_loop_inst0__0_
timestamp 1688980957
transform 1 0 8648 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM_IO_switch_matrix_inst_cus_mux81_buf_S4BEG1_cus_mux21_inst_break_comb_loop_inst1__0_
timestamp 1688980957
transform 1 0 9016 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix_inst_cus_mux81_buf_S4BEG1_cus_mux41_buf_inst0
timestamp 1688980957
transform 1 0 6532 0 -1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix_inst_cus_mux81_buf_S4BEG1_cus_mux41_buf_inst1
timestamp 1688980957
transform 1 0 6808 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_2  Inst_RAM_IO_switch_matrix_inst_cus_mux81_buf_S4BEG2_cus_mux21_inst__2_
timestamp 1688980957
transform 1 0 10672 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM_IO_switch_matrix_inst_cus_mux81_buf_S4BEG2_cus_mux21_inst__3_
timestamp 1688980957
transform 1 0 10396 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  Inst_RAM_IO_switch_matrix_inst_cus_mux81_buf_S4BEG2_cus_mux21_inst__4_
timestamp 1688980957
transform 1 0 10396 0 -1 28288
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM_IO_switch_matrix_inst_cus_mux81_buf_S4BEG2_cus_mux21_inst_break_comb_loop_inst0__0_
timestamp 1688980957
transform 1 0 9844 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM_IO_switch_matrix_inst_cus_mux81_buf_S4BEG2_cus_mux21_inst_break_comb_loop_inst1__0_
timestamp 1688980957
transform 1 0 10120 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix_inst_cus_mux81_buf_S4BEG2_cus_mux41_buf_inst0
timestamp 1688980957
transform 1 0 7728 0 -1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix_inst_cus_mux81_buf_S4BEG2_cus_mux41_buf_inst1
timestamp 1688980957
transform 1 0 7820 0 -1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_2  Inst_RAM_IO_switch_matrix_inst_cus_mux81_buf_S4BEG3_cus_mux21_inst__2_
timestamp 1688980957
transform 1 0 19228 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM_IO_switch_matrix_inst_cus_mux81_buf_S4BEG3_cus_mux21_inst__3_
timestamp 1688980957
transform 1 0 19504 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_RAM_IO_switch_matrix_inst_cus_mux81_buf_S4BEG3_cus_mux21_inst__4_
timestamp 1688980957
transform 1 0 18676 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM_IO_switch_matrix_inst_cus_mux81_buf_S4BEG3_cus_mux21_inst_break_comb_loop_inst0__0_
timestamp 1688980957
transform 1 0 18124 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM_IO_switch_matrix_inst_cus_mux81_buf_S4BEG3_cus_mux21_inst_break_comb_loop_inst1__0_
timestamp 1688980957
transform 1 0 18400 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix_inst_cus_mux81_buf_S4BEG3_cus_mux41_buf_inst0
timestamp 1688980957
transform 1 0 16652 0 -1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix_inst_cus_mux81_buf_S4BEG3_cus_mux41_buf_inst1
timestamp 1688980957
transform 1 0 16652 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_1  N4BEG_outbuf_0__0_
timestamp 1688980957
transform 1 0 5980 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  N4BEG_outbuf_1__0_
timestamp 1688980957
transform 1 0 5980 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  N4BEG_outbuf_2__0_
timestamp 1688980957
transform 1 0 7176 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  N4BEG_outbuf_3__0_
timestamp 1688980957
transform 1 0 6900 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  N4BEG_outbuf_4__0_
timestamp 1688980957
transform 1 0 10212 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  N4BEG_outbuf_5__0_
timestamp 1688980957
transform 1 0 3404 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  N4BEG_outbuf_6__0_
timestamp 1688980957
transform 1 0 8832 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  N4BEG_outbuf_7__0_
timestamp 1688980957
transform 1 0 9936 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  N4BEG_outbuf_8__0_
timestamp 1688980957
transform 1 0 3772 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  N4BEG_outbuf_9__0_
timestamp 1688980957
transform 1 0 8924 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  N4BEG_outbuf_10__0_
timestamp 1688980957
transform 1 0 9200 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  N4BEG_outbuf_11__0_
timestamp 1688980957
transform 1 0 9108 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  N4END_inbuf_0__0_
timestamp 1688980957
transform 1 0 5520 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  N4END_inbuf_1__0_
timestamp 1688980957
transform 1 0 5888 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  N4END_inbuf_2__0_
timestamp 1688980957
transform 1 0 5888 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  N4END_inbuf_3__0_
timestamp 1688980957
transform 1 0 6348 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  N4END_inbuf_4__0_
timestamp 1688980957
transform 1 0 6716 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  N4END_inbuf_5__0_
timestamp 1688980957
transform 1 0 7636 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  N4END_inbuf_6__0_
timestamp 1688980957
transform 1 0 7084 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  N4END_inbuf_7__0_
timestamp 1688980957
transform 1 0 7544 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  N4END_inbuf_8__0_
timestamp 1688980957
transform 1 0 7452 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  N4END_inbuf_9__0_
timestamp 1688980957
transform 1 0 7820 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  N4END_inbuf_10__0_
timestamp 1688980957
transform 1 0 8188 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  N4END_inbuf_11__0_
timestamp 1688980957
transform 1 0 8556 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output189
timestamp 1688980957
transform 1 0 23920 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output190
timestamp 1688980957
transform 1 0 23184 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output191
timestamp 1688980957
transform 1 0 22816 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output192
timestamp 1688980957
transform 1 0 23736 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output193
timestamp 1688980957
transform 1 0 23552 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output194
timestamp 1688980957
transform 1 0 23920 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output195
timestamp 1688980957
transform 1 0 23184 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output196
timestamp 1688980957
transform 1 0 23552 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output197
timestamp 1688980957
transform 1 0 23920 0 1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output198
timestamp 1688980957
transform 1 0 23184 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output199
timestamp 1688980957
transform 1 0 23920 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output200
timestamp 1688980957
transform 1 0 23736 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output201
timestamp 1688980957
transform 1 0 23552 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output202
timestamp 1688980957
transform 1 0 23184 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output203
timestamp 1688980957
transform 1 0 23552 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output204
timestamp 1688980957
transform 1 0 23184 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output205
timestamp 1688980957
transform 1 0 23368 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output206
timestamp 1688980957
transform 1 0 23920 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output207
timestamp 1688980957
transform 1 0 23552 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output208
timestamp 1688980957
transform 1 0 23736 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output209
timestamp 1688980957
transform 1 0 23552 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output210
timestamp 1688980957
transform 1 0 23920 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output211
timestamp 1688980957
transform 1 0 23736 0 -1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output212
timestamp 1688980957
transform 1 0 23920 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output213
timestamp 1688980957
transform 1 0 23368 0 1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output214
timestamp 1688980957
transform 1 0 23736 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output215
timestamp 1688980957
transform 1 0 23920 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output216
timestamp 1688980957
transform 1 0 23920 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output217
timestamp 1688980957
transform 1 0 23184 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output218
timestamp 1688980957
transform 1 0 23920 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output219
timestamp 1688980957
transform 1 0 23552 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output220
timestamp 1688980957
transform 1 0 23736 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output221
timestamp 1688980957
transform 1 0 23920 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output222
timestamp 1688980957
transform 1 0 23920 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output223
timestamp 1688980957
transform 1 0 23920 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output224
timestamp 1688980957
transform 1 0 23920 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output225
timestamp 1688980957
transform 1 0 23920 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output226
timestamp 1688980957
transform 1 0 23736 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output227
timestamp 1688980957
transform 1 0 23920 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output228
timestamp 1688980957
transform 1 0 23920 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output229
timestamp 1688980957
transform 1 0 23736 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output230
timestamp 1688980957
transform 1 0 23920 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output231
timestamp 1688980957
transform 1 0 23920 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output232
timestamp 1688980957
transform 1 0 23920 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output233
timestamp 1688980957
transform 1 0 23920 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output234
timestamp 1688980957
transform 1 0 23920 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output235
timestamp 1688980957
transform 1 0 23736 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output236
timestamp 1688980957
transform 1 0 23920 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output237
timestamp 1688980957
transform 1 0 23736 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output238
timestamp 1688980957
transform 1 0 23368 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output239
timestamp 1688980957
transform 1 0 22632 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output240
timestamp 1688980957
transform 1 0 23000 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output241
timestamp 1688980957
transform 1 0 23920 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output242
timestamp 1688980957
transform 1 0 23552 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output243
timestamp 1688980957
transform 1 0 23920 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output244
timestamp 1688980957
transform 1 0 22448 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output245
timestamp 1688980957
transform 1 0 21620 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output246
timestamp 1688980957
transform 1 0 23920 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output247
timestamp 1688980957
transform 1 0 23736 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output248
timestamp 1688980957
transform 1 0 23920 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output249
timestamp 1688980957
transform 1 0 23920 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output250
timestamp 1688980957
transform 1 0 23736 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output251
timestamp 1688980957
transform 1 0 23920 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output252
timestamp 1688980957
transform 1 0 23736 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output253
timestamp 1688980957
transform 1 0 20148 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output254
timestamp 1688980957
transform 1 0 21068 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output255
timestamp 1688980957
transform 1 0 22080 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output256
timestamp 1688980957
transform 1 0 23552 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output257
timestamp 1688980957
transform 1 0 23736 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output258
timestamp 1688980957
transform 1 0 23000 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output259
timestamp 1688980957
transform 1 0 23184 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output260
timestamp 1688980957
transform 1 0 23552 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output261
timestamp 1688980957
transform 1 0 22632 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output262
timestamp 1688980957
transform 1 0 23736 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output263
timestamp 1688980957
transform 1 0 21160 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output264
timestamp 1688980957
transform 1 0 20516 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output265
timestamp 1688980957
transform 1 0 21804 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output266
timestamp 1688980957
transform 1 0 21344 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output267
timestamp 1688980957
transform 1 0 22172 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output268
timestamp 1688980957
transform 1 0 22724 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output269
timestamp 1688980957
transform 1 0 22172 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output270
timestamp 1688980957
transform 1 0 22724 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output271
timestamp 1688980957
transform 1 0 23276 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output272
timestamp 1688980957
transform 1 0 21896 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output273
timestamp 1688980957
transform 1 0 9844 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output274
timestamp 1688980957
transform 1 0 6348 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output275
timestamp 1688980957
transform 1 0 8188 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output276
timestamp 1688980957
transform 1 0 6992 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output277
timestamp 1688980957
transform 1 0 5704 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output278
timestamp 1688980957
transform 1 0 1748 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output279
timestamp 1688980957
transform 1 0 6532 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output280
timestamp 1688980957
transform 1 0 3772 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output281
timestamp 1688980957
transform 1 0 5152 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output282
timestamp 1688980957
transform 1 0 1932 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output283
timestamp 1688980957
transform 1 0 4876 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output284
timestamp 1688980957
transform 1 0 1932 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output285
timestamp 1688980957
transform 1 0 1472 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output286
timestamp 1688980957
transform 1 0 2392 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output287
timestamp 1688980957
transform 1 0 4324 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output288
timestamp 1688980957
transform 1 0 5428 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output289
timestamp 1688980957
transform 1 0 2576 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output290
timestamp 1688980957
transform 1 0 3128 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output291
timestamp 1688980957
transform 1 0 1380 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output292
timestamp 1688980957
transform 1 0 3864 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output293
timestamp 1688980957
transform 1 0 2576 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output294
timestamp 1688980957
transform 1 0 8280 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output295
timestamp 1688980957
transform 1 0 7360 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output296
timestamp 1688980957
transform 1 0 8464 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output297
timestamp 1688980957
transform 1 0 9292 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output298
timestamp 1688980957
transform 1 0 8924 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output299
timestamp 1688980957
transform 1 0 9292 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output300
timestamp 1688980957
transform 1 0 3128 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output301
timestamp 1688980957
transform 1 0 7084 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output302
timestamp 1688980957
transform 1 0 1380 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output303
timestamp 1688980957
transform 1 0 5704 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output304
timestamp 1688980957
transform 1 0 6808 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output305
timestamp 1688980957
transform 1 0 6440 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output306
timestamp 1688980957
transform 1 0 6348 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output307
timestamp 1688980957
transform 1 0 7728 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output308
timestamp 1688980957
transform 1 0 8924 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output309
timestamp 1688980957
transform 1 0 8924 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output310
timestamp 1688980957
transform 1 0 10396 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output311
timestamp 1688980957
transform 1 0 9476 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output312
timestamp 1688980957
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output313
timestamp 1688980957
transform 1 0 13432 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output314
timestamp 1688980957
transform 1 0 14444 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output315
timestamp 1688980957
transform 1 0 14076 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output316
timestamp 1688980957
transform 1 0 14812 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output317
timestamp 1688980957
transform 1 0 15180 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output318
timestamp 1688980957
transform 1 0 15732 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output319
timestamp 1688980957
transform 1 0 16652 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output320
timestamp 1688980957
transform 1 0 15364 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output321
timestamp 1688980957
transform 1 0 8280 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output322
timestamp 1688980957
transform 1 0 7912 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output323
timestamp 1688980957
transform 1 0 11776 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output324
timestamp 1688980957
transform 1 0 11040 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output325
timestamp 1688980957
transform 1 0 11776 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output326
timestamp 1688980957
transform 1 0 12144 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output327
timestamp 1688980957
transform 1 0 12696 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output328
timestamp 1688980957
transform 1 0 13064 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output329
timestamp 1688980957
transform 1 0 15916 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output330
timestamp 1688980957
transform 1 0 17940 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output331
timestamp 1688980957
transform 1 0 18400 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output332
timestamp 1688980957
transform 1 0 18952 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output333
timestamp 1688980957
transform 1 0 19504 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output334
timestamp 1688980957
transform 1 0 19872 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output335
timestamp 1688980957
transform 1 0 20056 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output336
timestamp 1688980957
transform 1 0 17204 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output337
timestamp 1688980957
transform 1 0 18308 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output338
timestamp 1688980957
transform 1 0 16652 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output339
timestamp 1688980957
transform 1 0 18860 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output340
timestamp 1688980957
transform 1 0 17204 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output341
timestamp 1688980957
transform 1 0 17756 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output342
timestamp 1688980957
transform 1 0 17572 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output343
timestamp 1688980957
transform 1 0 20700 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output344
timestamp 1688980957
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  output345
timestamp 1688980957
transform 1 0 21344 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  output346
timestamp 1688980957
transform 1 0 3036 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output347
timestamp 1688980957
transform 1 0 4324 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output348
timestamp 1688980957
transform 1 0 1564 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output349
timestamp 1688980957
transform 1 0 1380 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output350
timestamp 1688980957
transform 1 0 3036 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output351
timestamp 1688980957
transform 1 0 3772 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output352
timestamp 1688980957
transform 1 0 2116 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output353
timestamp 1688980957
transform 1 0 4508 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output354
timestamp 1688980957
transform 1 0 3588 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output355
timestamp 1688980957
transform 1 0 5612 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output356
timestamp 1688980957
transform 1 0 5152 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output357
timestamp 1688980957
transform 1 0 1564 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output358
timestamp 1688980957
transform 1 0 3128 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output359
timestamp 1688980957
transform 1 0 1748 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output360
timestamp 1688980957
transform 1 0 5060 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output361
timestamp 1688980957
transform 1 0 3772 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output362
timestamp 1688980957
transform 1 0 4324 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output363
timestamp 1688980957
transform 1 0 4324 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output364
timestamp 1688980957
transform 1 0 1748 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output365
timestamp 1688980957
transform 1 0 5704 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output366
timestamp 1688980957
transform 1 0 2944 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output367
timestamp 1688980957
transform 1 0 3128 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output368
timestamp 1688980957
transform 1 0 3036 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output369
timestamp 1688980957
transform 1 0 2852 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output370
timestamp 1688980957
transform 1 0 3036 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output371
timestamp 1688980957
transform 1 0 2484 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output372
timestamp 1688980957
transform 1 0 1932 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output373
timestamp 1688980957
transform 1 0 1380 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output374
timestamp 1688980957
transform 1 0 3772 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output375
timestamp 1688980957
transform 1 0 3496 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output376
timestamp 1688980957
transform 1 0 1380 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output377
timestamp 1688980957
transform 1 0 3956 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output378
timestamp 1688980957
transform 1 0 4876 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output379
timestamp 1688980957
transform 1 0 2116 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output380
timestamp 1688980957
transform 1 0 1380 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output381
timestamp 1688980957
transform 1 0 4600 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output382
timestamp 1688980957
transform 1 0 1564 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output383
timestamp 1688980957
transform 1 0 1380 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output384
timestamp 1688980957
transform 1 0 3772 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output385
timestamp 1688980957
transform 1 0 5428 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output386
timestamp 1688980957
transform 1 0 3772 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output387
timestamp 1688980957
transform 1 0 2760 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output388
timestamp 1688980957
transform 1 0 1380 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output389
timestamp 1688980957
transform 1 0 3956 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output390
timestamp 1688980957
transform 1 0 3128 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output391
timestamp 1688980957
transform 1 0 4508 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output392
timestamp 1688980957
transform 1 0 1564 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output393
timestamp 1688980957
transform 1 0 4324 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1688980957
transform 1 0 1104 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1688980957
transform -1 0 24564 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1688980957
transform 1 0 1104 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1688980957
transform -1 0 24564 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1688980957
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1688980957
transform -1 0 24564 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1688980957
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1688980957
transform -1 0 24564 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1688980957
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1688980957
transform -1 0 24564 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1688980957
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1688980957
transform -1 0 24564 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1688980957
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1688980957
transform -1 0 24564 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1688980957
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1688980957
transform -1 0 24564 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1688980957
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1688980957
transform -1 0 24564 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1688980957
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1688980957
transform -1 0 24564 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1688980957
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1688980957
transform -1 0 24564 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1688980957
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1688980957
transform -1 0 24564 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1688980957
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1688980957
transform -1 0 24564 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1688980957
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1688980957
transform -1 0 24564 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1688980957
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1688980957
transform -1 0 24564 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1688980957
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1688980957
transform -1 0 24564 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1688980957
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1688980957
transform -1 0 24564 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1688980957
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1688980957
transform -1 0 24564 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1688980957
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1688980957
transform -1 0 24564 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1688980957
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1688980957
transform -1 0 24564 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1688980957
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1688980957
transform -1 0 24564 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1688980957
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1688980957
transform -1 0 24564 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1688980957
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1688980957
transform -1 0 24564 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1688980957
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1688980957
transform -1 0 24564 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1688980957
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1688980957
transform -1 0 24564 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1688980957
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1688980957
transform -1 0 24564 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1688980957
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1688980957
transform -1 0 24564 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1688980957
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1688980957
transform -1 0 24564 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1688980957
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1688980957
transform -1 0 24564 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1688980957
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1688980957
transform -1 0 24564 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1688980957
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1688980957
transform -1 0 24564 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1688980957
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1688980957
transform -1 0 24564 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1688980957
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1688980957
transform -1 0 24564 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1688980957
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1688980957
transform -1 0 24564 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1688980957
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1688980957
transform -1 0 24564 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1688980957
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1688980957
transform -1 0 24564 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1688980957
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1688980957
transform -1 0 24564 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1688980957
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1688980957
transform -1 0 24564 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1688980957
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1688980957
transform -1 0 24564 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1688980957
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1688980957
transform -1 0 24564 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1688980957
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1688980957
transform -1 0 24564 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1688980957
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1688980957
transform -1 0 24564 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1688980957
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1688980957
transform -1 0 24564 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1688980957
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1688980957
transform -1 0 24564 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1688980957
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1688980957
transform -1 0 24564 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1688980957
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1688980957
transform -1 0 24564 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1688980957
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1688980957
transform -1 0 24564 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1688980957
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1688980957
transform -1 0 24564 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1688980957
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1688980957
transform -1 0 24564 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1688980957
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1688980957
transform -1 0 24564 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1688980957
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1688980957
transform -1 0 24564 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1688980957
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1688980957
transform -1 0 24564 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1688980957
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1688980957
transform -1 0 24564 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1688980957
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1688980957
transform -1 0 24564 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1688980957
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1688980957
transform -1 0 24564 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1688980957
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1688980957
transform -1 0 24564 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1688980957
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1688980957
transform -1 0 24564 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1688980957
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1688980957
transform -1 0 24564 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1688980957
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1688980957
transform -1 0 24564 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1688980957
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1688980957
transform -1 0 24564 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1688980957
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1688980957
transform -1 0 24564 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1688980957
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1688980957
transform -1 0 24564 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1688980957
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1688980957
transform -1 0 24564 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1688980957
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1688980957
transform -1 0 24564 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1688980957
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1688980957
transform -1 0 24564 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1688980957
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1688980957
transform -1 0 24564 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1688980957
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1688980957
transform -1 0 24564 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1688980957
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1688980957
transform -1 0 24564 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1688980957
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1688980957
transform -1 0 24564 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1688980957
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1688980957
transform -1 0 24564 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1688980957
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1688980957
transform -1 0 24564 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1688980957
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1688980957
transform -1 0 24564 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1688980957
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1688980957
transform -1 0 24564 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1688980957
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1688980957
transform -1 0 24564 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1688980957
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1688980957
transform -1 0 24564 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1688980957
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1688980957
transform -1 0 24564 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1688980957
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1688980957
transform -1 0 24564 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1688980957
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1688980957
transform -1 0 24564 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  S4BEG_outbuf_0__0_
timestamp 1688980957
transform 1 0 16284 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  S4BEG_outbuf_1__0_
timestamp 1688980957
transform 1 0 16100 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  S4BEG_outbuf_2__0_
timestamp 1688980957
transform 1 0 16376 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  S4BEG_outbuf_3__0_
timestamp 1688980957
transform 1 0 16652 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  S4BEG_outbuf_4__0_
timestamp 1688980957
transform 1 0 16928 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  S4BEG_outbuf_5__0_
timestamp 1688980957
transform 1 0 24012 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  S4BEG_outbuf_6__0_
timestamp 1688980957
transform 1 0 17020 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  S4BEG_outbuf_7__0_
timestamp 1688980957
transform 1 0 19228 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  S4BEG_outbuf_8__0_
timestamp 1688980957
transform 1 0 18124 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  S4BEG_outbuf_9__0_
timestamp 1688980957
transform 1 0 18584 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  S4BEG_outbuf_10__0_
timestamp 1688980957
transform 1 0 21436 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  S4BEG_outbuf_11__0_
timestamp 1688980957
transform 1 0 24012 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  S4END_inbuf_0__0_
timestamp 1688980957
transform 1 0 16192 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  S4END_inbuf_1__0_
timestamp 1688980957
transform 1 0 16560 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  S4END_inbuf_2__0_
timestamp 1688980957
transform 1 0 16928 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  S4END_inbuf_3__0_
timestamp 1688980957
transform 1 0 17296 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  S4END_inbuf_4__0_
timestamp 1688980957
transform 1 0 17664 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  S4END_inbuf_5__0_
timestamp 1688980957
transform 1 0 18032 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  S4END_inbuf_6__0_
timestamp 1688980957
transform 1 0 18400 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  S4END_inbuf_7__0_
timestamp 1688980957
transform 1 0 18768 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  S4END_inbuf_8__0_
timestamp 1688980957
transform 1 0 18308 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  S4END_inbuf_9__0_
timestamp 1688980957
transform 1 0 19228 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  S4END_inbuf_10__0_
timestamp 1688980957
transform 1 0 19596 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  S4END_inbuf_11__0_
timestamp 1688980957
transform 1 0 19228 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_0__0_
timestamp 1688980957
transform 1 0 19872 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_1__0_
timestamp 1688980957
transform 1 0 20792 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_2__0_
timestamp 1688980957
transform 1 0 20332 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_3__0_
timestamp 1688980957
transform 1 0 20608 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_4__0_
timestamp 1688980957
transform 1 0 21620 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  strobe_inbuf_5__0_
timestamp 1688980957
transform 1 0 21160 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_6__0_
timestamp 1688980957
transform 1 0 21436 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_7__0_
timestamp 1688980957
transform 1 0 21068 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_8__0_
timestamp 1688980957
transform 1 0 22172 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_9__0_
timestamp 1688980957
transform 1 0 19596 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  strobe_inbuf_10__0_
timestamp 1688980957
transform 1 0 22816 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_11__0_
timestamp 1688980957
transform 1 0 22816 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_12__0_
timestamp 1688980957
transform 1 0 22632 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_13__0_
timestamp 1688980957
transform 1 0 20884 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_14__0_
timestamp 1688980957
transform 1 0 23460 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_15__0_
timestamp 1688980957
transform 1 0 23644 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_16__0_
timestamp 1688980957
transform 1 0 23644 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_17__0_
timestamp 1688980957
transform 1 0 23644 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_18__0_
timestamp 1688980957
transform 1 0 23184 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_19__0_
timestamp 1688980957
transform 1 0 23644 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_0__0_
timestamp 1688980957
transform 1 0 20240 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_1__0_
timestamp 1688980957
transform 1 0 20608 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_2__0_
timestamp 1688980957
transform 1 0 23276 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_3__0_
timestamp 1688980957
transform 1 0 20884 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_4__0_
timestamp 1688980957
transform 1 0 21436 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_5__0_
timestamp 1688980957
transform 1 0 20332 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_6__0_
timestamp 1688980957
transform 1 0 21804 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_7__0_
timestamp 1688980957
transform 1 0 22908 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_8__0_
timestamp 1688980957
transform 1 0 22264 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_9__0_
timestamp 1688980957
transform 1 0 22908 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_10__0_
timestamp 1688980957
transform 1 0 21988 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_11__0_
timestamp 1688980957
transform 1 0 21436 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_12__0_
timestamp 1688980957
transform 1 0 23184 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_13__0_
timestamp 1688980957
transform 1 0 21896 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_14__0_
timestamp 1688980957
transform 1 0 21160 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_15__0_
timestamp 1688980957
transform 1 0 23092 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_16__0_
timestamp 1688980957
transform 1 0 23368 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_17__0_
timestamp 1688980957
transform 1 0 23460 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  strobe_outbuf_18__0_
timestamp 1688980957
transform 1 0 23644 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_19__0_
timestamp 1688980957
transform 1 0 23368 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3680 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1688980957
transform 1 0 6256 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1688980957
transform 1 0 8832 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1688980957
transform 1 0 11408 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1688980957
transform 1 0 13984 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1688980957
transform 1 0 16560 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1688980957
transform 1 0 19136 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1688980957
transform 1 0 21712 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1688980957
transform 1 0 6256 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1688980957
transform 1 0 11408 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1688980957
transform 1 0 16560 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1688980957
transform 1 0 21712 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1688980957
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1688980957
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1688980957
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1688980957
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1688980957
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1688980957
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1688980957
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1688980957
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1688980957
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1688980957
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1688980957
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1688980957
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1688980957
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1688980957
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1688980957
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1688980957
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1688980957
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1688980957
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1688980957
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1688980957
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1688980957
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1688980957
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1688980957
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1688980957
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1688980957
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1688980957
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1688980957
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1688980957
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1688980957
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1688980957
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1688980957
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1688980957
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1688980957
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1688980957
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1688980957
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1688980957
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1688980957
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1688980957
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1688980957
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1688980957
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1688980957
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1688980957
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1688980957
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1688980957
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1688980957
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1688980957
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1688980957
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1688980957
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1688980957
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1688980957
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1688980957
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1688980957
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1688980957
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1688980957
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1688980957
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1688980957
transform 1 0 21712 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1688980957
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1688980957
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1688980957
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1688980957
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1688980957
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1688980957
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1688980957
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1688980957
transform 1 0 21712 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1688980957
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1688980957
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1688980957
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1688980957
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1688980957
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1688980957
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1688980957
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1688980957
transform 1 0 21712 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1688980957
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1688980957
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1688980957
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1688980957
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1688980957
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1688980957
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1688980957
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1688980957
transform 1 0 21712 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1688980957
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1688980957
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1688980957
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1688980957
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1688980957
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1688980957
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1688980957
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1688980957
transform 1 0 21712 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1688980957
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1688980957
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1688980957
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1688980957
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1688980957
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1688980957
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1688980957
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1688980957
transform 1 0 21712 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1688980957
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1688980957
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1688980957
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1688980957
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1688980957
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1688980957
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1688980957
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1688980957
transform 1 0 21712 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1688980957
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1688980957
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1688980957
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1688980957
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1688980957
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1688980957
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1688980957
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1688980957
transform 1 0 21712 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1688980957
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1688980957
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1688980957
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1688980957
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1688980957
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1688980957
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1688980957
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1688980957
transform 1 0 21712 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1688980957
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1688980957
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1688980957
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1688980957
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1688980957
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1688980957
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1688980957
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1688980957
transform 1 0 21712 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1688980957
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1688980957
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1688980957
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1688980957
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1688980957
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1688980957
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1688980957
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1688980957
transform 1 0 21712 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1688980957
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1688980957
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1688980957
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1688980957
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1688980957
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1688980957
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1688980957
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1688980957
transform 1 0 21712 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1688980957
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1688980957
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1688980957
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1688980957
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1688980957
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1688980957
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1688980957
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1688980957
transform 1 0 21712 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1688980957
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1688980957
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1688980957
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1688980957
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1688980957
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1688980957
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1688980957
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1688980957
transform 1 0 21712 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1688980957
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1688980957
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1688980957
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1688980957
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1688980957
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1688980957
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1688980957
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1688980957
transform 1 0 21712 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1688980957
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1688980957
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1688980957
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1688980957
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1688980957
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1688980957
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1688980957
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1688980957
transform 1 0 21712 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1688980957
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1688980957
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1688980957
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1688980957
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1688980957
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1688980957
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1688980957
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1688980957
transform 1 0 21712 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1688980957
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1688980957
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1688980957
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1688980957
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1688980957
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1688980957
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1688980957
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1688980957
transform 1 0 21712 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1688980957
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1688980957
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1688980957
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1688980957
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1688980957
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1688980957
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1688980957
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1688980957
transform 1 0 21712 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1688980957
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1688980957
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1688980957
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1688980957
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1688980957
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1688980957
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1688980957
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1688980957
transform 1 0 21712 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1688980957
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1688980957
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1688980957
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1688980957
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1688980957
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1688980957
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1688980957
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1688980957
transform 1 0 21712 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1688980957
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1688980957
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1688980957
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1688980957
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1688980957
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1688980957
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1688980957
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1688980957
transform 1 0 21712 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1688980957
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1688980957
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1688980957
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1688980957
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1688980957
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1688980957
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1688980957
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1688980957
transform 1 0 21712 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1688980957
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1688980957
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1688980957
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1688980957
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1688980957
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1688980957
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1688980957
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1688980957
transform 1 0 21712 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1688980957
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1688980957
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1688980957
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1688980957
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1688980957
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1688980957
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1688980957
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1688980957
transform 1 0 21712 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1688980957
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1688980957
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1688980957
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1688980957
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1688980957
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1688980957
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1688980957
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1688980957
transform 1 0 21712 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1688980957
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1688980957
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1688980957
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1688980957
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1688980957
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1688980957
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1688980957
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1688980957
transform 1 0 21712 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1688980957
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1688980957
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1688980957
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1688980957
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_436
timestamp 1688980957
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_437
timestamp 1688980957
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_438
timestamp 1688980957
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_439
timestamp 1688980957
transform 1 0 21712 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_440
timestamp 1688980957
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_441
timestamp 1688980957
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_442
timestamp 1688980957
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_443
timestamp 1688980957
transform 1 0 19136 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_444
timestamp 1688980957
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_445
timestamp 1688980957
transform 1 0 11408 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_446
timestamp 1688980957
transform 1 0 16560 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_447
timestamp 1688980957
transform 1 0 21712 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_448
timestamp 1688980957
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_449
timestamp 1688980957
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_450
timestamp 1688980957
transform 1 0 13984 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_451
timestamp 1688980957
transform 1 0 19136 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_452
timestamp 1688980957
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_453
timestamp 1688980957
transform 1 0 11408 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_454
timestamp 1688980957
transform 1 0 16560 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_455
timestamp 1688980957
transform 1 0 21712 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_456
timestamp 1688980957
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_457
timestamp 1688980957
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_458
timestamp 1688980957
transform 1 0 13984 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_459
timestamp 1688980957
transform 1 0 19136 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_460
timestamp 1688980957
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_461
timestamp 1688980957
transform 1 0 11408 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_462
timestamp 1688980957
transform 1 0 16560 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_463
timestamp 1688980957
transform 1 0 21712 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_464
timestamp 1688980957
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_465
timestamp 1688980957
transform 1 0 8832 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_466
timestamp 1688980957
transform 1 0 13984 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_467
timestamp 1688980957
transform 1 0 19136 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_468
timestamp 1688980957
transform 1 0 3680 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_469
timestamp 1688980957
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_470
timestamp 1688980957
transform 1 0 8832 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_471
timestamp 1688980957
transform 1 0 11408 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_472
timestamp 1688980957
transform 1 0 13984 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_473
timestamp 1688980957
transform 1 0 16560 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_474
timestamp 1688980957
transform 1 0 19136 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_475
timestamp 1688980957
transform 1 0 21712 0 -1 43520
box -38 -48 130 592
<< labels >>
flabel metal3 s 25540 9256 26000 9376 0 FreeSans 480 0 0 0 Config_accessC_bit0
port 0 nsew signal tristate
flabel metal3 s 25540 9800 26000 9920 0 FreeSans 480 0 0 0 Config_accessC_bit1
port 1 nsew signal tristate
flabel metal3 s 25540 10344 26000 10464 0 FreeSans 480 0 0 0 Config_accessC_bit2
port 2 nsew signal tristate
flabel metal3 s 25540 10888 26000 11008 0 FreeSans 480 0 0 0 Config_accessC_bit3
port 3 nsew signal tristate
flabel metal3 s -300 17960 160 18080 0 FreeSans 480 0 0 0 E1END[0]
port 4 nsew signal input
flabel metal3 s -300 18232 160 18352 0 FreeSans 480 0 0 0 E1END[1]
port 5 nsew signal input
flabel metal3 s -300 18504 160 18624 0 FreeSans 480 0 0 0 E1END[2]
port 6 nsew signal input
flabel metal3 s -300 18776 160 18896 0 FreeSans 480 0 0 0 E1END[3]
port 7 nsew signal input
flabel metal3 s -300 21224 160 21344 0 FreeSans 480 0 0 0 E2END[0]
port 8 nsew signal input
flabel metal3 s -300 21496 160 21616 0 FreeSans 480 0 0 0 E2END[1]
port 9 nsew signal input
flabel metal3 s -300 21768 160 21888 0 FreeSans 480 0 0 0 E2END[2]
port 10 nsew signal input
flabel metal3 s -300 22040 160 22160 0 FreeSans 480 0 0 0 E2END[3]
port 11 nsew signal input
flabel metal3 s -300 22312 160 22432 0 FreeSans 480 0 0 0 E2END[4]
port 12 nsew signal input
flabel metal3 s -300 22584 160 22704 0 FreeSans 480 0 0 0 E2END[5]
port 13 nsew signal input
flabel metal3 s -300 22856 160 22976 0 FreeSans 480 0 0 0 E2END[6]
port 14 nsew signal input
flabel metal3 s -300 23128 160 23248 0 FreeSans 480 0 0 0 E2END[7]
port 15 nsew signal input
flabel metal3 s -300 19048 160 19168 0 FreeSans 480 0 0 0 E2MID[0]
port 16 nsew signal input
flabel metal3 s -300 19320 160 19440 0 FreeSans 480 0 0 0 E2MID[1]
port 17 nsew signal input
flabel metal3 s -300 19592 160 19712 0 FreeSans 480 0 0 0 E2MID[2]
port 18 nsew signal input
flabel metal3 s -300 19864 160 19984 0 FreeSans 480 0 0 0 E2MID[3]
port 19 nsew signal input
flabel metal3 s -300 20136 160 20256 0 FreeSans 480 0 0 0 E2MID[4]
port 20 nsew signal input
flabel metal3 s -300 20408 160 20528 0 FreeSans 480 0 0 0 E2MID[5]
port 21 nsew signal input
flabel metal3 s -300 20680 160 20800 0 FreeSans 480 0 0 0 E2MID[6]
port 22 nsew signal input
flabel metal3 s -300 20952 160 21072 0 FreeSans 480 0 0 0 E2MID[7]
port 23 nsew signal input
flabel metal3 s -300 27752 160 27872 0 FreeSans 480 0 0 0 E6END[0]
port 24 nsew signal input
flabel metal3 s -300 30472 160 30592 0 FreeSans 480 0 0 0 E6END[10]
port 25 nsew signal input
flabel metal3 s -300 30744 160 30864 0 FreeSans 480 0 0 0 E6END[11]
port 26 nsew signal input
flabel metal3 s -300 28024 160 28144 0 FreeSans 480 0 0 0 E6END[1]
port 27 nsew signal input
flabel metal3 s -300 28296 160 28416 0 FreeSans 480 0 0 0 E6END[2]
port 28 nsew signal input
flabel metal3 s -300 28568 160 28688 0 FreeSans 480 0 0 0 E6END[3]
port 29 nsew signal input
flabel metal3 s -300 28840 160 28960 0 FreeSans 480 0 0 0 E6END[4]
port 30 nsew signal input
flabel metal3 s -300 29112 160 29232 0 FreeSans 480 0 0 0 E6END[5]
port 31 nsew signal input
flabel metal3 s -300 29384 160 29504 0 FreeSans 480 0 0 0 E6END[6]
port 32 nsew signal input
flabel metal3 s -300 29656 160 29776 0 FreeSans 480 0 0 0 E6END[7]
port 33 nsew signal input
flabel metal3 s -300 29928 160 30048 0 FreeSans 480 0 0 0 E6END[8]
port 34 nsew signal input
flabel metal3 s -300 30200 160 30320 0 FreeSans 480 0 0 0 E6END[9]
port 35 nsew signal input
flabel metal3 s -300 23400 160 23520 0 FreeSans 480 0 0 0 EE4END[0]
port 36 nsew signal input
flabel metal3 s -300 26120 160 26240 0 FreeSans 480 0 0 0 EE4END[10]
port 37 nsew signal input
flabel metal3 s -300 26392 160 26512 0 FreeSans 480 0 0 0 EE4END[11]
port 38 nsew signal input
flabel metal3 s -300 26664 160 26784 0 FreeSans 480 0 0 0 EE4END[12]
port 39 nsew signal input
flabel metal3 s -300 26936 160 27056 0 FreeSans 480 0 0 0 EE4END[13]
port 40 nsew signal input
flabel metal3 s -300 27208 160 27328 0 FreeSans 480 0 0 0 EE4END[14]
port 41 nsew signal input
flabel metal3 s -300 27480 160 27600 0 FreeSans 480 0 0 0 EE4END[15]
port 42 nsew signal input
flabel metal3 s -300 23672 160 23792 0 FreeSans 480 0 0 0 EE4END[1]
port 43 nsew signal input
flabel metal3 s -300 23944 160 24064 0 FreeSans 480 0 0 0 EE4END[2]
port 44 nsew signal input
flabel metal3 s -300 24216 160 24336 0 FreeSans 480 0 0 0 EE4END[3]
port 45 nsew signal input
flabel metal3 s -300 24488 160 24608 0 FreeSans 480 0 0 0 EE4END[4]
port 46 nsew signal input
flabel metal3 s -300 24760 160 24880 0 FreeSans 480 0 0 0 EE4END[5]
port 47 nsew signal input
flabel metal3 s -300 25032 160 25152 0 FreeSans 480 0 0 0 EE4END[6]
port 48 nsew signal input
flabel metal3 s -300 25304 160 25424 0 FreeSans 480 0 0 0 EE4END[7]
port 49 nsew signal input
flabel metal3 s -300 25576 160 25696 0 FreeSans 480 0 0 0 EE4END[8]
port 50 nsew signal input
flabel metal3 s -300 25848 160 25968 0 FreeSans 480 0 0 0 EE4END[9]
port 51 nsew signal input
flabel metal3 s 25540 15784 26000 15904 0 FreeSans 480 0 0 0 FAB2RAM_A0_O0
port 52 nsew signal tristate
flabel metal3 s 25540 16328 26000 16448 0 FreeSans 480 0 0 0 FAB2RAM_A0_O1
port 53 nsew signal tristate
flabel metal3 s 25540 16872 26000 16992 0 FreeSans 480 0 0 0 FAB2RAM_A0_O2
port 54 nsew signal tristate
flabel metal3 s 25540 17416 26000 17536 0 FreeSans 480 0 0 0 FAB2RAM_A0_O3
port 55 nsew signal tristate
flabel metal3 s 25540 13608 26000 13728 0 FreeSans 480 0 0 0 FAB2RAM_A1_O0
port 56 nsew signal tristate
flabel metal3 s 25540 14152 26000 14272 0 FreeSans 480 0 0 0 FAB2RAM_A1_O1
port 57 nsew signal tristate
flabel metal3 s 25540 14696 26000 14816 0 FreeSans 480 0 0 0 FAB2RAM_A1_O2
port 58 nsew signal tristate
flabel metal3 s 25540 15240 26000 15360 0 FreeSans 480 0 0 0 FAB2RAM_A1_O3
port 59 nsew signal tristate
flabel metal3 s 25540 11432 26000 11552 0 FreeSans 480 0 0 0 FAB2RAM_C_O0
port 60 nsew signal tristate
flabel metal3 s 25540 11976 26000 12096 0 FreeSans 480 0 0 0 FAB2RAM_C_O1
port 61 nsew signal tristate
flabel metal3 s 25540 12520 26000 12640 0 FreeSans 480 0 0 0 FAB2RAM_C_O2
port 62 nsew signal tristate
flabel metal3 s 25540 13064 26000 13184 0 FreeSans 480 0 0 0 FAB2RAM_C_O3
port 63 nsew signal tristate
flabel metal3 s 25540 24488 26000 24608 0 FreeSans 480 0 0 0 FAB2RAM_D0_O0
port 64 nsew signal tristate
flabel metal3 s 25540 25032 26000 25152 0 FreeSans 480 0 0 0 FAB2RAM_D0_O1
port 65 nsew signal tristate
flabel metal3 s 25540 25576 26000 25696 0 FreeSans 480 0 0 0 FAB2RAM_D0_O2
port 66 nsew signal tristate
flabel metal3 s 25540 26120 26000 26240 0 FreeSans 480 0 0 0 FAB2RAM_D0_O3
port 67 nsew signal tristate
flabel metal3 s 25540 22312 26000 22432 0 FreeSans 480 0 0 0 FAB2RAM_D1_O0
port 68 nsew signal tristate
flabel metal3 s 25540 22856 26000 22976 0 FreeSans 480 0 0 0 FAB2RAM_D1_O1
port 69 nsew signal tristate
flabel metal3 s 25540 23400 26000 23520 0 FreeSans 480 0 0 0 FAB2RAM_D1_O2
port 70 nsew signal tristate
flabel metal3 s 25540 23944 26000 24064 0 FreeSans 480 0 0 0 FAB2RAM_D1_O3
port 71 nsew signal tristate
flabel metal3 s 25540 20136 26000 20256 0 FreeSans 480 0 0 0 FAB2RAM_D2_O0
port 72 nsew signal tristate
flabel metal3 s 25540 20680 26000 20800 0 FreeSans 480 0 0 0 FAB2RAM_D2_O1
port 73 nsew signal tristate
flabel metal3 s 25540 21224 26000 21344 0 FreeSans 480 0 0 0 FAB2RAM_D2_O2
port 74 nsew signal tristate
flabel metal3 s 25540 21768 26000 21888 0 FreeSans 480 0 0 0 FAB2RAM_D2_O3
port 75 nsew signal tristate
flabel metal3 s 25540 17960 26000 18080 0 FreeSans 480 0 0 0 FAB2RAM_D3_O0
port 76 nsew signal tristate
flabel metal3 s 25540 18504 26000 18624 0 FreeSans 480 0 0 0 FAB2RAM_D3_O1
port 77 nsew signal tristate
flabel metal3 s 25540 19048 26000 19168 0 FreeSans 480 0 0 0 FAB2RAM_D3_O2
port 78 nsew signal tristate
flabel metal3 s 25540 19592 26000 19712 0 FreeSans 480 0 0 0 FAB2RAM_D3_O3
port 79 nsew signal tristate
flabel metal3 s -300 31016 160 31136 0 FreeSans 480 0 0 0 FrameData[0]
port 80 nsew signal input
flabel metal3 s -300 33736 160 33856 0 FreeSans 480 0 0 0 FrameData[10]
port 81 nsew signal input
flabel metal3 s -300 34008 160 34128 0 FreeSans 480 0 0 0 FrameData[11]
port 82 nsew signal input
flabel metal3 s -300 34280 160 34400 0 FreeSans 480 0 0 0 FrameData[12]
port 83 nsew signal input
flabel metal3 s -300 34552 160 34672 0 FreeSans 480 0 0 0 FrameData[13]
port 84 nsew signal input
flabel metal3 s -300 34824 160 34944 0 FreeSans 480 0 0 0 FrameData[14]
port 85 nsew signal input
flabel metal3 s -300 35096 160 35216 0 FreeSans 480 0 0 0 FrameData[15]
port 86 nsew signal input
flabel metal3 s -300 35368 160 35488 0 FreeSans 480 0 0 0 FrameData[16]
port 87 nsew signal input
flabel metal3 s -300 35640 160 35760 0 FreeSans 480 0 0 0 FrameData[17]
port 88 nsew signal input
flabel metal3 s -300 35912 160 36032 0 FreeSans 480 0 0 0 FrameData[18]
port 89 nsew signal input
flabel metal3 s -300 36184 160 36304 0 FreeSans 480 0 0 0 FrameData[19]
port 90 nsew signal input
flabel metal3 s -300 31288 160 31408 0 FreeSans 480 0 0 0 FrameData[1]
port 91 nsew signal input
flabel metal3 s -300 36456 160 36576 0 FreeSans 480 0 0 0 FrameData[20]
port 92 nsew signal input
flabel metal3 s -300 36728 160 36848 0 FreeSans 480 0 0 0 FrameData[21]
port 93 nsew signal input
flabel metal3 s -300 37000 160 37120 0 FreeSans 480 0 0 0 FrameData[22]
port 94 nsew signal input
flabel metal3 s -300 37272 160 37392 0 FreeSans 480 0 0 0 FrameData[23]
port 95 nsew signal input
flabel metal3 s -300 37544 160 37664 0 FreeSans 480 0 0 0 FrameData[24]
port 96 nsew signal input
flabel metal3 s -300 37816 160 37936 0 FreeSans 480 0 0 0 FrameData[25]
port 97 nsew signal input
flabel metal3 s -300 38088 160 38208 0 FreeSans 480 0 0 0 FrameData[26]
port 98 nsew signal input
flabel metal3 s -300 38360 160 38480 0 FreeSans 480 0 0 0 FrameData[27]
port 99 nsew signal input
flabel metal3 s -300 38632 160 38752 0 FreeSans 480 0 0 0 FrameData[28]
port 100 nsew signal input
flabel metal3 s -300 38904 160 39024 0 FreeSans 480 0 0 0 FrameData[29]
port 101 nsew signal input
flabel metal3 s -300 31560 160 31680 0 FreeSans 480 0 0 0 FrameData[2]
port 102 nsew signal input
flabel metal3 s -300 39176 160 39296 0 FreeSans 480 0 0 0 FrameData[30]
port 103 nsew signal input
flabel metal3 s -300 39448 160 39568 0 FreeSans 480 0 0 0 FrameData[31]
port 104 nsew signal input
flabel metal3 s -300 31832 160 31952 0 FreeSans 480 0 0 0 FrameData[3]
port 105 nsew signal input
flabel metal3 s -300 32104 160 32224 0 FreeSans 480 0 0 0 FrameData[4]
port 106 nsew signal input
flabel metal3 s -300 32376 160 32496 0 FreeSans 480 0 0 0 FrameData[5]
port 107 nsew signal input
flabel metal3 s -300 32648 160 32768 0 FreeSans 480 0 0 0 FrameData[6]
port 108 nsew signal input
flabel metal3 s -300 32920 160 33040 0 FreeSans 480 0 0 0 FrameData[7]
port 109 nsew signal input
flabel metal3 s -300 33192 160 33312 0 FreeSans 480 0 0 0 FrameData[8]
port 110 nsew signal input
flabel metal3 s -300 33464 160 33584 0 FreeSans 480 0 0 0 FrameData[9]
port 111 nsew signal input
flabel metal3 s 25540 26664 26000 26784 0 FreeSans 480 0 0 0 FrameData_O[0]
port 112 nsew signal tristate
flabel metal3 s 25540 32104 26000 32224 0 FreeSans 480 0 0 0 FrameData_O[10]
port 113 nsew signal tristate
flabel metal3 s 25540 32648 26000 32768 0 FreeSans 480 0 0 0 FrameData_O[11]
port 114 nsew signal tristate
flabel metal3 s 25540 33192 26000 33312 0 FreeSans 480 0 0 0 FrameData_O[12]
port 115 nsew signal tristate
flabel metal3 s 25540 33736 26000 33856 0 FreeSans 480 0 0 0 FrameData_O[13]
port 116 nsew signal tristate
flabel metal3 s 25540 34280 26000 34400 0 FreeSans 480 0 0 0 FrameData_O[14]
port 117 nsew signal tristate
flabel metal3 s 25540 34824 26000 34944 0 FreeSans 480 0 0 0 FrameData_O[15]
port 118 nsew signal tristate
flabel metal3 s 25540 35368 26000 35488 0 FreeSans 480 0 0 0 FrameData_O[16]
port 119 nsew signal tristate
flabel metal3 s 25540 35912 26000 36032 0 FreeSans 480 0 0 0 FrameData_O[17]
port 120 nsew signal tristate
flabel metal3 s 25540 36456 26000 36576 0 FreeSans 480 0 0 0 FrameData_O[18]
port 121 nsew signal tristate
flabel metal3 s 25540 37000 26000 37120 0 FreeSans 480 0 0 0 FrameData_O[19]
port 122 nsew signal tristate
flabel metal3 s 25540 27208 26000 27328 0 FreeSans 480 0 0 0 FrameData_O[1]
port 123 nsew signal tristate
flabel metal3 s 25540 37544 26000 37664 0 FreeSans 480 0 0 0 FrameData_O[20]
port 124 nsew signal tristate
flabel metal3 s 25540 38088 26000 38208 0 FreeSans 480 0 0 0 FrameData_O[21]
port 125 nsew signal tristate
flabel metal3 s 25540 38632 26000 38752 0 FreeSans 480 0 0 0 FrameData_O[22]
port 126 nsew signal tristate
flabel metal3 s 25540 39176 26000 39296 0 FreeSans 480 0 0 0 FrameData_O[23]
port 127 nsew signal tristate
flabel metal3 s 25540 39720 26000 39840 0 FreeSans 480 0 0 0 FrameData_O[24]
port 128 nsew signal tristate
flabel metal3 s 25540 40264 26000 40384 0 FreeSans 480 0 0 0 FrameData_O[25]
port 129 nsew signal tristate
flabel metal3 s 25540 40808 26000 40928 0 FreeSans 480 0 0 0 FrameData_O[26]
port 130 nsew signal tristate
flabel metal3 s 25540 41352 26000 41472 0 FreeSans 480 0 0 0 FrameData_O[27]
port 131 nsew signal tristate
flabel metal3 s 25540 41896 26000 42016 0 FreeSans 480 0 0 0 FrameData_O[28]
port 132 nsew signal tristate
flabel metal3 s 25540 42440 26000 42560 0 FreeSans 480 0 0 0 FrameData_O[29]
port 133 nsew signal tristate
flabel metal3 s 25540 27752 26000 27872 0 FreeSans 480 0 0 0 FrameData_O[2]
port 134 nsew signal tristate
flabel metal3 s 25540 42984 26000 43104 0 FreeSans 480 0 0 0 FrameData_O[30]
port 135 nsew signal tristate
flabel metal3 s 25540 43528 26000 43648 0 FreeSans 480 0 0 0 FrameData_O[31]
port 136 nsew signal tristate
flabel metal3 s 25540 28296 26000 28416 0 FreeSans 480 0 0 0 FrameData_O[3]
port 137 nsew signal tristate
flabel metal3 s 25540 28840 26000 28960 0 FreeSans 480 0 0 0 FrameData_O[4]
port 138 nsew signal tristate
flabel metal3 s 25540 29384 26000 29504 0 FreeSans 480 0 0 0 FrameData_O[5]
port 139 nsew signal tristate
flabel metal3 s 25540 29928 26000 30048 0 FreeSans 480 0 0 0 FrameData_O[6]
port 140 nsew signal tristate
flabel metal3 s 25540 30472 26000 30592 0 FreeSans 480 0 0 0 FrameData_O[7]
port 141 nsew signal tristate
flabel metal3 s 25540 31016 26000 31136 0 FreeSans 480 0 0 0 FrameData_O[8]
port 142 nsew signal tristate
flabel metal3 s 25540 31560 26000 31680 0 FreeSans 480 0 0 0 FrameData_O[9]
port 143 nsew signal tristate
flabel metal2 s 20258 -300 20314 160 0 FreeSans 224 90 0 0 FrameStrobe[0]
port 144 nsew signal input
flabel metal2 s 23018 -300 23074 160 0 FreeSans 224 90 0 0 FrameStrobe[10]
port 145 nsew signal input
flabel metal2 s 23294 -300 23350 160 0 FreeSans 224 90 0 0 FrameStrobe[11]
port 146 nsew signal input
flabel metal2 s 23570 -300 23626 160 0 FreeSans 224 90 0 0 FrameStrobe[12]
port 147 nsew signal input
flabel metal2 s 23846 -300 23902 160 0 FreeSans 224 90 0 0 FrameStrobe[13]
port 148 nsew signal input
flabel metal2 s 24122 -300 24178 160 0 FreeSans 224 90 0 0 FrameStrobe[14]
port 149 nsew signal input
flabel metal2 s 24398 -300 24454 160 0 FreeSans 224 90 0 0 FrameStrobe[15]
port 150 nsew signal input
flabel metal2 s 24674 -300 24730 160 0 FreeSans 224 90 0 0 FrameStrobe[16]
port 151 nsew signal input
flabel metal2 s 24950 -300 25006 160 0 FreeSans 224 90 0 0 FrameStrobe[17]
port 152 nsew signal input
flabel metal2 s 25226 -300 25282 160 0 FreeSans 224 90 0 0 FrameStrobe[18]
port 153 nsew signal input
flabel metal2 s 25502 -300 25558 160 0 FreeSans 224 90 0 0 FrameStrobe[19]
port 154 nsew signal input
flabel metal2 s 20534 -300 20590 160 0 FreeSans 224 90 0 0 FrameStrobe[1]
port 155 nsew signal input
flabel metal2 s 20810 -300 20866 160 0 FreeSans 224 90 0 0 FrameStrobe[2]
port 156 nsew signal input
flabel metal2 s 21086 -300 21142 160 0 FreeSans 224 90 0 0 FrameStrobe[3]
port 157 nsew signal input
flabel metal2 s 21362 -300 21418 160 0 FreeSans 224 90 0 0 FrameStrobe[4]
port 158 nsew signal input
flabel metal2 s 21638 -300 21694 160 0 FreeSans 224 90 0 0 FrameStrobe[5]
port 159 nsew signal input
flabel metal2 s 21914 -300 21970 160 0 FreeSans 224 90 0 0 FrameStrobe[6]
port 160 nsew signal input
flabel metal2 s 22190 -300 22246 160 0 FreeSans 224 90 0 0 FrameStrobe[7]
port 161 nsew signal input
flabel metal2 s 22466 -300 22522 160 0 FreeSans 224 90 0 0 FrameStrobe[8]
port 162 nsew signal input
flabel metal2 s 22742 -300 22798 160 0 FreeSans 224 90 0 0 FrameStrobe[9]
port 163 nsew signal input
flabel metal2 s 20258 44540 20314 45000 0 FreeSans 224 90 0 0 FrameStrobe_O[0]
port 164 nsew signal tristate
flabel metal2 s 23018 44540 23074 45000 0 FreeSans 224 90 0 0 FrameStrobe_O[10]
port 165 nsew signal tristate
flabel metal2 s 23294 44540 23350 45000 0 FreeSans 224 90 0 0 FrameStrobe_O[11]
port 166 nsew signal tristate
flabel metal2 s 23570 44540 23626 45000 0 FreeSans 224 90 0 0 FrameStrobe_O[12]
port 167 nsew signal tristate
flabel metal2 s 23846 44540 23902 45000 0 FreeSans 224 90 0 0 FrameStrobe_O[13]
port 168 nsew signal tristate
flabel metal2 s 24122 44540 24178 45000 0 FreeSans 224 90 0 0 FrameStrobe_O[14]
port 169 nsew signal tristate
flabel metal2 s 24398 44540 24454 45000 0 FreeSans 224 90 0 0 FrameStrobe_O[15]
port 170 nsew signal tristate
flabel metal2 s 24674 44540 24730 45000 0 FreeSans 224 90 0 0 FrameStrobe_O[16]
port 171 nsew signal tristate
flabel metal2 s 24950 44540 25006 45000 0 FreeSans 224 90 0 0 FrameStrobe_O[17]
port 172 nsew signal tristate
flabel metal2 s 25226 44540 25282 45000 0 FreeSans 224 90 0 0 FrameStrobe_O[18]
port 173 nsew signal tristate
flabel metal2 s 25502 44540 25558 45000 0 FreeSans 224 90 0 0 FrameStrobe_O[19]
port 174 nsew signal tristate
flabel metal2 s 20534 44540 20590 45000 0 FreeSans 224 90 0 0 FrameStrobe_O[1]
port 175 nsew signal tristate
flabel metal2 s 20810 44540 20866 45000 0 FreeSans 224 90 0 0 FrameStrobe_O[2]
port 176 nsew signal tristate
flabel metal2 s 21086 44540 21142 45000 0 FreeSans 224 90 0 0 FrameStrobe_O[3]
port 177 nsew signal tristate
flabel metal2 s 21362 44540 21418 45000 0 FreeSans 224 90 0 0 FrameStrobe_O[4]
port 178 nsew signal tristate
flabel metal2 s 21638 44540 21694 45000 0 FreeSans 224 90 0 0 FrameStrobe_O[5]
port 179 nsew signal tristate
flabel metal2 s 21914 44540 21970 45000 0 FreeSans 224 90 0 0 FrameStrobe_O[6]
port 180 nsew signal tristate
flabel metal2 s 22190 44540 22246 45000 0 FreeSans 224 90 0 0 FrameStrobe_O[7]
port 181 nsew signal tristate
flabel metal2 s 22466 44540 22522 45000 0 FreeSans 224 90 0 0 FrameStrobe_O[8]
port 182 nsew signal tristate
flabel metal2 s 22742 44540 22798 45000 0 FreeSans 224 90 0 0 FrameStrobe_O[9]
port 183 nsew signal tristate
flabel metal2 s 110 44540 166 45000 0 FreeSans 224 90 0 0 N1BEG[0]
port 184 nsew signal tristate
flabel metal2 s 386 44540 442 45000 0 FreeSans 224 90 0 0 N1BEG[1]
port 185 nsew signal tristate
flabel metal2 s 662 44540 718 45000 0 FreeSans 224 90 0 0 N1BEG[2]
port 186 nsew signal tristate
flabel metal2 s 938 44540 994 45000 0 FreeSans 224 90 0 0 N1BEG[3]
port 187 nsew signal tristate
flabel metal2 s 110 -300 166 160 0 FreeSans 224 90 0 0 N1END[0]
port 188 nsew signal input
flabel metal2 s 386 -300 442 160 0 FreeSans 224 90 0 0 N1END[1]
port 189 nsew signal input
flabel metal2 s 662 -300 718 160 0 FreeSans 224 90 0 0 N1END[2]
port 190 nsew signal input
flabel metal2 s 938 -300 994 160 0 FreeSans 224 90 0 0 N1END[3]
port 191 nsew signal input
flabel metal2 s 1214 44540 1270 45000 0 FreeSans 224 90 0 0 N2BEG[0]
port 192 nsew signal tristate
flabel metal2 s 1490 44540 1546 45000 0 FreeSans 224 90 0 0 N2BEG[1]
port 193 nsew signal tristate
flabel metal2 s 1766 44540 1822 45000 0 FreeSans 224 90 0 0 N2BEG[2]
port 194 nsew signal tristate
flabel metal2 s 2042 44540 2098 45000 0 FreeSans 224 90 0 0 N2BEG[3]
port 195 nsew signal tristate
flabel metal2 s 2318 44540 2374 45000 0 FreeSans 224 90 0 0 N2BEG[4]
port 196 nsew signal tristate
flabel metal2 s 2594 44540 2650 45000 0 FreeSans 224 90 0 0 N2BEG[5]
port 197 nsew signal tristate
flabel metal2 s 2870 44540 2926 45000 0 FreeSans 224 90 0 0 N2BEG[6]
port 198 nsew signal tristate
flabel metal2 s 3146 44540 3202 45000 0 FreeSans 224 90 0 0 N2BEG[7]
port 199 nsew signal tristate
flabel metal2 s 3422 44540 3478 45000 0 FreeSans 224 90 0 0 N2BEGb[0]
port 200 nsew signal tristate
flabel metal2 s 3698 44540 3754 45000 0 FreeSans 224 90 0 0 N2BEGb[1]
port 201 nsew signal tristate
flabel metal2 s 3974 44540 4030 45000 0 FreeSans 224 90 0 0 N2BEGb[2]
port 202 nsew signal tristate
flabel metal2 s 4250 44540 4306 45000 0 FreeSans 224 90 0 0 N2BEGb[3]
port 203 nsew signal tristate
flabel metal2 s 4526 44540 4582 45000 0 FreeSans 224 90 0 0 N2BEGb[4]
port 204 nsew signal tristate
flabel metal2 s 4802 44540 4858 45000 0 FreeSans 224 90 0 0 N2BEGb[5]
port 205 nsew signal tristate
flabel metal2 s 5078 44540 5134 45000 0 FreeSans 224 90 0 0 N2BEGb[6]
port 206 nsew signal tristate
flabel metal2 s 5354 44540 5410 45000 0 FreeSans 224 90 0 0 N2BEGb[7]
port 207 nsew signal tristate
flabel metal2 s 3422 -300 3478 160 0 FreeSans 224 90 0 0 N2END[0]
port 208 nsew signal input
flabel metal2 s 3698 -300 3754 160 0 FreeSans 224 90 0 0 N2END[1]
port 209 nsew signal input
flabel metal2 s 3974 -300 4030 160 0 FreeSans 224 90 0 0 N2END[2]
port 210 nsew signal input
flabel metal2 s 4250 -300 4306 160 0 FreeSans 224 90 0 0 N2END[3]
port 211 nsew signal input
flabel metal2 s 4526 -300 4582 160 0 FreeSans 224 90 0 0 N2END[4]
port 212 nsew signal input
flabel metal2 s 4802 -300 4858 160 0 FreeSans 224 90 0 0 N2END[5]
port 213 nsew signal input
flabel metal2 s 5078 -300 5134 160 0 FreeSans 224 90 0 0 N2END[6]
port 214 nsew signal input
flabel metal2 s 5354 -300 5410 160 0 FreeSans 224 90 0 0 N2END[7]
port 215 nsew signal input
flabel metal2 s 1214 -300 1270 160 0 FreeSans 224 90 0 0 N2MID[0]
port 216 nsew signal input
flabel metal2 s 1490 -300 1546 160 0 FreeSans 224 90 0 0 N2MID[1]
port 217 nsew signal input
flabel metal2 s 1766 -300 1822 160 0 FreeSans 224 90 0 0 N2MID[2]
port 218 nsew signal input
flabel metal2 s 2042 -300 2098 160 0 FreeSans 224 90 0 0 N2MID[3]
port 219 nsew signal input
flabel metal2 s 2318 -300 2374 160 0 FreeSans 224 90 0 0 N2MID[4]
port 220 nsew signal input
flabel metal2 s 2594 -300 2650 160 0 FreeSans 224 90 0 0 N2MID[5]
port 221 nsew signal input
flabel metal2 s 2870 -300 2926 160 0 FreeSans 224 90 0 0 N2MID[6]
port 222 nsew signal input
flabel metal2 s 3146 -300 3202 160 0 FreeSans 224 90 0 0 N2MID[7]
port 223 nsew signal input
flabel metal2 s 5630 44540 5686 45000 0 FreeSans 224 90 0 0 N4BEG[0]
port 224 nsew signal tristate
flabel metal2 s 8390 44540 8446 45000 0 FreeSans 224 90 0 0 N4BEG[10]
port 225 nsew signal tristate
flabel metal2 s 8666 44540 8722 45000 0 FreeSans 224 90 0 0 N4BEG[11]
port 226 nsew signal tristate
flabel metal2 s 8942 44540 8998 45000 0 FreeSans 224 90 0 0 N4BEG[12]
port 227 nsew signal tristate
flabel metal2 s 9218 44540 9274 45000 0 FreeSans 224 90 0 0 N4BEG[13]
port 228 nsew signal tristate
flabel metal2 s 9494 44540 9550 45000 0 FreeSans 224 90 0 0 N4BEG[14]
port 229 nsew signal tristate
flabel metal2 s 9770 44540 9826 45000 0 FreeSans 224 90 0 0 N4BEG[15]
port 230 nsew signal tristate
flabel metal2 s 5906 44540 5962 45000 0 FreeSans 224 90 0 0 N4BEG[1]
port 231 nsew signal tristate
flabel metal2 s 6182 44540 6238 45000 0 FreeSans 224 90 0 0 N4BEG[2]
port 232 nsew signal tristate
flabel metal2 s 6458 44540 6514 45000 0 FreeSans 224 90 0 0 N4BEG[3]
port 233 nsew signal tristate
flabel metal2 s 6734 44540 6790 45000 0 FreeSans 224 90 0 0 N4BEG[4]
port 234 nsew signal tristate
flabel metal2 s 7010 44540 7066 45000 0 FreeSans 224 90 0 0 N4BEG[5]
port 235 nsew signal tristate
flabel metal2 s 7286 44540 7342 45000 0 FreeSans 224 90 0 0 N4BEG[6]
port 236 nsew signal tristate
flabel metal2 s 7562 44540 7618 45000 0 FreeSans 224 90 0 0 N4BEG[7]
port 237 nsew signal tristate
flabel metal2 s 7838 44540 7894 45000 0 FreeSans 224 90 0 0 N4BEG[8]
port 238 nsew signal tristate
flabel metal2 s 8114 44540 8170 45000 0 FreeSans 224 90 0 0 N4BEG[9]
port 239 nsew signal tristate
flabel metal2 s 5630 -300 5686 160 0 FreeSans 224 90 0 0 N4END[0]
port 240 nsew signal input
flabel metal2 s 8390 -300 8446 160 0 FreeSans 224 90 0 0 N4END[10]
port 241 nsew signal input
flabel metal2 s 8666 -300 8722 160 0 FreeSans 224 90 0 0 N4END[11]
port 242 nsew signal input
flabel metal2 s 8942 -300 8998 160 0 FreeSans 224 90 0 0 N4END[12]
port 243 nsew signal input
flabel metal2 s 9218 -300 9274 160 0 FreeSans 224 90 0 0 N4END[13]
port 244 nsew signal input
flabel metal2 s 9494 -300 9550 160 0 FreeSans 224 90 0 0 N4END[14]
port 245 nsew signal input
flabel metal2 s 9770 -300 9826 160 0 FreeSans 224 90 0 0 N4END[15]
port 246 nsew signal input
flabel metal2 s 5906 -300 5962 160 0 FreeSans 224 90 0 0 N4END[1]
port 247 nsew signal input
flabel metal2 s 6182 -300 6238 160 0 FreeSans 224 90 0 0 N4END[2]
port 248 nsew signal input
flabel metal2 s 6458 -300 6514 160 0 FreeSans 224 90 0 0 N4END[3]
port 249 nsew signal input
flabel metal2 s 6734 -300 6790 160 0 FreeSans 224 90 0 0 N4END[4]
port 250 nsew signal input
flabel metal2 s 7010 -300 7066 160 0 FreeSans 224 90 0 0 N4END[5]
port 251 nsew signal input
flabel metal2 s 7286 -300 7342 160 0 FreeSans 224 90 0 0 N4END[6]
port 252 nsew signal input
flabel metal2 s 7562 -300 7618 160 0 FreeSans 224 90 0 0 N4END[7]
port 253 nsew signal input
flabel metal2 s 7838 -300 7894 160 0 FreeSans 224 90 0 0 N4END[8]
port 254 nsew signal input
flabel metal2 s 8114 -300 8170 160 0 FreeSans 224 90 0 0 N4END[9]
port 255 nsew signal input
flabel metal3 s 25540 7080 26000 7200 0 FreeSans 480 0 0 0 RAM2FAB_D0_I0
port 256 nsew signal input
flabel metal3 s 25540 7624 26000 7744 0 FreeSans 480 0 0 0 RAM2FAB_D0_I1
port 257 nsew signal input
flabel metal3 s 25540 8168 26000 8288 0 FreeSans 480 0 0 0 RAM2FAB_D0_I2
port 258 nsew signal input
flabel metal3 s 25540 8712 26000 8832 0 FreeSans 480 0 0 0 RAM2FAB_D0_I3
port 259 nsew signal input
flabel metal3 s 25540 4904 26000 5024 0 FreeSans 480 0 0 0 RAM2FAB_D1_I0
port 260 nsew signal input
flabel metal3 s 25540 5448 26000 5568 0 FreeSans 480 0 0 0 RAM2FAB_D1_I1
port 261 nsew signal input
flabel metal3 s 25540 5992 26000 6112 0 FreeSans 480 0 0 0 RAM2FAB_D1_I2
port 262 nsew signal input
flabel metal3 s 25540 6536 26000 6656 0 FreeSans 480 0 0 0 RAM2FAB_D1_I3
port 263 nsew signal input
flabel metal3 s 25540 2728 26000 2848 0 FreeSans 480 0 0 0 RAM2FAB_D2_I0
port 264 nsew signal input
flabel metal3 s 25540 3272 26000 3392 0 FreeSans 480 0 0 0 RAM2FAB_D2_I1
port 265 nsew signal input
flabel metal3 s 25540 3816 26000 3936 0 FreeSans 480 0 0 0 RAM2FAB_D2_I2
port 266 nsew signal input
flabel metal3 s 25540 4360 26000 4480 0 FreeSans 480 0 0 0 RAM2FAB_D2_I3
port 267 nsew signal input
flabel metal3 s 25540 552 26000 672 0 FreeSans 480 0 0 0 RAM2FAB_D3_I0
port 268 nsew signal input
flabel metal3 s 25540 1096 26000 1216 0 FreeSans 480 0 0 0 RAM2FAB_D3_I1
port 269 nsew signal input
flabel metal3 s 25540 1640 26000 1760 0 FreeSans 480 0 0 0 RAM2FAB_D3_I2
port 270 nsew signal input
flabel metal3 s 25540 2184 26000 2304 0 FreeSans 480 0 0 0 RAM2FAB_D3_I3
port 271 nsew signal input
flabel metal2 s 10046 -300 10102 160 0 FreeSans 224 90 0 0 S1BEG[0]
port 272 nsew signal tristate
flabel metal2 s 10322 -300 10378 160 0 FreeSans 224 90 0 0 S1BEG[1]
port 273 nsew signal tristate
flabel metal2 s 10598 -300 10654 160 0 FreeSans 224 90 0 0 S1BEG[2]
port 274 nsew signal tristate
flabel metal2 s 10874 -300 10930 160 0 FreeSans 224 90 0 0 S1BEG[3]
port 275 nsew signal tristate
flabel metal2 s 10046 44540 10102 45000 0 FreeSans 224 90 0 0 S1END[0]
port 276 nsew signal input
flabel metal2 s 10322 44540 10378 45000 0 FreeSans 224 90 0 0 S1END[1]
port 277 nsew signal input
flabel metal2 s 10598 44540 10654 45000 0 FreeSans 224 90 0 0 S1END[2]
port 278 nsew signal input
flabel metal2 s 10874 44540 10930 45000 0 FreeSans 224 90 0 0 S1END[3]
port 279 nsew signal input
flabel metal2 s 13358 -300 13414 160 0 FreeSans 224 90 0 0 S2BEG[0]
port 280 nsew signal tristate
flabel metal2 s 13634 -300 13690 160 0 FreeSans 224 90 0 0 S2BEG[1]
port 281 nsew signal tristate
flabel metal2 s 13910 -300 13966 160 0 FreeSans 224 90 0 0 S2BEG[2]
port 282 nsew signal tristate
flabel metal2 s 14186 -300 14242 160 0 FreeSans 224 90 0 0 S2BEG[3]
port 283 nsew signal tristate
flabel metal2 s 14462 -300 14518 160 0 FreeSans 224 90 0 0 S2BEG[4]
port 284 nsew signal tristate
flabel metal2 s 14738 -300 14794 160 0 FreeSans 224 90 0 0 S2BEG[5]
port 285 nsew signal tristate
flabel metal2 s 15014 -300 15070 160 0 FreeSans 224 90 0 0 S2BEG[6]
port 286 nsew signal tristate
flabel metal2 s 15290 -300 15346 160 0 FreeSans 224 90 0 0 S2BEG[7]
port 287 nsew signal tristate
flabel metal2 s 11150 -300 11206 160 0 FreeSans 224 90 0 0 S2BEGb[0]
port 288 nsew signal tristate
flabel metal2 s 11426 -300 11482 160 0 FreeSans 224 90 0 0 S2BEGb[1]
port 289 nsew signal tristate
flabel metal2 s 11702 -300 11758 160 0 FreeSans 224 90 0 0 S2BEGb[2]
port 290 nsew signal tristate
flabel metal2 s 11978 -300 12034 160 0 FreeSans 224 90 0 0 S2BEGb[3]
port 291 nsew signal tristate
flabel metal2 s 12254 -300 12310 160 0 FreeSans 224 90 0 0 S2BEGb[4]
port 292 nsew signal tristate
flabel metal2 s 12530 -300 12586 160 0 FreeSans 224 90 0 0 S2BEGb[5]
port 293 nsew signal tristate
flabel metal2 s 12806 -300 12862 160 0 FreeSans 224 90 0 0 S2BEGb[6]
port 294 nsew signal tristate
flabel metal2 s 13082 -300 13138 160 0 FreeSans 224 90 0 0 S2BEGb[7]
port 295 nsew signal tristate
flabel metal2 s 11150 44540 11206 45000 0 FreeSans 224 90 0 0 S2END[0]
port 296 nsew signal input
flabel metal2 s 11426 44540 11482 45000 0 FreeSans 224 90 0 0 S2END[1]
port 297 nsew signal input
flabel metal2 s 11702 44540 11758 45000 0 FreeSans 224 90 0 0 S2END[2]
port 298 nsew signal input
flabel metal2 s 11978 44540 12034 45000 0 FreeSans 224 90 0 0 S2END[3]
port 299 nsew signal input
flabel metal2 s 12254 44540 12310 45000 0 FreeSans 224 90 0 0 S2END[4]
port 300 nsew signal input
flabel metal2 s 12530 44540 12586 45000 0 FreeSans 224 90 0 0 S2END[5]
port 301 nsew signal input
flabel metal2 s 12806 44540 12862 45000 0 FreeSans 224 90 0 0 S2END[6]
port 302 nsew signal input
flabel metal2 s 13082 44540 13138 45000 0 FreeSans 224 90 0 0 S2END[7]
port 303 nsew signal input
flabel metal2 s 13358 44540 13414 45000 0 FreeSans 224 90 0 0 S2MID[0]
port 304 nsew signal input
flabel metal2 s 13634 44540 13690 45000 0 FreeSans 224 90 0 0 S2MID[1]
port 305 nsew signal input
flabel metal2 s 13910 44540 13966 45000 0 FreeSans 224 90 0 0 S2MID[2]
port 306 nsew signal input
flabel metal2 s 14186 44540 14242 45000 0 FreeSans 224 90 0 0 S2MID[3]
port 307 nsew signal input
flabel metal2 s 14462 44540 14518 45000 0 FreeSans 224 90 0 0 S2MID[4]
port 308 nsew signal input
flabel metal2 s 14738 44540 14794 45000 0 FreeSans 224 90 0 0 S2MID[5]
port 309 nsew signal input
flabel metal2 s 15014 44540 15070 45000 0 FreeSans 224 90 0 0 S2MID[6]
port 310 nsew signal input
flabel metal2 s 15290 44540 15346 45000 0 FreeSans 224 90 0 0 S2MID[7]
port 311 nsew signal input
flabel metal2 s 15566 -300 15622 160 0 FreeSans 224 90 0 0 S4BEG[0]
port 312 nsew signal tristate
flabel metal2 s 18326 -300 18382 160 0 FreeSans 224 90 0 0 S4BEG[10]
port 313 nsew signal tristate
flabel metal2 s 18602 -300 18658 160 0 FreeSans 224 90 0 0 S4BEG[11]
port 314 nsew signal tristate
flabel metal2 s 18878 -300 18934 160 0 FreeSans 224 90 0 0 S4BEG[12]
port 315 nsew signal tristate
flabel metal2 s 19154 -300 19210 160 0 FreeSans 224 90 0 0 S4BEG[13]
port 316 nsew signal tristate
flabel metal2 s 19430 -300 19486 160 0 FreeSans 224 90 0 0 S4BEG[14]
port 317 nsew signal tristate
flabel metal2 s 19706 -300 19762 160 0 FreeSans 224 90 0 0 S4BEG[15]
port 318 nsew signal tristate
flabel metal2 s 15842 -300 15898 160 0 FreeSans 224 90 0 0 S4BEG[1]
port 319 nsew signal tristate
flabel metal2 s 16118 -300 16174 160 0 FreeSans 224 90 0 0 S4BEG[2]
port 320 nsew signal tristate
flabel metal2 s 16394 -300 16450 160 0 FreeSans 224 90 0 0 S4BEG[3]
port 321 nsew signal tristate
flabel metal2 s 16670 -300 16726 160 0 FreeSans 224 90 0 0 S4BEG[4]
port 322 nsew signal tristate
flabel metal2 s 16946 -300 17002 160 0 FreeSans 224 90 0 0 S4BEG[5]
port 323 nsew signal tristate
flabel metal2 s 17222 -300 17278 160 0 FreeSans 224 90 0 0 S4BEG[6]
port 324 nsew signal tristate
flabel metal2 s 17498 -300 17554 160 0 FreeSans 224 90 0 0 S4BEG[7]
port 325 nsew signal tristate
flabel metal2 s 17774 -300 17830 160 0 FreeSans 224 90 0 0 S4BEG[8]
port 326 nsew signal tristate
flabel metal2 s 18050 -300 18106 160 0 FreeSans 224 90 0 0 S4BEG[9]
port 327 nsew signal tristate
flabel metal2 s 15566 44540 15622 45000 0 FreeSans 224 90 0 0 S4END[0]
port 328 nsew signal input
flabel metal2 s 18326 44540 18382 45000 0 FreeSans 224 90 0 0 S4END[10]
port 329 nsew signal input
flabel metal2 s 18602 44540 18658 45000 0 FreeSans 224 90 0 0 S4END[11]
port 330 nsew signal input
flabel metal2 s 18878 44540 18934 45000 0 FreeSans 224 90 0 0 S4END[12]
port 331 nsew signal input
flabel metal2 s 19154 44540 19210 45000 0 FreeSans 224 90 0 0 S4END[13]
port 332 nsew signal input
flabel metal2 s 19430 44540 19486 45000 0 FreeSans 224 90 0 0 S4END[14]
port 333 nsew signal input
flabel metal2 s 19706 44540 19762 45000 0 FreeSans 224 90 0 0 S4END[15]
port 334 nsew signal input
flabel metal2 s 15842 44540 15898 45000 0 FreeSans 224 90 0 0 S4END[1]
port 335 nsew signal input
flabel metal2 s 16118 44540 16174 45000 0 FreeSans 224 90 0 0 S4END[2]
port 336 nsew signal input
flabel metal2 s 16394 44540 16450 45000 0 FreeSans 224 90 0 0 S4END[3]
port 337 nsew signal input
flabel metal2 s 16670 44540 16726 45000 0 FreeSans 224 90 0 0 S4END[4]
port 338 nsew signal input
flabel metal2 s 16946 44540 17002 45000 0 FreeSans 224 90 0 0 S4END[5]
port 339 nsew signal input
flabel metal2 s 17222 44540 17278 45000 0 FreeSans 224 90 0 0 S4END[6]
port 340 nsew signal input
flabel metal2 s 17498 44540 17554 45000 0 FreeSans 224 90 0 0 S4END[7]
port 341 nsew signal input
flabel metal2 s 17774 44540 17830 45000 0 FreeSans 224 90 0 0 S4END[8]
port 342 nsew signal input
flabel metal2 s 18050 44540 18106 45000 0 FreeSans 224 90 0 0 S4END[9]
port 343 nsew signal input
flabel metal2 s 19982 -300 20038 160 0 FreeSans 224 90 0 0 UserCLK
port 344 nsew signal input
flabel metal2 s 19982 44540 20038 45000 0 FreeSans 224 90 0 0 UserCLKo
port 345 nsew signal tristate
flabel metal4 s 6808 1040 7128 43568 0 FreeSans 1920 90 0 0 VGND
port 346 nsew ground bidirectional
flabel metal4 s 12673 1040 12993 43568 0 FreeSans 1920 90 0 0 VGND
port 346 nsew ground bidirectional
flabel metal4 s 18538 1040 18858 43568 0 FreeSans 1920 90 0 0 VGND
port 346 nsew ground bidirectional
flabel metal4 s 24403 1040 24723 43568 0 FreeSans 1920 90 0 0 VGND
port 346 nsew ground bidirectional
flabel metal4 s 3876 1040 4196 43568 0 FreeSans 1920 90 0 0 VPWR
port 347 nsew power bidirectional
flabel metal4 s 9741 1040 10061 43568 0 FreeSans 1920 90 0 0 VPWR
port 347 nsew power bidirectional
flabel metal4 s 15606 1040 15926 43568 0 FreeSans 1920 90 0 0 VPWR
port 347 nsew power bidirectional
flabel metal4 s 21471 1040 21791 43568 0 FreeSans 1920 90 0 0 VPWR
port 347 nsew power bidirectional
flabel metal3 s -300 4904 160 5024 0 FreeSans 480 0 0 0 W1BEG[0]
port 348 nsew signal tristate
flabel metal3 s -300 5176 160 5296 0 FreeSans 480 0 0 0 W1BEG[1]
port 349 nsew signal tristate
flabel metal3 s -300 5448 160 5568 0 FreeSans 480 0 0 0 W1BEG[2]
port 350 nsew signal tristate
flabel metal3 s -300 5720 160 5840 0 FreeSans 480 0 0 0 W1BEG[3]
port 351 nsew signal tristate
flabel metal3 s -300 5992 160 6112 0 FreeSans 480 0 0 0 W2BEG[0]
port 352 nsew signal tristate
flabel metal3 s -300 6264 160 6384 0 FreeSans 480 0 0 0 W2BEG[1]
port 353 nsew signal tristate
flabel metal3 s -300 6536 160 6656 0 FreeSans 480 0 0 0 W2BEG[2]
port 354 nsew signal tristate
flabel metal3 s -300 6808 160 6928 0 FreeSans 480 0 0 0 W2BEG[3]
port 355 nsew signal tristate
flabel metal3 s -300 7080 160 7200 0 FreeSans 480 0 0 0 W2BEG[4]
port 356 nsew signal tristate
flabel metal3 s -300 7352 160 7472 0 FreeSans 480 0 0 0 W2BEG[5]
port 357 nsew signal tristate
flabel metal3 s -300 7624 160 7744 0 FreeSans 480 0 0 0 W2BEG[6]
port 358 nsew signal tristate
flabel metal3 s -300 7896 160 8016 0 FreeSans 480 0 0 0 W2BEG[7]
port 359 nsew signal tristate
flabel metal3 s -300 8168 160 8288 0 FreeSans 480 0 0 0 W2BEGb[0]
port 360 nsew signal tristate
flabel metal3 s -300 8440 160 8560 0 FreeSans 480 0 0 0 W2BEGb[1]
port 361 nsew signal tristate
flabel metal3 s -300 8712 160 8832 0 FreeSans 480 0 0 0 W2BEGb[2]
port 362 nsew signal tristate
flabel metal3 s -300 8984 160 9104 0 FreeSans 480 0 0 0 W2BEGb[3]
port 363 nsew signal tristate
flabel metal3 s -300 9256 160 9376 0 FreeSans 480 0 0 0 W2BEGb[4]
port 364 nsew signal tristate
flabel metal3 s -300 9528 160 9648 0 FreeSans 480 0 0 0 W2BEGb[5]
port 365 nsew signal tristate
flabel metal3 s -300 9800 160 9920 0 FreeSans 480 0 0 0 W2BEGb[6]
port 366 nsew signal tristate
flabel metal3 s -300 10072 160 10192 0 FreeSans 480 0 0 0 W2BEGb[7]
port 367 nsew signal tristate
flabel metal3 s -300 14696 160 14816 0 FreeSans 480 0 0 0 W6BEG[0]
port 368 nsew signal tristate
flabel metal3 s -300 17416 160 17536 0 FreeSans 480 0 0 0 W6BEG[10]
port 369 nsew signal tristate
flabel metal3 s -300 17688 160 17808 0 FreeSans 480 0 0 0 W6BEG[11]
port 370 nsew signal tristate
flabel metal3 s -300 14968 160 15088 0 FreeSans 480 0 0 0 W6BEG[1]
port 371 nsew signal tristate
flabel metal3 s -300 15240 160 15360 0 FreeSans 480 0 0 0 W6BEG[2]
port 372 nsew signal tristate
flabel metal3 s -300 15512 160 15632 0 FreeSans 480 0 0 0 W6BEG[3]
port 373 nsew signal tristate
flabel metal3 s -300 15784 160 15904 0 FreeSans 480 0 0 0 W6BEG[4]
port 374 nsew signal tristate
flabel metal3 s -300 16056 160 16176 0 FreeSans 480 0 0 0 W6BEG[5]
port 375 nsew signal tristate
flabel metal3 s -300 16328 160 16448 0 FreeSans 480 0 0 0 W6BEG[6]
port 376 nsew signal tristate
flabel metal3 s -300 16600 160 16720 0 FreeSans 480 0 0 0 W6BEG[7]
port 377 nsew signal tristate
flabel metal3 s -300 16872 160 16992 0 FreeSans 480 0 0 0 W6BEG[8]
port 378 nsew signal tristate
flabel metal3 s -300 17144 160 17264 0 FreeSans 480 0 0 0 W6BEG[9]
port 379 nsew signal tristate
flabel metal3 s -300 10344 160 10464 0 FreeSans 480 0 0 0 WW4BEG[0]
port 380 nsew signal tristate
flabel metal3 s -300 13064 160 13184 0 FreeSans 480 0 0 0 WW4BEG[10]
port 381 nsew signal tristate
flabel metal3 s -300 13336 160 13456 0 FreeSans 480 0 0 0 WW4BEG[11]
port 382 nsew signal tristate
flabel metal3 s -300 13608 160 13728 0 FreeSans 480 0 0 0 WW4BEG[12]
port 383 nsew signal tristate
flabel metal3 s -300 13880 160 14000 0 FreeSans 480 0 0 0 WW4BEG[13]
port 384 nsew signal tristate
flabel metal3 s -300 14152 160 14272 0 FreeSans 480 0 0 0 WW4BEG[14]
port 385 nsew signal tristate
flabel metal3 s -300 14424 160 14544 0 FreeSans 480 0 0 0 WW4BEG[15]
port 386 nsew signal tristate
flabel metal3 s -300 10616 160 10736 0 FreeSans 480 0 0 0 WW4BEG[1]
port 387 nsew signal tristate
flabel metal3 s -300 10888 160 11008 0 FreeSans 480 0 0 0 WW4BEG[2]
port 388 nsew signal tristate
flabel metal3 s -300 11160 160 11280 0 FreeSans 480 0 0 0 WW4BEG[3]
port 389 nsew signal tristate
flabel metal3 s -300 11432 160 11552 0 FreeSans 480 0 0 0 WW4BEG[4]
port 390 nsew signal tristate
flabel metal3 s -300 11704 160 11824 0 FreeSans 480 0 0 0 WW4BEG[5]
port 391 nsew signal tristate
flabel metal3 s -300 11976 160 12096 0 FreeSans 480 0 0 0 WW4BEG[6]
port 392 nsew signal tristate
flabel metal3 s -300 12248 160 12368 0 FreeSans 480 0 0 0 WW4BEG[7]
port 393 nsew signal tristate
flabel metal3 s -300 12520 160 12640 0 FreeSans 480 0 0 0 WW4BEG[8]
port 394 nsew signal tristate
flabel metal3 s -300 12792 160 12912 0 FreeSans 480 0 0 0 WW4BEG[9]
port 395 nsew signal tristate
rlabel via1 12913 43520 12913 43520 0 VGND
rlabel metal1 12834 42976 12834 42976 0 VPWR
rlabel metal1 17480 6426 17480 6426 0 ConfigBits\[0\]
rlabel metal2 13478 19924 13478 19924 0 ConfigBits\[100\]
rlabel metal1 13524 20026 13524 20026 0 ConfigBits\[101\]
rlabel metal1 8188 17510 8188 17510 0 ConfigBits\[102\]
rlabel metal1 8970 16218 8970 16218 0 ConfigBits\[103\]
rlabel metal1 11730 27574 11730 27574 0 ConfigBits\[104\]
rlabel metal2 12098 28356 12098 28356 0 ConfigBits\[105\]
rlabel metal1 13524 18122 13524 18122 0 ConfigBits\[106\]
rlabel metal1 14858 17850 14858 17850 0 ConfigBits\[107\]
rlabel metal1 13984 22474 13984 22474 0 ConfigBits\[108\]
rlabel via1 15318 22073 15318 22073 0 ConfigBits\[109\]
rlabel metal1 20056 12750 20056 12750 0 ConfigBits\[10\]
rlabel metal1 18170 22032 18170 22032 0 ConfigBits\[110\]
rlabel metal1 6900 22066 6900 22066 0 ConfigBits\[111\]
rlabel metal1 8004 21658 8004 21658 0 ConfigBits\[112\]
rlabel metal1 9568 21318 9568 21318 0 ConfigBits\[113\]
rlabel metal2 8418 29546 8418 29546 0 ConfigBits\[114\]
rlabel metal2 8970 29308 8970 29308 0 ConfigBits\[115\]
rlabel metal1 10442 29104 10442 29104 0 ConfigBits\[116\]
rlabel metal2 17342 18258 17342 18258 0 ConfigBits\[117\]
rlabel metal2 17894 18768 17894 18768 0 ConfigBits\[118\]
rlabel metal2 19550 18938 19550 18938 0 ConfigBits\[119\]
rlabel metal2 20838 10540 20838 10540 0 ConfigBits\[11\]
rlabel metal1 7590 4046 7590 4046 0 ConfigBits\[120\]
rlabel metal2 8326 4420 8326 4420 0 ConfigBits\[121\]
rlabel metal1 5060 13498 5060 13498 0 ConfigBits\[122\]
rlabel metal2 5566 14620 5566 14620 0 ConfigBits\[123\]
rlabel metal1 4692 8058 4692 8058 0 ConfigBits\[124\]
rlabel metal2 5106 8636 5106 8636 0 ConfigBits\[125\]
rlabel metal1 13524 3706 13524 3706 0 ConfigBits\[126\]
rlabel metal1 14076 4250 14076 4250 0 ConfigBits\[127\]
rlabel metal1 5152 5338 5152 5338 0 ConfigBits\[128\]
rlabel metal2 5658 6188 5658 6188 0 ConfigBits\[129\]
rlabel metal1 17756 4114 17756 4114 0 ConfigBits\[12\]
rlabel metal1 3404 6222 3404 6222 0 ConfigBits\[130\]
rlabel metal1 4186 6222 4186 6222 0 ConfigBits\[131\]
rlabel metal2 3358 12546 3358 12546 0 ConfigBits\[132\]
rlabel metal1 4186 12750 4186 12750 0 ConfigBits\[133\]
rlabel metal1 6118 6426 6118 6426 0 ConfigBits\[134\]
rlabel metal2 7406 6358 7406 6358 0 ConfigBits\[135\]
rlabel metal1 15502 5338 15502 5338 0 ConfigBits\[136\]
rlabel metal1 15916 4794 15916 4794 0 ConfigBits\[137\]
rlabel metal1 2300 10234 2300 10234 0 ConfigBits\[138\]
rlabel metal2 2714 11492 2714 11492 0 ConfigBits\[139\]
rlabel metal2 23138 6596 23138 6596 0 ConfigBits\[13\]
rlabel metal1 2300 4726 2300 4726 0 ConfigBits\[140\]
rlabel metal1 2576 5338 2576 5338 0 ConfigBits\[141\]
rlabel metal1 3082 3706 3082 3706 0 ConfigBits\[142\]
rlabel metal1 3542 2550 3542 2550 0 ConfigBits\[143\]
rlabel metal1 5106 2074 5106 2074 0 ConfigBits\[144\]
rlabel metal2 5014 3706 5014 3706 0 ConfigBits\[145\]
rlabel metal1 2990 9146 2990 9146 0 ConfigBits\[146\]
rlabel metal1 3496 8058 3496 8058 0 ConfigBits\[147\]
rlabel metal1 2070 16694 2070 16694 0 ConfigBits\[148\]
rlabel metal2 2806 16388 2806 16388 0 ConfigBits\[149\]
rlabel metal1 21114 6256 21114 6256 0 ConfigBits\[14\]
rlabel metal1 6072 9078 6072 9078 0 ConfigBits\[150\]
rlabel metal1 7084 8602 7084 8602 0 ConfigBits\[151\]
rlabel metal2 15226 7106 15226 7106 0 ConfigBits\[152\]
rlabel metal2 15686 7548 15686 7548 0 ConfigBits\[153\]
rlabel metal1 2208 13838 2208 13838 0 ConfigBits\[154\]
rlabel metal1 2622 13498 2622 13498 0 ConfigBits\[155\]
rlabel metal1 2300 6426 2300 6426 0 ConfigBits\[156\]
rlabel metal1 2622 7514 2622 7514 0 ConfigBits\[157\]
rlabel metal1 4140 2278 4140 2278 0 ConfigBits\[158\]
rlabel metal1 3864 2074 3864 2074 0 ConfigBits\[159\]
rlabel metal2 21114 3740 21114 3740 0 ConfigBits\[15\]
rlabel metal1 16284 8262 16284 8262 0 ConfigBits\[160\]
rlabel metal1 17296 8602 17296 8602 0 ConfigBits\[161\]
rlabel metal1 2392 18870 2392 18870 0 ConfigBits\[162\]
rlabel metal2 2898 18564 2898 18564 0 ConfigBits\[163\]
rlabel metal1 2300 21658 2300 21658 0 ConfigBits\[164\]
rlabel metal1 2576 22406 2576 22406 0 ConfigBits\[165\]
rlabel metal2 8326 5508 8326 5508 0 ConfigBits\[166\]
rlabel metal2 8878 5644 8878 5644 0 ConfigBits\[167\]
rlabel metal1 14720 10098 14720 10098 0 ConfigBits\[168\]
rlabel metal1 15226 9690 15226 9690 0 ConfigBits\[169\]
rlabel metal2 23690 25534 23690 25534 0 ConfigBits\[16\]
rlabel metal2 5750 10982 5750 10982 0 ConfigBits\[170\]
rlabel metal1 6394 11186 6394 11186 0 ConfigBits\[171\]
rlabel metal1 3772 16014 3772 16014 0 ConfigBits\[172\]
rlabel metal2 4462 16524 4462 16524 0 ConfigBits\[173\]
rlabel metal1 8372 7310 8372 7310 0 ConfigBits\[174\]
rlabel metal2 8970 7820 8970 7820 0 ConfigBits\[175\]
rlabel metal1 16284 10778 16284 10778 0 ConfigBits\[176\]
rlabel metal1 17296 10778 17296 10778 0 ConfigBits\[177\]
rlabel metal1 2898 10778 2898 10778 0 ConfigBits\[178\]
rlabel metal1 4600 10778 4600 10778 0 ConfigBits\[179\]
rlabel metal1 22586 30566 22586 30566 0 ConfigBits\[17\]
rlabel metal2 5566 16218 5566 16218 0 ConfigBits\[180\]
rlabel metal1 5704 16626 5704 16626 0 ConfigBits\[181\]
rlabel metal2 8510 9690 8510 9690 0 ConfigBits\[182\]
rlabel metal2 8326 9894 8326 9894 0 ConfigBits\[183\]
rlabel metal1 16192 13430 16192 13430 0 ConfigBits\[184\]
rlabel metal1 17204 13362 17204 13362 0 ConfigBits\[185\]
rlabel metal2 4278 18666 4278 18666 0 ConfigBits\[186\]
rlabel metal2 4830 18428 4830 18428 0 ConfigBits\[187\]
rlabel metal2 4416 21692 4416 21692 0 ConfigBits\[188\]
rlabel metal2 5014 21692 5014 21692 0 ConfigBits\[189\]
rlabel metal1 22908 27846 22908 27846 0 ConfigBits\[18\]
rlabel metal1 6164 3162 6164 3162 0 ConfigBits\[190\]
rlabel metal1 7130 2618 7130 2618 0 ConfigBits\[191\]
rlabel metal2 11086 10982 11086 10982 0 ConfigBits\[192\]
rlabel metal2 11638 10948 11638 10948 0 ConfigBits\[193\]
rlabel metal2 5750 34918 5750 34918 0 ConfigBits\[194\]
rlabel metal1 5796 35054 5796 35054 0 ConfigBits\[195\]
rlabel metal1 4324 26010 4324 26010 0 ConfigBits\[196\]
rlabel metal2 5014 26554 5014 26554 0 ConfigBits\[197\]
rlabel metal1 12662 12274 12662 12274 0 ConfigBits\[198\]
rlabel metal1 13386 11866 13386 11866 0 ConfigBits\[199\]
rlabel metal1 18584 28050 18584 28050 0 ConfigBits\[19\]
rlabel metal1 18124 9350 18124 9350 0 ConfigBits\[1\]
rlabel metal2 14950 12070 14950 12070 0 ConfigBits\[200\]
rlabel metal2 14766 12410 14766 12410 0 ConfigBits\[201\]
rlabel metal1 6210 13430 6210 13430 0 ConfigBits\[202\]
rlabel metal1 7222 13362 7222 13362 0 ConfigBits\[203\]
rlabel metal1 6854 16728 6854 16728 0 ConfigBits\[204\]
rlabel metal1 7544 16218 7544 16218 0 ConfigBits\[205\]
rlabel metal2 8510 11458 8510 11458 0 ConfigBits\[206\]
rlabel metal1 9522 11322 9522 11322 0 ConfigBits\[207\]
rlabel metal1 15042 14586 15042 14586 0 ConfigBits\[208\]
rlabel metal2 15502 15164 15502 15164 0 ConfigBits\[209\]
rlabel metal1 22034 22712 22034 22712 0 ConfigBits\[20\]
rlabel metal1 5980 18870 5980 18870 0 ConfigBits\[210\]
rlabel metal2 6808 19686 6808 19686 0 ConfigBits\[211\]
rlabel metal2 5796 21522 5796 21522 0 ConfigBits\[212\]
rlabel metal1 6670 20978 6670 20978 0 ConfigBits\[213\]
rlabel metal1 7820 12954 7820 12954 0 ConfigBits\[214\]
rlabel metal2 8326 14076 8326 14076 0 ConfigBits\[215\]
rlabel metal2 12558 25568 12558 25568 0 ConfigBits\[216\]
rlabel metal1 12926 25330 12926 25330 0 ConfigBits\[217\]
rlabel metal2 5934 32028 5934 32028 0 ConfigBits\[218\]
rlabel metal1 7038 31858 7038 31858 0 ConfigBits\[219\]
rlabel metal1 23552 22950 23552 22950 0 ConfigBits\[21\]
rlabel metal1 6033 27982 6033 27982 0 ConfigBits\[220\]
rlabel metal1 5980 27574 5980 27574 0 ConfigBits\[221\]
rlabel metal1 15364 27982 15364 27982 0 ConfigBits\[222\]
rlabel metal2 16514 27812 16514 27812 0 ConfigBits\[223\]
rlabel metal1 14766 25432 14766 25432 0 ConfigBits\[224\]
rlabel metal1 15410 25330 15410 25330 0 ConfigBits\[225\]
rlabel metal2 5934 25194 5934 25194 0 ConfigBits\[226\]
rlabel metal1 7084 24786 7084 24786 0 ConfigBits\[227\]
rlabel metal1 7176 26554 7176 26554 0 ConfigBits\[228\]
rlabel metal1 7728 27030 7728 27030 0 ConfigBits\[229\]
rlabel metal1 21620 25874 21620 25874 0 ConfigBits\[22\]
rlabel metal1 16928 25466 16928 25466 0 ConfigBits\[230\]
rlabel metal1 17480 26010 17480 26010 0 ConfigBits\[231\]
rlabel metal1 12558 23834 12558 23834 0 ConfigBits\[232\]
rlabel metal1 13110 24242 13110 24242 0 ConfigBits\[233\]
rlabel metal2 6762 34476 6762 34476 0 ConfigBits\[234\]
rlabel metal1 7314 33966 7314 33966 0 ConfigBits\[235\]
rlabel metal1 5934 29716 5934 29716 0 ConfigBits\[236\]
rlabel metal1 7360 29274 7360 29274 0 ConfigBits\[237\]
rlabel metal2 15962 31246 15962 31246 0 ConfigBits\[238\]
rlabel metal2 17342 31212 17342 31212 0 ConfigBits\[239\]
rlabel metal1 19918 26758 19918 26758 0 ConfigBits\[23\]
rlabel metal1 13800 24650 13800 24650 0 ConfigBits\[240\]
rlabel metal2 14858 25228 14858 25228 0 ConfigBits\[241\]
rlabel metal2 7406 23902 7406 23902 0 ConfigBits\[242\]
rlabel metal1 8326 24174 8326 24174 0 ConfigBits\[243\]
rlabel metal1 8740 26486 8740 26486 0 ConfigBits\[244\]
rlabel metal2 9522 26520 9522 26520 0 ConfigBits\[245\]
rlabel metal1 16790 23562 16790 23562 0 ConfigBits\[246\]
rlabel metal1 17526 23290 17526 23290 0 ConfigBits\[247\]
rlabel metal1 15364 16762 15364 16762 0 ConfigBits\[248\]
rlabel metal1 16100 16218 16100 16218 0 ConfigBits\[249\]
rlabel metal1 18906 24378 18906 24378 0 ConfigBits\[24\]
rlabel metal1 11684 17714 11684 17714 0 ConfigBits\[250\]
rlabel metal1 12512 17306 12512 17306 0 ConfigBits\[251\]
rlabel via1 9706 19125 9706 19125 0 ConfigBits\[252\]
rlabel metal1 10074 18394 10074 18394 0 ConfigBits\[253\]
rlabel metal1 15364 19958 15364 19958 0 ConfigBits\[254\]
rlabel metal1 15916 19482 15916 19482 0 ConfigBits\[255\]
rlabel metal2 13110 16218 13110 16218 0 ConfigBits\[256\]
rlabel metal2 13662 15878 13662 15878 0 ConfigBits\[257\]
rlabel metal1 8648 14858 8648 14858 0 ConfigBits\[258\]
rlabel metal1 10074 14586 10074 14586 0 ConfigBits\[259\]
rlabel metal1 22310 32878 22310 32878 0 ConfigBits\[25\]
rlabel metal1 10534 19958 10534 19958 0 ConfigBits\[260\]
rlabel metal1 11592 18938 11592 18938 0 ConfigBits\[261\]
rlabel metal1 16514 21046 16514 21046 0 ConfigBits\[262\]
rlabel metal1 17526 20978 17526 20978 0 ConfigBits\[263\]
rlabel metal1 12005 13838 12005 13838 0 ConfigBits\[264\]
rlabel metal1 12374 13498 12374 13498 0 ConfigBits\[265\]
rlabel metal2 7774 41219 7774 41219 0 ConfigBits\[266\]
rlabel metal1 8234 41174 8234 41174 0 ConfigBits\[267\]
rlabel metal1 12006 35598 12006 35598 0 ConfigBits\[268\]
rlabel metal2 12742 35428 12742 35428 0 ConfigBits\[269\]
rlabel metal1 20424 29138 20424 29138 0 ConfigBits\[26\]
rlabel metal2 17342 29308 17342 29308 0 ConfigBits\[270\]
rlabel metal2 17894 29308 17894 29308 0 ConfigBits\[271\]
rlabel metal1 8786 3162 8786 3162 0 ConfigBits\[272\]
rlabel metal1 9752 3162 9752 3162 0 ConfigBits\[273\]
rlabel metal2 5014 39644 5014 39644 0 ConfigBits\[274\]
rlabel metal1 5566 39066 5566 39066 0 ConfigBits\[275\]
rlabel metal1 3588 28662 3588 28662 0 ConfigBits\[276\]
rlabel metal2 4462 28730 4462 28730 0 ConfigBits\[277\]
rlabel metal2 13110 14042 13110 14042 0 ConfigBits\[278\]
rlabel metal1 13846 13498 13846 13498 0 ConfigBits\[279\]
rlabel metal1 19044 30702 19044 30702 0 ConfigBits\[27\]
rlabel metal1 9752 9894 9752 9894 0 ConfigBits\[280\]
rlabel metal1 10488 9146 10488 9146 0 ConfigBits\[281\]
rlabel metal2 5382 37553 5382 37553 0 ConfigBits\[282\]
rlabel metal1 5658 36890 5658 36890 0 ConfigBits\[283\]
rlabel metal2 3358 31450 3358 31450 0 ConfigBits\[284\]
rlabel metal1 4324 31994 4324 31994 0 ConfigBits\[285\]
rlabel metal2 12466 9622 12466 9622 0 ConfigBits\[286\]
rlabel metal1 12972 9690 12972 9690 0 ConfigBits\[287\]
rlabel metal1 10120 7718 10120 7718 0 ConfigBits\[288\]
rlabel metal1 10580 6970 10580 6970 0 ConfigBits\[289\]
rlabel metal1 20608 24174 20608 24174 0 ConfigBits\[28\]
rlabel metal2 5106 42092 5106 42092 0 ConfigBits\[290\]
rlabel metal1 5836 41582 5836 41582 0 ConfigBits\[291\]
rlabel metal1 4232 34374 4232 34374 0 ConfigBits\[292\]
rlabel metal1 5106 33626 5106 33626 0 ConfigBits\[293\]
rlabel metal1 13616 6970 13616 6970 0 ConfigBits\[294\]
rlabel metal2 14214 7072 14214 7072 0 ConfigBits\[295\]
rlabel metal1 10212 4794 10212 4794 0 ConfigBits\[296\]
rlabel metal2 10166 5372 10166 5372 0 ConfigBits\[297\]
rlabel metal1 4186 40970 4186 40970 0 ConfigBits\[298\]
rlabel metal1 5060 41174 5060 41174 0 ConfigBits\[299\]
rlabel metal1 23966 19856 23966 19856 0 ConfigBits\[29\]
rlabel metal1 22402 7990 22402 7990 0 ConfigBits\[2\]
rlabel metal1 3588 36278 3588 36278 0 ConfigBits\[300\]
rlabel metal1 4462 36142 4462 36142 0 ConfigBits\[301\]
rlabel metal1 11960 7718 11960 7718 0 ConfigBits\[302\]
rlabel metal1 12190 6970 12190 6970 0 ConfigBits\[303\]
rlabel metal1 10810 1530 10810 1530 0 ConfigBits\[304\]
rlabel metal1 10948 2074 10948 2074 0 ConfigBits\[305\]
rlabel metal2 10258 38692 10258 38692 0 ConfigBits\[306\]
rlabel metal1 10258 38998 10258 38998 0 ConfigBits\[307\]
rlabel metal1 4968 30362 4968 30362 0 ConfigBits\[308\]
rlabel metal1 5474 30702 5474 30702 0 ConfigBits\[309\]
rlabel metal1 21919 19958 21919 19958 0 ConfigBits\[30\]
rlabel metal1 11316 33354 11316 33354 0 ConfigBits\[310\]
rlabel metal1 12190 33558 12190 33558 0 ConfigBits\[311\]
rlabel metal2 11914 4182 11914 4182 0 ConfigBits\[312\]
rlabel metal2 12558 4420 12558 4420 0 ConfigBits\[313\]
rlabel metal2 7958 19686 7958 19686 0 ConfigBits\[314\]
rlabel metal1 8188 19822 8188 19822 0 ConfigBits\[315\]
rlabel metal2 11086 29852 11086 29852 0 ConfigBits\[316\]
rlabel metal1 11316 29614 11316 29614 0 ConfigBits\[317\]
rlabel metal2 12374 2652 12374 2652 0 ConfigBits\[318\]
rlabel metal1 12972 2074 12972 2074 0 ConfigBits\[319\]
rlabel metal1 19964 21862 19964 21862 0 ConfigBits\[31\]
rlabel metal2 9982 12954 9982 12954 0 ConfigBits\[320\]
rlabel metal1 10028 12818 10028 12818 0 ConfigBits\[321\]
rlabel metal2 2530 42636 2530 42636 0 ConfigBits\[322\]
rlabel metal1 3220 41786 3220 41786 0 ConfigBits\[323\]
rlabel metal2 3358 37434 3358 37434 0 ConfigBits\[324\]
rlabel metal2 3450 36686 3450 36686 0 ConfigBits\[325\]
rlabel metal1 13524 28730 13524 28730 0 ConfigBits\[326\]
rlabel metal1 14168 28186 14168 28186 0 ConfigBits\[327\]
rlabel metal1 19182 16218 19182 16218 0 ConfigBits\[32\]
rlabel metal1 21758 16524 21758 16524 0 ConfigBits\[33\]
rlabel metal1 23736 16762 23736 16762 0 ConfigBits\[34\]
rlabel metal1 23092 18598 23092 18598 0 ConfigBits\[35\]
rlabel metal2 18722 14790 18722 14790 0 ConfigBits\[36\]
rlabel metal1 23966 14008 23966 14008 0 ConfigBits\[37\]
rlabel metal2 20654 14790 20654 14790 0 ConfigBits\[38\]
rlabel metal2 21022 16762 21022 16762 0 ConfigBits\[39\]
rlabel metal1 19872 9486 19872 9486 0 ConfigBits\[3\]
rlabel metal1 22402 12818 22402 12818 0 ConfigBits\[40\]
rlabel metal1 20056 31450 20056 31450 0 ConfigBits\[41\]
rlabel metal1 20884 34578 20884 34578 0 ConfigBits\[42\]
rlabel metal1 20562 18700 20562 18700 0 ConfigBits\[43\]
rlabel metal1 23874 9044 23874 9044 0 ConfigBits\[44\]
rlabel metal1 22724 10030 22724 10030 0 ConfigBits\[45\]
rlabel metal1 22494 10064 22494 10064 0 ConfigBits\[46\]
rlabel metal1 24058 10642 24058 10642 0 ConfigBits\[47\]
rlabel metal2 10810 22236 10810 22236 0 ConfigBits\[48\]
rlabel metal1 10856 21658 10856 21658 0 ConfigBits\[49\]
rlabel metal2 18078 12517 18078 12517 0 ConfigBits\[4\]
rlabel metal1 2300 38794 2300 38794 0 ConfigBits\[50\]
rlabel metal1 2668 40154 2668 40154 0 ConfigBits\[51\]
rlabel metal1 2392 35190 2392 35190 0 ConfigBits\[52\]
rlabel metal2 2852 34714 2852 34714 0 ConfigBits\[53\]
rlabel metal2 15318 33473 15318 33473 0 ConfigBits\[54\]
rlabel metal1 16790 33082 16790 33082 0 ConfigBits\[55\]
rlabel metal1 3128 26486 3128 26486 0 ConfigBits\[56\]
rlabel metal1 3266 23290 3266 23290 0 ConfigBits\[57\]
rlabel metal1 2254 36890 2254 36890 0 ConfigBits\[58\]
rlabel metal2 2622 37468 2622 37468 0 ConfigBits\[59\]
rlabel metal2 21390 12517 21390 12517 0 ConfigBits\[5\]
rlabel metal1 2116 32334 2116 32334 0 ConfigBits\[60\]
rlabel metal2 2622 32572 2622 32572 0 ConfigBits\[61\]
rlabel metal1 2208 30158 2208 30158 0 ConfigBits\[62\]
rlabel metal2 2898 29988 2898 29988 0 ConfigBits\[63\]
rlabel metal1 4876 24310 4876 24310 0 ConfigBits\[64\]
rlabel metal2 5474 23834 5474 23834 0 ConfigBits\[65\]
rlabel metal2 2438 25500 2438 25500 0 ConfigBits\[66\]
rlabel metal1 2346 24922 2346 24922 0 ConfigBits\[67\]
rlabel metal1 2254 27098 2254 27098 0 ConfigBits\[68\]
rlabel metal2 2622 27812 2622 27812 0 ConfigBits\[69\]
rlabel metal2 20838 7004 20838 7004 0 ConfigBits\[6\]
rlabel metal2 2714 20502 2714 20502 0 ConfigBits\[70\]
rlabel metal2 2622 20706 2622 20706 0 ConfigBits\[71\]
rlabel metal2 9798 23902 9798 23902 0 ConfigBits\[72\]
rlabel metal1 10350 24208 10350 24208 0 ConfigBits\[73\]
rlabel metal1 10626 26316 10626 26316 0 ConfigBits\[74\]
rlabel metal2 7406 39338 7406 39338 0 ConfigBits\[75\]
rlabel metal2 7958 39100 7958 39100 0 ConfigBits\[76\]
rlabel metal1 9384 39406 9384 39406 0 ConfigBits\[77\]
rlabel metal1 8188 32334 8188 32334 0 ConfigBits\[78\]
rlabel metal2 8786 32844 8786 32844 0 ConfigBits\[79\]
rlabel metal2 19458 5984 19458 5984 0 ConfigBits\[7\]
rlabel metal2 10350 34374 10350 34374 0 ConfigBits\[80\]
rlabel metal1 14168 33082 14168 33082 0 ConfigBits\[81\]
rlabel via2 14398 32844 14398 32844 0 ConfigBits\[82\]
rlabel metal1 14536 35802 14536 35802 0 ConfigBits\[83\]
rlabel metal2 10212 16014 10212 16014 0 ConfigBits\[84\]
rlabel metal1 10810 16014 10810 16014 0 ConfigBits\[85\]
rlabel metal2 7958 36890 7958 36890 0 ConfigBits\[86\]
rlabel metal2 8418 36312 8418 36312 0 ConfigBits\[87\]
rlabel metal2 8510 35802 8510 35802 0 ConfigBits\[88\]
rlabel metal1 9568 35734 9568 35734 0 ConfigBits\[89\]
rlabel metal2 19274 3332 19274 3332 0 ConfigBits\[8\]
rlabel metal2 13846 30634 13846 30634 0 ConfigBits\[90\]
rlabel metal2 14490 30702 14490 30702 0 ConfigBits\[91\]
rlabel metal2 12466 21590 12466 21590 0 ConfigBits\[92\]
rlabel metal2 12374 21794 12374 21794 0 ConfigBits\[93\]
rlabel metal2 10994 37094 10994 37094 0 ConfigBits\[94\]
rlabel metal1 11822 37230 11822 37230 0 ConfigBits\[95\]
rlabel metal2 8878 31892 8878 31892 0 ConfigBits\[96\]
rlabel metal2 9522 31586 9522 31586 0 ConfigBits\[97\]
rlabel metal1 13018 30090 13018 30090 0 ConfigBits\[98\]
rlabel metal1 13294 31654 13294 31654 0 ConfigBits\[99\]
rlabel metal1 21482 5236 21482 5236 0 ConfigBits\[9\]
rlabel metal2 24150 9231 24150 9231 0 Config_accessC_bit0
rlabel metal3 25262 9860 25262 9860 0 Config_accessC_bit1
rlabel metal1 24104 9894 24104 9894 0 Config_accessC_bit2
rlabel metal1 24518 10234 24518 10234 0 Config_accessC_bit3
rlabel via2 3634 18037 3634 18037 0 E1END[0]
rlabel metal2 2806 17969 2806 17969 0 E1END[1]
rlabel metal2 3818 17561 3818 17561 0 E1END[2]
rlabel metal2 2806 19091 2806 19091 0 E1END[3]
rlabel metal3 636 21284 636 21284 0 E2END[0]
rlabel metal3 452 21556 452 21556 0 E2END[1]
rlabel metal3 544 21828 544 21828 0 E2END[2]
rlabel metal3 1050 22100 1050 22100 0 E2END[3]
rlabel metal3 728 22372 728 22372 0 E2END[4]
rlabel metal3 498 22644 498 22644 0 E2END[5]
rlabel metal3 452 22916 452 22916 0 E2END[6]
rlabel metal3 544 23188 544 23188 0 E2END[7]
rlabel metal3 452 19108 452 19108 0 E2MID[0]
rlabel metal3 636 19380 636 19380 0 E2MID[1]
rlabel metal3 728 19652 728 19652 0 E2MID[2]
rlabel metal3 774 19924 774 19924 0 E2MID[3]
rlabel metal3 452 20196 452 20196 0 E2MID[4]
rlabel metal3 544 20468 544 20468 0 E2MID[5]
rlabel metal3 820 20740 820 20740 0 E2MID[6]
rlabel metal3 728 21012 728 21012 0 E2MID[7]
rlabel metal3 728 27812 728 27812 0 E6END[0]
rlabel metal1 3680 32402 3680 32402 0 E6END[10]
rlabel metal3 1096 30804 1096 30804 0 E6END[11]
rlabel metal3 452 28084 452 28084 0 E6END[1]
rlabel metal3 475 28356 475 28356 0 E6END[2]
rlabel metal2 2806 29665 2806 29665 0 E6END[3]
rlabel metal3 1280 28900 1280 28900 0 E6END[4]
rlabel metal3 728 29172 728 29172 0 E6END[5]
rlabel metal3 728 29444 728 29444 0 E6END[6]
rlabel metal3 452 29716 452 29716 0 E6END[7]
rlabel metal3 728 29988 728 29988 0 E6END[8]
rlabel metal3 1602 30260 1602 30260 0 E6END[9]
rlabel metal3 452 23460 452 23460 0 EE4END[0]
rlabel metal2 2898 26571 2898 26571 0 EE4END[10]
rlabel metal3 728 26452 728 26452 0 EE4END[11]
rlabel metal3 682 26724 682 26724 0 EE4END[12]
rlabel metal3 728 26996 728 26996 0 EE4END[13]
rlabel metal3 498 27268 498 27268 0 EE4END[14]
rlabel metal2 3726 27795 3726 27795 0 EE4END[15]
rlabel metal3 498 23732 498 23732 0 EE4END[1]
rlabel metal3 728 24004 728 24004 0 EE4END[2]
rlabel metal3 452 24276 452 24276 0 EE4END[3]
rlabel metal3 682 24548 682 24548 0 EE4END[4]
rlabel metal3 728 24820 728 24820 0 EE4END[5]
rlabel metal3 475 25092 475 25092 0 EE4END[6]
rlabel metal3 498 25364 498 25364 0 EE4END[7]
rlabel metal3 728 25636 728 25636 0 EE4END[8]
rlabel metal2 2806 26435 2806 26435 0 EE4END[9]
rlabel metal1 16872 16558 16872 16558 0 FAB2RAM_A0_I0
rlabel metal1 19166 17578 19166 17578 0 FAB2RAM_A0_I1
rlabel metal2 20838 17952 20838 17952 0 FAB2RAM_A0_I2
rlabel metal1 19274 19720 19274 19720 0 FAB2RAM_A0_I3
rlabel metal3 24710 15844 24710 15844 0 FAB2RAM_A0_O0
rlabel metal1 24518 16218 24518 16218 0 FAB2RAM_A0_O1
rlabel metal3 24618 16932 24618 16932 0 FAB2RAM_A0_O2
rlabel metal3 25262 17476 25262 17476 0 FAB2RAM_A0_O3
rlabel metal1 16918 14994 16918 14994 0 FAB2RAM_A1_I0
rlabel metal1 17250 15096 17250 15096 0 FAB2RAM_A1_I1
rlabel metal1 19918 15470 19918 15470 0 FAB2RAM_A1_I2
rlabel metal1 18768 17646 18768 17646 0 FAB2RAM_A1_I3
rlabel metal2 24150 13583 24150 13583 0 FAB2RAM_A1_O0
rlabel metal3 25262 14212 25262 14212 0 FAB2RAM_A1_O1
rlabel metal3 24894 14756 24894 14756 0 FAB2RAM_A1_O2
rlabel metal3 25262 15300 25262 15300 0 FAB2RAM_A1_O3
rlabel metal1 21574 13872 21574 13872 0 FAB2RAM_C_I0
rlabel metal1 19080 32402 19080 32402 0 FAB2RAM_C_I1
rlabel metal2 17342 35258 17342 35258 0 FAB2RAM_C_I2
rlabel metal1 19310 19822 19310 19822 0 FAB2RAM_C_I3
rlabel metal3 24848 11492 24848 11492 0 FAB2RAM_C_O0
rlabel metal3 25262 12036 25262 12036 0 FAB2RAM_C_O1
rlabel metal3 24802 12580 24802 12580 0 FAB2RAM_C_O2
rlabel metal1 24150 12954 24150 12954 0 FAB2RAM_C_O3
rlabel metal1 14030 25466 14030 25466 0 FAB2RAM_D0_I0
rlabel metal1 13478 33014 13478 33014 0 FAB2RAM_D0_I1
rlabel metal1 21666 28084 21666 28084 0 FAB2RAM_D0_I2
rlabel metal1 17204 28050 17204 28050 0 FAB2RAM_D0_I3
rlabel metal1 23828 24378 23828 24378 0 FAB2RAM_D0_O0
rlabel metal3 25262 25092 25262 25092 0 FAB2RAM_D0_O1
rlabel metal3 24710 25636 24710 25636 0 FAB2RAM_D0_O2
rlabel metal3 25262 26180 25262 26180 0 FAB2RAM_D0_O3
rlabel metal1 19366 23086 19366 23086 0 FAB2RAM_D1_I0
rlabel via2 7866 24667 7866 24667 0 FAB2RAM_D1_I1
rlabel metal1 20930 26996 20930 26996 0 FAB2RAM_D1_I2
rlabel via1 18446 26350 18446 26350 0 FAB2RAM_D1_I3
rlabel metal3 24710 22372 24710 22372 0 FAB2RAM_D1_O0
rlabel metal1 24518 22406 24518 22406 0 FAB2RAM_D1_O1
rlabel metal3 24894 23460 24894 23460 0 FAB2RAM_D1_O2
rlabel metal3 25262 24004 25262 24004 0 FAB2RAM_D1_O3
rlabel metal1 15594 24174 15594 24174 0 FAB2RAM_D2_I0
rlabel metal1 21298 33490 21298 33490 0 FAB2RAM_D2_I1
rlabel metal1 19734 29580 19734 29580 0 FAB2RAM_D2_I2
rlabel metal1 17710 31790 17710 31790 0 FAB2RAM_D2_I3
rlabel metal2 23782 20111 23782 20111 0 FAB2RAM_D2_O0
rlabel metal3 25262 20740 25262 20740 0 FAB2RAM_D2_O1
rlabel metal3 24894 21284 24894 21284 0 FAB2RAM_D2_O2
rlabel metal1 24518 21862 24518 21862 0 FAB2RAM_D2_O3
rlabel via1 19550 24786 19550 24786 0 FAB2RAM_D3_I0
rlabel metal2 22034 21182 22034 21182 0 FAB2RAM_D3_I1
rlabel metal1 20132 20842 20132 20842 0 FAB2RAM_D3_I2
rlabel metal1 18676 21998 18676 21998 0 FAB2RAM_D3_I3
rlabel metal3 24618 18020 24618 18020 0 FAB2RAM_D3_O0
rlabel metal1 24518 17850 24518 17850 0 FAB2RAM_D3_O1
rlabel metal3 24802 19108 24802 19108 0 FAB2RAM_D3_O2
rlabel metal1 24656 18394 24656 18394 0 FAB2RAM_D3_O3
rlabel metal3 820 31076 820 31076 0 FrameData[0]
rlabel metal3 728 33796 728 33796 0 FrameData[10]
rlabel metal3 774 34068 774 34068 0 FrameData[11]
rlabel metal3 1441 34340 1441 34340 0 FrameData[12]
rlabel metal2 3910 34833 3910 34833 0 FrameData[13]
rlabel metal2 2806 35819 2806 35819 0 FrameData[14]
rlabel metal2 3082 35955 3082 35955 0 FrameData[15]
rlabel metal2 3634 36091 3634 36091 0 FrameData[16]
rlabel metal2 3266 36465 3266 36465 0 FrameData[17]
rlabel metal3 2752 35972 2752 35972 0 FrameData[18]
rlabel metal2 2898 36584 2898 36584 0 FrameData[19]
rlabel metal3 728 31348 728 31348 0 FrameData[1]
rlabel metal2 1748 42194 1748 42194 0 FrameData[20]
rlabel metal3 774 36788 774 36788 0 FrameData[21]
rlabel metal2 3082 37995 3082 37995 0 FrameData[22]
rlabel metal3 866 37332 866 37332 0 FrameData[23]
rlabel metal3 1441 37604 1441 37604 0 FrameData[24]
rlabel metal3 2568 37876 2568 37876 0 FrameData[25]
rlabel metal3 452 38148 452 38148 0 FrameData[26]
rlabel metal2 2806 38675 2806 38675 0 FrameData[27]
rlabel via2 3726 38709 3726 38709 0 FrameData[28]
rlabel metal1 2254 41548 2254 41548 0 FrameData[29]
rlabel metal3 2752 31620 2752 31620 0 FrameData[2]
rlabel metal3 774 39236 774 39236 0 FrameData[30]
rlabel metal2 2990 39797 2990 39797 0 FrameData[31]
rlabel metal3 728 31892 728 31892 0 FrameData[3]
rlabel metal3 843 32164 843 32164 0 FrameData[4]
rlabel metal3 774 32436 774 32436 0 FrameData[5]
rlabel metal3 1648 32708 1648 32708 0 FrameData[6]
rlabel metal3 567 32980 567 32980 0 FrameData[7]
rlabel metal3 728 33252 728 33252 0 FrameData[8]
rlabel metal3 636 33524 636 33524 0 FrameData[9]
rlabel metal3 24894 26724 24894 26724 0 FrameData_O[0]
rlabel metal3 24894 32164 24894 32164 0 FrameData_O[10]
rlabel metal3 25262 32708 25262 32708 0 FrameData_O[11]
rlabel metal3 24894 33252 24894 33252 0 FrameData_O[12]
rlabel metal3 25262 33796 25262 33796 0 FrameData_O[13]
rlabel metal3 25193 34340 25193 34340 0 FrameData_O[14]
rlabel metal3 25262 34884 25262 34884 0 FrameData_O[15]
rlabel metal3 24894 35428 24894 35428 0 FrameData_O[16]
rlabel metal3 25308 35972 25308 35972 0 FrameData_O[17]
rlabel metal3 24894 36516 24894 36516 0 FrameData_O[18]
rlabel metal3 25262 37060 25262 37060 0 FrameData_O[19]
rlabel metal3 25262 27268 25262 27268 0 FrameData_O[1]
rlabel metal3 24894 37604 24894 37604 0 FrameData_O[20]
rlabel metal3 25262 38148 25262 38148 0 FrameData_O[21]
rlabel metal3 24894 38692 24894 38692 0 FrameData_O[22]
rlabel metal3 25262 39236 25262 39236 0 FrameData_O[23]
rlabel metal3 24894 39780 24894 39780 0 FrameData_O[24]
rlabel metal3 25308 40324 25308 40324 0 FrameData_O[25]
rlabel metal3 24664 40868 24664 40868 0 FrameData_O[26]
rlabel metal3 24173 41548 24173 41548 0 FrameData_O[27]
rlabel metal3 24894 41956 24894 41956 0 FrameData_O[28]
rlabel metal1 24426 42330 24426 42330 0 FrameData_O[29]
rlabel metal3 24894 27812 24894 27812 0 FrameData_O[2]
rlabel metal1 22908 42330 22908 42330 0 FrameData_O[30]
rlabel metal2 22126 43146 22126 43146 0 FrameData_O[31]
rlabel metal3 25262 28356 25262 28356 0 FrameData_O[3]
rlabel metal3 24894 28900 24894 28900 0 FrameData_O[4]
rlabel metal3 25262 29444 25262 29444 0 FrameData_O[5]
rlabel metal3 24894 29988 24894 29988 0 FrameData_O[6]
rlabel metal3 25262 30532 25262 30532 0 FrameData_O[7]
rlabel metal3 24894 31076 24894 31076 0 FrameData_O[8]
rlabel metal1 24656 31790 24656 31790 0 FrameData_O[9]
rlabel metal1 23690 26962 23690 26962 0 FrameData_O_i\[0\]
rlabel metal1 23414 32436 23414 32436 0 FrameData_O_i\[10\]
rlabel metal1 23690 32878 23690 32878 0 FrameData_O_i\[11\]
rlabel metal1 23644 33490 23644 33490 0 FrameData_O_i\[12\]
rlabel metal1 23552 33626 23552 33626 0 FrameData_O_i\[13\]
rlabel metal1 23368 34578 23368 34578 0 FrameData_O_i\[14\]
rlabel metal1 23046 35258 23046 35258 0 FrameData_O_i\[15\]
rlabel metal2 22586 35734 22586 35734 0 FrameData_O_i\[16\]
rlabel metal1 23000 35802 23000 35802 0 FrameData_O_i\[17\]
rlabel metal1 21482 36108 21482 36108 0 FrameData_O_i\[18\]
rlabel metal1 21482 36618 21482 36618 0 FrameData_O_i\[19\]
rlabel metal1 23736 27438 23736 27438 0 FrameData_O_i\[1\]
rlabel metal1 20608 36890 20608 36890 0 FrameData_O_i\[20\]
rlabel metal2 23414 37604 23414 37604 0 FrameData_O_i\[21\]
rlabel metal2 22862 38148 22862 38148 0 FrameData_O_i\[22\]
rlabel metal1 20148 38522 20148 38522 0 FrameData_O_i\[23\]
rlabel metal1 19090 38522 19090 38522 0 FrameData_O_i\[24\]
rlabel metal2 22586 39236 22586 39236 0 FrameData_O_i\[25\]
rlabel metal1 22218 40052 22218 40052 0 FrameData_O_i\[26\]
rlabel metal2 21022 40018 21022 40018 0 FrameData_O_i\[27\]
rlabel metal1 18860 40698 18860 40698 0 FrameData_O_i\[28\]
rlabel metal1 23368 39406 23368 39406 0 FrameData_O_i\[29\]
rlabel metal1 23184 27438 23184 27438 0 FrameData_O_i\[2\]
rlabel metal1 21896 41582 21896 41582 0 FrameData_O_i\[30\]
rlabel metal1 21344 41582 21344 41582 0 FrameData_O_i\[31\]
rlabel metal1 23184 28526 23184 28526 0 FrameData_O_i\[3\]
rlabel metal2 23506 29444 23506 29444 0 FrameData_O_i\[4\]
rlabel metal1 23414 29818 23414 29818 0 FrameData_O_i\[5\]
rlabel metal1 23276 30226 23276 30226 0 FrameData_O_i\[6\]
rlabel metal1 23322 30362 23322 30362 0 FrameData_O_i\[7\]
rlabel metal1 23460 30906 23460 30906 0 FrameData_O_i\[8\]
rlabel metal1 23046 31858 23046 31858 0 FrameData_O_i\[9\]
rlabel metal2 20339 68 20339 68 0 FrameStrobe[0]
rlabel metal2 23046 1282 23046 1282 0 FrameStrobe[10]
rlabel metal1 23460 4114 23460 4114 0 FrameStrobe[11]
rlabel metal1 21482 4216 21482 4216 0 FrameStrobe[12]
rlabel metal2 23973 68 23973 68 0 FrameStrobe[13]
rlabel metal2 24150 1214 24150 1214 0 FrameStrobe[14]
rlabel metal2 24426 347 24426 347 0 FrameStrobe[15]
rlabel metal2 24755 68 24755 68 0 FrameStrobe[16]
rlabel metal2 24925 68 24925 68 0 FrameStrobe[17]
rlabel metal1 22862 2992 22862 2992 0 FrameStrobe[18]
rlabel metal1 24794 4522 24794 4522 0 FrameStrobe[19]
rlabel metal2 20615 68 20615 68 0 FrameStrobe[1]
rlabel metal1 20286 2414 20286 2414 0 FrameStrobe[2]
rlabel metal2 21167 68 21167 68 0 FrameStrobe[3]
rlabel metal2 21489 68 21489 68 0 FrameStrobe[4]
rlabel metal2 21765 68 21765 68 0 FrameStrobe[5]
rlabel metal1 21390 1326 21390 1326 0 FrameStrobe[6]
rlabel metal2 22218 636 22218 636 0 FrameStrobe[7]
rlabel metal1 22494 850 22494 850 0 FrameStrobe[8]
rlabel metal2 22770 1180 22770 1180 0 FrameStrobe[9]
rlabel metal1 20332 43418 20332 43418 0 FrameStrobe_O[0]
rlabel metal1 22126 42602 22126 42602 0 FrameStrobe_O[10]
rlabel metal1 22908 41718 22908 41718 0 FrameStrobe_O[11]
rlabel metal2 23598 43972 23598 43972 0 FrameStrobe_O[12]
rlabel metal2 23874 43802 23874 43802 0 FrameStrobe_O[13]
rlabel metal1 23782 42262 23782 42262 0 FrameStrobe_O[14]
rlabel metal1 23966 41718 23966 41718 0 FrameStrobe_O[15]
rlabel metal2 24748 43724 24748 43724 0 FrameStrobe_O[16]
rlabel metal1 24058 41582 24058 41582 0 FrameStrobe_O[17]
rlabel metal1 24702 40698 24702 40698 0 FrameStrobe_O[18]
rlabel metal1 25530 43384 25530 43384 0 FrameStrobe_O[19]
rlabel metal2 20562 43972 20562 43972 0 FrameStrobe_O[1]
rlabel metal1 21436 43146 21436 43146 0 FrameStrobe_O[2]
rlabel metal1 21344 42330 21344 42330 0 FrameStrobe_O[3]
rlabel metal2 21390 43972 21390 43972 0 FrameStrobe_O[4]
rlabel metal2 21666 43802 21666 43802 0 FrameStrobe_O[5]
rlabel metal2 21942 43938 21942 43938 0 FrameStrobe_O[6]
rlabel metal2 22218 43530 22218 43530 0 FrameStrobe_O[7]
rlabel metal2 22494 44057 22494 44057 0 FrameStrobe_O[8]
rlabel metal1 22540 42330 22540 42330 0 FrameStrobe_O[9]
rlabel metal1 20194 41786 20194 41786 0 FrameStrobe_O_i\[0\]
rlabel metal2 22540 17340 22540 17340 0 FrameStrobe_O_i\[10\]
rlabel metal2 21390 40358 21390 40358 0 FrameStrobe_O_i\[11\]
rlabel metal1 23414 40052 23414 40052 0 FrameStrobe_O_i\[12\]
rlabel metal1 20930 41480 20930 41480 0 FrameStrobe_O_i\[13\]
rlabel metal2 21298 40460 21298 40460 0 FrameStrobe_O_i\[14\]
rlabel metal1 23506 39610 23506 39610 0 FrameStrobe_O_i\[15\]
rlabel metal1 23644 35258 23644 35258 0 FrameStrobe_O_i\[16\]
rlabel metal2 23690 36278 23690 36278 0 FrameStrobe_O_i\[17\]
rlabel metal1 23460 31994 23460 31994 0 FrameStrobe_O_i\[18\]
rlabel metal1 23644 37434 23644 37434 0 FrameStrobe_O_i\[19\]
rlabel metal1 20884 41582 20884 41582 0 FrameStrobe_O_i\[1\]
rlabel metal1 23874 43214 23874 43214 0 FrameStrobe_O_i\[2\]
rlabel metal1 21022 41106 21022 41106 0 FrameStrobe_O_i\[3\]
rlabel metal1 21758 40698 21758 40698 0 FrameStrobe_O_i\[4\]
rlabel metal2 21390 21913 21390 21913 0 FrameStrobe_O_i\[5\]
rlabel metal1 21758 34170 21758 34170 0 FrameStrobe_O_i\[6\]
rlabel metal2 21114 39814 21114 39814 0 FrameStrobe_O_i\[7\]
rlabel metal1 22356 40698 22356 40698 0 FrameStrobe_O_i\[8\]
rlabel via1 21574 41429 21574 41429 0 FrameStrobe_O_i\[9\]
rlabel metal1 19228 16558 19228 16558 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux/Q\[0\]
rlabel metal1 21942 17170 21942 17170 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux/Q\[1\]
rlabel metal1 23046 17204 23046 17204 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux/Q\[2\]
rlabel metal1 23368 19346 23368 19346 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux/Q\[3\]
rlabel metal1 17434 16184 17434 16184 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux/cus_mux21_inst0/AIN\[0\]
rlabel metal1 19734 16524 19734 16524 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux/cus_mux21_inst0/AIN\[1\]
rlabel metal1 18814 16694 18814 16694 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux/cus_mux21_inst0/_0_
rlabel metal1 18998 16626 18998 16626 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux/cus_mux21_inst0/_1_
rlabel metal2 22126 17306 22126 17306 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux/cus_mux21_inst1/AIN\[0\]
rlabel viali 22577 16558 22577 16558 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux/cus_mux21_inst1/AIN\[1\]
rlabel metal1 22034 16762 22034 16762 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux/cus_mux21_inst1/_0_
rlabel metal1 22264 16626 22264 16626 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux/cus_mux21_inst1/_1_
rlabel metal1 22448 17170 22448 17170 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux/cus_mux21_inst2/AIN\[0\]
rlabel metal1 24242 16524 24242 16524 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux/cus_mux21_inst2/AIN\[1\]
rlabel metal1 23322 17034 23322 17034 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux/cus_mux21_inst2/_0_
rlabel metal1 24104 17102 24104 17102 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux/cus_mux21_inst2/_1_
rlabel metal1 22954 18292 22954 18292 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux/cus_mux21_inst3/AIN\[0\]
rlabel metal2 22862 18700 22862 18700 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux/cus_mux21_inst3/AIN\[1\]
rlabel metal1 23506 18394 23506 18394 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux/cus_mux21_inst3/_0_
rlabel metal1 22678 18394 22678 18394 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux/cus_mux21_inst3/_1_
rlabel metal1 18584 13906 18584 13906 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux/Q\[0\]
rlabel metal1 22770 14416 22770 14416 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux/Q\[1\]
rlabel metal1 21022 14994 21022 14994 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux/Q\[2\]
rlabel metal1 20838 16558 20838 16558 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux/Q\[3\]
rlabel metal1 18078 13974 18078 13974 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux/cus_mux21_inst0/AIN\[0\]
rlabel metal1 18768 14042 18768 14042 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux/cus_mux21_inst0/AIN\[1\]
rlabel metal2 18170 14178 18170 14178 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux/cus_mux21_inst0/_0_
rlabel metal1 19182 14450 19182 14450 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux/cus_mux21_inst0/_1_
rlabel metal1 22719 13896 22719 13896 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux/cus_mux21_inst1/AIN\[0\]
rlabel metal1 22540 14382 22540 14382 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux/cus_mux21_inst1/AIN\[1\]
rlabel metal1 23322 14042 23322 14042 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux/cus_mux21_inst1/_0_
rlabel metal1 24058 14484 24058 14484 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux/cus_mux21_inst1/_1_
rlabel viali 21018 14382 21018 14382 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux/cus_mux21_inst2/AIN\[0\]
rlabel metal1 21482 14450 21482 14450 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux/cus_mux21_inst2/AIN\[1\]
rlabel metal2 21114 14722 21114 14722 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux/cus_mux21_inst2/_0_
rlabel metal1 21160 14926 21160 14926 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux/cus_mux21_inst2/_1_
rlabel metal1 20010 16592 20010 16592 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux/cus_mux21_inst3/AIN\[0\]
rlabel metal1 21206 16524 21206 16524 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux/cus_mux21_inst3/AIN\[1\]
rlabel metal1 20286 16626 20286 16626 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux/cus_mux21_inst3/_0_
rlabel metal1 20884 16626 20884 16626 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux/cus_mux21_inst3/_1_
rlabel metal1 22402 13498 22402 13498 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux/Q\[0\]
rlabel metal1 21252 31790 21252 31790 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux/Q\[1\]
rlabel metal2 20286 34884 20286 34884 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux/Q\[2\]
rlabel metal1 20516 20026 20516 20026 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux/Q\[3\]
rlabel metal1 21712 12818 21712 12818 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux/cus_mux21_inst0/AIN\[0\]
rlabel metal2 22310 13974 22310 13974 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux/cus_mux21_inst0/AIN\[1\]
rlabel metal1 22356 12614 22356 12614 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux/cus_mux21_inst0/_0_
rlabel metal1 22494 12750 22494 12750 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux/cus_mux21_inst0/_1_
rlabel metal1 19918 31824 19918 31824 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux/cus_mux21_inst1/AIN\[0\]
rlabel metal1 21068 31790 21068 31790 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux/cus_mux21_inst1/AIN\[1\]
rlabel metal1 20378 31824 20378 31824 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux/cus_mux21_inst1/_0_
rlabel metal1 20746 31824 20746 31824 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux/cus_mux21_inst1/_1_
rlabel metal1 20010 35122 20010 35122 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux/cus_mux21_inst2/AIN\[0\]
rlabel metal1 21206 34646 21206 34646 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux/cus_mux21_inst2/AIN\[1\]
rlabel metal1 20332 34578 20332 34578 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux/cus_mux21_inst2/_0_
rlabel metal1 21022 34646 21022 34646 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux/cus_mux21_inst2/_1_
rlabel metal2 18906 20230 18906 20230 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux/cus_mux21_inst3/AIN\[0\]
rlabel metal1 20746 18802 20746 18802 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux/cus_mux21_inst3/AIN\[1\]
rlabel metal1 20056 18938 20056 18938 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux/cus_mux21_inst3/_0_
rlabel metal1 20562 18802 20562 18802 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux/cus_mux21_inst3/_1_
rlabel metal1 23874 24786 23874 24786 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux/Q\[0\]
rlabel metal2 23230 30906 23230 30906 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux/Q\[1\]
rlabel metal1 22402 27438 22402 27438 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux/Q\[2\]
rlabel metal1 18860 28526 18860 28526 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux/Q\[3\]
rlabel metal1 24058 25228 24058 25228 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux/cus_mux21_inst0/AIN\[0\]
rlabel metal2 24058 25432 24058 25432 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux/cus_mux21_inst0/AIN\[1\]
rlabel metal1 23966 25398 23966 25398 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux/cus_mux21_inst0/_0_
rlabel metal1 23690 25330 23690 25330 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux/cus_mux21_inst0/_1_
rlabel metal1 21482 30226 21482 30226 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux/cus_mux21_inst1/AIN\[0\]
rlabel metal1 23000 30702 23000 30702 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux/cus_mux21_inst1/AIN\[1\]
rlabel metal1 22126 30022 22126 30022 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux/cus_mux21_inst1/_0_
rlabel metal1 22545 30169 22545 30169 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux/cus_mux21_inst1/_1_
rlabel metal2 22126 28356 22126 28356 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux/cus_mux21_inst2/AIN\[0\]
rlabel metal1 22862 27472 22862 27472 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux/cus_mux21_inst2/AIN\[1\]
rlabel metal1 23506 28084 23506 28084 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux/cus_mux21_inst2/_0_
rlabel metal1 22770 27608 22770 27608 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux/cus_mux21_inst2/_1_
rlabel metal1 18262 28084 18262 28084 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux/cus_mux21_inst3/AIN\[0\]
rlabel metal1 19044 28050 19044 28050 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux/cus_mux21_inst3/AIN\[1\]
rlabel metal1 18492 27846 18492 27846 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux/cus_mux21_inst3/_0_
rlabel metal1 18906 27982 18906 27982 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux/cus_mux21_inst3/_1_
rlabel metal1 22034 22576 22034 22576 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux/Q\[0\]
rlabel metal1 23552 23698 23552 23698 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux/Q\[1\]
rlabel metal1 21804 26350 21804 26350 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux/Q\[2\]
rlabel metal1 19918 25874 19918 25874 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux/Q\[3\]
rlabel metal1 21068 23290 21068 23290 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux/cus_mux21_inst0/AIN\[0\]
rlabel metal1 22678 22542 22678 22542 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux/cus_mux21_inst0/AIN\[1\]
rlabel metal2 21942 23052 21942 23052 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux/cus_mux21_inst0/_0_
rlabel metal1 22356 22542 22356 22542 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux/cus_mux21_inst0/_1_
rlabel metal2 23230 23324 23230 23324 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux/cus_mux21_inst1/AIN\[0\]
rlabel metal1 23138 22644 23138 22644 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux/cus_mux21_inst1/AIN\[1\]
rlabel metal1 23414 22610 23414 22610 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux/cus_mux21_inst1/_0_
rlabel metal2 23138 22882 23138 22882 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux/cus_mux21_inst1/_1_
rlabel metal1 21022 25262 21022 25262 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux/cus_mux21_inst2/AIN\[0\]
rlabel metal2 22402 26180 22402 26180 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux/cus_mux21_inst2/AIN\[1\]
rlabel metal1 21666 25466 21666 25466 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux/cus_mux21_inst2/_0_
rlabel metal1 22218 25806 22218 25806 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux/cus_mux21_inst2/_1_
rlabel metal1 19458 26316 19458 26316 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux/cus_mux21_inst3/AIN\[0\]
rlabel metal1 20240 26010 20240 26010 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux/cus_mux21_inst3/AIN\[1\]
rlabel metal1 19734 26418 19734 26418 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux/cus_mux21_inst3/_0_
rlabel metal1 20148 26418 20148 26418 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux/cus_mux21_inst3/_1_
rlabel metal1 18952 24786 18952 24786 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux/Q\[0\]
rlabel metal1 22586 33558 22586 33558 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux/Q\[1\]
rlabel metal2 20378 29444 20378 29444 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux/Q\[2\]
rlabel metal1 18814 31450 18814 31450 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux/Q\[3\]
rlabel metal1 17848 24378 17848 24378 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux/cus_mux21_inst0/AIN\[0\]
rlabel metal1 19320 24786 19320 24786 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux/cus_mux21_inst0/AIN\[1\]
rlabel metal1 18768 23698 18768 23698 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux/cus_mux21_inst0/_0_
rlabel metal1 19090 23630 19090 23630 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux/cus_mux21_inst0/_1_
rlabel metal1 21850 33388 21850 33388 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux/cus_mux21_inst1/AIN\[0\]
rlabel metal2 23046 33082 23046 33082 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux/cus_mux21_inst1/AIN\[1\]
rlabel metal1 22402 33082 22402 33082 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux/cus_mux21_inst1/_0_
rlabel metal1 22862 32946 22862 32946 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux/cus_mux21_inst1/_1_
rlabel metal1 20838 29171 20838 29171 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux/cus_mux21_inst2/AIN\[0\]
rlabel metal1 21298 29172 21298 29172 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux/cus_mux21_inst2/AIN\[1\]
rlabel metal1 20562 29172 20562 29172 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux/cus_mux21_inst2/_0_
rlabel metal1 20746 29036 20746 29036 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux/cus_mux21_inst2/_1_
rlabel metal1 18354 31858 18354 31858 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux/cus_mux21_inst3/AIN\[0\]
rlabel metal1 19550 31994 19550 31994 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux/cus_mux21_inst3/AIN\[1\]
rlabel metal3 19090 31756 19090 31756 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux/cus_mux21_inst3/_0_
rlabel metal1 19642 30770 19642 30770 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux/cus_mux21_inst3/_1_
rlabel metal1 21574 24140 21574 24140 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux/Q\[0\]
rlabel metal1 23736 21114 23736 21114 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux/Q\[1\]
rlabel metal1 21758 20434 21758 20434 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux/Q\[2\]
rlabel metal1 19688 22610 19688 22610 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux/Q\[3\]
rlabel metal1 20102 24752 20102 24752 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux/cus_mux21_inst0/AIN\[0\]
rlabel metal1 21344 24174 21344 24174 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux/cus_mux21_inst0/AIN\[1\]
rlabel metal1 20516 24378 20516 24378 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux/cus_mux21_inst0/_0_
rlabel metal1 21114 24242 21114 24242 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux/cus_mux21_inst0/_1_
rlabel metal1 23414 21556 23414 21556 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux/cus_mux21_inst1/AIN\[0\]
rlabel metal1 23368 19822 23368 19822 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux/cus_mux21_inst1/AIN\[1\]
rlabel metal2 24058 20672 24058 20672 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux/cus_mux21_inst1/_0_
rlabel metal1 24242 19924 24242 19924 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux/cus_mux21_inst1/_1_
rlabel metal1 21206 20468 21206 20468 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux/cus_mux21_inst2/AIN\[0\]
rlabel metal1 22310 20502 22310 20502 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux/cus_mux21_inst2/AIN\[1\]
rlabel metal1 21390 19788 21390 19788 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux/cus_mux21_inst2/_0_
rlabel metal1 22356 19890 22356 19890 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux/cus_mux21_inst2/_1_
rlabel metal1 18768 21862 18768 21862 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux/cus_mux21_inst3/AIN\[0\]
rlabel metal2 20884 21964 20884 21964 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux/cus_mux21_inst3/AIN\[1\]
rlabel metal1 19734 21556 19734 21556 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux/cus_mux21_inst3/_0_
rlabel metal1 20332 21454 20332 21454 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux/cus_mux21_inst3/_1_
rlabel metal1 18630 6732 18630 6732 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux/Q\[0\]
rlabel metal1 19136 8466 19136 8466 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux/Q\[1\]
rlabel metal1 23828 8466 23828 8466 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux/Q\[2\]
rlabel metal1 20516 8466 20516 8466 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux/Q\[3\]
rlabel metal1 16560 6766 16560 6766 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux/cus_mux21_inst0/AIN\[0\]
rlabel metal1 18262 6358 18262 6358 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux/cus_mux21_inst0/AIN\[1\]
rlabel metal1 16744 6970 16744 6970 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux/cus_mux21_inst0/_0_
rlabel metal2 18170 6902 18170 6902 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux/cus_mux21_inst0/_1_
rlabel metal1 18078 8398 18078 8398 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux/cus_mux21_inst1/AIN\[0\]
rlabel metal1 18538 8432 18538 8432 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux/cus_mux21_inst1/AIN\[1\]
rlabel metal1 18216 8602 18216 8602 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux/cus_mux21_inst1/_0_
rlabel metal1 18400 8602 18400 8602 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux/cus_mux21_inst1/_1_
rlabel metal1 22540 8058 22540 8058 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux/cus_mux21_inst2/AIN\[0\]
rlabel metal1 23322 7888 23322 7888 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux/cus_mux21_inst2/AIN\[1\]
rlabel metal2 22126 8704 22126 8704 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux/cus_mux21_inst2/_0_
rlabel metal2 23046 8500 23046 8500 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux/cus_mux21_inst2/_1_
rlabel metal1 19688 8466 19688 8466 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux/cus_mux21_inst3/AIN\[0\]
rlabel metal1 20102 8602 20102 8602 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux/cus_mux21_inst3/AIN\[1\]
rlabel metal2 19642 9078 19642 9078 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux/cus_mux21_inst3/_0_
rlabel metal1 20792 9554 20792 9554 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux/cus_mux21_inst3/_1_
rlabel metal1 18952 11730 18952 11730 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux/Q\[0\]
rlabel metal1 22494 11322 22494 11322 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux/Q\[1\]
rlabel metal1 22264 5882 22264 5882 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux/Q\[2\]
rlabel metal1 20562 6256 20562 6256 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux/Q\[3\]
rlabel metal1 17710 11118 17710 11118 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux/cus_mux21_inst0/AIN\[0\]
rlabel metal1 18906 11628 18906 11628 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux/cus_mux21_inst0/AIN\[1\]
rlabel metal2 18078 11764 18078 11764 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux/cus_mux21_inst0/_0_
rlabel metal1 18446 12138 18446 12138 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux/cus_mux21_inst0/_1_
rlabel metal1 22126 10574 22126 10574 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux/cus_mux21_inst1/AIN\[0\]
rlabel metal1 22034 11695 22034 11695 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux/cus_mux21_inst1/AIN\[1\]
rlabel metal1 21896 10778 21896 10778 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux/cus_mux21_inst1/_0_
rlabel metal2 22126 12036 22126 12036 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux/cus_mux21_inst1/_1_
rlabel metal1 20792 6290 20792 6290 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux/cus_mux21_inst2/AIN\[0\]
rlabel metal1 22034 6698 22034 6698 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux/cus_mux21_inst2/AIN\[1\]
rlabel metal2 21022 6596 21022 6596 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux/cus_mux21_inst2/_0_
rlabel metal1 21574 6800 21574 6800 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux/cus_mux21_inst2/_1_
rlabel metal1 18814 6426 18814 6426 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux/cus_mux21_inst3/AIN\[0\]
rlabel metal1 20332 6290 20332 6290 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux/cus_mux21_inst3/AIN\[1\]
rlabel metal2 19642 6154 19642 6154 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux/cus_mux21_inst3/_0_
rlabel metal2 20194 5882 20194 5882 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux/cus_mux21_inst3/_1_
rlabel metal1 20378 2074 20378 2074 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux/Q\[0\]
rlabel metal1 19550 4556 19550 4556 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux/Q\[1\]
rlabel metal1 20700 11730 20700 11730 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux/Q\[2\]
rlabel metal2 22034 9350 22034 9350 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux/Q\[3\]
rlabel metal2 22126 1768 22126 1768 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux/cus_mux21_inst0/AIN\[0\]
rlabel metal1 17066 3026 17066 3026 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux/cus_mux21_inst0/AIN\[1\]
rlabel metal1 19412 1326 19412 1326 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux/cus_mux21_inst0/_0_
rlabel metal2 16974 3298 16974 3298 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux/cus_mux21_inst0/_1_
rlabel metal1 20194 4624 20194 4624 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux/cus_mux21_inst1/AIN\[0\]
rlabel metal1 19780 4794 19780 4794 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux/cus_mux21_inst1/AIN\[1\]
rlabel metal1 21114 4794 21114 4794 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux/cus_mux21_inst1/_0_
rlabel metal1 22678 5270 22678 5270 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux/cus_mux21_inst1/_1_
rlabel metal1 19228 11322 19228 11322 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux/cus_mux21_inst2/AIN\[0\]
rlabel metal1 20746 11866 20746 11866 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux/cus_mux21_inst2/AIN\[1\]
rlabel metal2 19642 12614 19642 12614 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux/cus_mux21_inst2/_0_
rlabel metal1 20378 12886 20378 12886 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux/cus_mux21_inst2/_1_
rlabel metal1 21022 8602 21022 8602 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux/cus_mux21_inst3/AIN\[0\]
rlabel metal1 21758 9554 21758 9554 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux/cus_mux21_inst3/AIN\[1\]
rlabel metal1 21114 9690 21114 9690 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux/cus_mux21_inst3/_0_
rlabel metal2 21574 9826 21574 9826 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux/cus_mux21_inst3/_1_
rlabel metal1 18722 2516 18722 2516 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux/Q\[0\]
rlabel metal1 24104 5882 24104 5882 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux/Q\[1\]
rlabel metal2 20194 1598 20194 1598 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux/Q\[2\]
rlabel metal1 20470 2006 20470 2006 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux/Q\[3\]
rlabel metal1 17526 3162 17526 3162 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux/cus_mux21_inst0/AIN\[0\]
rlabel metal1 19458 2890 19458 2890 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux/cus_mux21_inst0/AIN\[1\]
rlabel metal1 17848 3706 17848 3706 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux/cus_mux21_inst0/_0_
rlabel metal1 17894 3638 17894 3638 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux/cus_mux21_inst0/_1_
rlabel metal1 23552 6290 23552 6290 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux/cus_mux21_inst1/AIN\[0\]
rlabel metal1 23966 6324 23966 6324 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux/cus_mux21_inst1/AIN\[1\]
rlabel metal1 23552 6426 23552 6426 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux/cus_mux21_inst1/_0_
rlabel metal2 23874 6596 23874 6596 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux/cus_mux21_inst1/_1_
rlabel metal1 19182 4590 19182 4590 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux/cus_mux21_inst2/AIN\[0\]
rlabel metal1 16054 2618 16054 2618 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux/cus_mux21_inst2/AIN\[1\]
rlabel metal1 20562 3502 20562 3502 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux/cus_mux21_inst2/_0_
rlabel metal2 23506 4522 23506 4522 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux/cus_mux21_inst2/_1_
rlabel metal1 17158 3604 17158 3604 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux/cus_mux21_inst3/AIN\[0\]
rlabel metal1 19964 4726 19964 4726 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux/cus_mux21_inst3/AIN\[1\]
rlabel via2 17250 3587 17250 3587 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux/cus_mux21_inst3/_0_
rlabel metal1 21689 6154 21689 6154 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux/cus_mux21_inst3/_1_
rlabel metal1 10902 25466 10902 25466 0 Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_N4BEG0/cus_mux21_inst/AIN\[0\]
rlabel metal1 11270 26010 11270 26010 0 Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_N4BEG0/cus_mux21_inst/AIN\[1\]
rlabel metal1 10902 26486 10902 26486 0 Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_N4BEG0/cus_mux21_inst/_0_
rlabel metal1 11132 26418 11132 26418 0 Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_N4BEG0/cus_mux21_inst/_1_
rlabel metal2 10994 24548 10994 24548 0 Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_N4BEG0/cus_mux41_buf_out0
rlabel metal1 10948 24378 10948 24378 0 Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_N4BEG0/cus_mux41_buf_out1
rlabel metal1 9200 39066 9200 39066 0 Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_N4BEG1/cus_mux21_inst/AIN\[0\]
rlabel metal1 9108 38182 9108 38182 0 Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_N4BEG1/cus_mux21_inst/AIN\[1\]
rlabel metal1 9384 39542 9384 39542 0 Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_N4BEG1/cus_mux21_inst/_0_
rlabel metal1 9338 39474 9338 39474 0 Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_N4BEG1/cus_mux21_inst/_1_
rlabel metal1 8648 38522 8648 38522 0 Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_N4BEG1/cus_mux41_buf_out0
rlabel metal1 8878 38318 8878 38318 0 Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_N4BEG1/cus_mux41_buf_out1
rlabel metal1 8832 33966 8832 33966 0 Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_N4BEG2/cus_mux21_inst/AIN\[0\]
rlabel metal1 10258 33626 10258 33626 0 Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_N4BEG2/cus_mux21_inst/AIN\[1\]
rlabel metal2 8694 34272 8694 34272 0 Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_N4BEG2/cus_mux21_inst/_0_
rlabel metal1 10350 34510 10350 34510 0 Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_N4BEG2/cus_mux21_inst/_1_
rlabel metal1 8970 31994 8970 31994 0 Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_N4BEG2/cus_mux41_buf_out0
rlabel metal2 9430 33014 9430 33014 0 Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_N4BEG2/cus_mux41_buf_out1
rlabel metal1 14858 35258 14858 35258 0 Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_N4BEG3/cus_mux21_inst/AIN\[0\]
rlabel metal2 15042 35700 15042 35700 0 Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_N4BEG3/cus_mux21_inst/AIN\[1\]
rlabel metal1 15134 35530 15134 35530 0 Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_N4BEG3/cus_mux21_inst/_0_
rlabel metal1 14950 35598 14950 35598 0 Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_N4BEG3/cus_mux21_inst/_1_
rlabel metal1 14996 32538 14996 32538 0 Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_N4BEG3/cus_mux41_buf_out0
rlabel metal1 15594 33082 15594 33082 0 Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_N4BEG3/cus_mux41_buf_out1
rlabel metal1 17434 21998 17434 21998 0 Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_S4BEG0/cus_mux21_inst/AIN\[0\]
rlabel metal1 17802 21896 17802 21896 0 Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_S4BEG0/cus_mux21_inst/AIN\[1\]
rlabel metal1 18032 21114 18032 21114 0 Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_S4BEG0/cus_mux21_inst/_0_
rlabel metal1 18354 21046 18354 21046 0 Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_S4BEG0/cus_mux21_inst/_1_
rlabel metal1 16284 22610 16284 22610 0 Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_S4BEG0/cus_mux41_buf_out0
rlabel metal1 17986 22032 17986 22032 0 Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_S4BEG0/cus_mux41_buf_out1
rlabel metal1 8924 20910 8924 20910 0 Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_S4BEG1/cus_mux21_inst/AIN\[0\]
rlabel metal1 9062 21896 9062 21896 0 Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_S4BEG1/cus_mux21_inst/AIN\[1\]
rlabel metal1 9614 20944 9614 20944 0 Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_S4BEG1/cus_mux21_inst/_0_
rlabel metal1 9982 20978 9982 20978 0 Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_S4BEG1/cus_mux21_inst/_1_
rlabel metal1 8648 22610 8648 22610 0 Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_S4BEG1/cus_mux41_buf_out0
rlabel metal1 8970 21998 8970 21998 0 Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_S4BEG1/cus_mux41_buf_out1
rlabel metal1 10718 29070 10718 29070 0 Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_S4BEG2/cus_mux21_inst/AIN\[0\]
rlabel metal1 10626 29172 10626 29172 0 Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_S4BEG2/cus_mux21_inst/AIN\[1\]
rlabel metal1 10718 28050 10718 28050 0 Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_S4BEG2/cus_mux21_inst/_0_
rlabel metal1 10764 28118 10764 28118 0 Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_S4BEG2/cus_mux21_inst/_1_
rlabel metal1 9844 29138 9844 29138 0 Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_S4BEG2/cus_mux41_buf_out0
rlabel metal1 9936 28186 9936 28186 0 Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_S4BEG2/cus_mux41_buf_out1
rlabel metal1 19044 18734 19044 18734 0 Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_S4BEG3/cus_mux21_inst/AIN\[0\]
rlabel metal1 19734 18802 19734 18802 0 Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_S4BEG3/cus_mux21_inst/AIN\[1\]
rlabel metal1 19090 18870 19090 18870 0 Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_S4BEG3/cus_mux21_inst/_0_
rlabel metal1 19320 18802 19320 18802 0 Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_S4BEG3/cus_mux21_inst/_1_
rlabel metal1 18354 18768 18354 18768 0 Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_S4BEG3/cus_mux41_buf_out0
rlabel metal1 18492 18394 18492 18394 0 Inst_RAM_IO_switch_matrix/inst_cus_mux81_buf_S4BEG3/cus_mux41_buf_out1
rlabel metal1 10442 21930 10442 21930 0 J_NS1_BEG\[0\]
rlabel metal1 7682 36822 7682 36822 0 J_NS1_BEG\[1\]
rlabel metal2 12558 35156 12558 35156 0 J_NS1_BEG\[2\]
rlabel metal1 15778 29206 15778 29206 0 J_NS1_BEG\[3\]
rlabel metal1 15376 17102 15376 17102 0 J_NS2_BEG\[0\]
rlabel metal2 2346 37604 2346 37604 0 J_NS2_BEG\[1\]
rlabel metal2 2346 32470 2346 32470 0 J_NS2_BEG\[2\]
rlabel via1 15698 19822 15698 19822 0 J_NS2_BEG\[3\]
rlabel metal1 13248 20434 13248 20434 0 J_NS2_BEG\[4\]
rlabel metal1 8740 20026 8740 20026 0 J_NS2_BEG\[5\]
rlabel metal2 2346 28118 2346 28118 0 J_NS2_BEG\[6\]
rlabel metal2 966 16116 966 16116 0 J_NS2_BEG\[7\]
rlabel via1 6831 3570 6831 3570 0 J_NS4_BEG\[0\]
rlabel metal3 5681 15844 5681 15844 0 J_NS4_BEG\[10\]
rlabel metal1 15134 32742 15134 32742 0 J_NS4_BEG\[11\]
rlabel metal1 11040 4998 11040 4998 0 J_NS4_BEG\[12\]
rlabel metal1 7314 36822 7314 36822 0 J_NS4_BEG\[13\]
rlabel metal1 1622 18802 1622 18802 0 J_NS4_BEG\[14\]
rlabel via1 17722 18190 17722 18190 0 J_NS4_BEG\[15\]
rlabel metal1 5221 21454 5221 21454 0 J_NS4_BEG\[1\]
rlabel metal1 5336 18802 5336 18802 0 J_NS4_BEG\[2\]
rlabel metal2 16468 19482 16468 19482 0 J_NS4_BEG\[3\]
rlabel metal1 14260 22066 14260 22066 0 J_NS4_BEG\[4\]
rlabel metal2 6210 16830 6210 16830 0 J_NS4_BEG\[5\]
rlabel metal1 8050 27948 8050 27948 0 J_NS4_BEG\[6\]
rlabel metal3 15548 32300 15548 32300 0 J_NS4_BEG\[7\]
rlabel metal1 13340 13702 13340 13702 0 J_NS4_BEG\[8\]
rlabel metal1 6866 16626 6866 16626 0 J_NS4_BEG\[9\]
rlabel metal2 138 44142 138 44142 0 N1BEG[0]
rlabel metal2 414 42306 414 42306 0 N1BEG[1]
rlabel metal2 690 44414 690 44414 0 N1BEG[2]
rlabel metal2 966 43598 966 43598 0 N1BEG[3]
rlabel metal2 138 262 138 262 0 N1END[0]
rlabel metal2 513 68 513 68 0 N1END[1]
rlabel metal1 1058 3502 1058 3502 0 N1END[2]
rlabel metal2 966 976 966 976 0 N1END[3]
rlabel metal2 1242 43530 1242 43530 0 N2BEG[0]
rlabel metal1 1794 39542 1794 39542 0 N2BEG[1]
rlabel metal2 1794 43853 1794 43853 0 N2BEG[2]
rlabel metal2 2070 43513 2070 43513 0 N2BEG[3]
rlabel metal2 2346 44074 2346 44074 0 N2BEG[4]
rlabel metal1 2484 42330 2484 42330 0 N2BEG[5]
rlabel metal2 2944 40358 2944 40358 0 N2BEG[6]
rlabel metal2 3174 43972 3174 43972 0 N2BEG[7]
rlabel metal2 3450 43632 3450 43632 0 N2BEGb[0]
rlabel metal1 3266 41242 3266 41242 0 N2BEGb[1]
rlabel metal2 3956 40698 3956 40698 0 N2BEGb[2]
rlabel metal2 4646 40698 4646 40698 0 N2BEGb[3]
rlabel metal1 3036 42874 3036 42874 0 N2BEGb[4]
rlabel metal1 4186 42534 4186 42534 0 N2BEGb[5]
rlabel metal1 3312 41446 3312 41446 0 N2BEGb[6]
rlabel metal1 4508 41786 4508 41786 0 N2BEGb[7]
rlabel metal2 3450 432 3450 432 0 N2END[0]
rlabel metal2 3726 704 3726 704 0 N2END[1]
rlabel metal2 4002 704 4002 704 0 N2END[2]
rlabel metal2 4278 670 4278 670 0 N2END[3]
rlabel metal2 4653 68 4653 68 0 N2END[4]
rlabel metal2 4830 636 4830 636 0 N2END[5]
rlabel metal2 5205 68 5205 68 0 N2END[6]
rlabel metal2 5382 1010 5382 1010 0 N2END[7]
rlabel metal2 1242 2540 1242 2540 0 N2MID[0]
rlabel metal2 1518 1095 1518 1095 0 N2MID[1]
rlabel metal2 1794 347 1794 347 0 N2MID[2]
rlabel metal1 2254 4182 2254 4182 0 N2MID[3]
rlabel metal2 2346 1724 2346 1724 0 N2MID[4]
rlabel metal2 2622 2336 2622 2336 0 N2MID[5]
rlabel metal1 2254 1292 2254 1292 0 N2MID[6]
rlabel metal1 4232 4658 4232 4658 0 N2MID[7]
rlabel metal1 3312 43350 3312 43350 0 N4BEG[0]
rlabel metal2 8418 44057 8418 44057 0 N4BEG[10]
rlabel metal1 8234 43146 8234 43146 0 N4BEG[11]
rlabel metal1 8832 43418 8832 43418 0 N4BEG[12]
rlabel metal2 9246 43921 9246 43921 0 N4BEG[13]
rlabel metal1 9338 43418 9338 43418 0 N4BEG[14]
rlabel metal1 9752 43418 9752 43418 0 N4BEG[15]
rlabel metal1 4784 43350 4784 43350 0 N4BEG[1]
rlabel metal1 6946 41786 6946 41786 0 N4BEG[2]
rlabel metal2 1610 43554 1610 43554 0 N4BEG[3]
rlabel metal1 6440 43418 6440 43418 0 N4BEG[4]
rlabel metal2 7038 44176 7038 44176 0 N4BEG[5]
rlabel metal1 6992 42330 6992 42330 0 N4BEG[6]
rlabel metal1 7084 43146 7084 43146 0 N4BEG[7]
rlabel metal2 7866 44057 7866 44057 0 N4BEG[8]
rlabel metal1 8740 42534 8740 42534 0 N4BEG[9]
rlabel metal2 6210 40545 6210 40545 0 N4BEG_i\[0\]
rlabel via2 8418 1819 8418 1819 0 N4BEG_i\[10\]
rlabel metal1 8832 2074 8832 2074 0 N4BEG_i\[11\]
rlabel metal2 506 1703 506 1703 0 N4BEG_i\[1\]
rlabel metal2 6118 1802 6118 1802 0 N4BEG_i\[2\]
rlabel metal2 1104 12420 1104 12420 0 N4BEG_i\[3\]
rlabel metal1 7130 2074 7130 2074 0 N4BEG_i\[4\]
rlabel metal4 644 21284 644 21284 0 N4BEG_i\[5\]
rlabel metal1 7728 1938 7728 1938 0 N4BEG_i\[6\]
rlabel metal4 828 19652 828 19652 0 N4BEG_i\[7\]
rlabel metal4 1012 22372 1012 22372 0 N4BEG_i\[8\]
rlabel metal1 8096 2074 8096 2074 0 N4BEG_i\[9\]
rlabel metal2 5658 500 5658 500 0 N4END[0]
rlabel metal2 8418 636 8418 636 0 N4END[10]
rlabel metal2 8694 636 8694 636 0 N4END[11]
rlabel metal2 9069 68 9069 68 0 N4END[12]
rlabel metal2 9345 68 9345 68 0 N4END[13]
rlabel metal2 9614 2465 9614 2465 0 N4END[14]
rlabel metal1 13202 1768 13202 1768 0 N4END[15]
rlabel metal2 5934 279 5934 279 0 N4END[1]
rlabel metal2 6210 347 6210 347 0 N4END[2]
rlabel metal2 6486 636 6486 636 0 N4END[3]
rlabel metal2 6663 68 6663 68 0 N4END[4]
rlabel metal2 7137 68 7137 68 0 N4END[5]
rlabel metal2 7314 619 7314 619 0 N4END[6]
rlabel metal2 7590 1421 7590 1421 0 N4END[7]
rlabel metal2 7912 3468 7912 3468 0 N4END[8]
rlabel metal2 8195 68 8195 68 0 N4END[9]
rlabel metal3 24848 7140 24848 7140 0 RAM2FAB_D0_I0
rlabel metal3 25285 7684 25285 7684 0 RAM2FAB_D0_I1
rlabel metal3 24940 8228 24940 8228 0 RAM2FAB_D0_I2
rlabel metal3 25285 8772 25285 8772 0 RAM2FAB_D0_I3
rlabel metal1 15088 13362 15088 13362 0 RAM2FAB_D0_O0
rlabel metal1 1840 18734 1840 18734 0 RAM2FAB_D0_O1
rlabel metal1 19734 8568 19734 8568 0 RAM2FAB_D0_O2
rlabel metal1 20838 9384 20838 9384 0 RAM2FAB_D0_O3
rlabel metal3 24848 4964 24848 4964 0 RAM2FAB_D1_I0
rlabel metal3 25285 5508 25285 5508 0 RAM2FAB_D1_I1
rlabel metal3 24917 6052 24917 6052 0 RAM2FAB_D1_I2
rlabel metal3 25262 6596 25262 6596 0 RAM2FAB_D1_I3
rlabel metal1 14490 7378 14490 7378 0 RAM2FAB_D1_O0
rlabel metal1 1886 13804 1886 13804 0 RAM2FAB_D1_O1
rlabel metal2 2346 15215 2346 15215 0 RAM2FAB_D1_O2
rlabel metal1 19320 5814 19320 5814 0 RAM2FAB_D1_O3
rlabel metal2 21022 4063 21022 4063 0 RAM2FAB_D2_I0
rlabel metal3 25285 3332 25285 3332 0 RAM2FAB_D2_I1
rlabel metal2 20930 4607 20930 4607 0 RAM2FAB_D2_I2
rlabel metal3 25285 4420 25285 4420 0 RAM2FAB_D2_I3
rlabel metal3 16100 3672 16100 3672 0 RAM2FAB_D2_O0
rlabel metal2 11638 5984 11638 5984 0 RAM2FAB_D2_O1
rlabel metal1 10074 13192 10074 13192 0 RAM2FAB_D2_O2
rlabel metal1 6992 10098 6992 10098 0 RAM2FAB_D2_O3
rlabel metal3 24020 612 24020 612 0 RAM2FAB_D3_I0
rlabel metal3 25285 1156 25285 1156 0 RAM2FAB_D3_I1
rlabel metal3 23836 1700 23836 1700 0 RAM2FAB_D3_I2
rlabel metal3 25285 2244 25285 2244 0 RAM2FAB_D3_I3
rlabel metal1 15410 13294 15410 13294 0 RAM2FAB_D3_O0
rlabel metal1 1656 18734 1656 18734 0 RAM2FAB_D3_O1
rlabel metal2 1518 21369 1518 21369 0 RAM2FAB_D3_O2
rlabel metal2 22310 3553 22310 3553 0 RAM2FAB_D3_O3
rlabel metal2 9522 1411 9522 1411 0 S1BEG[0]
rlabel metal2 10403 68 10403 68 0 S1BEG[1]
rlabel metal2 10626 483 10626 483 0 S1BEG[2]
rlabel metal2 10948 2788 10948 2788 0 S1BEG[3]
rlabel metal2 10074 44074 10074 44074 0 S1END[0]
rlabel metal2 10350 43598 10350 43598 0 S1END[1]
rlabel metal2 10626 43598 10626 43598 0 S1END[2]
rlabel metal2 10902 44193 10902 44193 0 S1END[3]
rlabel metal2 13386 636 13386 636 0 S2BEG[0]
rlabel metal2 13662 772 13662 772 0 S2BEG[1]
rlabel metal2 13938 636 13938 636 0 S2BEG[2]
rlabel metal2 14214 908 14214 908 0 S2BEG[3]
rlabel metal2 14490 806 14490 806 0 S2BEG[4]
rlabel metal2 14865 68 14865 68 0 S2BEG[5]
rlabel metal2 15095 68 15095 68 0 S2BEG[6]
rlabel metal2 15318 908 15318 908 0 S2BEG[7]
rlabel metal2 11178 772 11178 772 0 S2BEGb[0]
rlabel metal2 11454 466 11454 466 0 S2BEGb[1]
rlabel metal2 11730 483 11730 483 0 S2BEGb[2]
rlabel metal2 12006 330 12006 330 0 S2BEGb[3]
rlabel metal2 12282 636 12282 636 0 S2BEGb[4]
rlabel metal2 12558 738 12558 738 0 S2BEGb[5]
rlabel metal2 12933 68 12933 68 0 S2BEGb[6]
rlabel metal2 13110 143 13110 143 0 S2BEGb[7]
rlabel metal2 11178 43904 11178 43904 0 S2END[0]
rlabel metal2 11454 43598 11454 43598 0 S2END[1]
rlabel metal2 11730 43598 11730 43598 0 S2END[2]
rlabel metal2 12006 44193 12006 44193 0 S2END[3]
rlabel metal2 12282 43938 12282 43938 0 S2END[4]
rlabel metal2 12558 43972 12558 43972 0 S2END[5]
rlabel metal2 12834 44193 12834 44193 0 S2END[6]
rlabel metal2 13110 44261 13110 44261 0 S2END[7]
rlabel metal2 13386 43938 13386 43938 0 S2MID[0]
rlabel metal2 13662 44057 13662 44057 0 S2MID[1]
rlabel metal2 13938 43904 13938 43904 0 S2MID[2]
rlabel metal2 14214 44057 14214 44057 0 S2MID[3]
rlabel metal2 14490 43904 14490 43904 0 S2MID[4]
rlabel metal2 14766 43904 14766 43904 0 S2MID[5]
rlabel metal2 15042 44057 15042 44057 0 S2MID[6]
rlabel metal2 15318 43938 15318 43938 0 S2MID[7]
rlabel metal2 15693 68 15693 68 0 S4BEG[0]
rlabel metal2 18255 68 18255 68 0 S4BEG[10]
rlabel metal2 18729 68 18729 68 0 S4BEG[11]
rlabel metal2 18906 211 18906 211 0 S4BEG[12]
rlabel metal2 19235 68 19235 68 0 S4BEG[13]
rlabel metal2 19458 432 19458 432 0 S4BEG[14]
rlabel metal1 20010 3910 20010 3910 0 S4BEG[15]
rlabel metal2 15870 738 15870 738 0 S4BEG[1]
rlabel metal2 16245 68 16245 68 0 S4BEG[2]
rlabel metal2 16422 908 16422 908 0 S4BEG[3]
rlabel metal2 16698 942 16698 942 0 S4BEG[4]
rlabel metal2 16974 908 16974 908 0 S4BEG[5]
rlabel metal2 17349 68 17349 68 0 S4BEG[6]
rlabel metal1 17664 2822 17664 2822 0 S4BEG[7]
rlabel metal3 19182 3060 19182 3060 0 S4BEG[8]
rlabel metal2 18170 3468 18170 3468 0 S4BEG[9]
rlabel metal2 16514 918 16514 918 0 S4BEG_i\[0\]
rlabel metal3 20424 8364 20424 8364 0 S4BEG_i\[10\]
rlabel metal1 24012 1938 24012 1938 0 S4BEG_i\[11\]
rlabel metal1 22218 1972 22218 1972 0 S4BEG_i\[1\]
rlabel metal1 16836 2482 16836 2482 0 S4BEG_i\[2\]
rlabel metal3 16951 2652 16951 2652 0 S4BEG_i\[3\]
rlabel via3 17181 2652 17181 2652 0 S4BEG_i\[4\]
rlabel via3 22195 2652 22195 2652 0 S4BEG_i\[5\]
rlabel metal3 17871 5508 17871 5508 0 S4BEG_i\[6\]
rlabel via3 19619 2652 19619 2652 0 S4BEG_i\[7\]
rlabel metal1 18584 11050 18584 11050 0 S4BEG_i\[8\]
rlabel metal3 19389 8500 19389 8500 0 S4BEG_i\[9\]
rlabel metal2 15594 43904 15594 43904 0 S4END[0]
rlabel metal2 18354 43853 18354 43853 0 S4END[10]
rlabel metal2 18630 44193 18630 44193 0 S4END[11]
rlabel metal2 18906 44261 18906 44261 0 S4END[12]
rlabel metal2 19182 44397 19182 44397 0 S4END[13]
rlabel metal2 19458 44057 19458 44057 0 S4END[14]
rlabel metal1 20562 40086 20562 40086 0 S4END[15]
rlabel metal2 15870 43938 15870 43938 0 S4END[1]
rlabel metal2 16146 43972 16146 43972 0 S4END[2]
rlabel metal2 16422 43904 16422 43904 0 S4END[3]
rlabel metal2 16698 43870 16698 43870 0 S4END[4]
rlabel metal2 16974 43938 16974 43938 0 S4END[5]
rlabel metal2 17250 44193 17250 44193 0 S4END[6]
rlabel metal2 17526 44261 17526 44261 0 S4END[7]
rlabel metal2 17802 44329 17802 44329 0 S4END[8]
rlabel metal2 18078 44312 18078 44312 0 S4END[9]
rlabel metal1 16974 14858 16974 14858 0 UserCLK
rlabel metal1 20792 40698 20792 40698 0 UserCLKo
rlabel metal3 728 4964 728 4964 0 W1BEG[0]
rlabel metal2 3726 5015 3726 5015 0 W1BEG[1]
rlabel metal3 567 5508 567 5508 0 W1BEG[2]
rlabel metal1 2346 2006 2346 2006 0 W1BEG[3]
rlabel metal2 3266 5695 3266 5695 0 W2BEG[0]
rlabel metal3 1372 6324 1372 6324 0 W2BEG[1]
rlabel metal2 2898 4811 2898 4811 0 W2BEG[2]
rlabel metal2 4738 7021 4738 7021 0 W2BEG[3]
rlabel metal2 3542 6239 3542 6239 0 W2BEG[4]
rlabel metal2 4094 7463 4094 7463 0 W2BEG[5]
rlabel via2 4094 7701 4094 7701 0 W2BEG[6]
rlabel metal3 1004 7956 1004 7956 0 W2BEG[7]
rlabel metal2 3082 5933 3082 5933 0 W2BEGb[0]
rlabel metal3 1050 8500 1050 8500 0 W2BEGb[1]
rlabel metal2 3542 8075 3542 8075 0 W2BEGb[2]
rlabel metal3 2223 9044 2223 9044 0 W2BEGb[3]
rlabel metal3 1441 9316 1441 9316 0 W2BEGb[4]
rlabel metal2 4140 9588 4140 9588 0 W2BEGb[5]
rlabel metal2 2944 9860 2944 9860 0 W2BEGb[6]
rlabel metal2 4094 9911 4094 9911 0 W2BEGb[7]
rlabel metal3 728 14756 728 14756 0 W6BEG[0]
rlabel metal3 728 17476 728 17476 0 W6BEG[10]
rlabel metal2 3266 17901 3266 17901 0 W6BEG[11]
rlabel metal3 636 15028 636 15028 0 W6BEG[1]
rlabel metal3 682 15300 682 15300 0 W6BEG[2]
rlabel metal3 728 15572 728 15572 0 W6BEG[3]
rlabel metal3 636 15844 636 15844 0 W6BEG[4]
rlabel metal3 866 16116 866 16116 0 W6BEG[5]
rlabel metal2 3358 16031 3358 16031 0 W6BEG[6]
rlabel metal2 3726 15895 3726 15895 0 W6BEG[7]
rlabel metal3 498 16932 498 16932 0 W6BEG[8]
rlabel metal2 3450 17357 3450 17357 0 W6BEG[9]
rlabel metal2 3634 10319 3634 10319 0 WW4BEG[0]
rlabel metal3 682 13124 682 13124 0 WW4BEG[10]
rlabel metal3 406 13396 406 13396 0 WW4BEG[11]
rlabel metal2 3634 13311 3634 13311 0 WW4BEG[12]
rlabel metal3 567 13940 567 13940 0 WW4BEG[13]
rlabel metal3 659 14212 659 14212 0 WW4BEG[14]
rlabel metal2 4002 14535 4002 14535 0 WW4BEG[15]
rlabel metal2 3726 10421 3726 10421 0 WW4BEG[1]
rlabel via2 4002 10965 4002 10965 0 WW4BEG[2]
rlabel metal2 2990 10727 2990 10727 0 WW4BEG[3]
rlabel metal3 866 11492 866 11492 0 WW4BEG[4]
rlabel metal2 3450 11917 3450 11917 0 WW4BEG[5]
rlabel metal3 728 12036 728 12036 0 WW4BEG[6]
rlabel metal2 3726 12359 3726 12359 0 WW4BEG[7]
rlabel metal3 958 12580 958 12580 0 WW4BEG[8]
rlabel metal3 1878 12852 1878 12852 0 WW4BEG[9]
rlabel metal2 11638 14722 11638 14722 0 net1
rlabel via2 1426 32317 1426 32317 0 net10
rlabel metal2 20700 20298 20700 20298 0 net100
rlabel metal1 10902 7446 10902 7446 0 net101
rlabel metal1 1380 1190 1380 1190 0 net102
rlabel metal2 1610 3859 1610 3859 0 net103
rlabel metal1 2530 1768 2530 1768 0 net104
rlabel metal2 9430 4046 9430 4046 0 net105
rlabel metal4 19412 20196 19412 20196 0 net106
rlabel metal2 414 21148 414 21148 0 net107
rlabel metal1 17066 884 17066 884 0 net108
rlabel metal1 7360 3910 7360 3910 0 net109
rlabel metal2 2438 37808 2438 37808 0 net11
rlabel via2 7498 1173 7498 1173 0 net110
rlabel metal3 17963 19380 17963 19380 0 net111
rlabel metal1 6762 1768 6762 1768 0 net112
rlabel metal2 11086 1853 11086 1853 0 net113
rlabel metal1 1794 3910 1794 3910 0 net114
rlabel metal1 2116 1190 2116 1190 0 net115
rlabel metal2 12834 33405 12834 33405 0 net116
rlabel metal2 11454 4352 11454 4352 0 net117
rlabel metal1 1058 16422 1058 16422 0 net118
rlabel metal2 2438 884 2438 884 0 net119
rlabel metal1 3588 23698 3588 23698 0 net12
rlabel metal1 5382 2346 5382 2346 0 net120
rlabel metal2 6670 1020 6670 1020 0 net121
rlabel metal1 7222 1904 7222 1904 0 net122
rlabel metal1 7590 1292 7590 1292 0 net123
rlabel metal1 7682 2006 7682 2006 0 net124
rlabel metal1 8602 2006 8602 2006 0 net125
rlabel metal1 8326 1938 8326 1938 0 net126
rlabel metal1 9522 2006 9522 2006 0 net127
rlabel metal3 16169 8364 16169 8364 0 net128
rlabel metal2 5704 21658 5704 21658 0 net129
rlabel metal1 2622 18088 2622 18088 0 net13
rlabel metal1 8372 2482 8372 2482 0 net130
rlabel metal1 6992 2414 6992 2414 0 net131
rlabel metal2 6026 1802 6026 1802 0 net132
rlabel metal1 6394 1938 6394 1938 0 net133
rlabel metal1 6900 2890 6900 2890 0 net134
rlabel metal1 7406 1802 7406 1802 0 net135
rlabel metal1 8004 2346 8004 2346 0 net136
rlabel metal2 20746 7191 20746 7191 0 net137
rlabel metal1 18906 8466 18906 8466 0 net138
rlabel metal1 23046 7820 23046 7820 0 net139
rlabel metal1 2300 20570 2300 20570 0 net14
rlabel metal1 20010 8432 20010 8432 0 net140
rlabel metal1 17342 11798 17342 11798 0 net141
rlabel metal1 22448 10642 22448 10642 0 net142
rlabel metal1 20608 6766 20608 6766 0 net143
rlabel metal1 19407 6358 19407 6358 0 net144
rlabel metal1 22678 2380 22678 2380 0 net145
rlabel metal1 21707 4522 21707 4522 0 net146
rlabel metal1 21022 5338 21022 5338 0 net147
rlabel metal1 21436 8466 21436 8466 0 net148
rlabel metal1 17418 2346 17418 2346 0 net149
rlabel metal1 8648 17170 8648 17170 0 net15
rlabel metal1 17986 748 17986 748 0 net150
rlabel metal1 21712 3910 21712 3910 0 net151
rlabel metal1 20424 3366 20424 3366 0 net152
rlabel metal4 21068 26112 21068 26112 0 net153
rlabel metal1 4416 14382 4416 14382 0 net154
rlabel metal1 3588 36006 3588 36006 0 net155
rlabel metal2 13248 36550 13248 36550 0 net156
rlabel metal3 10327 2516 10327 2516 0 net157
rlabel metal2 10074 39049 10074 39049 0 net158
rlabel metal3 8464 30804 8464 30804 0 net159
rlabel metal1 3220 18938 3220 18938 0 net16
rlabel metal1 12144 43078 12144 43078 0 net160
rlabel via2 12558 43061 12558 43061 0 net161
rlabel metal2 12466 41973 12466 41973 0 net162
rlabel metal1 11316 33014 11316 33014 0 net163
rlabel metal2 13340 20604 13340 20604 0 net164
rlabel metal3 13455 20740 13455 20740 0 net165
rlabel metal1 13938 42568 13938 42568 0 net166
rlabel metal2 12144 37468 12144 37468 0 net167
rlabel metal1 13800 42738 13800 42738 0 net168
rlabel metal2 14674 40936 14674 40936 0 net169
rlabel metal2 1702 20009 1702 20009 0 net17
rlabel via3 15019 42908 15019 42908 0 net170
rlabel metal1 13340 30294 13340 30294 0 net171
rlabel metal1 13892 2414 13892 2414 0 net172
rlabel metal1 13570 18394 13570 18394 0 net173
rlabel metal1 18998 42602 18998 42602 0 net174
rlabel metal1 18906 42704 18906 42704 0 net175
rlabel metal1 18446 42296 18446 42296 0 net176
rlabel metal1 19688 42670 19688 42670 0 net177
rlabel metal1 20194 42602 20194 42602 0 net178
rlabel metal1 20424 40154 20424 40154 0 net179
rlabel metal1 2024 20570 2024 20570 0 net18
rlabel metal2 16882 43486 16882 43486 0 net180
rlabel metal2 14122 42364 14122 42364 0 net181
rlabel metal2 13938 14535 13938 14535 0 net182
rlabel metal1 16652 42670 16652 42670 0 net183
rlabel metal1 17158 42602 17158 42602 0 net184
rlabel metal1 17204 42670 17204 42670 0 net185
rlabel metal1 17434 42704 17434 42704 0 net186
rlabel metal1 17848 42670 17848 42670 0 net187
rlabel metal1 18170 42738 18170 42738 0 net188
rlabel metal1 23966 8908 23966 8908 0 net189
rlabel metal1 1150 20570 1150 20570 0 net19
rlabel metal1 23213 9962 23213 9962 0 net190
rlabel viali 22862 10027 22862 10027 0 net191
rlabel metal1 23966 10030 23966 10030 0 net192
rlabel metal2 21482 16456 21482 16456 0 net193
rlabel metal1 23966 16116 23966 16116 0 net194
rlabel metal1 23460 17170 23460 17170 0 net195
rlabel metal1 23736 17646 23736 17646 0 net196
rlabel metal1 23966 13260 23966 13260 0 net197
rlabel metal1 23690 14314 23690 14314 0 net198
rlabel metal1 23966 15062 23966 15062 0 net199
rlabel via2 1702 40477 1702 40477 0 net2
rlabel metal1 3496 21318 3496 21318 0 net20
rlabel metal2 20654 16779 20654 16779 0 net200
rlabel metal2 23414 12852 23414 12852 0 net201
rlabel metal2 20700 21964 20700 21964 0 net202
rlabel metal2 20424 19346 20424 19346 0 net203
rlabel metal1 21298 12648 21298 12648 0 net204
rlabel metal1 23598 24174 23598 24174 0 net205
rlabel metal1 23874 25874 23874 25874 0 net206
rlabel metal2 23598 26860 23598 26860 0 net207
rlabel metal2 22034 27098 22034 27098 0 net208
rlabel metal1 23598 22508 23598 22508 0 net209
rlabel via1 12570 25330 12570 25330 0 net21
rlabel metal1 24380 22610 24380 22610 0 net210
rlabel metal1 23920 23766 23920 23766 0 net211
rlabel metal1 20654 26248 20654 26248 0 net212
rlabel metal2 20608 19482 20608 19482 0 net213
rlabel metal1 25392 21998 25392 21998 0 net214
rlabel metal2 21942 21767 21942 21767 0 net215
rlabel metal1 24748 22066 24748 22066 0 net216
rlabel metal1 21436 24038 21436 24038 0 net217
rlabel metal1 24104 17646 24104 17646 0 net218
rlabel metal1 23644 19414 23644 19414 0 net219
rlabel metal2 10166 32470 10166 32470 0 net22
rlabel metal1 23644 18258 23644 18258 0 net220
rlabel metal1 23966 26928 23966 26928 0 net221
rlabel metal1 23966 32470 23966 32470 0 net222
rlabel metal1 23966 32912 23966 32912 0 net223
rlabel metal1 23966 33456 23966 33456 0 net224
rlabel metal1 23966 34000 23966 34000 0 net225
rlabel metal1 23644 34646 23644 34646 0 net226
rlabel metal1 23966 35088 23966 35088 0 net227
rlabel metal1 23966 35632 23966 35632 0 net228
rlabel metal1 23506 36074 23506 36074 0 net229
rlabel metal1 9520 31144 9520 31144 0 net23
rlabel metal2 23966 36550 23966 36550 0 net230
rlabel metal1 22034 37230 22034 37230 0 net231
rlabel metal1 23966 27404 23966 27404 0 net232
rlabel metal1 21850 37128 21850 37128 0 net233
rlabel metal1 23828 37978 23828 37978 0 net234
rlabel metal1 22954 38522 22954 38522 0 net235
rlabel metal2 20378 39270 20378 39270 0 net236
rlabel metal1 20654 39542 20654 39542 0 net237
rlabel metal1 22816 39542 22816 39542 0 net238
rlabel metal2 22034 40630 22034 40630 0 net239
rlabel via1 2450 28050 2450 28050 0 net24
rlabel metal1 23184 38794 23184 38794 0 net240
rlabel metal1 23874 42670 23874 42670 0 net241
rlabel metal1 23644 42194 23644 42194 0 net242
rlabel metal1 23460 27574 23460 27574 0 net243
rlabel metal2 22586 41990 22586 41990 0 net244
rlabel metal1 21252 41786 21252 41786 0 net245
rlabel metal1 23966 28492 23966 28492 0 net246
rlabel metal1 23782 29206 23782 29206 0 net247
rlabel metal1 23966 29648 23966 29648 0 net248
rlabel metal1 23966 30192 23966 30192 0 net249
rlabel metal1 11546 35734 11546 35734 0 net25
rlabel metal1 23782 30702 23782 30702 0 net250
rlabel metal1 23966 31348 23966 31348 0 net251
rlabel metal1 23874 31824 23874 31824 0 net252
rlabel metal1 20240 42874 20240 42874 0 net253
rlabel metal1 21988 40970 21988 40970 0 net254
rlabel metal1 21850 41242 21850 41242 0 net255
rlabel metal1 23414 40154 23414 40154 0 net256
rlabel metal2 21942 40783 21942 40783 0 net257
rlabel metal1 21206 41208 21206 41208 0 net258
rlabel metal1 23230 40698 23230 40698 0 net259
rlabel via1 15755 28050 15755 28050 0 net26
rlabel metal1 23644 36278 23644 36278 0 net260
rlabel metal1 23414 41446 23414 41446 0 net261
rlabel metal1 23828 32266 23828 32266 0 net262
rlabel metal3 21643 43180 21643 43180 0 net263
rlabel metal1 20654 41718 20654 41718 0 net264
rlabel viali 21850 43284 21850 43284 0 net265
rlabel metal1 21022 41242 21022 41242 0 net266
rlabel metal1 21942 41718 21942 41718 0 net267
rlabel metal2 22862 43044 22862 43044 0 net268
rlabel metal2 21850 37315 21850 37315 0 net269
rlabel metal1 2668 29002 2668 29002 0 net27
rlabel metal1 23184 42670 23184 42670 0 net270
rlabel metal1 23046 42602 23046 42602 0 net271
rlabel metal1 22034 42160 22034 42160 0 net272
rlabel metal1 12282 34102 12282 34102 0 net273
rlabel metal1 4554 40562 4554 40562 0 net274
rlabel metal2 3542 37434 3542 37434 0 net275
rlabel metal1 16468 33626 16468 33626 0 net276
rlabel metal2 16606 36023 16606 36023 0 net277
rlabel metal2 1886 38386 1886 38386 0 net278
rlabel metal1 3634 32198 3634 32198 0 net279
rlabel metal2 2714 32572 2714 32572 0 net28
rlabel metal4 2668 35904 2668 35904 0 net280
rlabel metal2 6118 24599 6118 24599 0 net281
rlabel metal2 14030 35972 14030 35972 0 net282
rlabel metal1 1840 28526 1840 28526 0 net283
rlabel metal4 2668 28152 2668 28152 0 net284
rlabel metal1 1794 42602 1794 42602 0 net285
rlabel via1 2622 39627 2622 39627 0 net286
rlabel metal1 3818 31450 3818 31450 0 net287
rlabel metal1 4278 33626 4278 33626 0 net288
rlabel via2 2714 42619 2714 42619 0 net289
rlabel metal1 1748 35054 1748 35054 0 net29
rlabel metal3 4899 20604 4899 20604 0 net290
rlabel metal3 1495 41412 1495 41412 0 net291
rlabel via2 5382 2635 5382 2635 0 net292
rlabel metal2 2714 43588 2714 43588 0 net293
rlabel metal2 9246 42194 9246 42194 0 net294
rlabel metal2 9154 42772 9154 42772 0 net295
rlabel metal1 8648 43282 8648 43282 0 net296
rlabel metal1 9292 39610 9292 39610 0 net297
rlabel metal1 10120 34714 10120 34714 0 net298
rlabel metal1 15042 35802 15042 35802 0 net299
rlabel metal2 13110 26979 13110 26979 0 net3
rlabel via1 17722 19278 17722 19278 0 net30
rlabel metal1 4646 43826 4646 43826 0 net300
rlabel metal2 7176 41582 7176 41582 0 net301
rlabel metal1 1426 43928 1426 43928 0 net302
rlabel metal1 10258 42296 10258 42296 0 net303
rlabel metal2 3450 41208 3450 41208 0 net304
rlabel metal1 6486 42228 6486 42228 0 net305
rlabel metal1 6394 43180 6394 43180 0 net306
rlabel metal1 6854 42670 6854 42670 0 net307
rlabel metal2 8970 42228 8970 42228 0 net308
rlabel metal1 10258 15878 10258 15878 0 net309
rlabel metal1 10488 16422 10488 16422 0 net31
rlabel metal1 9660 17306 9660 17306 0 net310
rlabel metal1 9614 1904 9614 1904 0 net311
rlabel metal3 18699 29036 18699 29036 0 net312
rlabel via3 13501 1292 13501 1292 0 net313
rlabel via3 14605 1292 14605 1292 0 net314
rlabel metal3 14191 1292 14191 1292 0 net315
rlabel via2 14490 2091 14490 2091 0 net316
rlabel metal1 15272 1326 15272 1326 0 net317
rlabel metal1 12098 1360 12098 1360 0 net318
rlabel metal2 16882 7548 16882 7548 0 net319
rlabel metal1 6394 33830 6394 33830 0 net32
rlabel metal2 15318 17170 15318 17170 0 net320
rlabel metal1 8832 1258 8832 1258 0 net321
rlabel metal3 8349 1292 8349 1292 0 net322
rlabel metal3 11983 2380 11983 2380 0 net323
rlabel via3 11109 1292 11109 1292 0 net324
rlabel metal2 11822 1530 11822 1530 0 net325
rlabel metal2 12236 1326 12236 1326 0 net326
rlabel via2 12742 1309 12742 1309 0 net327
rlabel metal1 13248 1326 13248 1326 0 net328
rlabel metal1 16192 1530 16192 1530 0 net329
rlabel metal1 9154 23732 9154 23732 0 net33
rlabel metal1 20424 3162 20424 3162 0 net330
rlabel metal1 19182 3978 19182 3978 0 net331
rlabel metal2 18952 20604 18952 20604 0 net332
rlabel metal2 12466 19040 12466 19040 0 net333
rlabel metal3 20079 4012 20079 4012 0 net334
rlabel metal1 19136 18598 19136 18598 0 net335
rlabel metal1 16744 1258 16744 1258 0 net336
rlabel metal1 18216 2006 18216 2006 0 net337
rlabel metal1 16744 2006 16744 2006 0 net338
rlabel metal1 18906 2006 18906 2006 0 net339
rlabel metal1 5612 28050 5612 28050 0 net34
rlabel metal1 23184 1190 23184 1190 0 net340
rlabel metal1 17664 2006 17664 2006 0 net341
rlabel metal1 19228 2278 19228 2278 0 net342
rlabel metal1 18630 2822 18630 2822 0 net343
rlabel metal1 18538 3502 18538 3502 0 net344
rlabel metal1 21114 40562 21114 40562 0 net345
rlabel metal2 8970 4386 8970 4386 0 net346
rlabel metal1 5658 14246 5658 14246 0 net347
rlabel metal1 1932 2414 1932 2414 0 net348
rlabel metal1 1610 2006 1610 2006 0 net349
rlabel metal1 14674 28118 14674 28118 0 net35
rlabel metal1 4738 5270 4738 5270 0 net350
rlabel metal1 4278 4590 4278 4590 0 net351
rlabel metal2 2254 3638 2254 3638 0 net352
rlabel metal2 7498 7208 7498 7208 0 net353
rlabel metal1 14375 5542 14375 5542 0 net354
rlabel metal1 5750 7344 5750 7344 0 net355
rlabel metal1 3910 5882 3910 5882 0 net356
rlabel metal1 2231 3094 2231 3094 0 net357
rlabel metal1 3634 3434 3634 3434 0 net358
rlabel metal1 3128 7786 3128 7786 0 net359
rlabel metal1 14030 25262 14030 25262 0 net36
rlabel metal1 5336 7378 5336 7378 0 net360
rlabel metal1 3864 9962 3864 9962 0 net361
rlabel metal1 14904 7514 14904 7514 0 net362
rlabel metal1 3864 10030 3864 10030 0 net363
rlabel metal2 2070 8109 2070 8109 0 net364
rlabel metal1 4922 3162 4922 3162 0 net365
rlabel metal2 10672 12988 10672 12988 0 net366
rlabel metal1 3496 17646 3496 17646 0 net367
rlabel metal1 8372 14042 8372 14042 0 net368
rlabel metal2 2714 16949 2714 16949 0 net369
rlabel metal1 7314 24888 7314 24888 0 net37
rlabel metal3 5727 17884 5727 17884 0 net370
rlabel metal1 13202 12410 13202 12410 0 net371
rlabel metal1 1886 15470 1886 15470 0 net372
rlabel metal2 1518 14178 1518 14178 0 net373
rlabel metal1 5980 15402 5980 15402 0 net374
rlabel metal2 7498 12818 7498 12818 0 net375
rlabel metal2 1518 16575 1518 16575 0 net376
rlabel metal1 4830 17578 4830 17578 0 net377
rlabel metal1 14950 9112 14950 9112 0 net378
rlabel metal2 2254 13022 2254 13022 0 net379
rlabel metal1 7636 29070 7636 29070 0 net38
rlabel metal1 2070 10472 2070 10472 0 net380
rlabel metal2 17342 13056 17342 13056 0 net381
rlabel metal2 2162 15368 2162 15368 0 net382
rlabel via3 1541 12172 1541 12172 0 net383
rlabel metal2 7590 5440 7590 5440 0 net384
rlabel metal1 5612 10030 5612 10030 0 net385
rlabel metal2 3266 21862 3266 21862 0 net386
rlabel metal2 9522 6052 9522 6052 0 net387
rlabel via2 1518 6715 1518 6715 0 net388
rlabel metal1 6256 11322 6256 11322 0 net389
rlabel metal1 9522 28152 9522 28152 0 net39
rlabel metal2 4186 12852 4186 12852 0 net390
rlabel metal1 8648 7174 8648 7174 0 net391
rlabel metal2 17434 10863 17434 10863 0 net392
rlabel metal1 4462 11152 4462 11152 0 net393
rlabel metal1 14076 28730 14076 28730 0 net394
rlabel metal2 15594 17408 15594 17408 0 net395
rlabel metal1 12098 17714 12098 17714 0 net396
rlabel metal2 9430 19006 9430 19006 0 net397
rlabel metal1 15824 19890 15824 19890 0 net398
rlabel metal2 13386 16320 13386 16320 0 net399
rlabel metal1 16744 19278 16744 19278 0 net4
rlabel via2 1610 24667 1610 24667 0 net40
rlabel metal2 9430 15232 9430 15232 0 net400
rlabel metal2 11178 20026 11178 20026 0 net401
rlabel metal2 17066 21488 17066 21488 0 net402
rlabel metal2 12466 14076 12466 14076 0 net403
rlabel metal1 7314 41140 7314 41140 0 net404
rlabel metal1 12282 35564 12282 35564 0 net405
rlabel metal1 10166 12886 10166 12886 0 net406
rlabel metal1 2438 42262 2438 42262 0 net407
rlabel metal1 3358 35768 3358 35768 0 net408
rlabel viali 16514 29141 16514 29141 0 net409
rlabel metal1 6992 31790 6992 31790 0 net41
rlabel metal1 13754 32198 13754 32198 0 net42
rlabel metal1 13754 24786 13754 24786 0 net43
rlabel metal1 7590 24922 7590 24922 0 net44
rlabel metal1 8142 27064 8142 27064 0 net45
rlabel metal1 6210 25976 6210 25976 0 net46
rlabel metal1 3266 25160 3266 25160 0 net47
rlabel metal1 3266 26758 3266 26758 0 net48
rlabel metal2 1748 31790 1748 31790 0 net49
rlabel via1 14410 18258 14410 18258 0 net5
rlabel metal1 1702 39013 1702 39013 0 net50
rlabel metal2 2484 8228 2484 8228 0 net51
rlabel metal1 17986 33388 17986 33388 0 net52
rlabel metal1 17250 34408 17250 34408 0 net53
rlabel via1 16973 17646 16973 17646 0 net54
rlabel metal1 7865 14382 7865 14382 0 net55
rlabel metal1 17250 35190 17250 35190 0 net56
rlabel metal2 2714 23205 2714 23205 0 net57
rlabel metal1 20654 36176 20654 36176 0 net58
rlabel metal1 21206 36720 21206 36720 0 net59
rlabel metal1 8878 17850 8878 17850 0 net6
rlabel metal1 15087 4590 15087 4590 0 net60
rlabel metal2 1656 40052 1656 40052 0 net61
rlabel metal2 19366 36329 19366 36329 0 net62
rlabel metal1 20637 19822 20637 19822 0 net63
rlabel metal2 2024 32164 2024 32164 0 net64
rlabel via1 15501 8466 15501 8466 0 net65
rlabel metal2 22034 38658 22034 38658 0 net66
rlabel metal3 2461 6460 2461 6460 0 net67
rlabel metal1 2575 41582 2575 41582 0 net68
rlabel metal2 2392 17068 2392 17068 0 net69
rlabel metal1 2070 20774 2070 20774 0 net7
rlabel metal3 2277 41412 2277 41412 0 net70
rlabel metal1 19687 33966 19687 33966 0 net71
rlabel metal1 1518 41038 1518 41038 0 net72
rlabel metal1 19642 20808 19642 20808 0 net73
rlabel metal2 19964 14212 19964 14212 0 net74
rlabel via1 2253 17170 2253 17170 0 net75
rlabel metal3 1817 5508 1817 5508 0 net76
rlabel metal1 18537 21522 18537 21522 0 net77
rlabel metal1 16651 31790 16651 31790 0 net78
rlabel metal1 20286 24174 20286 24174 0 net79
rlabel metal1 13294 19992 13294 19992 0 net8
rlabel metal1 15042 32198 15042 32198 0 net80
rlabel metal2 2622 35071 2622 35071 0 net81
rlabel metal2 20378 13294 20378 13294 0 net82
rlabel metal2 23644 16796 23644 16796 0 net83
rlabel metal1 22678 40494 22678 40494 0 net84
rlabel metal2 25070 35836 25070 35836 0 net85
rlabel metal1 24610 2618 24610 2618 0 net86
rlabel metal2 25300 35564 25300 35564 0 net87
rlabel metal3 21183 2380 21183 2380 0 net88
rlabel metal2 23322 35037 23322 35037 0 net89
rlabel metal2 12466 16218 12466 16218 0 net9
rlabel metal2 23000 13804 23000 13804 0 net90
rlabel metal2 25530 34476 25530 34476 0 net91
rlabel metal1 21298 2550 21298 2550 0 net92
rlabel metal2 19918 2278 19918 2278 0 net93
rlabel metal1 18446 41038 18446 41038 0 net94
rlabel metal2 20838 15062 20838 15062 0 net95
rlabel metal1 23368 2482 23368 2482 0 net96
rlabel metal1 21252 1258 21252 1258 0 net97
rlabel metal1 19918 1428 19918 1428 0 net98
rlabel metal1 1564 32878 1564 32878 0 net99
<< properties >>
string FIXED_BBOX 0 0 25700 44700
<< end >>
