magic
tech sky130A
magscale 1 2
timestamp 1733615923
<< obsli1 >>
rect 1104 1071 45540 43537
<< obsm1 >>
rect 198 620 46630 43988
<< metal2 >>
rect 478 44540 534 45000
rect 846 44540 902 45000
rect 1214 44540 1270 45000
rect 1582 44540 1638 45000
rect 1950 44540 2006 45000
rect 2318 44540 2374 45000
rect 2686 44540 2742 45000
rect 3054 44540 3110 45000
rect 3422 44540 3478 45000
rect 3790 44540 3846 45000
rect 4158 44540 4214 45000
rect 4526 44540 4582 45000
rect 4894 44540 4950 45000
rect 5262 44540 5318 45000
rect 5630 44540 5686 45000
rect 5998 44540 6054 45000
rect 6366 44540 6422 45000
rect 6734 44540 6790 45000
rect 7102 44540 7158 45000
rect 7470 44540 7526 45000
rect 7838 44540 7894 45000
rect 8206 44540 8262 45000
rect 8574 44540 8630 45000
rect 8942 44540 8998 45000
rect 9310 44540 9366 45000
rect 9678 44540 9734 45000
rect 10046 44540 10102 45000
rect 10414 44540 10470 45000
rect 10782 44540 10838 45000
rect 11150 44540 11206 45000
rect 11518 44540 11574 45000
rect 11886 44540 11942 45000
rect 12254 44540 12310 45000
rect 12622 44540 12678 45000
rect 12990 44540 13046 45000
rect 13358 44540 13414 45000
rect 13726 44540 13782 45000
rect 14094 44540 14150 45000
rect 14462 44540 14518 45000
rect 14830 44540 14886 45000
rect 15198 44540 15254 45000
rect 15566 44540 15622 45000
rect 15934 44540 15990 45000
rect 16302 44540 16358 45000
rect 16670 44540 16726 45000
rect 17038 44540 17094 45000
rect 17406 44540 17462 45000
rect 17774 44540 17830 45000
rect 18142 44540 18198 45000
rect 18510 44540 18566 45000
rect 18878 44540 18934 45000
rect 19246 44540 19302 45000
rect 19614 44540 19670 45000
rect 19982 44540 20038 45000
rect 20350 44540 20406 45000
rect 20718 44540 20774 45000
rect 21086 44540 21142 45000
rect 21454 44540 21510 45000
rect 21822 44540 21878 45000
rect 22190 44540 22246 45000
rect 22558 44540 22614 45000
rect 22926 44540 22982 45000
rect 23294 44540 23350 45000
rect 23662 44540 23718 45000
rect 24030 44540 24086 45000
rect 24398 44540 24454 45000
rect 24766 44540 24822 45000
rect 25134 44540 25190 45000
rect 25502 44540 25558 45000
rect 25870 44540 25926 45000
rect 26238 44540 26294 45000
rect 26606 44540 26662 45000
rect 26974 44540 27030 45000
rect 27342 44540 27398 45000
rect 27710 44540 27766 45000
rect 28078 44540 28134 45000
rect 28446 44540 28502 45000
rect 28814 44540 28870 45000
rect 29182 44540 29238 45000
rect 29550 44540 29606 45000
rect 29918 44540 29974 45000
rect 30286 44540 30342 45000
rect 30654 44540 30710 45000
rect 31022 44540 31078 45000
rect 31390 44540 31446 45000
rect 31758 44540 31814 45000
rect 32126 44540 32182 45000
rect 32494 44540 32550 45000
rect 32862 44540 32918 45000
rect 33230 44540 33286 45000
rect 33598 44540 33654 45000
rect 33966 44540 34022 45000
rect 34334 44540 34390 45000
rect 34702 44540 34758 45000
rect 35070 44540 35126 45000
rect 35438 44540 35494 45000
rect 35806 44540 35862 45000
rect 36174 44540 36230 45000
rect 36542 44540 36598 45000
rect 36910 44540 36966 45000
rect 37278 44540 37334 45000
rect 37646 44540 37702 45000
rect 38014 44540 38070 45000
rect 38382 44540 38438 45000
rect 38750 44540 38806 45000
rect 39118 44540 39174 45000
rect 39486 44540 39542 45000
rect 39854 44540 39910 45000
rect 40222 44540 40278 45000
rect 40590 44540 40646 45000
rect 40958 44540 41014 45000
rect 41326 44540 41382 45000
rect 41694 44540 41750 45000
rect 42062 44540 42118 45000
rect 42430 44540 42486 45000
rect 42798 44540 42854 45000
rect 43166 44540 43222 45000
rect 43534 44540 43590 45000
rect 43902 44540 43958 45000
rect 44270 44540 44326 45000
rect 44638 44540 44694 45000
rect 45006 44540 45062 45000
rect 45374 44540 45430 45000
rect 45742 44540 45798 45000
rect 46110 44540 46166 45000
rect 478 -300 534 160
rect 846 -300 902 160
rect 1214 -300 1270 160
rect 1582 -300 1638 160
rect 1950 -300 2006 160
rect 2318 -300 2374 160
rect 2686 -300 2742 160
rect 3054 -300 3110 160
rect 3422 -300 3478 160
rect 3790 -300 3846 160
rect 4158 -300 4214 160
rect 4526 -300 4582 160
rect 4894 -300 4950 160
rect 5262 -300 5318 160
rect 5630 -300 5686 160
rect 5998 -300 6054 160
rect 6366 -300 6422 160
rect 6734 -300 6790 160
rect 7102 -300 7158 160
rect 7470 -300 7526 160
rect 7838 -300 7894 160
rect 8206 -300 8262 160
rect 8574 -300 8630 160
rect 8942 -300 8998 160
rect 9310 -300 9366 160
rect 9678 -300 9734 160
rect 10046 -300 10102 160
rect 10414 -300 10470 160
rect 10782 -300 10838 160
rect 11150 -300 11206 160
rect 11518 -300 11574 160
rect 11886 -300 11942 160
rect 12254 -300 12310 160
rect 12622 -300 12678 160
rect 12990 -300 13046 160
rect 13358 -300 13414 160
rect 13726 -300 13782 160
rect 14094 -300 14150 160
rect 14462 -300 14518 160
rect 14830 -300 14886 160
rect 15198 -300 15254 160
rect 15566 -300 15622 160
rect 15934 -300 15990 160
rect 16302 -300 16358 160
rect 16670 -300 16726 160
rect 17038 -300 17094 160
rect 17406 -300 17462 160
rect 17774 -300 17830 160
rect 18142 -300 18198 160
rect 18510 -300 18566 160
rect 18878 -300 18934 160
rect 19246 -300 19302 160
rect 19614 -300 19670 160
rect 19982 -300 20038 160
rect 20350 -300 20406 160
rect 20718 -300 20774 160
rect 21086 -300 21142 160
rect 21454 -300 21510 160
rect 21822 -300 21878 160
rect 22190 -300 22246 160
rect 22558 -300 22614 160
rect 22926 -300 22982 160
rect 23294 -300 23350 160
rect 23662 -300 23718 160
rect 24030 -300 24086 160
rect 24398 -300 24454 160
rect 24766 -300 24822 160
rect 25134 -300 25190 160
rect 25502 -300 25558 160
rect 25870 -300 25926 160
rect 26238 -300 26294 160
rect 26606 -300 26662 160
rect 26974 -300 27030 160
rect 27342 -300 27398 160
rect 27710 -300 27766 160
rect 28078 -300 28134 160
rect 28446 -300 28502 160
rect 28814 -300 28870 160
rect 29182 -300 29238 160
rect 29550 -300 29606 160
rect 29918 -300 29974 160
rect 30286 -300 30342 160
rect 30654 -300 30710 160
rect 31022 -300 31078 160
rect 31390 -300 31446 160
rect 31758 -300 31814 160
rect 32126 -300 32182 160
rect 32494 -300 32550 160
rect 32862 -300 32918 160
rect 33230 -300 33286 160
rect 33598 -300 33654 160
rect 33966 -300 34022 160
rect 34334 -300 34390 160
rect 34702 -300 34758 160
rect 35070 -300 35126 160
rect 35438 -300 35494 160
rect 35806 -300 35862 160
rect 36174 -300 36230 160
rect 36542 -300 36598 160
rect 36910 -300 36966 160
rect 37278 -300 37334 160
rect 37646 -300 37702 160
rect 38014 -300 38070 160
rect 38382 -300 38438 160
rect 38750 -300 38806 160
rect 39118 -300 39174 160
rect 39486 -300 39542 160
rect 39854 -300 39910 160
rect 40222 -300 40278 160
rect 40590 -300 40646 160
rect 40958 -300 41014 160
rect 41326 -300 41382 160
rect 41694 -300 41750 160
rect 42062 -300 42118 160
rect 42430 -300 42486 160
rect 42798 -300 42854 160
rect 43166 -300 43222 160
rect 43534 -300 43590 160
rect 43902 -300 43958 160
rect 44270 -300 44326 160
rect 44638 -300 44694 160
rect 45006 -300 45062 160
rect 45374 -300 45430 160
rect 45742 -300 45798 160
rect 46110 -300 46166 160
<< obsm2 >>
rect 204 44484 422 44554
rect 590 44484 790 44554
rect 958 44484 1158 44554
rect 1326 44484 1526 44554
rect 1694 44484 1894 44554
rect 2062 44484 2262 44554
rect 2430 44484 2630 44554
rect 2798 44484 2998 44554
rect 3166 44484 3366 44554
rect 3534 44484 3734 44554
rect 3902 44484 4102 44554
rect 4270 44484 4470 44554
rect 4638 44484 4838 44554
rect 5006 44484 5206 44554
rect 5374 44484 5574 44554
rect 5742 44484 5942 44554
rect 6110 44484 6310 44554
rect 6478 44484 6678 44554
rect 6846 44484 7046 44554
rect 7214 44484 7414 44554
rect 7582 44484 7782 44554
rect 7950 44484 8150 44554
rect 8318 44484 8518 44554
rect 8686 44484 8886 44554
rect 9054 44484 9254 44554
rect 9422 44484 9622 44554
rect 9790 44484 9990 44554
rect 10158 44484 10358 44554
rect 10526 44484 10726 44554
rect 10894 44484 11094 44554
rect 11262 44484 11462 44554
rect 11630 44484 11830 44554
rect 11998 44484 12198 44554
rect 12366 44484 12566 44554
rect 12734 44484 12934 44554
rect 13102 44484 13302 44554
rect 13470 44484 13670 44554
rect 13838 44484 14038 44554
rect 14206 44484 14406 44554
rect 14574 44484 14774 44554
rect 14942 44484 15142 44554
rect 15310 44484 15510 44554
rect 15678 44484 15878 44554
rect 16046 44484 16246 44554
rect 16414 44484 16614 44554
rect 16782 44484 16982 44554
rect 17150 44484 17350 44554
rect 17518 44484 17718 44554
rect 17886 44484 18086 44554
rect 18254 44484 18454 44554
rect 18622 44484 18822 44554
rect 18990 44484 19190 44554
rect 19358 44484 19558 44554
rect 19726 44484 19926 44554
rect 20094 44484 20294 44554
rect 20462 44484 20662 44554
rect 20830 44484 21030 44554
rect 21198 44484 21398 44554
rect 21566 44484 21766 44554
rect 21934 44484 22134 44554
rect 22302 44484 22502 44554
rect 22670 44484 22870 44554
rect 23038 44484 23238 44554
rect 23406 44484 23606 44554
rect 23774 44484 23974 44554
rect 24142 44484 24342 44554
rect 24510 44484 24710 44554
rect 24878 44484 25078 44554
rect 25246 44484 25446 44554
rect 25614 44484 25814 44554
rect 25982 44484 26182 44554
rect 26350 44484 26550 44554
rect 26718 44484 26918 44554
rect 27086 44484 27286 44554
rect 27454 44484 27654 44554
rect 27822 44484 28022 44554
rect 28190 44484 28390 44554
rect 28558 44484 28758 44554
rect 28926 44484 29126 44554
rect 29294 44484 29494 44554
rect 29662 44484 29862 44554
rect 30030 44484 30230 44554
rect 30398 44484 30598 44554
rect 30766 44484 30966 44554
rect 31134 44484 31334 44554
rect 31502 44484 31702 44554
rect 31870 44484 32070 44554
rect 32238 44484 32438 44554
rect 32606 44484 32806 44554
rect 32974 44484 33174 44554
rect 33342 44484 33542 44554
rect 33710 44484 33910 44554
rect 34078 44484 34278 44554
rect 34446 44484 34646 44554
rect 34814 44484 35014 44554
rect 35182 44484 35382 44554
rect 35550 44484 35750 44554
rect 35918 44484 36118 44554
rect 36286 44484 36486 44554
rect 36654 44484 36854 44554
rect 37022 44484 37222 44554
rect 37390 44484 37590 44554
rect 37758 44484 37958 44554
rect 38126 44484 38326 44554
rect 38494 44484 38694 44554
rect 38862 44484 39062 44554
rect 39230 44484 39430 44554
rect 39598 44484 39798 44554
rect 39966 44484 40166 44554
rect 40334 44484 40534 44554
rect 40702 44484 40902 44554
rect 41070 44484 41270 44554
rect 41438 44484 41638 44554
rect 41806 44484 42006 44554
rect 42174 44484 42374 44554
rect 42542 44484 42742 44554
rect 42910 44484 43110 44554
rect 43278 44484 43478 44554
rect 43646 44484 43846 44554
rect 44014 44484 44214 44554
rect 44382 44484 44582 44554
rect 44750 44484 44950 44554
rect 45118 44484 45318 44554
rect 45486 44484 45686 44554
rect 45854 44484 46054 44554
rect 46222 44484 46626 44554
rect 204 216 46626 44484
rect 204 54 422 216
rect 590 54 790 216
rect 958 54 1158 216
rect 1326 54 1526 216
rect 1694 54 1894 216
rect 2062 54 2262 216
rect 2430 54 2630 216
rect 2798 54 2998 216
rect 3166 54 3366 216
rect 3534 54 3734 216
rect 3902 54 4102 216
rect 4270 54 4470 216
rect 4638 54 4838 216
rect 5006 54 5206 216
rect 5374 54 5574 216
rect 5742 54 5942 216
rect 6110 54 6310 216
rect 6478 54 6678 216
rect 6846 54 7046 216
rect 7214 54 7414 216
rect 7582 54 7782 216
rect 7950 54 8150 216
rect 8318 54 8518 216
rect 8686 54 8886 216
rect 9054 54 9254 216
rect 9422 54 9622 216
rect 9790 54 9990 216
rect 10158 54 10358 216
rect 10526 54 10726 216
rect 10894 54 11094 216
rect 11262 54 11462 216
rect 11630 54 11830 216
rect 11998 54 12198 216
rect 12366 54 12566 216
rect 12734 54 12934 216
rect 13102 54 13302 216
rect 13470 54 13670 216
rect 13838 54 14038 216
rect 14206 54 14406 216
rect 14574 54 14774 216
rect 14942 54 15142 216
rect 15310 54 15510 216
rect 15678 54 15878 216
rect 16046 54 16246 216
rect 16414 54 16614 216
rect 16782 54 16982 216
rect 17150 54 17350 216
rect 17518 54 17718 216
rect 17886 54 18086 216
rect 18254 54 18454 216
rect 18622 54 18822 216
rect 18990 54 19190 216
rect 19358 54 19558 216
rect 19726 54 19926 216
rect 20094 54 20294 216
rect 20462 54 20662 216
rect 20830 54 21030 216
rect 21198 54 21398 216
rect 21566 54 21766 216
rect 21934 54 22134 216
rect 22302 54 22502 216
rect 22670 54 22870 216
rect 23038 54 23238 216
rect 23406 54 23606 216
rect 23774 54 23974 216
rect 24142 54 24342 216
rect 24510 54 24710 216
rect 24878 54 25078 216
rect 25246 54 25446 216
rect 25614 54 25814 216
rect 25982 54 26182 216
rect 26350 54 26550 216
rect 26718 54 26918 216
rect 27086 54 27286 216
rect 27454 54 27654 216
rect 27822 54 28022 216
rect 28190 54 28390 216
rect 28558 54 28758 216
rect 28926 54 29126 216
rect 29294 54 29494 216
rect 29662 54 29862 216
rect 30030 54 30230 216
rect 30398 54 30598 216
rect 30766 54 30966 216
rect 31134 54 31334 216
rect 31502 54 31702 216
rect 31870 54 32070 216
rect 32238 54 32438 216
rect 32606 54 32806 216
rect 32974 54 33174 216
rect 33342 54 33542 216
rect 33710 54 33910 216
rect 34078 54 34278 216
rect 34446 54 34646 216
rect 34814 54 35014 216
rect 35182 54 35382 216
rect 35550 54 35750 216
rect 35918 54 36118 216
rect 36286 54 36486 216
rect 36654 54 36854 216
rect 37022 54 37222 216
rect 37390 54 37590 216
rect 37758 54 37958 216
rect 38126 54 38326 216
rect 38494 54 38694 216
rect 38862 54 39062 216
rect 39230 54 39430 216
rect 39598 54 39798 216
rect 39966 54 40166 216
rect 40334 54 40534 216
rect 40702 54 40902 216
rect 41070 54 41270 216
rect 41438 54 41638 216
rect 41806 54 42006 216
rect 42174 54 42374 216
rect 42542 54 42742 216
rect 42910 54 43110 216
rect 43278 54 43478 216
rect 43646 54 43846 216
rect 44014 54 44214 216
rect 44382 54 44582 216
rect 44750 54 44950 216
rect 45118 54 45318 216
rect 45486 54 45686 216
rect 45854 54 46054 216
rect 46222 54 46626 216
<< metal3 >>
rect -300 39448 160 39568
rect -300 39176 160 39296
rect -300 38904 160 39024
rect -300 38632 160 38752
rect -300 38360 160 38480
rect -300 38088 160 38208
rect -300 37816 160 37936
rect -300 37544 160 37664
rect -300 37272 160 37392
rect -300 37000 160 37120
rect -300 36728 160 36848
rect -300 36456 160 36576
rect -300 36184 160 36304
rect -300 35912 160 36032
rect -300 35640 160 35760
rect -300 35368 160 35488
rect -300 35096 160 35216
rect -300 34824 160 34944
rect -300 34552 160 34672
rect -300 34280 160 34400
rect -300 34008 160 34128
rect -300 33736 160 33856
rect -300 33464 160 33584
rect -300 33192 160 33312
rect -300 32920 160 33040
rect -300 32648 160 32768
rect -300 32376 160 32496
rect -300 32104 160 32224
rect -300 31832 160 31952
rect -300 31560 160 31680
rect -300 31288 160 31408
rect -300 31016 160 31136
rect -300 30744 160 30864
rect -300 30472 160 30592
rect -300 30200 160 30320
rect -300 29928 160 30048
rect -300 29656 160 29776
rect -300 29384 160 29504
rect -300 29112 160 29232
rect -300 28840 160 28960
rect -300 28568 160 28688
rect -300 28296 160 28416
rect -300 28024 160 28144
rect -300 27752 160 27872
rect -300 27480 160 27600
rect -300 27208 160 27328
rect -300 26936 160 27056
rect -300 26664 160 26784
rect -300 26392 160 26512
rect -300 26120 160 26240
rect -300 25848 160 25968
rect -300 25576 160 25696
rect -300 25304 160 25424
rect -300 25032 160 25152
rect -300 24760 160 24880
rect -300 24488 160 24608
rect -300 24216 160 24336
rect -300 23944 160 24064
rect -300 23672 160 23792
rect -300 23400 160 23520
rect -300 23128 160 23248
rect -300 22856 160 22976
rect -300 22584 160 22704
rect -300 22312 160 22432
rect -300 22040 160 22160
rect -300 21768 160 21888
rect -300 21496 160 21616
rect -300 21224 160 21344
rect -300 20952 160 21072
rect -300 20680 160 20800
rect -300 20408 160 20528
rect -300 20136 160 20256
rect -300 19864 160 19984
rect -300 19592 160 19712
rect -300 19320 160 19440
rect -300 19048 160 19168
rect -300 18776 160 18896
rect -300 18504 160 18624
rect -300 18232 160 18352
rect -300 17960 160 18080
rect -300 17688 160 17808
rect -300 17416 160 17536
rect -300 17144 160 17264
rect -300 16872 160 16992
rect -300 16600 160 16720
rect -300 16328 160 16448
rect -300 16056 160 16176
rect -300 15784 160 15904
rect -300 15512 160 15632
rect -300 15240 160 15360
rect -300 14968 160 15088
rect -300 14696 160 14816
rect -300 14424 160 14544
rect -300 14152 160 14272
rect -300 13880 160 14000
rect -300 13608 160 13728
rect -300 13336 160 13456
rect -300 13064 160 13184
rect -300 12792 160 12912
rect -300 12520 160 12640
rect -300 12248 160 12368
rect -300 11976 160 12096
rect -300 11704 160 11824
rect -300 11432 160 11552
rect -300 11160 160 11280
rect -300 10888 160 11008
rect -300 10616 160 10736
rect -300 10344 160 10464
rect -300 10072 160 10192
rect -300 9800 160 9920
rect -300 9528 160 9648
rect -300 9256 160 9376
rect -300 8984 160 9104
rect -300 8712 160 8832
rect -300 8440 160 8560
rect -300 8168 160 8288
rect -300 7896 160 8016
rect -300 7624 160 7744
rect -300 7352 160 7472
rect -300 7080 160 7200
rect -300 6808 160 6928
rect -300 6536 160 6656
rect -300 6264 160 6384
rect -300 5992 160 6112
rect -300 5720 160 5840
rect -300 5448 160 5568
rect -300 5176 160 5296
rect -300 4904 160 5024
rect 46540 39448 47000 39568
rect 46540 39176 47000 39296
rect 46540 38904 47000 39024
rect 46540 38632 47000 38752
rect 46540 38360 47000 38480
rect 46540 38088 47000 38208
rect 46540 37816 47000 37936
rect 46540 37544 47000 37664
rect 46540 37272 47000 37392
rect 46540 37000 47000 37120
rect 46540 36728 47000 36848
rect 46540 36456 47000 36576
rect 46540 36184 47000 36304
rect 46540 35912 47000 36032
rect 46540 35640 47000 35760
rect 46540 35368 47000 35488
rect 46540 35096 47000 35216
rect 46540 34824 47000 34944
rect 46540 34552 47000 34672
rect 46540 34280 47000 34400
rect 46540 34008 47000 34128
rect 46540 33736 47000 33856
rect 46540 33464 47000 33584
rect 46540 33192 47000 33312
rect 46540 32920 47000 33040
rect 46540 32648 47000 32768
rect 46540 32376 47000 32496
rect 46540 32104 47000 32224
rect 46540 31832 47000 31952
rect 46540 31560 47000 31680
rect 46540 31288 47000 31408
rect 46540 31016 47000 31136
rect 46540 30744 47000 30864
rect 46540 30472 47000 30592
rect 46540 30200 47000 30320
rect 46540 29928 47000 30048
rect 46540 29656 47000 29776
rect 46540 29384 47000 29504
rect 46540 29112 47000 29232
rect 46540 28840 47000 28960
rect 46540 28568 47000 28688
rect 46540 28296 47000 28416
rect 46540 28024 47000 28144
rect 46540 27752 47000 27872
rect 46540 27480 47000 27600
rect 46540 27208 47000 27328
rect 46540 26936 47000 27056
rect 46540 26664 47000 26784
rect 46540 26392 47000 26512
rect 46540 26120 47000 26240
rect 46540 25848 47000 25968
rect 46540 25576 47000 25696
rect 46540 25304 47000 25424
rect 46540 25032 47000 25152
rect 46540 24760 47000 24880
rect 46540 24488 47000 24608
rect 46540 24216 47000 24336
rect 46540 23944 47000 24064
rect 46540 23672 47000 23792
rect 46540 23400 47000 23520
rect 46540 23128 47000 23248
rect 46540 22856 47000 22976
rect 46540 22584 47000 22704
rect 46540 22312 47000 22432
rect 46540 22040 47000 22160
rect 46540 21768 47000 21888
rect 46540 21496 47000 21616
rect 46540 21224 47000 21344
rect 46540 20952 47000 21072
rect 46540 20680 47000 20800
rect 46540 20408 47000 20528
rect 46540 20136 47000 20256
rect 46540 19864 47000 19984
rect 46540 19592 47000 19712
rect 46540 19320 47000 19440
rect 46540 19048 47000 19168
rect 46540 18776 47000 18896
rect 46540 18504 47000 18624
rect 46540 18232 47000 18352
rect 46540 17960 47000 18080
rect 46540 17688 47000 17808
rect 46540 17416 47000 17536
rect 46540 17144 47000 17264
rect 46540 16872 47000 16992
rect 46540 16600 47000 16720
rect 46540 16328 47000 16448
rect 46540 16056 47000 16176
rect 46540 15784 47000 15904
rect 46540 15512 47000 15632
rect 46540 15240 47000 15360
rect 46540 14968 47000 15088
rect 46540 14696 47000 14816
rect 46540 14424 47000 14544
rect 46540 14152 47000 14272
rect 46540 13880 47000 14000
rect 46540 13608 47000 13728
rect 46540 13336 47000 13456
rect 46540 13064 47000 13184
rect 46540 12792 47000 12912
rect 46540 12520 47000 12640
rect 46540 12248 47000 12368
rect 46540 11976 47000 12096
rect 46540 11704 47000 11824
rect 46540 11432 47000 11552
rect 46540 11160 47000 11280
rect 46540 10888 47000 11008
rect 46540 10616 47000 10736
rect 46540 10344 47000 10464
rect 46540 10072 47000 10192
rect 46540 9800 47000 9920
rect 46540 9528 47000 9648
rect 46540 9256 47000 9376
rect 46540 8984 47000 9104
rect 46540 8712 47000 8832
rect 46540 8440 47000 8560
rect 46540 8168 47000 8288
rect 46540 7896 47000 8016
rect 46540 7624 47000 7744
rect 46540 7352 47000 7472
rect 46540 7080 47000 7200
rect 46540 6808 47000 6928
rect 46540 6536 47000 6656
rect 46540 6264 47000 6384
rect 46540 5992 47000 6112
rect 46540 5720 47000 5840
rect 46540 5448 47000 5568
rect 46540 5176 47000 5296
rect 46540 4904 47000 5024
<< obsm3 >>
rect 160 39648 46631 43553
rect 240 4824 46460 39648
rect 160 851 46631 4824
<< metal4 >>
rect 4208 1040 4528 43568
rect 19568 1040 19888 43568
rect 34928 1040 35248 43568
<< obsm4 >>
rect 611 960 4128 42941
rect 4608 960 19488 42941
rect 19968 960 34848 42941
rect 35328 960 45573 42941
rect 611 851 45573 960
<< labels >>
rlabel metal3 s 46540 17960 47000 18080 6 E1BEG[0]
port 1 nsew signal output
rlabel metal3 s 46540 18232 47000 18352 6 E1BEG[1]
port 2 nsew signal output
rlabel metal3 s 46540 18504 47000 18624 6 E1BEG[2]
port 3 nsew signal output
rlabel metal3 s 46540 18776 47000 18896 6 E1BEG[3]
port 4 nsew signal output
rlabel metal3 s -300 17960 160 18080 4 E1END[0]
port 5 nsew signal input
rlabel metal3 s -300 18232 160 18352 4 E1END[1]
port 6 nsew signal input
rlabel metal3 s -300 18504 160 18624 4 E1END[2]
port 7 nsew signal input
rlabel metal3 s -300 18776 160 18896 4 E1END[3]
port 8 nsew signal input
rlabel metal3 s 46540 19048 47000 19168 6 E2BEG[0]
port 9 nsew signal output
rlabel metal3 s 46540 19320 47000 19440 6 E2BEG[1]
port 10 nsew signal output
rlabel metal3 s 46540 19592 47000 19712 6 E2BEG[2]
port 11 nsew signal output
rlabel metal3 s 46540 19864 47000 19984 6 E2BEG[3]
port 12 nsew signal output
rlabel metal3 s 46540 20136 47000 20256 6 E2BEG[4]
port 13 nsew signal output
rlabel metal3 s 46540 20408 47000 20528 6 E2BEG[5]
port 14 nsew signal output
rlabel metal3 s 46540 20680 47000 20800 6 E2BEG[6]
port 15 nsew signal output
rlabel metal3 s 46540 20952 47000 21072 6 E2BEG[7]
port 16 nsew signal output
rlabel metal3 s 46540 21224 47000 21344 6 E2BEGb[0]
port 17 nsew signal output
rlabel metal3 s 46540 21496 47000 21616 6 E2BEGb[1]
port 18 nsew signal output
rlabel metal3 s 46540 21768 47000 21888 6 E2BEGb[2]
port 19 nsew signal output
rlabel metal3 s 46540 22040 47000 22160 6 E2BEGb[3]
port 20 nsew signal output
rlabel metal3 s 46540 22312 47000 22432 6 E2BEGb[4]
port 21 nsew signal output
rlabel metal3 s 46540 22584 47000 22704 6 E2BEGb[5]
port 22 nsew signal output
rlabel metal3 s 46540 22856 47000 22976 6 E2BEGb[6]
port 23 nsew signal output
rlabel metal3 s 46540 23128 47000 23248 6 E2BEGb[7]
port 24 nsew signal output
rlabel metal3 s -300 21224 160 21344 4 E2END[0]
port 25 nsew signal input
rlabel metal3 s -300 21496 160 21616 4 E2END[1]
port 26 nsew signal input
rlabel metal3 s -300 21768 160 21888 4 E2END[2]
port 27 nsew signal input
rlabel metal3 s -300 22040 160 22160 4 E2END[3]
port 28 nsew signal input
rlabel metal3 s -300 22312 160 22432 4 E2END[4]
port 29 nsew signal input
rlabel metal3 s -300 22584 160 22704 4 E2END[5]
port 30 nsew signal input
rlabel metal3 s -300 22856 160 22976 4 E2END[6]
port 31 nsew signal input
rlabel metal3 s -300 23128 160 23248 4 E2END[7]
port 32 nsew signal input
rlabel metal3 s -300 19048 160 19168 4 E2MID[0]
port 33 nsew signal input
rlabel metal3 s -300 19320 160 19440 4 E2MID[1]
port 34 nsew signal input
rlabel metal3 s -300 19592 160 19712 4 E2MID[2]
port 35 nsew signal input
rlabel metal3 s -300 19864 160 19984 4 E2MID[3]
port 36 nsew signal input
rlabel metal3 s -300 20136 160 20256 4 E2MID[4]
port 37 nsew signal input
rlabel metal3 s -300 20408 160 20528 4 E2MID[5]
port 38 nsew signal input
rlabel metal3 s -300 20680 160 20800 4 E2MID[6]
port 39 nsew signal input
rlabel metal3 s -300 20952 160 21072 4 E2MID[7]
port 40 nsew signal input
rlabel metal3 s 46540 27752 47000 27872 6 E6BEG[0]
port 41 nsew signal output
rlabel metal3 s 46540 30472 47000 30592 6 E6BEG[10]
port 42 nsew signal output
rlabel metal3 s 46540 30744 47000 30864 6 E6BEG[11]
port 43 nsew signal output
rlabel metal3 s 46540 28024 47000 28144 6 E6BEG[1]
port 44 nsew signal output
rlabel metal3 s 46540 28296 47000 28416 6 E6BEG[2]
port 45 nsew signal output
rlabel metal3 s 46540 28568 47000 28688 6 E6BEG[3]
port 46 nsew signal output
rlabel metal3 s 46540 28840 47000 28960 6 E6BEG[4]
port 47 nsew signal output
rlabel metal3 s 46540 29112 47000 29232 6 E6BEG[5]
port 48 nsew signal output
rlabel metal3 s 46540 29384 47000 29504 6 E6BEG[6]
port 49 nsew signal output
rlabel metal3 s 46540 29656 47000 29776 6 E6BEG[7]
port 50 nsew signal output
rlabel metal3 s 46540 29928 47000 30048 6 E6BEG[8]
port 51 nsew signal output
rlabel metal3 s 46540 30200 47000 30320 6 E6BEG[9]
port 52 nsew signal output
rlabel metal3 s -300 27752 160 27872 4 E6END[0]
port 53 nsew signal input
rlabel metal3 s -300 30472 160 30592 4 E6END[10]
port 54 nsew signal input
rlabel metal3 s -300 30744 160 30864 4 E6END[11]
port 55 nsew signal input
rlabel metal3 s -300 28024 160 28144 4 E6END[1]
port 56 nsew signal input
rlabel metal3 s -300 28296 160 28416 4 E6END[2]
port 57 nsew signal input
rlabel metal3 s -300 28568 160 28688 4 E6END[3]
port 58 nsew signal input
rlabel metal3 s -300 28840 160 28960 4 E6END[4]
port 59 nsew signal input
rlabel metal3 s -300 29112 160 29232 4 E6END[5]
port 60 nsew signal input
rlabel metal3 s -300 29384 160 29504 4 E6END[6]
port 61 nsew signal input
rlabel metal3 s -300 29656 160 29776 4 E6END[7]
port 62 nsew signal input
rlabel metal3 s -300 29928 160 30048 4 E6END[8]
port 63 nsew signal input
rlabel metal3 s -300 30200 160 30320 4 E6END[9]
port 64 nsew signal input
rlabel metal3 s 46540 23400 47000 23520 6 EE4BEG[0]
port 65 nsew signal output
rlabel metal3 s 46540 26120 47000 26240 6 EE4BEG[10]
port 66 nsew signal output
rlabel metal3 s 46540 26392 47000 26512 6 EE4BEG[11]
port 67 nsew signal output
rlabel metal3 s 46540 26664 47000 26784 6 EE4BEG[12]
port 68 nsew signal output
rlabel metal3 s 46540 26936 47000 27056 6 EE4BEG[13]
port 69 nsew signal output
rlabel metal3 s 46540 27208 47000 27328 6 EE4BEG[14]
port 70 nsew signal output
rlabel metal3 s 46540 27480 47000 27600 6 EE4BEG[15]
port 71 nsew signal output
rlabel metal3 s 46540 23672 47000 23792 6 EE4BEG[1]
port 72 nsew signal output
rlabel metal3 s 46540 23944 47000 24064 6 EE4BEG[2]
port 73 nsew signal output
rlabel metal3 s 46540 24216 47000 24336 6 EE4BEG[3]
port 74 nsew signal output
rlabel metal3 s 46540 24488 47000 24608 6 EE4BEG[4]
port 75 nsew signal output
rlabel metal3 s 46540 24760 47000 24880 6 EE4BEG[5]
port 76 nsew signal output
rlabel metal3 s 46540 25032 47000 25152 6 EE4BEG[6]
port 77 nsew signal output
rlabel metal3 s 46540 25304 47000 25424 6 EE4BEG[7]
port 78 nsew signal output
rlabel metal3 s 46540 25576 47000 25696 6 EE4BEG[8]
port 79 nsew signal output
rlabel metal3 s 46540 25848 47000 25968 6 EE4BEG[9]
port 80 nsew signal output
rlabel metal3 s -300 23400 160 23520 4 EE4END[0]
port 81 nsew signal input
rlabel metal3 s -300 26120 160 26240 4 EE4END[10]
port 82 nsew signal input
rlabel metal3 s -300 26392 160 26512 4 EE4END[11]
port 83 nsew signal input
rlabel metal3 s -300 26664 160 26784 4 EE4END[12]
port 84 nsew signal input
rlabel metal3 s -300 26936 160 27056 4 EE4END[13]
port 85 nsew signal input
rlabel metal3 s -300 27208 160 27328 4 EE4END[14]
port 86 nsew signal input
rlabel metal3 s -300 27480 160 27600 4 EE4END[15]
port 87 nsew signal input
rlabel metal3 s -300 23672 160 23792 4 EE4END[1]
port 88 nsew signal input
rlabel metal3 s -300 23944 160 24064 4 EE4END[2]
port 89 nsew signal input
rlabel metal3 s -300 24216 160 24336 4 EE4END[3]
port 90 nsew signal input
rlabel metal3 s -300 24488 160 24608 4 EE4END[4]
port 91 nsew signal input
rlabel metal3 s -300 24760 160 24880 4 EE4END[5]
port 92 nsew signal input
rlabel metal3 s -300 25032 160 25152 4 EE4END[6]
port 93 nsew signal input
rlabel metal3 s -300 25304 160 25424 4 EE4END[7]
port 94 nsew signal input
rlabel metal3 s -300 25576 160 25696 4 EE4END[8]
port 95 nsew signal input
rlabel metal3 s -300 25848 160 25968 4 EE4END[9]
port 96 nsew signal input
rlabel metal3 s -300 31016 160 31136 4 FrameData[0]
port 97 nsew signal input
rlabel metal3 s -300 33736 160 33856 4 FrameData[10]
port 98 nsew signal input
rlabel metal3 s -300 34008 160 34128 4 FrameData[11]
port 99 nsew signal input
rlabel metal3 s -300 34280 160 34400 4 FrameData[12]
port 100 nsew signal input
rlabel metal3 s -300 34552 160 34672 4 FrameData[13]
port 101 nsew signal input
rlabel metal3 s -300 34824 160 34944 4 FrameData[14]
port 102 nsew signal input
rlabel metal3 s -300 35096 160 35216 4 FrameData[15]
port 103 nsew signal input
rlabel metal3 s -300 35368 160 35488 4 FrameData[16]
port 104 nsew signal input
rlabel metal3 s -300 35640 160 35760 4 FrameData[17]
port 105 nsew signal input
rlabel metal3 s -300 35912 160 36032 4 FrameData[18]
port 106 nsew signal input
rlabel metal3 s -300 36184 160 36304 4 FrameData[19]
port 107 nsew signal input
rlabel metal3 s -300 31288 160 31408 4 FrameData[1]
port 108 nsew signal input
rlabel metal3 s -300 36456 160 36576 4 FrameData[20]
port 109 nsew signal input
rlabel metal3 s -300 36728 160 36848 4 FrameData[21]
port 110 nsew signal input
rlabel metal3 s -300 37000 160 37120 4 FrameData[22]
port 111 nsew signal input
rlabel metal3 s -300 37272 160 37392 4 FrameData[23]
port 112 nsew signal input
rlabel metal3 s -300 37544 160 37664 4 FrameData[24]
port 113 nsew signal input
rlabel metal3 s -300 37816 160 37936 4 FrameData[25]
port 114 nsew signal input
rlabel metal3 s -300 38088 160 38208 4 FrameData[26]
port 115 nsew signal input
rlabel metal3 s -300 38360 160 38480 4 FrameData[27]
port 116 nsew signal input
rlabel metal3 s -300 38632 160 38752 4 FrameData[28]
port 117 nsew signal input
rlabel metal3 s -300 38904 160 39024 4 FrameData[29]
port 118 nsew signal input
rlabel metal3 s -300 31560 160 31680 4 FrameData[2]
port 119 nsew signal input
rlabel metal3 s -300 39176 160 39296 4 FrameData[30]
port 120 nsew signal input
rlabel metal3 s -300 39448 160 39568 4 FrameData[31]
port 121 nsew signal input
rlabel metal3 s -300 31832 160 31952 4 FrameData[3]
port 122 nsew signal input
rlabel metal3 s -300 32104 160 32224 4 FrameData[4]
port 123 nsew signal input
rlabel metal3 s -300 32376 160 32496 4 FrameData[5]
port 124 nsew signal input
rlabel metal3 s -300 32648 160 32768 4 FrameData[6]
port 125 nsew signal input
rlabel metal3 s -300 32920 160 33040 4 FrameData[7]
port 126 nsew signal input
rlabel metal3 s -300 33192 160 33312 4 FrameData[8]
port 127 nsew signal input
rlabel metal3 s -300 33464 160 33584 4 FrameData[9]
port 128 nsew signal input
rlabel metal3 s 46540 31016 47000 31136 6 FrameData_O[0]
port 129 nsew signal output
rlabel metal3 s 46540 33736 47000 33856 6 FrameData_O[10]
port 130 nsew signal output
rlabel metal3 s 46540 34008 47000 34128 6 FrameData_O[11]
port 131 nsew signal output
rlabel metal3 s 46540 34280 47000 34400 6 FrameData_O[12]
port 132 nsew signal output
rlabel metal3 s 46540 34552 47000 34672 6 FrameData_O[13]
port 133 nsew signal output
rlabel metal3 s 46540 34824 47000 34944 6 FrameData_O[14]
port 134 nsew signal output
rlabel metal3 s 46540 35096 47000 35216 6 FrameData_O[15]
port 135 nsew signal output
rlabel metal3 s 46540 35368 47000 35488 6 FrameData_O[16]
port 136 nsew signal output
rlabel metal3 s 46540 35640 47000 35760 6 FrameData_O[17]
port 137 nsew signal output
rlabel metal3 s 46540 35912 47000 36032 6 FrameData_O[18]
port 138 nsew signal output
rlabel metal3 s 46540 36184 47000 36304 6 FrameData_O[19]
port 139 nsew signal output
rlabel metal3 s 46540 31288 47000 31408 6 FrameData_O[1]
port 140 nsew signal output
rlabel metal3 s 46540 36456 47000 36576 6 FrameData_O[20]
port 141 nsew signal output
rlabel metal3 s 46540 36728 47000 36848 6 FrameData_O[21]
port 142 nsew signal output
rlabel metal3 s 46540 37000 47000 37120 6 FrameData_O[22]
port 143 nsew signal output
rlabel metal3 s 46540 37272 47000 37392 6 FrameData_O[23]
port 144 nsew signal output
rlabel metal3 s 46540 37544 47000 37664 6 FrameData_O[24]
port 145 nsew signal output
rlabel metal3 s 46540 37816 47000 37936 6 FrameData_O[25]
port 146 nsew signal output
rlabel metal3 s 46540 38088 47000 38208 6 FrameData_O[26]
port 147 nsew signal output
rlabel metal3 s 46540 38360 47000 38480 6 FrameData_O[27]
port 148 nsew signal output
rlabel metal3 s 46540 38632 47000 38752 6 FrameData_O[28]
port 149 nsew signal output
rlabel metal3 s 46540 38904 47000 39024 6 FrameData_O[29]
port 150 nsew signal output
rlabel metal3 s 46540 31560 47000 31680 6 FrameData_O[2]
port 151 nsew signal output
rlabel metal3 s 46540 39176 47000 39296 6 FrameData_O[30]
port 152 nsew signal output
rlabel metal3 s 46540 39448 47000 39568 6 FrameData_O[31]
port 153 nsew signal output
rlabel metal3 s 46540 31832 47000 31952 6 FrameData_O[3]
port 154 nsew signal output
rlabel metal3 s 46540 32104 47000 32224 6 FrameData_O[4]
port 155 nsew signal output
rlabel metal3 s 46540 32376 47000 32496 6 FrameData_O[5]
port 156 nsew signal output
rlabel metal3 s 46540 32648 47000 32768 6 FrameData_O[6]
port 157 nsew signal output
rlabel metal3 s 46540 32920 47000 33040 6 FrameData_O[7]
port 158 nsew signal output
rlabel metal3 s 46540 33192 47000 33312 6 FrameData_O[8]
port 159 nsew signal output
rlabel metal3 s 46540 33464 47000 33584 6 FrameData_O[9]
port 160 nsew signal output
rlabel metal2 s 39118 -300 39174 160 8 FrameStrobe[0]
port 161 nsew signal input
rlabel metal2 s 42798 -300 42854 160 8 FrameStrobe[10]
port 162 nsew signal input
rlabel metal2 s 43166 -300 43222 160 8 FrameStrobe[11]
port 163 nsew signal input
rlabel metal2 s 43534 -300 43590 160 8 FrameStrobe[12]
port 164 nsew signal input
rlabel metal2 s 43902 -300 43958 160 8 FrameStrobe[13]
port 165 nsew signal input
rlabel metal2 s 44270 -300 44326 160 8 FrameStrobe[14]
port 166 nsew signal input
rlabel metal2 s 44638 -300 44694 160 8 FrameStrobe[15]
port 167 nsew signal input
rlabel metal2 s 45006 -300 45062 160 8 FrameStrobe[16]
port 168 nsew signal input
rlabel metal2 s 45374 -300 45430 160 8 FrameStrobe[17]
port 169 nsew signal input
rlabel metal2 s 45742 -300 45798 160 8 FrameStrobe[18]
port 170 nsew signal input
rlabel metal2 s 46110 -300 46166 160 8 FrameStrobe[19]
port 171 nsew signal input
rlabel metal2 s 39486 -300 39542 160 8 FrameStrobe[1]
port 172 nsew signal input
rlabel metal2 s 39854 -300 39910 160 8 FrameStrobe[2]
port 173 nsew signal input
rlabel metal2 s 40222 -300 40278 160 8 FrameStrobe[3]
port 174 nsew signal input
rlabel metal2 s 40590 -300 40646 160 8 FrameStrobe[4]
port 175 nsew signal input
rlabel metal2 s 40958 -300 41014 160 8 FrameStrobe[5]
port 176 nsew signal input
rlabel metal2 s 41326 -300 41382 160 8 FrameStrobe[6]
port 177 nsew signal input
rlabel metal2 s 41694 -300 41750 160 8 FrameStrobe[7]
port 178 nsew signal input
rlabel metal2 s 42062 -300 42118 160 8 FrameStrobe[8]
port 179 nsew signal input
rlabel metal2 s 42430 -300 42486 160 8 FrameStrobe[9]
port 180 nsew signal input
rlabel metal2 s 39118 44540 39174 45000 6 FrameStrobe_O[0]
port 181 nsew signal output
rlabel metal2 s 42798 44540 42854 45000 6 FrameStrobe_O[10]
port 182 nsew signal output
rlabel metal2 s 43166 44540 43222 45000 6 FrameStrobe_O[11]
port 183 nsew signal output
rlabel metal2 s 43534 44540 43590 45000 6 FrameStrobe_O[12]
port 184 nsew signal output
rlabel metal2 s 43902 44540 43958 45000 6 FrameStrobe_O[13]
port 185 nsew signal output
rlabel metal2 s 44270 44540 44326 45000 6 FrameStrobe_O[14]
port 186 nsew signal output
rlabel metal2 s 44638 44540 44694 45000 6 FrameStrobe_O[15]
port 187 nsew signal output
rlabel metal2 s 45006 44540 45062 45000 6 FrameStrobe_O[16]
port 188 nsew signal output
rlabel metal2 s 45374 44540 45430 45000 6 FrameStrobe_O[17]
port 189 nsew signal output
rlabel metal2 s 45742 44540 45798 45000 6 FrameStrobe_O[18]
port 190 nsew signal output
rlabel metal2 s 46110 44540 46166 45000 6 FrameStrobe_O[19]
port 191 nsew signal output
rlabel metal2 s 39486 44540 39542 45000 6 FrameStrobe_O[1]
port 192 nsew signal output
rlabel metal2 s 39854 44540 39910 45000 6 FrameStrobe_O[2]
port 193 nsew signal output
rlabel metal2 s 40222 44540 40278 45000 6 FrameStrobe_O[3]
port 194 nsew signal output
rlabel metal2 s 40590 44540 40646 45000 6 FrameStrobe_O[4]
port 195 nsew signal output
rlabel metal2 s 40958 44540 41014 45000 6 FrameStrobe_O[5]
port 196 nsew signal output
rlabel metal2 s 41326 44540 41382 45000 6 FrameStrobe_O[6]
port 197 nsew signal output
rlabel metal2 s 41694 44540 41750 45000 6 FrameStrobe_O[7]
port 198 nsew signal output
rlabel metal2 s 42062 44540 42118 45000 6 FrameStrobe_O[8]
port 199 nsew signal output
rlabel metal2 s 42430 44540 42486 45000 6 FrameStrobe_O[9]
port 200 nsew signal output
rlabel metal2 s 478 44540 534 45000 6 N1BEG[0]
port 201 nsew signal output
rlabel metal2 s 846 44540 902 45000 6 N1BEG[1]
port 202 nsew signal output
rlabel metal2 s 1214 44540 1270 45000 6 N1BEG[2]
port 203 nsew signal output
rlabel metal2 s 1582 44540 1638 45000 6 N1BEG[3]
port 204 nsew signal output
rlabel metal2 s 478 -300 534 160 8 N1END[0]
port 205 nsew signal input
rlabel metal2 s 846 -300 902 160 8 N1END[1]
port 206 nsew signal input
rlabel metal2 s 1214 -300 1270 160 8 N1END[2]
port 207 nsew signal input
rlabel metal2 s 1582 -300 1638 160 8 N1END[3]
port 208 nsew signal input
rlabel metal2 s 1950 44540 2006 45000 6 N2BEG[0]
port 209 nsew signal output
rlabel metal2 s 2318 44540 2374 45000 6 N2BEG[1]
port 210 nsew signal output
rlabel metal2 s 2686 44540 2742 45000 6 N2BEG[2]
port 211 nsew signal output
rlabel metal2 s 3054 44540 3110 45000 6 N2BEG[3]
port 212 nsew signal output
rlabel metal2 s 3422 44540 3478 45000 6 N2BEG[4]
port 213 nsew signal output
rlabel metal2 s 3790 44540 3846 45000 6 N2BEG[5]
port 214 nsew signal output
rlabel metal2 s 4158 44540 4214 45000 6 N2BEG[6]
port 215 nsew signal output
rlabel metal2 s 4526 44540 4582 45000 6 N2BEG[7]
port 216 nsew signal output
rlabel metal2 s 4894 44540 4950 45000 6 N2BEGb[0]
port 217 nsew signal output
rlabel metal2 s 5262 44540 5318 45000 6 N2BEGb[1]
port 218 nsew signal output
rlabel metal2 s 5630 44540 5686 45000 6 N2BEGb[2]
port 219 nsew signal output
rlabel metal2 s 5998 44540 6054 45000 6 N2BEGb[3]
port 220 nsew signal output
rlabel metal2 s 6366 44540 6422 45000 6 N2BEGb[4]
port 221 nsew signal output
rlabel metal2 s 6734 44540 6790 45000 6 N2BEGb[5]
port 222 nsew signal output
rlabel metal2 s 7102 44540 7158 45000 6 N2BEGb[6]
port 223 nsew signal output
rlabel metal2 s 7470 44540 7526 45000 6 N2BEGb[7]
port 224 nsew signal output
rlabel metal2 s 4894 -300 4950 160 8 N2END[0]
port 225 nsew signal input
rlabel metal2 s 5262 -300 5318 160 8 N2END[1]
port 226 nsew signal input
rlabel metal2 s 5630 -300 5686 160 8 N2END[2]
port 227 nsew signal input
rlabel metal2 s 5998 -300 6054 160 8 N2END[3]
port 228 nsew signal input
rlabel metal2 s 6366 -300 6422 160 8 N2END[4]
port 229 nsew signal input
rlabel metal2 s 6734 -300 6790 160 8 N2END[5]
port 230 nsew signal input
rlabel metal2 s 7102 -300 7158 160 8 N2END[6]
port 231 nsew signal input
rlabel metal2 s 7470 -300 7526 160 8 N2END[7]
port 232 nsew signal input
rlabel metal2 s 1950 -300 2006 160 8 N2MID[0]
port 233 nsew signal input
rlabel metal2 s 2318 -300 2374 160 8 N2MID[1]
port 234 nsew signal input
rlabel metal2 s 2686 -300 2742 160 8 N2MID[2]
port 235 nsew signal input
rlabel metal2 s 3054 -300 3110 160 8 N2MID[3]
port 236 nsew signal input
rlabel metal2 s 3422 -300 3478 160 8 N2MID[4]
port 237 nsew signal input
rlabel metal2 s 3790 -300 3846 160 8 N2MID[5]
port 238 nsew signal input
rlabel metal2 s 4158 -300 4214 160 8 N2MID[6]
port 239 nsew signal input
rlabel metal2 s 4526 -300 4582 160 8 N2MID[7]
port 240 nsew signal input
rlabel metal2 s 7838 44540 7894 45000 6 N4BEG[0]
port 241 nsew signal output
rlabel metal2 s 11518 44540 11574 45000 6 N4BEG[10]
port 242 nsew signal output
rlabel metal2 s 11886 44540 11942 45000 6 N4BEG[11]
port 243 nsew signal output
rlabel metal2 s 12254 44540 12310 45000 6 N4BEG[12]
port 244 nsew signal output
rlabel metal2 s 12622 44540 12678 45000 6 N4BEG[13]
port 245 nsew signal output
rlabel metal2 s 12990 44540 13046 45000 6 N4BEG[14]
port 246 nsew signal output
rlabel metal2 s 13358 44540 13414 45000 6 N4BEG[15]
port 247 nsew signal output
rlabel metal2 s 8206 44540 8262 45000 6 N4BEG[1]
port 248 nsew signal output
rlabel metal2 s 8574 44540 8630 45000 6 N4BEG[2]
port 249 nsew signal output
rlabel metal2 s 8942 44540 8998 45000 6 N4BEG[3]
port 250 nsew signal output
rlabel metal2 s 9310 44540 9366 45000 6 N4BEG[4]
port 251 nsew signal output
rlabel metal2 s 9678 44540 9734 45000 6 N4BEG[5]
port 252 nsew signal output
rlabel metal2 s 10046 44540 10102 45000 6 N4BEG[6]
port 253 nsew signal output
rlabel metal2 s 10414 44540 10470 45000 6 N4BEG[7]
port 254 nsew signal output
rlabel metal2 s 10782 44540 10838 45000 6 N4BEG[8]
port 255 nsew signal output
rlabel metal2 s 11150 44540 11206 45000 6 N4BEG[9]
port 256 nsew signal output
rlabel metal2 s 7838 -300 7894 160 8 N4END[0]
port 257 nsew signal input
rlabel metal2 s 11518 -300 11574 160 8 N4END[10]
port 258 nsew signal input
rlabel metal2 s 11886 -300 11942 160 8 N4END[11]
port 259 nsew signal input
rlabel metal2 s 12254 -300 12310 160 8 N4END[12]
port 260 nsew signal input
rlabel metal2 s 12622 -300 12678 160 8 N4END[13]
port 261 nsew signal input
rlabel metal2 s 12990 -300 13046 160 8 N4END[14]
port 262 nsew signal input
rlabel metal2 s 13358 -300 13414 160 8 N4END[15]
port 263 nsew signal input
rlabel metal2 s 8206 -300 8262 160 8 N4END[1]
port 264 nsew signal input
rlabel metal2 s 8574 -300 8630 160 8 N4END[2]
port 265 nsew signal input
rlabel metal2 s 8942 -300 8998 160 8 N4END[3]
port 266 nsew signal input
rlabel metal2 s 9310 -300 9366 160 8 N4END[4]
port 267 nsew signal input
rlabel metal2 s 9678 -300 9734 160 8 N4END[5]
port 268 nsew signal input
rlabel metal2 s 10046 -300 10102 160 8 N4END[6]
port 269 nsew signal input
rlabel metal2 s 10414 -300 10470 160 8 N4END[7]
port 270 nsew signal input
rlabel metal2 s 10782 -300 10838 160 8 N4END[8]
port 271 nsew signal input
rlabel metal2 s 11150 -300 11206 160 8 N4END[9]
port 272 nsew signal input
rlabel metal2 s 13726 44540 13782 45000 6 NN4BEG[0]
port 273 nsew signal output
rlabel metal2 s 17406 44540 17462 45000 6 NN4BEG[10]
port 274 nsew signal output
rlabel metal2 s 17774 44540 17830 45000 6 NN4BEG[11]
port 275 nsew signal output
rlabel metal2 s 18142 44540 18198 45000 6 NN4BEG[12]
port 276 nsew signal output
rlabel metal2 s 18510 44540 18566 45000 6 NN4BEG[13]
port 277 nsew signal output
rlabel metal2 s 18878 44540 18934 45000 6 NN4BEG[14]
port 278 nsew signal output
rlabel metal2 s 19246 44540 19302 45000 6 NN4BEG[15]
port 279 nsew signal output
rlabel metal2 s 14094 44540 14150 45000 6 NN4BEG[1]
port 280 nsew signal output
rlabel metal2 s 14462 44540 14518 45000 6 NN4BEG[2]
port 281 nsew signal output
rlabel metal2 s 14830 44540 14886 45000 6 NN4BEG[3]
port 282 nsew signal output
rlabel metal2 s 15198 44540 15254 45000 6 NN4BEG[4]
port 283 nsew signal output
rlabel metal2 s 15566 44540 15622 45000 6 NN4BEG[5]
port 284 nsew signal output
rlabel metal2 s 15934 44540 15990 45000 6 NN4BEG[6]
port 285 nsew signal output
rlabel metal2 s 16302 44540 16358 45000 6 NN4BEG[7]
port 286 nsew signal output
rlabel metal2 s 16670 44540 16726 45000 6 NN4BEG[8]
port 287 nsew signal output
rlabel metal2 s 17038 44540 17094 45000 6 NN4BEG[9]
port 288 nsew signal output
rlabel metal2 s 13726 -300 13782 160 8 NN4END[0]
port 289 nsew signal input
rlabel metal2 s 17406 -300 17462 160 8 NN4END[10]
port 290 nsew signal input
rlabel metal2 s 17774 -300 17830 160 8 NN4END[11]
port 291 nsew signal input
rlabel metal2 s 18142 -300 18198 160 8 NN4END[12]
port 292 nsew signal input
rlabel metal2 s 18510 -300 18566 160 8 NN4END[13]
port 293 nsew signal input
rlabel metal2 s 18878 -300 18934 160 8 NN4END[14]
port 294 nsew signal input
rlabel metal2 s 19246 -300 19302 160 8 NN4END[15]
port 295 nsew signal input
rlabel metal2 s 14094 -300 14150 160 8 NN4END[1]
port 296 nsew signal input
rlabel metal2 s 14462 -300 14518 160 8 NN4END[2]
port 297 nsew signal input
rlabel metal2 s 14830 -300 14886 160 8 NN4END[3]
port 298 nsew signal input
rlabel metal2 s 15198 -300 15254 160 8 NN4END[4]
port 299 nsew signal input
rlabel metal2 s 15566 -300 15622 160 8 NN4END[5]
port 300 nsew signal input
rlabel metal2 s 15934 -300 15990 160 8 NN4END[6]
port 301 nsew signal input
rlabel metal2 s 16302 -300 16358 160 8 NN4END[7]
port 302 nsew signal input
rlabel metal2 s 16670 -300 16726 160 8 NN4END[8]
port 303 nsew signal input
rlabel metal2 s 17038 -300 17094 160 8 NN4END[9]
port 304 nsew signal input
rlabel metal2 s 19614 -300 19670 160 8 S1BEG[0]
port 305 nsew signal output
rlabel metal2 s 19982 -300 20038 160 8 S1BEG[1]
port 306 nsew signal output
rlabel metal2 s 20350 -300 20406 160 8 S1BEG[2]
port 307 nsew signal output
rlabel metal2 s 20718 -300 20774 160 8 S1BEG[3]
port 308 nsew signal output
rlabel metal2 s 19614 44540 19670 45000 6 S1END[0]
port 309 nsew signal input
rlabel metal2 s 19982 44540 20038 45000 6 S1END[1]
port 310 nsew signal input
rlabel metal2 s 20350 44540 20406 45000 6 S1END[2]
port 311 nsew signal input
rlabel metal2 s 20718 44540 20774 45000 6 S1END[3]
port 312 nsew signal input
rlabel metal2 s 24030 -300 24086 160 8 S2BEG[0]
port 313 nsew signal output
rlabel metal2 s 24398 -300 24454 160 8 S2BEG[1]
port 314 nsew signal output
rlabel metal2 s 24766 -300 24822 160 8 S2BEG[2]
port 315 nsew signal output
rlabel metal2 s 25134 -300 25190 160 8 S2BEG[3]
port 316 nsew signal output
rlabel metal2 s 25502 -300 25558 160 8 S2BEG[4]
port 317 nsew signal output
rlabel metal2 s 25870 -300 25926 160 8 S2BEG[5]
port 318 nsew signal output
rlabel metal2 s 26238 -300 26294 160 8 S2BEG[6]
port 319 nsew signal output
rlabel metal2 s 26606 -300 26662 160 8 S2BEG[7]
port 320 nsew signal output
rlabel metal2 s 21086 -300 21142 160 8 S2BEGb[0]
port 321 nsew signal output
rlabel metal2 s 21454 -300 21510 160 8 S2BEGb[1]
port 322 nsew signal output
rlabel metal2 s 21822 -300 21878 160 8 S2BEGb[2]
port 323 nsew signal output
rlabel metal2 s 22190 -300 22246 160 8 S2BEGb[3]
port 324 nsew signal output
rlabel metal2 s 22558 -300 22614 160 8 S2BEGb[4]
port 325 nsew signal output
rlabel metal2 s 22926 -300 22982 160 8 S2BEGb[5]
port 326 nsew signal output
rlabel metal2 s 23294 -300 23350 160 8 S2BEGb[6]
port 327 nsew signal output
rlabel metal2 s 23662 -300 23718 160 8 S2BEGb[7]
port 328 nsew signal output
rlabel metal2 s 21086 44540 21142 45000 6 S2END[0]
port 329 nsew signal input
rlabel metal2 s 21454 44540 21510 45000 6 S2END[1]
port 330 nsew signal input
rlabel metal2 s 21822 44540 21878 45000 6 S2END[2]
port 331 nsew signal input
rlabel metal2 s 22190 44540 22246 45000 6 S2END[3]
port 332 nsew signal input
rlabel metal2 s 22558 44540 22614 45000 6 S2END[4]
port 333 nsew signal input
rlabel metal2 s 22926 44540 22982 45000 6 S2END[5]
port 334 nsew signal input
rlabel metal2 s 23294 44540 23350 45000 6 S2END[6]
port 335 nsew signal input
rlabel metal2 s 23662 44540 23718 45000 6 S2END[7]
port 336 nsew signal input
rlabel metal2 s 24030 44540 24086 45000 6 S2MID[0]
port 337 nsew signal input
rlabel metal2 s 24398 44540 24454 45000 6 S2MID[1]
port 338 nsew signal input
rlabel metal2 s 24766 44540 24822 45000 6 S2MID[2]
port 339 nsew signal input
rlabel metal2 s 25134 44540 25190 45000 6 S2MID[3]
port 340 nsew signal input
rlabel metal2 s 25502 44540 25558 45000 6 S2MID[4]
port 341 nsew signal input
rlabel metal2 s 25870 44540 25926 45000 6 S2MID[5]
port 342 nsew signal input
rlabel metal2 s 26238 44540 26294 45000 6 S2MID[6]
port 343 nsew signal input
rlabel metal2 s 26606 44540 26662 45000 6 S2MID[7]
port 344 nsew signal input
rlabel metal2 s 26974 -300 27030 160 8 S4BEG[0]
port 345 nsew signal output
rlabel metal2 s 30654 -300 30710 160 8 S4BEG[10]
port 346 nsew signal output
rlabel metal2 s 31022 -300 31078 160 8 S4BEG[11]
port 347 nsew signal output
rlabel metal2 s 31390 -300 31446 160 8 S4BEG[12]
port 348 nsew signal output
rlabel metal2 s 31758 -300 31814 160 8 S4BEG[13]
port 349 nsew signal output
rlabel metal2 s 32126 -300 32182 160 8 S4BEG[14]
port 350 nsew signal output
rlabel metal2 s 32494 -300 32550 160 8 S4BEG[15]
port 351 nsew signal output
rlabel metal2 s 27342 -300 27398 160 8 S4BEG[1]
port 352 nsew signal output
rlabel metal2 s 27710 -300 27766 160 8 S4BEG[2]
port 353 nsew signal output
rlabel metal2 s 28078 -300 28134 160 8 S4BEG[3]
port 354 nsew signal output
rlabel metal2 s 28446 -300 28502 160 8 S4BEG[4]
port 355 nsew signal output
rlabel metal2 s 28814 -300 28870 160 8 S4BEG[5]
port 356 nsew signal output
rlabel metal2 s 29182 -300 29238 160 8 S4BEG[6]
port 357 nsew signal output
rlabel metal2 s 29550 -300 29606 160 8 S4BEG[7]
port 358 nsew signal output
rlabel metal2 s 29918 -300 29974 160 8 S4BEG[8]
port 359 nsew signal output
rlabel metal2 s 30286 -300 30342 160 8 S4BEG[9]
port 360 nsew signal output
rlabel metal2 s 26974 44540 27030 45000 6 S4END[0]
port 361 nsew signal input
rlabel metal2 s 30654 44540 30710 45000 6 S4END[10]
port 362 nsew signal input
rlabel metal2 s 31022 44540 31078 45000 6 S4END[11]
port 363 nsew signal input
rlabel metal2 s 31390 44540 31446 45000 6 S4END[12]
port 364 nsew signal input
rlabel metal2 s 31758 44540 31814 45000 6 S4END[13]
port 365 nsew signal input
rlabel metal2 s 32126 44540 32182 45000 6 S4END[14]
port 366 nsew signal input
rlabel metal2 s 32494 44540 32550 45000 6 S4END[15]
port 367 nsew signal input
rlabel metal2 s 27342 44540 27398 45000 6 S4END[1]
port 368 nsew signal input
rlabel metal2 s 27710 44540 27766 45000 6 S4END[2]
port 369 nsew signal input
rlabel metal2 s 28078 44540 28134 45000 6 S4END[3]
port 370 nsew signal input
rlabel metal2 s 28446 44540 28502 45000 6 S4END[4]
port 371 nsew signal input
rlabel metal2 s 28814 44540 28870 45000 6 S4END[5]
port 372 nsew signal input
rlabel metal2 s 29182 44540 29238 45000 6 S4END[6]
port 373 nsew signal input
rlabel metal2 s 29550 44540 29606 45000 6 S4END[7]
port 374 nsew signal input
rlabel metal2 s 29918 44540 29974 45000 6 S4END[8]
port 375 nsew signal input
rlabel metal2 s 30286 44540 30342 45000 6 S4END[9]
port 376 nsew signal input
rlabel metal2 s 32862 -300 32918 160 8 SS4BEG[0]
port 377 nsew signal output
rlabel metal2 s 36542 -300 36598 160 8 SS4BEG[10]
port 378 nsew signal output
rlabel metal2 s 36910 -300 36966 160 8 SS4BEG[11]
port 379 nsew signal output
rlabel metal2 s 37278 -300 37334 160 8 SS4BEG[12]
port 380 nsew signal output
rlabel metal2 s 37646 -300 37702 160 8 SS4BEG[13]
port 381 nsew signal output
rlabel metal2 s 38014 -300 38070 160 8 SS4BEG[14]
port 382 nsew signal output
rlabel metal2 s 38382 -300 38438 160 8 SS4BEG[15]
port 383 nsew signal output
rlabel metal2 s 33230 -300 33286 160 8 SS4BEG[1]
port 384 nsew signal output
rlabel metal2 s 33598 -300 33654 160 8 SS4BEG[2]
port 385 nsew signal output
rlabel metal2 s 33966 -300 34022 160 8 SS4BEG[3]
port 386 nsew signal output
rlabel metal2 s 34334 -300 34390 160 8 SS4BEG[4]
port 387 nsew signal output
rlabel metal2 s 34702 -300 34758 160 8 SS4BEG[5]
port 388 nsew signal output
rlabel metal2 s 35070 -300 35126 160 8 SS4BEG[6]
port 389 nsew signal output
rlabel metal2 s 35438 -300 35494 160 8 SS4BEG[7]
port 390 nsew signal output
rlabel metal2 s 35806 -300 35862 160 8 SS4BEG[8]
port 391 nsew signal output
rlabel metal2 s 36174 -300 36230 160 8 SS4BEG[9]
port 392 nsew signal output
rlabel metal2 s 32862 44540 32918 45000 6 SS4END[0]
port 393 nsew signal input
rlabel metal2 s 36542 44540 36598 45000 6 SS4END[10]
port 394 nsew signal input
rlabel metal2 s 36910 44540 36966 45000 6 SS4END[11]
port 395 nsew signal input
rlabel metal2 s 37278 44540 37334 45000 6 SS4END[12]
port 396 nsew signal input
rlabel metal2 s 37646 44540 37702 45000 6 SS4END[13]
port 397 nsew signal input
rlabel metal2 s 38014 44540 38070 45000 6 SS4END[14]
port 398 nsew signal input
rlabel metal2 s 38382 44540 38438 45000 6 SS4END[15]
port 399 nsew signal input
rlabel metal2 s 33230 44540 33286 45000 6 SS4END[1]
port 400 nsew signal input
rlabel metal2 s 33598 44540 33654 45000 6 SS4END[2]
port 401 nsew signal input
rlabel metal2 s 33966 44540 34022 45000 6 SS4END[3]
port 402 nsew signal input
rlabel metal2 s 34334 44540 34390 45000 6 SS4END[4]
port 403 nsew signal input
rlabel metal2 s 34702 44540 34758 45000 6 SS4END[5]
port 404 nsew signal input
rlabel metal2 s 35070 44540 35126 45000 6 SS4END[6]
port 405 nsew signal input
rlabel metal2 s 35438 44540 35494 45000 6 SS4END[7]
port 406 nsew signal input
rlabel metal2 s 35806 44540 35862 45000 6 SS4END[8]
port 407 nsew signal input
rlabel metal2 s 36174 44540 36230 45000 6 SS4END[9]
port 408 nsew signal input
rlabel metal2 s 38750 -300 38806 160 8 UserCLK
port 409 nsew signal input
rlabel metal2 s 38750 44540 38806 45000 6 UserCLKo
port 410 nsew signal output
rlabel metal4 s 19568 1040 19888 43568 6 VGND
port 411 nsew ground bidirectional
rlabel metal4 s 4208 1040 4528 43568 6 VPWR
port 412 nsew power bidirectional
rlabel metal4 s 34928 1040 35248 43568 6 VPWR
port 412 nsew power bidirectional
rlabel metal3 s -300 4904 160 5024 4 W1BEG[0]
port 413 nsew signal output
rlabel metal3 s -300 5176 160 5296 4 W1BEG[1]
port 414 nsew signal output
rlabel metal3 s -300 5448 160 5568 4 W1BEG[2]
port 415 nsew signal output
rlabel metal3 s -300 5720 160 5840 4 W1BEG[3]
port 416 nsew signal output
rlabel metal3 s 46540 4904 47000 5024 6 W1END[0]
port 417 nsew signal input
rlabel metal3 s 46540 5176 47000 5296 6 W1END[1]
port 418 nsew signal input
rlabel metal3 s 46540 5448 47000 5568 6 W1END[2]
port 419 nsew signal input
rlabel metal3 s 46540 5720 47000 5840 6 W1END[3]
port 420 nsew signal input
rlabel metal3 s -300 5992 160 6112 4 W2BEG[0]
port 421 nsew signal output
rlabel metal3 s -300 6264 160 6384 4 W2BEG[1]
port 422 nsew signal output
rlabel metal3 s -300 6536 160 6656 4 W2BEG[2]
port 423 nsew signal output
rlabel metal3 s -300 6808 160 6928 4 W2BEG[3]
port 424 nsew signal output
rlabel metal3 s -300 7080 160 7200 4 W2BEG[4]
port 425 nsew signal output
rlabel metal3 s -300 7352 160 7472 4 W2BEG[5]
port 426 nsew signal output
rlabel metal3 s -300 7624 160 7744 4 W2BEG[6]
port 427 nsew signal output
rlabel metal3 s -300 7896 160 8016 4 W2BEG[7]
port 428 nsew signal output
rlabel metal3 s -300 8168 160 8288 4 W2BEGb[0]
port 429 nsew signal output
rlabel metal3 s -300 8440 160 8560 4 W2BEGb[1]
port 430 nsew signal output
rlabel metal3 s -300 8712 160 8832 4 W2BEGb[2]
port 431 nsew signal output
rlabel metal3 s -300 8984 160 9104 4 W2BEGb[3]
port 432 nsew signal output
rlabel metal3 s -300 9256 160 9376 4 W2BEGb[4]
port 433 nsew signal output
rlabel metal3 s -300 9528 160 9648 4 W2BEGb[5]
port 434 nsew signal output
rlabel metal3 s -300 9800 160 9920 4 W2BEGb[6]
port 435 nsew signal output
rlabel metal3 s -300 10072 160 10192 4 W2BEGb[7]
port 436 nsew signal output
rlabel metal3 s 46540 8168 47000 8288 6 W2END[0]
port 437 nsew signal input
rlabel metal3 s 46540 8440 47000 8560 6 W2END[1]
port 438 nsew signal input
rlabel metal3 s 46540 8712 47000 8832 6 W2END[2]
port 439 nsew signal input
rlabel metal3 s 46540 8984 47000 9104 6 W2END[3]
port 440 nsew signal input
rlabel metal3 s 46540 9256 47000 9376 6 W2END[4]
port 441 nsew signal input
rlabel metal3 s 46540 9528 47000 9648 6 W2END[5]
port 442 nsew signal input
rlabel metal3 s 46540 9800 47000 9920 6 W2END[6]
port 443 nsew signal input
rlabel metal3 s 46540 10072 47000 10192 6 W2END[7]
port 444 nsew signal input
rlabel metal3 s 46540 5992 47000 6112 6 W2MID[0]
port 445 nsew signal input
rlabel metal3 s 46540 6264 47000 6384 6 W2MID[1]
port 446 nsew signal input
rlabel metal3 s 46540 6536 47000 6656 6 W2MID[2]
port 447 nsew signal input
rlabel metal3 s 46540 6808 47000 6928 6 W2MID[3]
port 448 nsew signal input
rlabel metal3 s 46540 7080 47000 7200 6 W2MID[4]
port 449 nsew signal input
rlabel metal3 s 46540 7352 47000 7472 6 W2MID[5]
port 450 nsew signal input
rlabel metal3 s 46540 7624 47000 7744 6 W2MID[6]
port 451 nsew signal input
rlabel metal3 s 46540 7896 47000 8016 6 W2MID[7]
port 452 nsew signal input
rlabel metal3 s -300 14696 160 14816 4 W6BEG[0]
port 453 nsew signal output
rlabel metal3 s -300 17416 160 17536 4 W6BEG[10]
port 454 nsew signal output
rlabel metal3 s -300 17688 160 17808 4 W6BEG[11]
port 455 nsew signal output
rlabel metal3 s -300 14968 160 15088 4 W6BEG[1]
port 456 nsew signal output
rlabel metal3 s -300 15240 160 15360 4 W6BEG[2]
port 457 nsew signal output
rlabel metal3 s -300 15512 160 15632 4 W6BEG[3]
port 458 nsew signal output
rlabel metal3 s -300 15784 160 15904 4 W6BEG[4]
port 459 nsew signal output
rlabel metal3 s -300 16056 160 16176 4 W6BEG[5]
port 460 nsew signal output
rlabel metal3 s -300 16328 160 16448 4 W6BEG[6]
port 461 nsew signal output
rlabel metal3 s -300 16600 160 16720 4 W6BEG[7]
port 462 nsew signal output
rlabel metal3 s -300 16872 160 16992 4 W6BEG[8]
port 463 nsew signal output
rlabel metal3 s -300 17144 160 17264 4 W6BEG[9]
port 464 nsew signal output
rlabel metal3 s 46540 14696 47000 14816 6 W6END[0]
port 465 nsew signal input
rlabel metal3 s 46540 17416 47000 17536 6 W6END[10]
port 466 nsew signal input
rlabel metal3 s 46540 17688 47000 17808 6 W6END[11]
port 467 nsew signal input
rlabel metal3 s 46540 14968 47000 15088 6 W6END[1]
port 468 nsew signal input
rlabel metal3 s 46540 15240 47000 15360 6 W6END[2]
port 469 nsew signal input
rlabel metal3 s 46540 15512 47000 15632 6 W6END[3]
port 470 nsew signal input
rlabel metal3 s 46540 15784 47000 15904 6 W6END[4]
port 471 nsew signal input
rlabel metal3 s 46540 16056 47000 16176 6 W6END[5]
port 472 nsew signal input
rlabel metal3 s 46540 16328 47000 16448 6 W6END[6]
port 473 nsew signal input
rlabel metal3 s 46540 16600 47000 16720 6 W6END[7]
port 474 nsew signal input
rlabel metal3 s 46540 16872 47000 16992 6 W6END[8]
port 475 nsew signal input
rlabel metal3 s 46540 17144 47000 17264 6 W6END[9]
port 476 nsew signal input
rlabel metal3 s -300 10344 160 10464 4 WW4BEG[0]
port 477 nsew signal output
rlabel metal3 s -300 13064 160 13184 4 WW4BEG[10]
port 478 nsew signal output
rlabel metal3 s -300 13336 160 13456 4 WW4BEG[11]
port 479 nsew signal output
rlabel metal3 s -300 13608 160 13728 4 WW4BEG[12]
port 480 nsew signal output
rlabel metal3 s -300 13880 160 14000 4 WW4BEG[13]
port 481 nsew signal output
rlabel metal3 s -300 14152 160 14272 4 WW4BEG[14]
port 482 nsew signal output
rlabel metal3 s -300 14424 160 14544 4 WW4BEG[15]
port 483 nsew signal output
rlabel metal3 s -300 10616 160 10736 4 WW4BEG[1]
port 484 nsew signal output
rlabel metal3 s -300 10888 160 11008 4 WW4BEG[2]
port 485 nsew signal output
rlabel metal3 s -300 11160 160 11280 4 WW4BEG[3]
port 486 nsew signal output
rlabel metal3 s -300 11432 160 11552 4 WW4BEG[4]
port 487 nsew signal output
rlabel metal3 s -300 11704 160 11824 4 WW4BEG[5]
port 488 nsew signal output
rlabel metal3 s -300 11976 160 12096 4 WW4BEG[6]
port 489 nsew signal output
rlabel metal3 s -300 12248 160 12368 4 WW4BEG[7]
port 490 nsew signal output
rlabel metal3 s -300 12520 160 12640 4 WW4BEG[8]
port 491 nsew signal output
rlabel metal3 s -300 12792 160 12912 4 WW4BEG[9]
port 492 nsew signal output
rlabel metal3 s 46540 10344 47000 10464 6 WW4END[0]
port 493 nsew signal input
rlabel metal3 s 46540 13064 47000 13184 6 WW4END[10]
port 494 nsew signal input
rlabel metal3 s 46540 13336 47000 13456 6 WW4END[11]
port 495 nsew signal input
rlabel metal3 s 46540 13608 47000 13728 6 WW4END[12]
port 496 nsew signal input
rlabel metal3 s 46540 13880 47000 14000 6 WW4END[13]
port 497 nsew signal input
rlabel metal3 s 46540 14152 47000 14272 6 WW4END[14]
port 498 nsew signal input
rlabel metal3 s 46540 14424 47000 14544 6 WW4END[15]
port 499 nsew signal input
rlabel metal3 s 46540 10616 47000 10736 6 WW4END[1]
port 500 nsew signal input
rlabel metal3 s 46540 10888 47000 11008 6 WW4END[2]
port 501 nsew signal input
rlabel metal3 s 46540 11160 47000 11280 6 WW4END[3]
port 502 nsew signal input
rlabel metal3 s 46540 11432 47000 11552 6 WW4END[4]
port 503 nsew signal input
rlabel metal3 s 46540 11704 47000 11824 6 WW4END[5]
port 504 nsew signal input
rlabel metal3 s 46540 11976 47000 12096 6 WW4END[6]
port 505 nsew signal input
rlabel metal3 s 46540 12248 47000 12368 6 WW4END[7]
port 506 nsew signal input
rlabel metal3 s 46540 12520 47000 12640 6 WW4END[8]
port 507 nsew signal input
rlabel metal3 s 46540 12792 47000 12912 6 WW4END[9]
port 508 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 46700 44700
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 7709022
string GDS_FILE /home/asma/Desktop/open_eFPGA/openlane/RegFile/runs/24_12_07_23_54/results/signoff/RegFile.magic.gds
string GDS_START 287328
<< end >>

