magic
tech sky130A
magscale 1 2
timestamp 1733618660
<< viali >>
rect 2145 8585 2179 8619
rect 2789 8585 2823 8619
rect 3525 8585 3559 8619
rect 4537 8585 4571 8619
rect 4997 8585 5031 8619
rect 5549 8585 5583 8619
rect 6561 8585 6595 8619
rect 7021 8585 7055 8619
rect 7757 8585 7791 8619
rect 8125 8585 8159 8619
rect 8677 8585 8711 8619
rect 9229 8585 9263 8619
rect 9781 8585 9815 8619
rect 10333 8585 10367 8619
rect 10701 8585 10735 8619
rect 11253 8585 11287 8619
rect 11989 8585 12023 8619
rect 12541 8585 12575 8619
rect 13277 8585 13311 8619
rect 13645 8585 13679 8619
rect 14381 8585 14415 8619
rect 14749 8585 14783 8619
rect 15301 8585 15335 8619
rect 15669 8585 15703 8619
rect 16037 8585 16071 8619
rect 16405 8585 16439 8619
rect 16865 8585 16899 8619
rect 17509 8585 17543 8619
rect 18061 8585 18095 8619
rect 18429 8585 18463 8619
rect 18797 8585 18831 8619
rect 19901 8585 19935 8619
rect 20637 8585 20671 8619
rect 22845 8585 22879 8619
rect 22937 8585 22971 8619
rect 23397 8585 23431 8619
rect 31493 8585 31527 8619
rect 32321 8585 32355 8619
rect 32413 8585 32447 8619
rect 33149 8585 33183 8619
rect 33517 8585 33551 8619
rect 33885 8585 33919 8619
rect 34253 8585 34287 8619
rect 35449 8585 35483 8619
rect 35725 8585 35759 8619
rect 38301 8585 38335 8619
rect 38669 8585 38703 8619
rect 39037 8585 39071 8619
rect 39589 8585 39623 8619
rect 40049 8585 40083 8619
rect 40601 8585 40635 8619
rect 41521 8585 41555 8619
rect 42625 8585 42659 8619
rect 44281 8585 44315 8619
rect 3249 8517 3283 8551
rect 5825 8517 5859 8551
rect 6193 8517 6227 8551
rect 6929 8517 6963 8551
rect 10977 8517 11011 8551
rect 11897 8517 11931 8551
rect 12449 8517 12483 8551
rect 43085 8517 43119 8551
rect 44189 8517 44223 8551
rect 2329 8449 2363 8483
rect 2697 8449 2731 8483
rect 4169 8449 4203 8483
rect 4721 8449 4755 8483
rect 4813 8449 4847 8483
rect 5273 8449 5307 8483
rect 6377 8449 6411 8483
rect 7573 8449 7607 8483
rect 8033 8449 8067 8483
rect 8493 8449 8527 8483
rect 9045 8449 9079 8483
rect 9505 8449 9539 8483
rect 10149 8449 10183 8483
rect 10517 8449 10551 8483
rect 13093 8449 13127 8483
rect 13553 8449 13587 8483
rect 14197 8449 14231 8483
rect 14565 8449 14599 8483
rect 15025 8449 15059 8483
rect 15485 8449 15519 8483
rect 15853 8449 15887 8483
rect 16221 8449 16255 8483
rect 16773 8449 16807 8483
rect 17325 8449 17359 8483
rect 17785 8449 17819 8483
rect 18245 8449 18279 8483
rect 18613 8449 18647 8483
rect 19625 8449 19659 8483
rect 19809 8449 19843 8483
rect 20545 8449 20579 8483
rect 20821 8449 20855 8483
rect 21097 8449 21131 8483
rect 21373 8449 21407 8483
rect 21649 8449 21683 8483
rect 22017 8449 22051 8483
rect 22293 8449 22327 8483
rect 22569 8449 22603 8483
rect 22661 8449 22695 8483
rect 23121 8449 23155 8483
rect 23581 8449 23615 8483
rect 23765 8449 23799 8483
rect 24225 8449 24259 8483
rect 24685 8449 24719 8483
rect 24961 8449 24995 8483
rect 25237 8449 25271 8483
rect 25513 8449 25547 8483
rect 25789 8449 25823 8483
rect 26157 8449 26191 8483
rect 26525 8449 26559 8483
rect 27169 8449 27203 8483
rect 27445 8449 27479 8483
rect 27721 8449 27755 8483
rect 27997 8449 28031 8483
rect 28365 8449 28399 8483
rect 28733 8449 28767 8483
rect 29101 8449 29135 8483
rect 29745 8449 29779 8483
rect 30021 8449 30055 8483
rect 30297 8449 30331 8483
rect 30573 8473 30607 8507
rect 30941 8449 30975 8483
rect 31309 8449 31343 8483
rect 31677 8449 31711 8483
rect 32137 8449 32171 8483
rect 32597 8449 32631 8483
rect 32689 8449 32723 8483
rect 32965 8449 32999 8483
rect 33333 8449 33367 8483
rect 33701 8449 33735 8483
rect 34069 8449 34103 8483
rect 34713 8449 34747 8483
rect 34989 8449 35023 8483
rect 35265 8449 35299 8483
rect 35541 8449 35575 8483
rect 35909 8449 35943 8483
rect 36277 8449 36311 8483
rect 36645 8449 36679 8483
rect 37289 8449 37323 8483
rect 37565 8449 37599 8483
rect 37841 8449 37875 8483
rect 38117 8449 38151 8483
rect 38485 8449 38519 8483
rect 38945 8449 38979 8483
rect 39405 8449 39439 8483
rect 39957 8449 39991 8483
rect 40509 8449 40543 8483
rect 40969 8449 41003 8483
rect 41429 8449 41463 8483
rect 42533 8449 42567 8483
rect 43637 8449 43671 8483
rect 1777 8313 1811 8347
rect 20913 8313 20947 8347
rect 22109 8313 22143 8347
rect 22385 8313 22419 8347
rect 23949 8313 23983 8347
rect 24041 8313 24075 8347
rect 26341 8313 26375 8347
rect 26985 8313 27019 8347
rect 28181 8313 28215 8347
rect 34897 8313 34931 8347
rect 35173 8313 35207 8347
rect 36093 8313 36127 8347
rect 36461 8313 36495 8347
rect 36829 8313 36863 8347
rect 37473 8313 37507 8347
rect 37749 8313 37783 8347
rect 38025 8313 38059 8347
rect 41153 8313 41187 8347
rect 43269 8313 43303 8347
rect 43821 8313 43855 8347
rect 19441 8245 19475 8279
rect 20361 8245 20395 8279
rect 21189 8245 21223 8279
rect 21465 8245 21499 8279
rect 21833 8245 21867 8279
rect 24501 8245 24535 8279
rect 24777 8245 24811 8279
rect 25053 8245 25087 8279
rect 25329 8245 25363 8279
rect 25605 8245 25639 8279
rect 25973 8245 26007 8279
rect 27261 8245 27295 8279
rect 27537 8245 27571 8279
rect 27813 8245 27847 8279
rect 28549 8245 28583 8279
rect 28917 8245 28951 8279
rect 29561 8245 29595 8279
rect 29837 8245 29871 8279
rect 30113 8245 30147 8279
rect 30389 8245 30423 8279
rect 30757 8245 30791 8279
rect 31125 8245 31159 8279
rect 32873 8245 32907 8279
rect 2053 8041 2087 8075
rect 2789 8041 2823 8075
rect 3157 8041 3191 8075
rect 3525 8041 3559 8075
rect 4169 8041 4203 8075
rect 4629 8041 4663 8075
rect 6469 8041 6503 8075
rect 7573 8041 7607 8075
rect 9137 8041 9171 8075
rect 10149 8041 10183 8075
rect 11621 8041 11655 8075
rect 12173 8041 12207 8075
rect 13093 8041 13127 8075
rect 14289 8041 14323 8075
rect 17325 8041 17359 8075
rect 17785 8041 17819 8075
rect 18061 8041 18095 8075
rect 19533 8041 19567 8075
rect 20453 8041 20487 8075
rect 20913 8041 20947 8075
rect 21557 8041 21591 8075
rect 22385 8041 22419 8075
rect 24593 8041 24627 8075
rect 27261 8041 27295 8075
rect 27629 8041 27663 8075
rect 27905 8041 27939 8075
rect 41153 8041 41187 8075
rect 43269 8041 43303 8075
rect 43821 8041 43855 8075
rect 44373 8041 44407 8075
rect 23949 7973 23983 8007
rect 24869 7973 24903 8007
rect 26525 7973 26559 8007
rect 42901 7973 42935 8007
rect 2973 7837 3007 7871
rect 3341 7837 3375 7871
rect 4445 7837 4479 7871
rect 7389 7837 7423 7871
rect 9965 7837 9999 7871
rect 11529 7837 11563 7871
rect 11989 7837 12023 7871
rect 12909 7837 12943 7871
rect 17141 7837 17175 7871
rect 17693 7837 17727 7871
rect 17969 7837 18003 7871
rect 18245 7837 18279 7871
rect 18337 7837 18371 7871
rect 18797 7837 18831 7871
rect 18889 7837 18923 7871
rect 19901 7837 19935 7871
rect 20177 7837 20211 7871
rect 20637 7837 20671 7871
rect 20729 7837 20763 7871
rect 21005 7837 21039 7871
rect 21281 7837 21315 7871
rect 21741 7837 21775 7871
rect 22017 7837 22051 7871
rect 22293 7837 22327 7871
rect 22569 7837 22603 7871
rect 22845 7837 22879 7871
rect 22937 7837 22971 7871
rect 23213 7837 23247 7871
rect 23489 7837 23523 7871
rect 23765 7837 23799 7871
rect 24041 7837 24075 7871
rect 24409 7837 24443 7871
rect 24685 7837 24719 7871
rect 24961 7837 24995 7871
rect 25237 7837 25271 7871
rect 25513 7837 25547 7871
rect 25789 7837 25823 7871
rect 26065 7837 26099 7871
rect 26341 7837 26375 7871
rect 26709 7837 26743 7871
rect 27077 7837 27111 7871
rect 27445 7837 27479 7871
rect 27721 7837 27755 7871
rect 27997 7837 28031 7871
rect 28273 7837 28307 7871
rect 28549 7837 28583 7871
rect 40969 7837 41003 7871
rect 1961 7769 1995 7803
rect 2513 7769 2547 7803
rect 3893 7769 3927 7803
rect 6377 7769 6411 7803
rect 9045 7769 9079 7803
rect 14197 7769 14231 7803
rect 19441 7769 19475 7803
rect 42625 7769 42659 7803
rect 43177 7769 43211 7803
rect 43729 7769 43763 7803
rect 44281 7769 44315 7803
rect 17509 7701 17543 7735
rect 18521 7701 18555 7735
rect 18613 7701 18647 7735
rect 19073 7701 19107 7735
rect 20085 7701 20119 7735
rect 20361 7701 20395 7735
rect 21189 7701 21223 7735
rect 21465 7701 21499 7735
rect 21833 7701 21867 7735
rect 22109 7701 22143 7735
rect 22661 7701 22695 7735
rect 23121 7701 23155 7735
rect 23397 7701 23431 7735
rect 23673 7701 23707 7735
rect 24225 7701 24259 7735
rect 25145 7701 25179 7735
rect 25421 7701 25455 7735
rect 25697 7701 25731 7735
rect 25973 7701 26007 7735
rect 26249 7701 26283 7735
rect 26893 7701 26927 7735
rect 28181 7701 28215 7735
rect 28457 7701 28491 7735
rect 28733 7701 28767 7735
rect 1777 7497 1811 7531
rect 2329 7497 2363 7531
rect 17509 7497 17543 7531
rect 18797 7497 18831 7531
rect 18889 7497 18923 7531
rect 19257 7497 19291 7531
rect 19717 7497 19751 7531
rect 22109 7497 22143 7531
rect 22477 7497 22511 7531
rect 43453 7497 43487 7531
rect 44741 7497 44775 7531
rect 2237 7429 2271 7463
rect 44281 7429 44315 7463
rect 1685 7361 1719 7395
rect 17693 7361 17727 7395
rect 18613 7361 18647 7395
rect 19073 7361 19107 7395
rect 19441 7361 19475 7395
rect 19901 7361 19935 7395
rect 21925 7361 21959 7395
rect 22201 7361 22235 7395
rect 22661 7361 22695 7395
rect 22937 7361 22971 7395
rect 23029 7361 23063 7395
rect 23397 7361 23431 7395
rect 23765 7361 23799 7395
rect 24041 7361 24075 7395
rect 43361 7361 43395 7395
rect 43913 7361 43947 7395
rect 44465 7361 44499 7395
rect 22385 7157 22419 7191
rect 22753 7157 22787 7191
rect 23213 7157 23247 7191
rect 23581 7157 23615 7191
rect 23949 7157 23983 7191
rect 24225 7157 24259 7191
rect 1777 6817 1811 6851
rect 44741 6817 44775 6851
rect 44281 6749 44315 6783
rect 1501 6681 1535 6715
rect 43913 6681 43947 6715
rect 44465 6681 44499 6715
rect 44925 6409 44959 6443
rect 44833 6273 44867 6307
rect 20453 2601 20487 2635
rect 22385 2601 22419 2635
rect 23397 2601 23431 2635
rect 23673 2601 23707 2635
rect 23949 2601 23983 2635
rect 24225 2601 24259 2635
rect 24869 2601 24903 2635
rect 27077 2601 27111 2635
rect 29285 2601 29319 2635
rect 43913 2601 43947 2635
rect 44189 2601 44223 2635
rect 44465 2601 44499 2635
rect 45017 2601 45051 2635
rect 22753 2533 22787 2567
rect 31493 2533 31527 2567
rect 33701 2533 33735 2567
rect 35909 2533 35943 2567
rect 22201 2397 22235 2431
rect 22937 2397 22971 2431
rect 23213 2397 23247 2431
rect 23489 2397 23523 2431
rect 23765 2397 23799 2431
rect 24041 2397 24075 2431
rect 24685 2397 24719 2431
rect 26893 2397 26927 2431
rect 29101 2397 29135 2431
rect 31309 2397 31343 2431
rect 33517 2397 33551 2431
rect 35725 2397 35759 2431
rect 37933 2397 37967 2431
rect 44097 2397 44131 2431
rect 44373 2397 44407 2431
rect 44649 2397 44683 2431
rect 45201 2397 45235 2431
rect 20361 2329 20395 2363
rect 22569 2329 22603 2363
rect 23121 2261 23155 2295
rect 38117 2261 38151 2295
rect 19441 2057 19475 2091
rect 21189 2057 21223 2091
rect 22293 2057 22327 2091
rect 22569 2057 22603 2091
rect 23121 2057 23155 2091
rect 23397 2057 23431 2091
rect 23857 2057 23891 2091
rect 26065 2057 26099 2091
rect 28273 2057 28307 2091
rect 30481 2057 30515 2091
rect 32689 2057 32723 2091
rect 34897 2057 34931 2091
rect 37289 2057 37323 2091
rect 41613 2057 41647 2091
rect 43453 2057 43487 2091
rect 43913 2057 43947 2091
rect 44373 2057 44407 2091
rect 20269 1989 20303 2023
rect 19625 1921 19659 1955
rect 20085 1921 20119 1955
rect 21373 1921 21407 1955
rect 21649 1921 21683 1955
rect 22201 1921 22235 1955
rect 22477 1921 22511 1955
rect 22753 1921 22787 1955
rect 22845 1921 22879 1955
rect 23305 1921 23339 1955
rect 23581 1921 23615 1955
rect 24041 1921 24075 1955
rect 26249 1921 26283 1955
rect 28457 1921 28491 1955
rect 30665 1921 30699 1955
rect 32873 1921 32907 1955
rect 35081 1921 35115 1955
rect 37473 1921 37507 1955
rect 41797 1921 41831 1955
rect 43637 1921 43671 1955
rect 44097 1921 44131 1955
rect 44557 1921 44591 1955
rect 22017 1785 22051 1819
rect 21465 1717 21499 1751
rect 23029 1717 23063 1751
rect 1593 1513 1627 1547
rect 19257 1513 19291 1547
rect 21189 1513 21223 1547
rect 22109 1513 22143 1547
rect 23397 1513 23431 1547
rect 27813 1513 27847 1547
rect 32229 1513 32263 1547
rect 34713 1513 34747 1547
rect 43269 1513 43303 1547
rect 45017 1513 45051 1547
rect 1409 1309 1443 1343
rect 3801 1309 3835 1343
rect 5733 1309 5767 1343
rect 7941 1309 7975 1343
rect 10149 1309 10183 1343
rect 12357 1309 12391 1343
rect 14749 1309 14783 1343
rect 16957 1309 16991 1343
rect 19441 1309 19475 1343
rect 21373 1309 21407 1343
rect 22293 1309 22327 1343
rect 23581 1309 23615 1343
rect 25789 1309 25823 1343
rect 27997 1309 28031 1343
rect 30205 1309 30239 1343
rect 32413 1309 32447 1343
rect 34897 1309 34931 1343
rect 36829 1309 36863 1343
rect 39037 1309 39071 1343
rect 41245 1309 41279 1343
rect 43453 1309 43487 1343
rect 45201 1309 45235 1343
rect 3985 1173 4019 1207
rect 5917 1173 5951 1207
rect 8125 1173 8159 1207
rect 10333 1173 10367 1207
rect 12541 1173 12575 1207
rect 14565 1173 14599 1207
rect 16773 1173 16807 1207
rect 25605 1173 25639 1207
rect 30021 1173 30055 1207
rect 36645 1173 36679 1207
rect 38853 1173 38887 1207
rect 41061 1173 41095 1207
<< metal1 >>
rect 13630 9976 13636 9988
rect 6886 9948 13636 9976
rect 6886 9908 6914 9948
rect 13630 9936 13636 9948
rect 13688 9936 13694 9988
rect 14918 9936 14924 9988
rect 14976 9976 14982 9988
rect 18322 9976 18328 9988
rect 14976 9948 18328 9976
rect 14976 9936 14982 9948
rect 18322 9936 18328 9948
rect 18380 9936 18386 9988
rect 18414 9936 18420 9988
rect 18472 9976 18478 9988
rect 19518 9976 19524 9988
rect 18472 9948 19524 9976
rect 18472 9936 18478 9948
rect 19518 9936 19524 9948
rect 19576 9936 19582 9988
rect 20622 9936 20628 9988
rect 20680 9976 20686 9988
rect 35710 9976 35716 9988
rect 20680 9948 35716 9976
rect 20680 9936 20686 9948
rect 35710 9936 35716 9948
rect 35768 9936 35774 9988
rect 5368 9880 6914 9908
rect 5368 9784 5396 9880
rect 8754 9868 8760 9920
rect 8812 9908 8818 9920
rect 14642 9908 14648 9920
rect 8812 9880 14648 9908
rect 8812 9868 8818 9880
rect 14642 9868 14648 9880
rect 14700 9868 14706 9920
rect 16482 9868 16488 9920
rect 16540 9908 16546 9920
rect 19886 9908 19892 9920
rect 16540 9880 19892 9908
rect 16540 9868 16546 9880
rect 19886 9868 19892 9880
rect 19944 9868 19950 9920
rect 9490 9800 9496 9852
rect 9548 9840 9554 9852
rect 14366 9840 14372 9852
rect 9548 9812 14372 9840
rect 9548 9800 9554 9812
rect 14366 9800 14372 9812
rect 14424 9800 14430 9852
rect 17678 9800 17684 9852
rect 17736 9840 17742 9852
rect 28902 9840 28908 9852
rect 17736 9812 28908 9840
rect 17736 9800 17742 9812
rect 28902 9800 28908 9812
rect 28960 9800 28966 9852
rect 5350 9732 5356 9784
rect 5408 9732 5414 9784
rect 8018 9732 8024 9784
rect 8076 9772 8082 9784
rect 14550 9772 14556 9784
rect 8076 9744 14556 9772
rect 8076 9732 8082 9744
rect 14550 9732 14556 9744
rect 14608 9732 14614 9784
rect 16390 9732 16396 9784
rect 16448 9772 16454 9784
rect 20070 9772 20076 9784
rect 16448 9744 20076 9772
rect 16448 9732 16454 9744
rect 20070 9732 20076 9744
rect 20128 9732 20134 9784
rect 22738 9732 22744 9784
rect 22796 9772 22802 9784
rect 22796 9744 28396 9772
rect 22796 9732 22802 9744
rect 7558 9664 7564 9716
rect 7616 9704 7622 9716
rect 17218 9704 17224 9716
rect 7616 9676 17224 9704
rect 7616 9664 7622 9676
rect 17218 9664 17224 9676
rect 17276 9664 17282 9716
rect 17310 9664 17316 9716
rect 17368 9704 17374 9716
rect 24118 9704 24124 9716
rect 17368 9676 24124 9704
rect 17368 9664 17374 9676
rect 24118 9664 24124 9676
rect 24176 9664 24182 9716
rect 5810 9596 5816 9648
rect 5868 9636 5874 9648
rect 14918 9636 14924 9648
rect 5868 9608 14924 9636
rect 5868 9596 5874 9608
rect 14918 9596 14924 9608
rect 14976 9596 14982 9648
rect 15010 9596 15016 9648
rect 15068 9636 15074 9648
rect 19334 9636 19340 9648
rect 15068 9608 19340 9636
rect 15068 9596 15074 9608
rect 19334 9596 19340 9608
rect 19392 9596 19398 9648
rect 19518 9596 19524 9648
rect 19576 9636 19582 9648
rect 28368 9636 28396 9744
rect 28534 9664 28540 9716
rect 28592 9704 28598 9716
rect 32306 9704 32312 9716
rect 28592 9676 32312 9704
rect 28592 9664 28598 9676
rect 32306 9664 32312 9676
rect 32364 9664 32370 9716
rect 36814 9636 36820 9648
rect 19576 9608 24348 9636
rect 28368 9608 36820 9636
rect 19576 9596 19582 9608
rect 19978 9568 19984 9580
rect 6886 9540 19984 9568
rect 4798 9188 4804 9240
rect 4856 9228 4862 9240
rect 6886 9228 6914 9540
rect 19978 9528 19984 9540
rect 20036 9528 20042 9580
rect 7374 9460 7380 9512
rect 7432 9500 7438 9512
rect 22370 9500 22376 9512
rect 7432 9472 22376 9500
rect 7432 9460 7438 9472
rect 22370 9460 22376 9472
rect 22428 9460 22434 9512
rect 17126 9432 17132 9444
rect 8864 9404 17132 9432
rect 8864 9240 8892 9404
rect 17126 9392 17132 9404
rect 17184 9392 17190 9444
rect 17218 9392 17224 9444
rect 17276 9432 17282 9444
rect 24026 9432 24032 9444
rect 17276 9404 24032 9432
rect 17276 9392 17282 9404
rect 24026 9392 24032 9404
rect 24084 9392 24090 9444
rect 24320 9432 24348 9608
rect 36814 9596 36820 9608
rect 36872 9596 36878 9648
rect 27430 9460 27436 9512
rect 27488 9500 27494 9512
rect 38654 9500 38660 9512
rect 27488 9472 38660 9500
rect 27488 9460 27494 9472
rect 38654 9460 38660 9472
rect 38712 9460 38718 9512
rect 34882 9432 34888 9444
rect 24320 9404 34888 9432
rect 34882 9392 34888 9404
rect 34940 9392 34946 9444
rect 36078 9392 36084 9444
rect 36136 9432 36142 9444
rect 36136 9404 41414 9432
rect 36136 9392 36142 9404
rect 26234 9364 26240 9376
rect 13096 9336 26240 9364
rect 13096 9308 13124 9336
rect 26234 9324 26240 9336
rect 26292 9324 26298 9376
rect 26326 9324 26332 9376
rect 26384 9364 26390 9376
rect 33502 9364 33508 9376
rect 26384 9336 33508 9364
rect 26384 9324 26390 9336
rect 33502 9324 33508 9336
rect 33560 9324 33566 9376
rect 33778 9324 33784 9376
rect 33836 9364 33842 9376
rect 33836 9336 41276 9364
rect 33836 9324 33842 9336
rect 13078 9256 13084 9308
rect 13136 9256 13142 9308
rect 13170 9256 13176 9308
rect 13228 9296 13234 9308
rect 16758 9296 16764 9308
rect 13228 9268 16764 9296
rect 13228 9256 13234 9268
rect 16758 9256 16764 9268
rect 16816 9256 16822 9308
rect 17310 9296 17316 9308
rect 17144 9268 17316 9296
rect 4856 9200 6914 9228
rect 4856 9188 4862 9200
rect 8846 9188 8852 9240
rect 8904 9188 8910 9240
rect 9030 9188 9036 9240
rect 9088 9228 9094 9240
rect 16942 9228 16948 9240
rect 9088 9200 16948 9228
rect 9088 9188 9094 9200
rect 16942 9188 16948 9200
rect 17000 9188 17006 9240
rect 17144 9160 17172 9268
rect 17310 9256 17316 9268
rect 17368 9256 17374 9308
rect 19334 9256 19340 9308
rect 19392 9296 19398 9308
rect 19886 9296 19892 9308
rect 19392 9268 19892 9296
rect 19392 9256 19398 9268
rect 19886 9256 19892 9268
rect 19944 9256 19950 9308
rect 28902 9256 28908 9308
rect 28960 9296 28966 9308
rect 35158 9296 35164 9308
rect 28960 9268 35164 9296
rect 28960 9256 28966 9268
rect 35158 9256 35164 9268
rect 35216 9256 35222 9308
rect 35342 9256 35348 9308
rect 35400 9296 35406 9308
rect 41046 9296 41052 9308
rect 35400 9268 41052 9296
rect 35400 9256 35406 9268
rect 41046 9256 41052 9268
rect 41104 9256 41110 9308
rect 6886 9132 17172 9160
rect 17236 9200 22876 9228
rect 6886 9024 6914 9132
rect 10502 9052 10508 9104
rect 10560 9092 10566 9104
rect 17236 9092 17264 9200
rect 18322 9120 18328 9172
rect 18380 9160 18386 9172
rect 22848 9160 22876 9200
rect 22922 9188 22928 9240
rect 22980 9228 22986 9240
rect 27430 9228 27436 9240
rect 22980 9200 27436 9228
rect 22980 9188 22986 9200
rect 27430 9188 27436 9200
rect 27488 9188 27494 9240
rect 27890 9228 27896 9240
rect 27540 9200 27896 9228
rect 27540 9160 27568 9200
rect 27890 9188 27896 9200
rect 27948 9188 27954 9240
rect 28092 9200 31754 9228
rect 18380 9132 22784 9160
rect 22848 9132 27568 9160
rect 18380 9120 18386 9132
rect 10560 9064 17264 9092
rect 10560 9052 10566 9064
rect 17770 9052 17776 9104
rect 17828 9092 17834 9104
rect 22756 9092 22784 9132
rect 17828 9064 22692 9092
rect 22756 9064 22876 9092
rect 17828 9052 17834 9064
rect 13170 9024 13176 9036
rect 3252 8996 6914 9024
rect 7300 8996 13176 9024
rect 3252 8832 3280 8996
rect 5442 8916 5448 8968
rect 5500 8956 5506 8968
rect 7300 8956 7328 8996
rect 13170 8984 13176 8996
rect 13228 8984 13234 9036
rect 22186 9024 22192 9036
rect 14016 8996 22192 9024
rect 14016 8956 14044 8996
rect 22186 8984 22192 8996
rect 22244 8984 22250 9036
rect 22664 9024 22692 9064
rect 22848 9024 22876 9064
rect 23014 9052 23020 9104
rect 23072 9092 23078 9104
rect 28092 9092 28120 9200
rect 31726 9160 31754 9200
rect 32766 9188 32772 9240
rect 32824 9228 32830 9240
rect 32824 9200 34744 9228
rect 32824 9188 32830 9200
rect 34606 9160 34612 9172
rect 31726 9132 34612 9160
rect 34606 9120 34612 9132
rect 34664 9120 34670 9172
rect 34716 9160 34744 9200
rect 41248 9160 41276 9336
rect 41386 9228 41414 9404
rect 43622 9228 43628 9240
rect 41386 9200 43628 9228
rect 43622 9188 43628 9200
rect 43680 9188 43686 9240
rect 42886 9160 42892 9172
rect 34716 9132 36860 9160
rect 41248 9132 42892 9160
rect 34054 9092 34060 9104
rect 23072 9064 28120 9092
rect 28966 9064 34060 9092
rect 23072 9052 23078 9064
rect 28966 9024 28994 9064
rect 34054 9052 34060 9064
rect 34112 9052 34118 9104
rect 22664 8996 22784 9024
rect 22848 8996 28994 9024
rect 36832 9024 36860 9132
rect 42886 9120 42892 9132
rect 42944 9120 42950 9172
rect 36832 8996 41414 9024
rect 20162 8956 20168 8968
rect 5500 8928 7328 8956
rect 8496 8928 14044 8956
rect 14108 8928 20168 8956
rect 5500 8916 5506 8928
rect 8496 8832 8524 8928
rect 14108 8888 14136 8928
rect 20162 8916 20168 8928
rect 20220 8916 20226 8968
rect 22756 8956 22784 8996
rect 22922 8956 22928 8968
rect 22756 8928 22928 8956
rect 22922 8916 22928 8928
rect 22980 8916 22986 8968
rect 27246 8916 27252 8968
rect 27304 8956 27310 8968
rect 33410 8956 33416 8968
rect 27304 8928 33416 8956
rect 27304 8916 27310 8928
rect 33410 8916 33416 8928
rect 33468 8916 33474 8968
rect 33870 8916 33876 8968
rect 33928 8956 33934 8968
rect 41386 8956 41414 8996
rect 43254 8956 43260 8968
rect 33928 8928 40724 8956
rect 41386 8928 43260 8956
rect 33928 8916 33934 8928
rect 11808 8860 14136 8888
rect 11808 8832 11836 8860
rect 14182 8848 14188 8900
rect 14240 8888 14246 8900
rect 16666 8888 16672 8900
rect 14240 8860 16672 8888
rect 14240 8848 14246 8860
rect 16666 8848 16672 8860
rect 16724 8848 16730 8900
rect 16758 8848 16764 8900
rect 16816 8888 16822 8900
rect 20254 8888 20260 8900
rect 16816 8860 20260 8888
rect 16816 8848 16822 8860
rect 20254 8848 20260 8860
rect 20312 8848 20318 8900
rect 23658 8848 23664 8900
rect 23716 8888 23722 8900
rect 31478 8888 31484 8900
rect 23716 8860 31484 8888
rect 23716 8848 23722 8860
rect 31478 8848 31484 8860
rect 31536 8848 31542 8900
rect 35618 8848 35624 8900
rect 35676 8888 35682 8900
rect 39942 8888 39948 8900
rect 35676 8860 39948 8888
rect 35676 8848 35682 8860
rect 39942 8848 39948 8860
rect 40000 8848 40006 8900
rect 40696 8832 40724 8928
rect 43254 8916 43260 8928
rect 43312 8916 43318 8968
rect 3234 8780 3240 8832
rect 3292 8780 3298 8832
rect 8478 8780 8484 8832
rect 8536 8780 8542 8832
rect 11790 8780 11796 8832
rect 11848 8780 11854 8832
rect 13538 8780 13544 8832
rect 13596 8820 13602 8832
rect 17770 8820 17776 8832
rect 13596 8792 17776 8820
rect 13596 8780 13602 8792
rect 17770 8780 17776 8792
rect 17828 8780 17834 8832
rect 19058 8780 19064 8832
rect 19116 8820 19122 8832
rect 22462 8820 22468 8832
rect 19116 8792 22468 8820
rect 19116 8780 19122 8792
rect 22462 8780 22468 8792
rect 22520 8780 22526 8832
rect 23750 8780 23756 8832
rect 23808 8820 23814 8832
rect 32398 8820 32404 8832
rect 23808 8792 32404 8820
rect 23808 8780 23814 8792
rect 32398 8780 32404 8792
rect 32456 8780 32462 8832
rect 35986 8780 35992 8832
rect 36044 8820 36050 8832
rect 40494 8820 40500 8832
rect 36044 8792 40500 8820
rect 36044 8780 36050 8792
rect 40494 8780 40500 8792
rect 40552 8780 40558 8832
rect 40678 8780 40684 8832
rect 40736 8780 40742 8832
rect 1104 8730 45696 8752
rect 1104 8678 12058 8730
rect 12110 8678 12122 8730
rect 12174 8678 12186 8730
rect 12238 8678 12250 8730
rect 12302 8678 12314 8730
rect 12366 8678 23166 8730
rect 23218 8678 23230 8730
rect 23282 8678 23294 8730
rect 23346 8678 23358 8730
rect 23410 8678 23422 8730
rect 23474 8678 34274 8730
rect 34326 8678 34338 8730
rect 34390 8678 34402 8730
rect 34454 8678 34466 8730
rect 34518 8678 34530 8730
rect 34582 8678 45382 8730
rect 45434 8678 45446 8730
rect 45498 8678 45510 8730
rect 45562 8678 45574 8730
rect 45626 8678 45638 8730
rect 45690 8678 45696 8730
rect 1104 8656 45696 8678
rect 2133 8619 2191 8625
rect 2133 8585 2145 8619
rect 2179 8616 2191 8619
rect 2314 8616 2320 8628
rect 2179 8588 2320 8616
rect 2179 8585 2191 8588
rect 2133 8579 2191 8585
rect 2314 8576 2320 8588
rect 2372 8576 2378 8628
rect 2777 8619 2835 8625
rect 2777 8585 2789 8619
rect 2823 8585 2835 8619
rect 2777 8579 2835 8585
rect 3513 8619 3571 8625
rect 3513 8585 3525 8619
rect 3559 8616 3571 8619
rect 4154 8616 4160 8628
rect 3559 8588 4160 8616
rect 3559 8585 3571 8588
rect 3513 8579 3571 8585
rect 750 8508 756 8560
rect 808 8548 814 8560
rect 2792 8548 2820 8579
rect 4154 8576 4160 8588
rect 4212 8576 4218 8628
rect 4525 8619 4583 8625
rect 4525 8585 4537 8619
rect 4571 8616 4583 8619
rect 4890 8616 4896 8628
rect 4571 8588 4896 8616
rect 4571 8585 4583 8588
rect 4525 8579 4583 8585
rect 4890 8576 4896 8588
rect 4948 8576 4954 8628
rect 4985 8619 5043 8625
rect 4985 8585 4997 8619
rect 5031 8616 5043 8619
rect 5258 8616 5264 8628
rect 5031 8588 5264 8616
rect 5031 8585 5043 8588
rect 4985 8579 5043 8585
rect 5258 8576 5264 8588
rect 5316 8576 5322 8628
rect 5442 8576 5448 8628
rect 5500 8576 5506 8628
rect 5537 8619 5595 8625
rect 5537 8585 5549 8619
rect 5583 8616 5595 8619
rect 5626 8616 5632 8628
rect 5583 8588 5632 8616
rect 5583 8585 5595 8588
rect 5537 8579 5595 8585
rect 5626 8576 5632 8588
rect 5684 8576 5690 8628
rect 5994 8576 6000 8628
rect 6052 8616 6058 8628
rect 6549 8619 6607 8625
rect 6549 8616 6561 8619
rect 6052 8588 6561 8616
rect 6052 8576 6058 8588
rect 6549 8585 6561 8588
rect 6595 8585 6607 8619
rect 6549 8579 6607 8585
rect 6730 8576 6736 8628
rect 6788 8576 6794 8628
rect 7006 8576 7012 8628
rect 7064 8576 7070 8628
rect 7745 8619 7803 8625
rect 7745 8585 7757 8619
rect 7791 8616 7803 8619
rect 7834 8616 7840 8628
rect 7791 8588 7840 8616
rect 7791 8585 7803 8588
rect 7745 8579 7803 8585
rect 7834 8576 7840 8588
rect 7892 8576 7898 8628
rect 8110 8576 8116 8628
rect 8168 8576 8174 8628
rect 8570 8576 8576 8628
rect 8628 8616 8634 8628
rect 8665 8619 8723 8625
rect 8665 8616 8677 8619
rect 8628 8588 8677 8616
rect 8628 8576 8634 8588
rect 8665 8585 8677 8588
rect 8711 8585 8723 8619
rect 8665 8579 8723 8585
rect 9217 8619 9275 8625
rect 9217 8585 9229 8619
rect 9263 8616 9275 8619
rect 9306 8616 9312 8628
rect 9263 8588 9312 8616
rect 9263 8585 9275 8588
rect 9217 8579 9275 8585
rect 9306 8576 9312 8588
rect 9364 8576 9370 8628
rect 9766 8576 9772 8628
rect 9824 8576 9830 8628
rect 10321 8619 10379 8625
rect 10321 8585 10333 8619
rect 10367 8616 10379 8619
rect 10410 8616 10416 8628
rect 10367 8588 10416 8616
rect 10367 8585 10379 8588
rect 10321 8579 10379 8585
rect 10410 8576 10416 8588
rect 10468 8576 10474 8628
rect 10689 8619 10747 8625
rect 10689 8585 10701 8619
rect 10735 8616 10747 8619
rect 10778 8616 10784 8628
rect 10735 8588 10784 8616
rect 10735 8585 10747 8588
rect 10689 8579 10747 8585
rect 10778 8576 10784 8588
rect 10836 8576 10842 8628
rect 10888 8588 11100 8616
rect 808 8520 2820 8548
rect 808 8508 814 8520
rect 3234 8508 3240 8560
rect 3292 8508 3298 8560
rect 5460 8548 5488 8576
rect 4724 8520 5488 8548
rect 4724 8489 4752 8520
rect 5810 8508 5816 8560
rect 5868 8508 5874 8560
rect 6181 8551 6239 8557
rect 6181 8517 6193 8551
rect 6227 8548 6239 8551
rect 6748 8548 6776 8576
rect 6227 8520 6776 8548
rect 6917 8551 6975 8557
rect 6227 8517 6239 8520
rect 6181 8511 6239 8517
rect 6917 8517 6929 8551
rect 6963 8548 6975 8551
rect 8846 8548 8852 8560
rect 6963 8520 8852 8548
rect 6963 8517 6975 8520
rect 6917 8511 6975 8517
rect 8846 8508 8852 8520
rect 8904 8508 8910 8560
rect 10888 8548 10916 8588
rect 8956 8520 10916 8548
rect 10965 8551 11023 8557
rect 2317 8483 2375 8489
rect 2317 8449 2329 8483
rect 2363 8449 2375 8483
rect 2317 8443 2375 8449
rect 2685 8483 2743 8489
rect 2685 8449 2697 8483
rect 2731 8449 2743 8483
rect 2685 8443 2743 8449
rect 4157 8483 4215 8489
rect 4157 8449 4169 8483
rect 4203 8480 4215 8483
rect 4709 8483 4767 8489
rect 4709 8480 4721 8483
rect 4203 8452 4721 8480
rect 4203 8449 4215 8452
rect 4157 8443 4215 8449
rect 4709 8449 4721 8452
rect 4755 8449 4767 8483
rect 4709 8443 4767 8449
rect 1765 8347 1823 8353
rect 1765 8313 1777 8347
rect 1811 8344 1823 8347
rect 2332 8344 2360 8443
rect 2700 8412 2728 8443
rect 4798 8440 4804 8492
rect 4856 8440 4862 8492
rect 5261 8483 5319 8489
rect 5261 8449 5273 8483
rect 5307 8480 5319 8483
rect 5350 8480 5356 8492
rect 5307 8452 5356 8480
rect 5307 8449 5319 8452
rect 5261 8443 5319 8449
rect 5350 8440 5356 8452
rect 5408 8440 5414 8492
rect 6365 8483 6423 8489
rect 6365 8449 6377 8483
rect 6411 8480 6423 8483
rect 7374 8480 7380 8492
rect 6411 8452 7380 8480
rect 6411 8449 6423 8452
rect 6365 8443 6423 8449
rect 7374 8440 7380 8452
rect 7432 8440 7438 8492
rect 7558 8440 7564 8492
rect 7616 8440 7622 8492
rect 8018 8440 8024 8492
rect 8076 8440 8082 8492
rect 8478 8440 8484 8492
rect 8536 8440 8542 8492
rect 8754 8440 8760 8492
rect 8812 8440 8818 8492
rect 8772 8412 8800 8440
rect 2700 8384 8800 8412
rect 8956 8344 8984 8520
rect 10965 8517 10977 8551
rect 11011 8517 11023 8551
rect 11072 8548 11100 8588
rect 11238 8576 11244 8628
rect 11296 8576 11302 8628
rect 11974 8576 11980 8628
rect 12032 8576 12038 8628
rect 12526 8576 12532 8628
rect 12584 8576 12590 8628
rect 13265 8619 13323 8625
rect 13265 8585 13277 8619
rect 13311 8616 13323 8619
rect 13354 8616 13360 8628
rect 13311 8588 13360 8616
rect 13311 8585 13323 8588
rect 13265 8579 13323 8585
rect 13354 8576 13360 8588
rect 13412 8576 13418 8628
rect 13630 8576 13636 8628
rect 13688 8576 13694 8628
rect 14369 8619 14427 8625
rect 14369 8585 14381 8619
rect 14415 8616 14427 8619
rect 14458 8616 14464 8628
rect 14415 8588 14464 8616
rect 14415 8585 14427 8588
rect 14369 8579 14427 8585
rect 14458 8576 14464 8588
rect 14516 8576 14522 8628
rect 14737 8619 14795 8625
rect 14737 8585 14749 8619
rect 14783 8616 14795 8619
rect 14826 8616 14832 8628
rect 14783 8588 14832 8616
rect 14783 8585 14795 8588
rect 14737 8579 14795 8585
rect 14826 8576 14832 8588
rect 14884 8576 14890 8628
rect 15286 8576 15292 8628
rect 15344 8576 15350 8628
rect 15562 8576 15568 8628
rect 15620 8616 15626 8628
rect 15657 8619 15715 8625
rect 15657 8616 15669 8619
rect 15620 8588 15669 8616
rect 15620 8576 15626 8588
rect 15657 8585 15669 8588
rect 15703 8585 15715 8619
rect 15657 8579 15715 8585
rect 15930 8576 15936 8628
rect 15988 8616 15994 8628
rect 16025 8619 16083 8625
rect 16025 8616 16037 8619
rect 15988 8588 16037 8616
rect 15988 8576 15994 8588
rect 16025 8585 16037 8588
rect 16071 8585 16083 8619
rect 16025 8579 16083 8585
rect 16298 8576 16304 8628
rect 16356 8616 16362 8628
rect 16393 8619 16451 8625
rect 16393 8616 16405 8619
rect 16356 8588 16405 8616
rect 16356 8576 16362 8588
rect 16393 8585 16405 8588
rect 16439 8585 16451 8619
rect 16393 8579 16451 8585
rect 16850 8576 16856 8628
rect 16908 8576 16914 8628
rect 17402 8576 17408 8628
rect 17460 8616 17466 8628
rect 17497 8619 17555 8625
rect 17497 8616 17509 8619
rect 17460 8588 17509 8616
rect 17460 8576 17466 8588
rect 17497 8585 17509 8588
rect 17543 8585 17555 8619
rect 17497 8579 17555 8585
rect 18046 8576 18052 8628
rect 18104 8576 18110 8628
rect 18138 8576 18144 8628
rect 18196 8616 18202 8628
rect 18417 8619 18475 8625
rect 18417 8616 18429 8619
rect 18196 8588 18429 8616
rect 18196 8576 18202 8588
rect 18417 8585 18429 8588
rect 18463 8585 18475 8619
rect 18417 8579 18475 8585
rect 18506 8576 18512 8628
rect 18564 8616 18570 8628
rect 18785 8619 18843 8625
rect 18785 8616 18797 8619
rect 18564 8588 18797 8616
rect 18564 8576 18570 8588
rect 18785 8585 18797 8588
rect 18831 8585 18843 8619
rect 18785 8579 18843 8585
rect 19150 8576 19156 8628
rect 19208 8616 19214 8628
rect 19889 8619 19947 8625
rect 19889 8616 19901 8619
rect 19208 8588 19901 8616
rect 19208 8576 19214 8588
rect 19889 8585 19901 8588
rect 19935 8585 19947 8619
rect 19889 8579 19947 8585
rect 20254 8576 20260 8628
rect 20312 8616 20318 8628
rect 20625 8619 20683 8625
rect 20625 8616 20637 8619
rect 20312 8588 20637 8616
rect 20312 8576 20318 8588
rect 20625 8585 20637 8588
rect 20671 8585 20683 8619
rect 22833 8619 22891 8625
rect 22833 8616 22845 8619
rect 20625 8579 20683 8585
rect 20732 8588 22845 8616
rect 11072 8520 11192 8548
rect 10965 8511 11023 8517
rect 9030 8440 9036 8492
rect 9088 8440 9094 8492
rect 9490 8440 9496 8492
rect 9548 8440 9554 8492
rect 10137 8483 10195 8489
rect 10137 8449 10149 8483
rect 10183 8480 10195 8483
rect 10410 8480 10416 8492
rect 10183 8452 10416 8480
rect 10183 8449 10195 8452
rect 10137 8443 10195 8449
rect 10410 8440 10416 8452
rect 10468 8440 10474 8492
rect 10502 8440 10508 8492
rect 10560 8440 10566 8492
rect 10980 8412 11008 8511
rect 11164 8480 11192 8520
rect 11790 8508 11796 8560
rect 11848 8548 11854 8560
rect 11885 8551 11943 8557
rect 11885 8548 11897 8551
rect 11848 8520 11897 8548
rect 11848 8508 11854 8520
rect 11885 8517 11897 8520
rect 11931 8517 11943 8551
rect 11885 8511 11943 8517
rect 12434 8508 12440 8560
rect 12492 8508 12498 8560
rect 14568 8520 19932 8548
rect 12618 8480 12624 8492
rect 11164 8452 12624 8480
rect 12618 8440 12624 8452
rect 12676 8440 12682 8492
rect 13078 8440 13084 8492
rect 13136 8440 13142 8492
rect 13538 8440 13544 8492
rect 13596 8440 13602 8492
rect 14182 8440 14188 8492
rect 14240 8440 14246 8492
rect 14568 8489 14596 8520
rect 14553 8483 14611 8489
rect 14553 8449 14565 8483
rect 14599 8449 14611 8483
rect 14553 8443 14611 8449
rect 15010 8440 15016 8492
rect 15068 8440 15074 8492
rect 15470 8440 15476 8492
rect 15528 8440 15534 8492
rect 15841 8483 15899 8489
rect 15841 8449 15853 8483
rect 15887 8480 15899 8483
rect 16114 8480 16120 8492
rect 15887 8452 16120 8480
rect 15887 8449 15899 8452
rect 15841 8443 15899 8449
rect 16114 8440 16120 8452
rect 16172 8440 16178 8492
rect 16209 8483 16267 8489
rect 16209 8449 16221 8483
rect 16255 8449 16267 8483
rect 16209 8443 16267 8449
rect 14366 8412 14372 8424
rect 10980 8384 14372 8412
rect 14366 8372 14372 8384
rect 14424 8372 14430 8424
rect 1811 8316 8984 8344
rect 16224 8344 16252 8443
rect 16758 8440 16764 8492
rect 16816 8440 16822 8492
rect 17310 8440 17316 8492
rect 17368 8440 17374 8492
rect 17494 8440 17500 8492
rect 17552 8480 17558 8492
rect 17773 8483 17831 8489
rect 17773 8480 17785 8483
rect 17552 8452 17785 8480
rect 17552 8440 17558 8452
rect 17773 8449 17785 8452
rect 17819 8449 17831 8483
rect 17773 8443 17831 8449
rect 18230 8440 18236 8492
rect 18288 8440 18294 8492
rect 18601 8483 18659 8489
rect 18601 8449 18613 8483
rect 18647 8480 18659 8483
rect 18874 8480 18880 8492
rect 18647 8452 18880 8480
rect 18647 8449 18659 8452
rect 18601 8443 18659 8449
rect 18874 8440 18880 8452
rect 18932 8440 18938 8492
rect 19610 8440 19616 8492
rect 19668 8440 19674 8492
rect 19797 8483 19855 8489
rect 19797 8449 19809 8483
rect 19843 8449 19855 8483
rect 19797 8443 19855 8449
rect 19150 8372 19156 8424
rect 19208 8412 19214 8424
rect 19812 8412 19840 8443
rect 19208 8384 19840 8412
rect 19904 8412 19932 8520
rect 19978 8508 19984 8560
rect 20036 8548 20042 8560
rect 20732 8548 20760 8588
rect 22833 8585 22845 8588
rect 22879 8585 22891 8619
rect 22833 8579 22891 8585
rect 22922 8576 22928 8628
rect 22980 8576 22986 8628
rect 23385 8619 23443 8625
rect 23385 8585 23397 8619
rect 23431 8585 23443 8619
rect 23385 8579 23443 8585
rect 23400 8548 23428 8579
rect 23474 8576 23480 8628
rect 23532 8616 23538 8628
rect 23532 8588 30236 8616
rect 23532 8576 23538 8588
rect 20036 8520 20760 8548
rect 22664 8520 23428 8548
rect 23492 8520 24072 8548
rect 20036 8508 20042 8520
rect 20530 8440 20536 8492
rect 20588 8440 20594 8492
rect 20806 8440 20812 8492
rect 20864 8440 20870 8492
rect 21082 8440 21088 8492
rect 21140 8440 21146 8492
rect 21358 8440 21364 8492
rect 21416 8440 21422 8492
rect 21634 8440 21640 8492
rect 21692 8440 21698 8492
rect 22002 8440 22008 8492
rect 22060 8440 22066 8492
rect 22094 8440 22100 8492
rect 22152 8440 22158 8492
rect 22278 8440 22284 8492
rect 22336 8440 22342 8492
rect 22370 8440 22376 8492
rect 22428 8440 22434 8492
rect 22554 8440 22560 8492
rect 22612 8440 22618 8492
rect 22664 8489 22692 8520
rect 22649 8483 22707 8489
rect 22649 8449 22661 8483
rect 22695 8449 22707 8483
rect 22649 8443 22707 8449
rect 22830 8440 22836 8492
rect 22888 8480 22894 8492
rect 23109 8483 23167 8489
rect 23109 8480 23121 8483
rect 22888 8452 23121 8480
rect 22888 8440 22894 8452
rect 23109 8449 23121 8452
rect 23155 8449 23167 8483
rect 23492 8480 23520 8520
rect 23109 8443 23167 8449
rect 23216 8452 23520 8480
rect 22112 8412 22140 8440
rect 22388 8412 22416 8440
rect 19904 8384 22140 8412
rect 22296 8384 22416 8412
rect 19208 8372 19214 8384
rect 22296 8356 22324 8384
rect 23014 8372 23020 8424
rect 23072 8412 23078 8424
rect 23216 8412 23244 8452
rect 23566 8440 23572 8492
rect 23624 8440 23630 8492
rect 23750 8440 23756 8492
rect 23808 8440 23814 8492
rect 23072 8384 23244 8412
rect 23072 8372 23078 8384
rect 16224 8316 20484 8344
rect 1811 8313 1823 8316
rect 1765 8307 1823 8313
rect 19426 8236 19432 8288
rect 19484 8236 19490 8288
rect 20346 8236 20352 8288
rect 20404 8236 20410 8288
rect 20456 8276 20484 8316
rect 20530 8304 20536 8356
rect 20588 8344 20594 8356
rect 20901 8347 20959 8353
rect 20901 8344 20913 8347
rect 20588 8316 20913 8344
rect 20588 8304 20594 8316
rect 20901 8313 20913 8316
rect 20947 8313 20959 8347
rect 21542 8344 21548 8356
rect 20901 8307 20959 8313
rect 21100 8316 21548 8344
rect 21100 8276 21128 8316
rect 21542 8304 21548 8316
rect 21600 8304 21606 8356
rect 21910 8304 21916 8356
rect 21968 8344 21974 8356
rect 22097 8347 22155 8353
rect 22097 8344 22109 8347
rect 21968 8316 22109 8344
rect 21968 8304 21974 8316
rect 22097 8313 22109 8316
rect 22143 8313 22155 8347
rect 22097 8307 22155 8313
rect 22186 8304 22192 8356
rect 22244 8304 22250 8356
rect 22278 8304 22284 8356
rect 22336 8304 22342 8356
rect 22370 8304 22376 8356
rect 22428 8304 22434 8356
rect 22830 8304 22836 8356
rect 22888 8344 22894 8356
rect 23842 8344 23848 8356
rect 22888 8316 23848 8344
rect 22888 8304 22894 8316
rect 23842 8304 23848 8316
rect 23900 8304 23906 8356
rect 23934 8304 23940 8356
rect 23992 8304 23998 8356
rect 24044 8353 24072 8520
rect 24394 8508 24400 8560
rect 24452 8548 24458 8560
rect 24452 8520 24808 8548
rect 24452 8508 24458 8520
rect 24213 8483 24271 8489
rect 24213 8449 24225 8483
rect 24259 8480 24271 8483
rect 24302 8480 24308 8492
rect 24259 8452 24308 8480
rect 24259 8449 24271 8452
rect 24213 8443 24271 8449
rect 24302 8440 24308 8452
rect 24360 8440 24366 8492
rect 24670 8440 24676 8492
rect 24728 8440 24734 8492
rect 24780 8480 24808 8520
rect 24854 8508 24860 8560
rect 24912 8548 24918 8560
rect 24912 8520 25268 8548
rect 24912 8508 24918 8520
rect 25240 8489 25268 8520
rect 26970 8508 26976 8560
rect 27028 8548 27034 8560
rect 27028 8520 27476 8548
rect 27028 8508 27034 8520
rect 24949 8483 25007 8489
rect 24949 8480 24961 8483
rect 24780 8452 24961 8480
rect 24949 8449 24961 8452
rect 24995 8449 25007 8483
rect 24949 8443 25007 8449
rect 25225 8483 25283 8489
rect 25225 8449 25237 8483
rect 25271 8449 25283 8483
rect 25225 8443 25283 8449
rect 25498 8440 25504 8492
rect 25556 8440 25562 8492
rect 25774 8440 25780 8492
rect 25832 8440 25838 8492
rect 26142 8440 26148 8492
rect 26200 8440 26206 8492
rect 26510 8440 26516 8492
rect 26568 8440 26574 8492
rect 26602 8440 26608 8492
rect 26660 8480 26666 8492
rect 27448 8489 27476 8520
rect 29546 8508 29552 8560
rect 29604 8548 29610 8560
rect 30208 8548 30236 8588
rect 30282 8576 30288 8628
rect 30340 8616 30346 8628
rect 30340 8588 30604 8616
rect 30340 8576 30346 8588
rect 29604 8520 30052 8548
rect 30208 8520 30512 8548
rect 29604 8508 29610 8520
rect 27157 8483 27215 8489
rect 27157 8480 27169 8483
rect 26660 8452 27169 8480
rect 26660 8440 26666 8452
rect 27157 8449 27169 8452
rect 27203 8449 27215 8483
rect 27157 8443 27215 8449
rect 27433 8483 27491 8489
rect 27433 8449 27445 8483
rect 27479 8449 27491 8483
rect 27433 8443 27491 8449
rect 27522 8440 27528 8492
rect 27580 8480 27586 8492
rect 27709 8483 27767 8489
rect 27709 8480 27721 8483
rect 27580 8452 27721 8480
rect 27580 8440 27586 8452
rect 27709 8449 27721 8452
rect 27755 8449 27767 8483
rect 27709 8443 27767 8449
rect 27982 8440 27988 8492
rect 28040 8440 28046 8492
rect 28350 8440 28356 8492
rect 28408 8440 28414 8492
rect 28718 8440 28724 8492
rect 28776 8440 28782 8492
rect 28810 8440 28816 8492
rect 28868 8480 28874 8492
rect 29089 8483 29147 8489
rect 29089 8480 29101 8483
rect 28868 8452 29101 8480
rect 28868 8440 28874 8452
rect 29089 8449 29101 8452
rect 29135 8449 29147 8483
rect 29089 8443 29147 8449
rect 29178 8440 29184 8492
rect 29236 8480 29242 8492
rect 30024 8489 30052 8520
rect 29733 8483 29791 8489
rect 29733 8480 29745 8483
rect 29236 8452 29745 8480
rect 29236 8440 29242 8452
rect 29733 8449 29745 8452
rect 29779 8449 29791 8483
rect 29733 8443 29791 8449
rect 30009 8483 30067 8489
rect 30009 8449 30021 8483
rect 30055 8449 30067 8483
rect 30009 8443 30067 8449
rect 30282 8440 30288 8492
rect 30340 8440 30346 8492
rect 24486 8372 24492 8424
rect 24544 8412 24550 8424
rect 30374 8412 30380 8424
rect 24544 8384 30380 8412
rect 24544 8372 24550 8384
rect 30374 8372 30380 8384
rect 30432 8372 30438 8424
rect 30484 8412 30512 8520
rect 30576 8513 30604 8588
rect 31478 8576 31484 8628
rect 31536 8576 31542 8628
rect 32306 8576 32312 8628
rect 32364 8576 32370 8628
rect 32398 8576 32404 8628
rect 32456 8576 32462 8628
rect 32490 8576 32496 8628
rect 32548 8616 32554 8628
rect 33137 8619 33195 8625
rect 33137 8616 33149 8619
rect 32548 8588 33149 8616
rect 32548 8576 32554 8588
rect 33137 8585 33149 8588
rect 33183 8585 33195 8619
rect 33137 8579 33195 8585
rect 33502 8576 33508 8628
rect 33560 8576 33566 8628
rect 33873 8619 33931 8625
rect 33873 8585 33885 8619
rect 33919 8585 33931 8619
rect 33873 8579 33931 8585
rect 30561 8507 30619 8513
rect 30650 8508 30656 8560
rect 30708 8548 30714 8560
rect 33888 8548 33916 8579
rect 34054 8576 34060 8628
rect 34112 8616 34118 8628
rect 34241 8619 34299 8625
rect 34241 8616 34253 8619
rect 34112 8588 34253 8616
rect 34112 8576 34118 8588
rect 34241 8585 34253 8588
rect 34287 8585 34299 8619
rect 34241 8579 34299 8585
rect 34606 8576 34612 8628
rect 34664 8576 34670 8628
rect 34790 8576 34796 8628
rect 34848 8616 34854 8628
rect 35437 8619 35495 8625
rect 35437 8616 35449 8619
rect 34848 8588 35449 8616
rect 34848 8576 34854 8588
rect 35437 8585 35449 8588
rect 35483 8585 35495 8619
rect 35437 8579 35495 8585
rect 35710 8576 35716 8628
rect 35768 8576 35774 8628
rect 35894 8576 35900 8628
rect 35952 8616 35958 8628
rect 38289 8619 38347 8625
rect 38289 8616 38301 8619
rect 35952 8588 38301 8616
rect 35952 8576 35958 8588
rect 38289 8585 38301 8588
rect 38335 8585 38347 8619
rect 38289 8579 38347 8585
rect 38654 8576 38660 8628
rect 38712 8576 38718 8628
rect 39022 8576 39028 8628
rect 39080 8576 39086 8628
rect 39114 8576 39120 8628
rect 39172 8616 39178 8628
rect 39577 8619 39635 8625
rect 39577 8616 39589 8619
rect 39172 8588 39589 8616
rect 39172 8576 39178 8588
rect 39577 8585 39589 8588
rect 39623 8585 39635 8619
rect 39577 8579 39635 8585
rect 39758 8576 39764 8628
rect 39816 8616 39822 8628
rect 40037 8619 40095 8625
rect 40037 8616 40049 8619
rect 39816 8588 40049 8616
rect 39816 8576 39822 8588
rect 40037 8585 40049 8588
rect 40083 8585 40095 8619
rect 40037 8579 40095 8585
rect 40589 8619 40647 8625
rect 40589 8585 40601 8619
rect 40635 8585 40647 8619
rect 40589 8579 40647 8585
rect 30708 8520 33916 8548
rect 34624 8548 34652 8576
rect 34624 8520 36492 8548
rect 30708 8508 30714 8520
rect 30561 8473 30573 8507
rect 30607 8473 30619 8507
rect 30561 8467 30619 8473
rect 30926 8440 30932 8492
rect 30984 8440 30990 8492
rect 31294 8440 31300 8492
rect 31352 8440 31358 8492
rect 31662 8440 31668 8492
rect 31720 8440 31726 8492
rect 31754 8440 31760 8492
rect 31812 8480 31818 8492
rect 32125 8483 32183 8489
rect 32125 8480 32137 8483
rect 31812 8452 32137 8480
rect 31812 8440 31818 8452
rect 32125 8449 32137 8452
rect 32171 8449 32183 8483
rect 32125 8443 32183 8449
rect 32306 8440 32312 8492
rect 32364 8480 32370 8492
rect 32585 8483 32643 8489
rect 32585 8480 32597 8483
rect 32364 8452 32597 8480
rect 32364 8440 32370 8452
rect 32585 8449 32597 8452
rect 32631 8449 32643 8483
rect 32585 8443 32643 8449
rect 32674 8440 32680 8492
rect 32732 8440 32738 8492
rect 32953 8483 33011 8489
rect 32953 8449 32965 8483
rect 32999 8449 33011 8483
rect 32953 8443 33011 8449
rect 32968 8412 32996 8443
rect 33318 8440 33324 8492
rect 33376 8440 33382 8492
rect 33686 8440 33692 8492
rect 33744 8440 33750 8492
rect 34054 8440 34060 8492
rect 34112 8440 34118 8492
rect 34146 8440 34152 8492
rect 34204 8480 34210 8492
rect 34701 8483 34759 8489
rect 34701 8480 34713 8483
rect 34204 8452 34713 8480
rect 34204 8440 34210 8452
rect 34701 8449 34713 8452
rect 34747 8449 34759 8483
rect 34701 8443 34759 8449
rect 34974 8440 34980 8492
rect 35032 8440 35038 8492
rect 35250 8440 35256 8492
rect 35308 8440 35314 8492
rect 35526 8440 35532 8492
rect 35584 8440 35590 8492
rect 35802 8440 35808 8492
rect 35860 8480 35866 8492
rect 35897 8483 35955 8489
rect 35897 8480 35909 8483
rect 35860 8452 35909 8480
rect 35860 8440 35866 8452
rect 35897 8449 35909 8452
rect 35943 8449 35955 8483
rect 35897 8443 35955 8449
rect 36262 8440 36268 8492
rect 36320 8440 36326 8492
rect 33042 8412 33048 8424
rect 30484 8384 32904 8412
rect 32968 8384 33048 8412
rect 24029 8347 24087 8353
rect 24029 8313 24041 8347
rect 24075 8313 24087 8347
rect 24029 8307 24087 8313
rect 25866 8304 25872 8356
rect 25924 8344 25930 8356
rect 26329 8347 26387 8353
rect 26329 8344 26341 8347
rect 25924 8316 26341 8344
rect 25924 8304 25930 8316
rect 26329 8313 26341 8316
rect 26375 8313 26387 8347
rect 26973 8347 27031 8353
rect 26973 8344 26985 8347
rect 26329 8307 26387 8313
rect 26436 8316 26985 8344
rect 20456 8248 21128 8276
rect 21174 8236 21180 8288
rect 21232 8236 21238 8288
rect 21450 8236 21456 8288
rect 21508 8236 21514 8288
rect 21818 8236 21824 8288
rect 21876 8236 21882 8288
rect 22204 8276 22232 8304
rect 23382 8276 23388 8288
rect 22204 8248 23388 8276
rect 23382 8236 23388 8248
rect 23440 8236 23446 8288
rect 23474 8236 23480 8288
rect 23532 8276 23538 8288
rect 24302 8276 24308 8288
rect 23532 8248 24308 8276
rect 23532 8236 23538 8248
rect 24302 8236 24308 8248
rect 24360 8236 24366 8288
rect 24486 8236 24492 8288
rect 24544 8236 24550 8288
rect 24762 8236 24768 8288
rect 24820 8236 24826 8288
rect 25038 8236 25044 8288
rect 25096 8236 25102 8288
rect 25130 8236 25136 8288
rect 25188 8276 25194 8288
rect 25317 8279 25375 8285
rect 25317 8276 25329 8279
rect 25188 8248 25329 8276
rect 25188 8236 25194 8248
rect 25317 8245 25329 8248
rect 25363 8245 25375 8279
rect 25317 8239 25375 8245
rect 25406 8236 25412 8288
rect 25464 8276 25470 8288
rect 25593 8279 25651 8285
rect 25593 8276 25605 8279
rect 25464 8248 25605 8276
rect 25464 8236 25470 8248
rect 25593 8245 25605 8248
rect 25639 8245 25651 8279
rect 25593 8239 25651 8245
rect 25682 8236 25688 8288
rect 25740 8276 25746 8288
rect 25961 8279 26019 8285
rect 25961 8276 25973 8279
rect 25740 8248 25973 8276
rect 25740 8236 25746 8248
rect 25961 8245 25973 8248
rect 26007 8245 26019 8279
rect 25961 8239 26019 8245
rect 26142 8236 26148 8288
rect 26200 8276 26206 8288
rect 26436 8276 26464 8316
rect 26973 8313 26985 8316
rect 27019 8313 27031 8347
rect 26973 8307 27031 8313
rect 27614 8304 27620 8356
rect 27672 8344 27678 8356
rect 28169 8347 28227 8353
rect 28169 8344 28181 8347
rect 27672 8316 28181 8344
rect 27672 8304 27678 8316
rect 28169 8313 28181 8316
rect 28215 8313 28227 8347
rect 28169 8307 28227 8313
rect 28258 8304 28264 8356
rect 28316 8344 28322 8356
rect 32490 8344 32496 8356
rect 28316 8316 32496 8344
rect 28316 8304 28322 8316
rect 32490 8304 32496 8316
rect 32548 8304 32554 8356
rect 26200 8248 26464 8276
rect 26200 8236 26206 8248
rect 26602 8236 26608 8288
rect 26660 8276 26666 8288
rect 27249 8279 27307 8285
rect 27249 8276 27261 8279
rect 26660 8248 27261 8276
rect 26660 8236 26666 8248
rect 27249 8245 27261 8248
rect 27295 8245 27307 8279
rect 27249 8239 27307 8245
rect 27522 8236 27528 8288
rect 27580 8236 27586 8288
rect 27798 8236 27804 8288
rect 27856 8236 27862 8288
rect 28534 8236 28540 8288
rect 28592 8236 28598 8288
rect 28626 8236 28632 8288
rect 28684 8276 28690 8288
rect 28905 8279 28963 8285
rect 28905 8276 28917 8279
rect 28684 8248 28917 8276
rect 28684 8236 28690 8248
rect 28905 8245 28917 8248
rect 28951 8245 28963 8279
rect 28905 8239 28963 8245
rect 29546 8236 29552 8288
rect 29604 8236 29610 8288
rect 29822 8236 29828 8288
rect 29880 8236 29886 8288
rect 30098 8236 30104 8288
rect 30156 8236 30162 8288
rect 30374 8236 30380 8288
rect 30432 8236 30438 8288
rect 30742 8236 30748 8288
rect 30800 8236 30806 8288
rect 31110 8236 31116 8288
rect 31168 8236 31174 8288
rect 32876 8285 32904 8384
rect 33042 8372 33048 8384
rect 33100 8372 33106 8424
rect 33244 8384 36124 8412
rect 32861 8279 32919 8285
rect 32861 8245 32873 8279
rect 32907 8245 32919 8279
rect 32861 8239 32919 8245
rect 33042 8236 33048 8288
rect 33100 8276 33106 8288
rect 33244 8276 33272 8384
rect 33410 8304 33416 8356
rect 33468 8304 33474 8356
rect 34882 8304 34888 8356
rect 34940 8304 34946 8356
rect 35158 8304 35164 8356
rect 35216 8304 35222 8356
rect 36096 8353 36124 8384
rect 36464 8353 36492 8520
rect 39850 8508 39856 8560
rect 39908 8548 39914 8560
rect 40604 8548 40632 8579
rect 40954 8576 40960 8628
rect 41012 8616 41018 8628
rect 41509 8619 41567 8625
rect 41509 8616 41521 8619
rect 41012 8588 41521 8616
rect 41012 8576 41018 8588
rect 41509 8585 41521 8588
rect 41555 8585 41567 8619
rect 41509 8579 41567 8585
rect 42613 8619 42671 8625
rect 42613 8585 42625 8619
rect 42659 8585 42671 8619
rect 42613 8579 42671 8585
rect 39908 8520 40632 8548
rect 39908 8508 39914 8520
rect 41322 8508 41328 8560
rect 41380 8548 41386 8560
rect 42628 8548 42656 8579
rect 42702 8576 42708 8628
rect 42760 8616 42766 8628
rect 44269 8619 44327 8625
rect 44269 8616 44281 8619
rect 42760 8588 44281 8616
rect 42760 8576 42766 8588
rect 44269 8585 44281 8588
rect 44315 8585 44327 8619
rect 44269 8579 44327 8585
rect 41380 8520 42656 8548
rect 41380 8508 41386 8520
rect 42886 8508 42892 8560
rect 42944 8548 42950 8560
rect 43073 8551 43131 8557
rect 43073 8548 43085 8551
rect 42944 8520 43085 8548
rect 42944 8508 42950 8520
rect 43073 8517 43085 8520
rect 43119 8517 43131 8551
rect 43073 8511 43131 8517
rect 43254 8508 43260 8560
rect 43312 8548 43318 8560
rect 44177 8551 44235 8557
rect 44177 8548 44189 8551
rect 43312 8520 44189 8548
rect 43312 8508 43318 8520
rect 44177 8517 44189 8520
rect 44223 8517 44235 8551
rect 44177 8511 44235 8517
rect 36630 8440 36636 8492
rect 36688 8440 36694 8492
rect 36814 8440 36820 8492
rect 36872 8440 36878 8492
rect 36906 8440 36912 8492
rect 36964 8480 36970 8492
rect 37277 8483 37335 8489
rect 37277 8480 37289 8483
rect 36964 8452 37289 8480
rect 36964 8440 36970 8452
rect 37277 8449 37289 8452
rect 37323 8449 37335 8483
rect 37277 8443 37335 8449
rect 37550 8440 37556 8492
rect 37608 8440 37614 8492
rect 37826 8440 37832 8492
rect 37884 8440 37890 8492
rect 38102 8440 38108 8492
rect 38160 8440 38166 8492
rect 38470 8440 38476 8492
rect 38528 8440 38534 8492
rect 38562 8440 38568 8492
rect 38620 8480 38626 8492
rect 38933 8483 38991 8489
rect 38933 8480 38945 8483
rect 38620 8452 38945 8480
rect 38620 8440 38626 8452
rect 38933 8449 38945 8452
rect 38979 8449 38991 8483
rect 38933 8443 38991 8449
rect 39393 8483 39451 8489
rect 39393 8449 39405 8483
rect 39439 8449 39451 8483
rect 39393 8443 39451 8449
rect 36832 8353 36860 8440
rect 36924 8384 38056 8412
rect 36081 8347 36139 8353
rect 36081 8313 36093 8347
rect 36127 8313 36139 8347
rect 36081 8307 36139 8313
rect 36449 8347 36507 8353
rect 36449 8313 36461 8347
rect 36495 8313 36507 8347
rect 36449 8307 36507 8313
rect 36817 8347 36875 8353
rect 36817 8313 36829 8347
rect 36863 8313 36875 8347
rect 36817 8307 36875 8313
rect 33100 8248 33272 8276
rect 33428 8276 33456 8304
rect 36924 8276 36952 8384
rect 37458 8304 37464 8356
rect 37516 8304 37522 8356
rect 37734 8304 37740 8356
rect 37792 8304 37798 8356
rect 38028 8353 38056 8384
rect 38013 8347 38071 8353
rect 38013 8313 38025 8347
rect 38059 8313 38071 8347
rect 39408 8344 39436 8443
rect 39942 8440 39948 8492
rect 40000 8440 40006 8492
rect 40218 8440 40224 8492
rect 40276 8440 40282 8492
rect 40494 8440 40500 8492
rect 40552 8440 40558 8492
rect 40678 8440 40684 8492
rect 40736 8480 40742 8492
rect 40957 8483 41015 8489
rect 40957 8480 40969 8483
rect 40736 8452 40969 8480
rect 40736 8440 40742 8452
rect 40957 8449 40969 8452
rect 41003 8449 41015 8483
rect 40957 8443 41015 8449
rect 41046 8440 41052 8492
rect 41104 8480 41110 8492
rect 41417 8483 41475 8489
rect 41417 8480 41429 8483
rect 41104 8452 41429 8480
rect 41104 8440 41110 8452
rect 41417 8449 41429 8452
rect 41463 8449 41475 8483
rect 41417 8443 41475 8449
rect 42518 8440 42524 8492
rect 42576 8440 42582 8492
rect 43622 8440 43628 8492
rect 43680 8440 43686 8492
rect 38013 8307 38071 8313
rect 38120 8316 39436 8344
rect 40236 8344 40264 8440
rect 42058 8372 42064 8424
rect 42116 8412 42122 8424
rect 42116 8384 43852 8412
rect 42116 8372 42122 8384
rect 41141 8347 41199 8353
rect 41141 8344 41153 8347
rect 40236 8316 41153 8344
rect 33428 8248 36952 8276
rect 33100 8236 33106 8248
rect 37182 8236 37188 8288
rect 37240 8276 37246 8288
rect 38120 8276 38148 8316
rect 41141 8313 41153 8316
rect 41187 8313 41199 8347
rect 41141 8307 41199 8313
rect 41690 8304 41696 8356
rect 41748 8344 41754 8356
rect 43824 8353 43852 8384
rect 43257 8347 43315 8353
rect 43257 8344 43269 8347
rect 41748 8316 43269 8344
rect 41748 8304 41754 8316
rect 43257 8313 43269 8316
rect 43303 8313 43315 8347
rect 43257 8307 43315 8313
rect 43809 8347 43867 8353
rect 43809 8313 43821 8347
rect 43855 8313 43867 8347
rect 43809 8307 43867 8313
rect 37240 8248 38148 8276
rect 37240 8236 37246 8248
rect 1104 8186 45540 8208
rect 1104 8134 6504 8186
rect 6556 8134 6568 8186
rect 6620 8134 6632 8186
rect 6684 8134 6696 8186
rect 6748 8134 6760 8186
rect 6812 8134 17612 8186
rect 17664 8134 17676 8186
rect 17728 8134 17740 8186
rect 17792 8134 17804 8186
rect 17856 8134 17868 8186
rect 17920 8134 28720 8186
rect 28772 8134 28784 8186
rect 28836 8134 28848 8186
rect 28900 8134 28912 8186
rect 28964 8134 28976 8186
rect 29028 8134 39828 8186
rect 39880 8134 39892 8186
rect 39944 8134 39956 8186
rect 40008 8134 40020 8186
rect 40072 8134 40084 8186
rect 40136 8134 45540 8186
rect 1104 8112 45540 8134
rect 2038 8032 2044 8084
rect 2096 8032 2102 8084
rect 2774 8032 2780 8084
rect 2832 8032 2838 8084
rect 3050 8032 3056 8084
rect 3108 8072 3114 8084
rect 3145 8075 3203 8081
rect 3145 8072 3157 8075
rect 3108 8044 3157 8072
rect 3108 8032 3114 8044
rect 3145 8041 3157 8044
rect 3191 8041 3203 8075
rect 3145 8035 3203 8041
rect 3418 8032 3424 8084
rect 3476 8072 3482 8084
rect 3513 8075 3571 8081
rect 3513 8072 3525 8075
rect 3476 8044 3525 8072
rect 3476 8032 3482 8044
rect 3513 8041 3525 8044
rect 3559 8041 3571 8075
rect 3513 8035 3571 8041
rect 4154 8032 4160 8084
rect 4212 8032 4218 8084
rect 4522 8032 4528 8084
rect 4580 8072 4586 8084
rect 4617 8075 4675 8081
rect 4617 8072 4629 8075
rect 4580 8044 4629 8072
rect 4580 8032 4586 8044
rect 4617 8041 4629 8044
rect 4663 8041 4675 8075
rect 4617 8035 4675 8041
rect 6362 8032 6368 8084
rect 6420 8072 6426 8084
rect 6457 8075 6515 8081
rect 6457 8072 6469 8075
rect 6420 8044 6469 8072
rect 6420 8032 6426 8044
rect 6457 8041 6469 8044
rect 6503 8041 6515 8075
rect 6457 8035 6515 8041
rect 7466 8032 7472 8084
rect 7524 8072 7530 8084
rect 7561 8075 7619 8081
rect 7561 8072 7573 8075
rect 7524 8044 7573 8072
rect 7524 8032 7530 8044
rect 7561 8041 7573 8044
rect 7607 8041 7619 8075
rect 7561 8035 7619 8041
rect 9122 8032 9128 8084
rect 9180 8032 9186 8084
rect 10042 8032 10048 8084
rect 10100 8072 10106 8084
rect 10137 8075 10195 8081
rect 10137 8072 10149 8075
rect 10100 8044 10149 8072
rect 10100 8032 10106 8044
rect 10137 8041 10149 8044
rect 10183 8041 10195 8075
rect 10137 8035 10195 8041
rect 11606 8032 11612 8084
rect 11664 8032 11670 8084
rect 11882 8032 11888 8084
rect 11940 8072 11946 8084
rect 12161 8075 12219 8081
rect 12161 8072 12173 8075
rect 11940 8044 12173 8072
rect 11940 8032 11946 8044
rect 12161 8041 12173 8044
rect 12207 8041 12219 8075
rect 12161 8035 12219 8041
rect 12986 8032 12992 8084
rect 13044 8072 13050 8084
rect 13081 8075 13139 8081
rect 13081 8072 13093 8075
rect 13044 8044 13093 8072
rect 13044 8032 13050 8044
rect 13081 8041 13093 8044
rect 13127 8041 13139 8075
rect 13081 8035 13139 8041
rect 14274 8032 14280 8084
rect 14332 8032 14338 8084
rect 17034 8032 17040 8084
rect 17092 8072 17098 8084
rect 17313 8075 17371 8081
rect 17313 8072 17325 8075
rect 17092 8044 17325 8072
rect 17092 8032 17098 8044
rect 17313 8041 17325 8044
rect 17359 8041 17371 8075
rect 17313 8035 17371 8041
rect 17494 8032 17500 8084
rect 17552 8072 17558 8084
rect 17773 8075 17831 8081
rect 17773 8072 17785 8075
rect 17552 8044 17785 8072
rect 17552 8032 17558 8044
rect 17773 8041 17785 8044
rect 17819 8041 17831 8075
rect 17773 8035 17831 8041
rect 18049 8075 18107 8081
rect 18049 8041 18061 8075
rect 18095 8072 18107 8075
rect 18230 8072 18236 8084
rect 18095 8044 18236 8072
rect 18095 8041 18107 8044
rect 18049 8035 18107 8041
rect 18230 8032 18236 8044
rect 18288 8032 18294 8084
rect 19242 8032 19248 8084
rect 19300 8072 19306 8084
rect 19521 8075 19579 8081
rect 19521 8072 19533 8075
rect 19300 8044 19533 8072
rect 19300 8032 19306 8044
rect 19521 8041 19533 8044
rect 19567 8041 19579 8075
rect 19521 8035 19579 8041
rect 20438 8032 20444 8084
rect 20496 8032 20502 8084
rect 20898 8032 20904 8084
rect 20956 8032 20962 8084
rect 21174 8032 21180 8084
rect 21232 8032 21238 8084
rect 21542 8032 21548 8084
rect 21600 8032 21606 8084
rect 21818 8032 21824 8084
rect 21876 8032 21882 8084
rect 22186 8032 22192 8084
rect 22244 8072 22250 8084
rect 22373 8075 22431 8081
rect 22373 8072 22385 8075
rect 22244 8044 22385 8072
rect 22244 8032 22250 8044
rect 22373 8041 22385 8044
rect 22419 8041 22431 8075
rect 22373 8035 22431 8041
rect 24302 8032 24308 8084
rect 24360 8072 24366 8084
rect 24360 8044 24440 8072
rect 24360 8032 24366 8044
rect 10410 7964 10416 8016
rect 10468 8004 10474 8016
rect 10468 7976 16712 8004
rect 10468 7964 10474 7976
rect 16684 7936 16712 7976
rect 17218 7964 17224 8016
rect 17276 8004 17282 8016
rect 19334 8004 19340 8016
rect 17276 7976 19340 8004
rect 17276 7964 17282 7976
rect 19334 7964 19340 7976
rect 19392 7964 19398 8016
rect 19426 7964 19432 8016
rect 19484 7964 19490 8016
rect 20346 8004 20352 8016
rect 19628 7976 20352 8004
rect 18046 7936 18052 7948
rect 11624 7908 15240 7936
rect 16684 7908 18052 7936
rect 2958 7828 2964 7880
rect 3016 7828 3022 7880
rect 3326 7828 3332 7880
rect 3384 7828 3390 7880
rect 4430 7828 4436 7880
rect 4488 7828 4494 7880
rect 7377 7871 7435 7877
rect 7377 7837 7389 7871
rect 7423 7868 7435 7871
rect 7423 7840 9674 7868
rect 7423 7837 7435 7840
rect 7377 7831 7435 7837
rect 1949 7803 2007 7809
rect 1949 7769 1961 7803
rect 1995 7769 2007 7803
rect 1949 7763 2007 7769
rect 1964 7732 1992 7763
rect 2498 7760 2504 7812
rect 2556 7760 2562 7812
rect 3878 7760 3884 7812
rect 3936 7760 3942 7812
rect 6362 7760 6368 7812
rect 6420 7760 6426 7812
rect 9033 7803 9091 7809
rect 9033 7769 9045 7803
rect 9079 7769 9091 7803
rect 9646 7800 9674 7840
rect 9950 7828 9956 7880
rect 10008 7828 10014 7880
rect 11514 7828 11520 7880
rect 11572 7828 11578 7880
rect 11624 7800 11652 7908
rect 11977 7871 12035 7877
rect 11977 7837 11989 7871
rect 12023 7837 12035 7871
rect 11977 7831 12035 7837
rect 9646 7772 11652 7800
rect 11992 7800 12020 7831
rect 12894 7828 12900 7880
rect 12952 7828 12958 7880
rect 14108 7840 15148 7868
rect 14108 7800 14136 7840
rect 15120 7812 15148 7840
rect 11992 7772 14136 7800
rect 9033 7763 9091 7769
rect 5442 7732 5448 7744
rect 1964 7704 5448 7732
rect 5442 7692 5448 7704
rect 5500 7692 5506 7744
rect 9048 7732 9076 7763
rect 14182 7760 14188 7812
rect 14240 7760 14246 7812
rect 15102 7760 15108 7812
rect 15160 7760 15166 7812
rect 15212 7800 15240 7908
rect 18046 7896 18052 7908
rect 18104 7896 18110 7948
rect 19444 7936 19472 7964
rect 18340 7908 19472 7936
rect 17126 7828 17132 7880
rect 17184 7828 17190 7880
rect 17218 7828 17224 7880
rect 17276 7828 17282 7880
rect 17310 7828 17316 7880
rect 17368 7828 17374 7880
rect 17681 7871 17739 7877
rect 17681 7837 17693 7871
rect 17727 7868 17739 7871
rect 17862 7868 17868 7880
rect 17727 7840 17868 7868
rect 17727 7837 17739 7840
rect 17681 7831 17739 7837
rect 17862 7828 17868 7840
rect 17920 7828 17926 7880
rect 17957 7871 18015 7877
rect 17957 7837 17969 7871
rect 18003 7837 18015 7871
rect 17957 7831 18015 7837
rect 17236 7800 17264 7828
rect 15212 7772 17264 7800
rect 17328 7800 17356 7828
rect 17972 7800 18000 7831
rect 18230 7828 18236 7880
rect 18288 7828 18294 7880
rect 18340 7877 18368 7908
rect 18325 7871 18383 7877
rect 18325 7837 18337 7871
rect 18371 7837 18383 7871
rect 18325 7831 18383 7837
rect 18782 7828 18788 7880
rect 18840 7828 18846 7880
rect 18877 7871 18935 7877
rect 18877 7837 18889 7871
rect 18923 7868 18935 7871
rect 19628 7868 19656 7976
rect 20346 7964 20352 7976
rect 20404 7964 20410 8016
rect 20254 7936 20260 7948
rect 19904 7908 20260 7936
rect 19904 7877 19932 7908
rect 20254 7896 20260 7908
rect 20312 7896 20318 7948
rect 21192 7936 21220 8032
rect 21836 7936 21864 8032
rect 22094 7964 22100 8016
rect 22152 8004 22158 8016
rect 23937 8007 23995 8013
rect 23937 8004 23949 8007
rect 22152 7976 23949 8004
rect 22152 7964 22158 7976
rect 23937 7973 23949 7976
rect 23983 7973 23995 8007
rect 24412 8004 24440 8044
rect 24578 8032 24584 8084
rect 24636 8032 24642 8084
rect 25038 8032 25044 8084
rect 25096 8032 25102 8084
rect 25222 8032 25228 8084
rect 25280 8072 25286 8084
rect 27249 8075 27307 8081
rect 27249 8072 27261 8075
rect 25280 8044 27261 8072
rect 25280 8032 25286 8044
rect 27249 8041 27261 8044
rect 27295 8041 27307 8075
rect 27249 8035 27307 8041
rect 27522 8032 27528 8084
rect 27580 8032 27586 8084
rect 27617 8075 27675 8081
rect 27617 8041 27629 8075
rect 27663 8072 27675 8075
rect 27706 8072 27712 8084
rect 27663 8044 27712 8072
rect 27663 8041 27675 8044
rect 27617 8035 27675 8041
rect 27706 8032 27712 8044
rect 27764 8032 27770 8084
rect 27798 8032 27804 8084
rect 27856 8032 27862 8084
rect 27890 8032 27896 8084
rect 27948 8032 27954 8084
rect 28534 8032 28540 8084
rect 28592 8032 28598 8084
rect 28626 8032 28632 8084
rect 28684 8032 28690 8084
rect 40586 8032 40592 8084
rect 40644 8072 40650 8084
rect 41141 8075 41199 8081
rect 41141 8072 41153 8075
rect 40644 8044 41153 8072
rect 40644 8032 40650 8044
rect 41141 8041 41153 8044
rect 41187 8041 41199 8075
rect 41141 8035 41199 8041
rect 42794 8032 42800 8084
rect 42852 8072 42858 8084
rect 43257 8075 43315 8081
rect 43257 8072 43269 8075
rect 42852 8044 43269 8072
rect 42852 8032 42858 8044
rect 43257 8041 43269 8044
rect 43303 8041 43315 8075
rect 43257 8035 43315 8041
rect 43530 8032 43536 8084
rect 43588 8072 43594 8084
rect 43809 8075 43867 8081
rect 43809 8072 43821 8075
rect 43588 8044 43821 8072
rect 43588 8032 43594 8044
rect 43809 8041 43821 8044
rect 43855 8041 43867 8075
rect 43809 8035 43867 8041
rect 43898 8032 43904 8084
rect 43956 8072 43962 8084
rect 44361 8075 44419 8081
rect 44361 8072 44373 8075
rect 43956 8044 44373 8072
rect 43956 8032 43962 8044
rect 44361 8041 44373 8044
rect 44407 8041 44419 8075
rect 44361 8035 44419 8041
rect 24857 8007 24915 8013
rect 24857 8004 24869 8007
rect 24412 7976 24869 8004
rect 23937 7967 23995 7973
rect 24857 7973 24869 7976
rect 24903 7973 24915 8007
rect 24857 7967 24915 7973
rect 20732 7908 21220 7936
rect 21284 7908 21864 7936
rect 22204 7908 22416 7936
rect 18923 7840 19656 7868
rect 19889 7871 19947 7877
rect 18923 7837 18935 7840
rect 18877 7831 18935 7837
rect 19889 7837 19901 7871
rect 19935 7837 19947 7871
rect 19889 7831 19947 7837
rect 20165 7871 20223 7877
rect 20165 7837 20177 7871
rect 20211 7868 20223 7871
rect 20530 7868 20536 7880
rect 20211 7840 20536 7868
rect 20211 7837 20223 7840
rect 20165 7831 20223 7837
rect 20530 7828 20536 7840
rect 20588 7828 20594 7880
rect 20622 7828 20628 7880
rect 20680 7828 20686 7880
rect 20732 7877 20760 7908
rect 21284 7877 21312 7908
rect 20717 7871 20775 7877
rect 20717 7837 20729 7871
rect 20763 7837 20775 7871
rect 20717 7831 20775 7837
rect 20993 7871 21051 7877
rect 20993 7837 21005 7871
rect 21039 7837 21051 7871
rect 20993 7831 21051 7837
rect 21269 7871 21327 7877
rect 21269 7837 21281 7871
rect 21315 7837 21327 7871
rect 21269 7831 21327 7837
rect 18414 7800 18420 7812
rect 17328 7772 17540 7800
rect 17972 7772 18420 7800
rect 17218 7732 17224 7744
rect 9048 7704 17224 7732
rect 17218 7692 17224 7704
rect 17276 7692 17282 7744
rect 17512 7741 17540 7772
rect 18414 7760 18420 7772
rect 18472 7760 18478 7812
rect 19429 7803 19487 7809
rect 19429 7800 19441 7803
rect 18616 7772 19441 7800
rect 17497 7735 17555 7741
rect 17497 7701 17509 7735
rect 17543 7701 17555 7735
rect 17497 7695 17555 7701
rect 18506 7692 18512 7744
rect 18564 7692 18570 7744
rect 18616 7741 18644 7772
rect 19429 7769 19441 7772
rect 19475 7769 19487 7803
rect 21008 7800 21036 7831
rect 21450 7828 21456 7880
rect 21508 7828 21514 7880
rect 21726 7828 21732 7880
rect 21784 7828 21790 7880
rect 22002 7828 22008 7880
rect 22060 7828 22066 7880
rect 21468 7800 21496 7828
rect 19429 7763 19487 7769
rect 19536 7772 20392 7800
rect 21008 7772 21496 7800
rect 18601 7735 18659 7741
rect 18601 7701 18613 7735
rect 18647 7701 18659 7735
rect 18601 7695 18659 7701
rect 18690 7692 18696 7744
rect 18748 7732 18754 7744
rect 19061 7735 19119 7741
rect 19061 7732 19073 7735
rect 18748 7704 19073 7732
rect 18748 7692 18754 7704
rect 19061 7701 19073 7704
rect 19107 7701 19119 7735
rect 19061 7695 19119 7701
rect 19334 7692 19340 7744
rect 19392 7732 19398 7744
rect 19536 7732 19564 7772
rect 19392 7704 19564 7732
rect 19392 7692 19398 7704
rect 20070 7692 20076 7744
rect 20128 7692 20134 7744
rect 20364 7741 20392 7772
rect 21634 7760 21640 7812
rect 21692 7800 21698 7812
rect 22204 7800 22232 7908
rect 22281 7871 22339 7877
rect 22281 7837 22293 7871
rect 22327 7837 22339 7871
rect 22281 7831 22339 7837
rect 21692 7772 22232 7800
rect 21692 7760 21698 7772
rect 20349 7735 20407 7741
rect 20349 7701 20361 7735
rect 20395 7701 20407 7735
rect 20349 7695 20407 7701
rect 21177 7735 21235 7741
rect 21177 7701 21189 7735
rect 21223 7732 21235 7735
rect 21358 7732 21364 7744
rect 21223 7704 21364 7732
rect 21223 7701 21235 7704
rect 21177 7695 21235 7701
rect 21358 7692 21364 7704
rect 21416 7692 21422 7744
rect 21450 7692 21456 7744
rect 21508 7692 21514 7744
rect 21818 7692 21824 7744
rect 21876 7692 21882 7744
rect 22002 7692 22008 7744
rect 22060 7732 22066 7744
rect 22097 7735 22155 7741
rect 22097 7732 22109 7735
rect 22060 7704 22109 7732
rect 22060 7692 22066 7704
rect 22097 7701 22109 7704
rect 22143 7701 22155 7735
rect 22296 7732 22324 7831
rect 22388 7800 22416 7908
rect 22462 7896 22468 7948
rect 22520 7936 22526 7948
rect 25056 7936 25084 8032
rect 26234 7964 26240 8016
rect 26292 8004 26298 8016
rect 26513 8007 26571 8013
rect 26513 8004 26525 8007
rect 26292 7976 26525 8004
rect 26292 7964 26298 7976
rect 26513 7973 26525 7976
rect 26559 7973 26571 8007
rect 27540 8004 27568 8032
rect 26513 7967 26571 7973
rect 26712 7976 27568 8004
rect 22520 7908 22876 7936
rect 22520 7896 22526 7908
rect 22557 7871 22615 7877
rect 22557 7837 22569 7871
rect 22603 7868 22615 7871
rect 22738 7868 22744 7880
rect 22603 7840 22744 7868
rect 22603 7837 22615 7840
rect 22557 7831 22615 7837
rect 22738 7828 22744 7840
rect 22796 7828 22802 7880
rect 22848 7877 22876 7908
rect 22940 7908 23980 7936
rect 22940 7877 22968 7908
rect 23952 7880 23980 7908
rect 24320 7908 25084 7936
rect 22833 7871 22891 7877
rect 22833 7837 22845 7871
rect 22879 7837 22891 7871
rect 22833 7831 22891 7837
rect 22925 7871 22983 7877
rect 22925 7837 22937 7871
rect 22971 7837 22983 7871
rect 22925 7831 22983 7837
rect 23198 7828 23204 7880
rect 23256 7828 23262 7880
rect 23477 7871 23535 7877
rect 23477 7837 23489 7871
rect 23523 7868 23535 7871
rect 23658 7868 23664 7880
rect 23523 7840 23664 7868
rect 23523 7837 23535 7840
rect 23477 7831 23535 7837
rect 23658 7828 23664 7840
rect 23716 7828 23722 7880
rect 23753 7871 23811 7877
rect 23753 7837 23765 7871
rect 23799 7837 23811 7871
rect 23753 7831 23811 7837
rect 23768 7800 23796 7831
rect 23934 7828 23940 7880
rect 23992 7828 23998 7880
rect 24029 7871 24087 7877
rect 24029 7837 24041 7871
rect 24075 7868 24087 7871
rect 24320 7868 24348 7908
rect 24075 7840 24348 7868
rect 24397 7871 24455 7877
rect 24075 7837 24087 7840
rect 24029 7831 24087 7837
rect 24397 7837 24409 7871
rect 24443 7837 24455 7871
rect 24397 7831 24455 7837
rect 24673 7871 24731 7877
rect 24673 7837 24685 7871
rect 24719 7837 24731 7871
rect 24673 7831 24731 7837
rect 24949 7871 25007 7877
rect 24949 7837 24961 7871
rect 24995 7868 25007 7871
rect 25130 7868 25136 7880
rect 24995 7840 25136 7868
rect 24995 7837 25007 7840
rect 24949 7831 25007 7837
rect 22388 7772 23704 7800
rect 23768 7772 24348 7800
rect 22554 7732 22560 7744
rect 22296 7704 22560 7732
rect 22097 7695 22155 7701
rect 22554 7692 22560 7704
rect 22612 7692 22618 7744
rect 22646 7692 22652 7744
rect 22704 7692 22710 7744
rect 22830 7692 22836 7744
rect 22888 7732 22894 7744
rect 23109 7735 23167 7741
rect 23109 7732 23121 7735
rect 22888 7704 23121 7732
rect 22888 7692 22894 7704
rect 23109 7701 23121 7704
rect 23155 7701 23167 7735
rect 23109 7695 23167 7701
rect 23382 7692 23388 7744
rect 23440 7692 23446 7744
rect 23676 7741 23704 7772
rect 24320 7744 24348 7772
rect 23661 7735 23719 7741
rect 23661 7701 23673 7735
rect 23707 7701 23719 7735
rect 23661 7695 23719 7701
rect 24210 7692 24216 7744
rect 24268 7692 24274 7744
rect 24302 7692 24308 7744
rect 24360 7692 24366 7744
rect 24412 7732 24440 7831
rect 24688 7800 24716 7831
rect 25130 7828 25136 7840
rect 25188 7828 25194 7880
rect 25225 7871 25283 7877
rect 25225 7837 25237 7871
rect 25271 7868 25283 7871
rect 25406 7868 25412 7880
rect 25271 7840 25412 7868
rect 25271 7837 25283 7840
rect 25225 7831 25283 7837
rect 25406 7828 25412 7840
rect 25464 7828 25470 7880
rect 25501 7871 25559 7877
rect 25501 7837 25513 7871
rect 25547 7868 25559 7871
rect 25682 7868 25688 7880
rect 25547 7840 25688 7868
rect 25547 7837 25559 7840
rect 25501 7831 25559 7837
rect 25682 7828 25688 7840
rect 25740 7828 25746 7880
rect 25777 7871 25835 7877
rect 25777 7837 25789 7871
rect 25823 7868 25835 7871
rect 25866 7868 25872 7880
rect 25823 7840 25872 7868
rect 25823 7837 25835 7840
rect 25777 7831 25835 7837
rect 25866 7828 25872 7840
rect 25924 7828 25930 7880
rect 26053 7871 26111 7877
rect 26053 7837 26065 7871
rect 26099 7868 26111 7871
rect 26142 7868 26148 7880
rect 26099 7840 26148 7868
rect 26099 7837 26111 7840
rect 26053 7831 26111 7837
rect 26142 7828 26148 7840
rect 26200 7828 26206 7880
rect 26329 7871 26387 7877
rect 26329 7837 26341 7871
rect 26375 7868 26387 7871
rect 26602 7868 26608 7880
rect 26375 7840 26608 7868
rect 26375 7837 26387 7840
rect 26329 7831 26387 7837
rect 26602 7828 26608 7840
rect 26660 7828 26666 7880
rect 26712 7877 26740 7976
rect 27816 7936 27844 8032
rect 28552 8004 28580 8032
rect 27080 7908 27844 7936
rect 28000 7976 28580 8004
rect 27080 7877 27108 7908
rect 26697 7871 26755 7877
rect 26697 7837 26709 7871
rect 26743 7837 26755 7871
rect 26697 7831 26755 7837
rect 27065 7871 27123 7877
rect 27065 7837 27077 7871
rect 27111 7837 27123 7871
rect 27065 7831 27123 7837
rect 27433 7871 27491 7877
rect 27433 7837 27445 7871
rect 27479 7868 27491 7871
rect 27614 7868 27620 7880
rect 27479 7840 27620 7868
rect 27479 7837 27491 7840
rect 27433 7831 27491 7837
rect 27614 7828 27620 7840
rect 27672 7828 27678 7880
rect 28000 7877 28028 7976
rect 28644 7936 28672 8032
rect 42889 8007 42947 8013
rect 42889 7973 42901 8007
rect 42935 8004 42947 8007
rect 44266 8004 44272 8016
rect 42935 7976 44272 8004
rect 42935 7973 42947 7976
rect 42889 7967 42947 7973
rect 44266 7964 44272 7976
rect 44324 7964 44330 8016
rect 28276 7908 28672 7936
rect 28276 7877 28304 7908
rect 27709 7871 27767 7877
rect 27709 7837 27721 7871
rect 27755 7837 27767 7871
rect 27709 7831 27767 7837
rect 27985 7871 28043 7877
rect 27985 7837 27997 7871
rect 28031 7837 28043 7871
rect 27985 7831 28043 7837
rect 28261 7871 28319 7877
rect 28261 7837 28273 7871
rect 28307 7837 28319 7871
rect 28261 7831 28319 7837
rect 28537 7871 28595 7877
rect 28537 7837 28549 7871
rect 28583 7868 28595 7871
rect 29546 7868 29552 7880
rect 28583 7840 29552 7868
rect 28583 7837 28595 7840
rect 28537 7831 28595 7837
rect 27724 7800 27752 7831
rect 29546 7828 29552 7840
rect 29604 7828 29610 7880
rect 29822 7828 29828 7880
rect 29880 7828 29886 7880
rect 33042 7828 33048 7880
rect 33100 7868 33106 7880
rect 40957 7871 41015 7877
rect 40957 7868 40969 7871
rect 33100 7840 40969 7868
rect 33100 7828 33106 7840
rect 40957 7837 40969 7840
rect 41003 7837 41015 7871
rect 40957 7831 41015 7837
rect 29840 7800 29868 7828
rect 24688 7772 27016 7800
rect 27724 7772 29868 7800
rect 25038 7732 25044 7744
rect 24412 7704 25044 7732
rect 25038 7692 25044 7704
rect 25096 7692 25102 7744
rect 25130 7692 25136 7744
rect 25188 7692 25194 7744
rect 25406 7692 25412 7744
rect 25464 7692 25470 7744
rect 25682 7692 25688 7744
rect 25740 7692 25746 7744
rect 25958 7692 25964 7744
rect 26016 7692 26022 7744
rect 26234 7692 26240 7744
rect 26292 7692 26298 7744
rect 26878 7692 26884 7744
rect 26936 7692 26942 7744
rect 26988 7732 27016 7772
rect 39666 7760 39672 7812
rect 39724 7800 39730 7812
rect 42613 7803 42671 7809
rect 42613 7800 42625 7803
rect 39724 7772 42625 7800
rect 39724 7760 39730 7772
rect 42613 7769 42625 7772
rect 42659 7769 42671 7803
rect 42613 7763 42671 7769
rect 42794 7760 42800 7812
rect 42852 7800 42858 7812
rect 43165 7803 43223 7809
rect 43165 7800 43177 7803
rect 42852 7772 43177 7800
rect 42852 7760 42858 7772
rect 43165 7769 43177 7772
rect 43211 7769 43223 7803
rect 43165 7763 43223 7769
rect 43438 7760 43444 7812
rect 43496 7800 43502 7812
rect 43717 7803 43775 7809
rect 43717 7800 43729 7803
rect 43496 7772 43729 7800
rect 43496 7760 43502 7772
rect 43717 7769 43729 7772
rect 43763 7769 43775 7803
rect 43717 7763 43775 7769
rect 44266 7760 44272 7812
rect 44324 7760 44330 7812
rect 27338 7732 27344 7744
rect 26988 7704 27344 7732
rect 27338 7692 27344 7704
rect 27396 7692 27402 7744
rect 28166 7692 28172 7744
rect 28224 7692 28230 7744
rect 28442 7692 28448 7744
rect 28500 7692 28506 7744
rect 28534 7692 28540 7744
rect 28592 7732 28598 7744
rect 28721 7735 28779 7741
rect 28721 7732 28733 7735
rect 28592 7704 28733 7732
rect 28592 7692 28598 7704
rect 28721 7701 28733 7704
rect 28767 7701 28779 7735
rect 28721 7695 28779 7701
rect 1104 7642 45696 7664
rect 1104 7590 12058 7642
rect 12110 7590 12122 7642
rect 12174 7590 12186 7642
rect 12238 7590 12250 7642
rect 12302 7590 12314 7642
rect 12366 7590 23166 7642
rect 23218 7590 23230 7642
rect 23282 7590 23294 7642
rect 23346 7590 23358 7642
rect 23410 7590 23422 7642
rect 23474 7590 34274 7642
rect 34326 7590 34338 7642
rect 34390 7590 34402 7642
rect 34454 7590 34466 7642
rect 34518 7590 34530 7642
rect 34582 7590 45382 7642
rect 45434 7590 45446 7642
rect 45498 7590 45510 7642
rect 45562 7590 45574 7642
rect 45626 7590 45638 7642
rect 45690 7590 45696 7642
rect 1104 7568 45696 7590
rect 842 7488 848 7540
rect 900 7528 906 7540
rect 1765 7531 1823 7537
rect 1765 7528 1777 7531
rect 900 7500 1777 7528
rect 900 7488 906 7500
rect 1765 7497 1777 7500
rect 1811 7497 1823 7531
rect 2317 7531 2375 7537
rect 2317 7528 2329 7531
rect 1765 7491 1823 7497
rect 1872 7500 2329 7528
rect 1578 7420 1584 7472
rect 1636 7460 1642 7472
rect 1872 7460 1900 7500
rect 2317 7497 2329 7500
rect 2363 7497 2375 7531
rect 2317 7491 2375 7497
rect 3878 7488 3884 7540
rect 3936 7528 3942 7540
rect 11054 7528 11060 7540
rect 3936 7500 11060 7528
rect 3936 7488 3942 7500
rect 11054 7488 11060 7500
rect 11112 7488 11118 7540
rect 15102 7528 15108 7540
rect 11624 7500 15108 7528
rect 1636 7432 1900 7460
rect 2225 7463 2283 7469
rect 1636 7420 1642 7432
rect 2225 7429 2237 7463
rect 2271 7460 2283 7463
rect 11624 7460 11652 7500
rect 15102 7488 15108 7500
rect 15160 7488 15166 7540
rect 17126 7488 17132 7540
rect 17184 7528 17190 7540
rect 17497 7531 17555 7537
rect 17497 7528 17509 7531
rect 17184 7500 17509 7528
rect 17184 7488 17190 7500
rect 17497 7497 17509 7500
rect 17543 7497 17555 7531
rect 18690 7528 18696 7540
rect 17497 7491 17555 7497
rect 17604 7500 18696 7528
rect 17604 7460 17632 7500
rect 18690 7488 18696 7500
rect 18748 7488 18754 7540
rect 18782 7488 18788 7540
rect 18840 7488 18846 7540
rect 18874 7488 18880 7540
rect 18932 7488 18938 7540
rect 19150 7488 19156 7540
rect 19208 7528 19214 7540
rect 19245 7531 19303 7537
rect 19245 7528 19257 7531
rect 19208 7500 19257 7528
rect 19208 7488 19214 7500
rect 19245 7497 19257 7500
rect 19291 7497 19303 7531
rect 19245 7491 19303 7497
rect 19705 7531 19763 7537
rect 19705 7497 19717 7531
rect 19751 7497 19763 7531
rect 19705 7491 19763 7497
rect 19720 7460 19748 7491
rect 19886 7488 19892 7540
rect 19944 7528 19950 7540
rect 21818 7528 21824 7540
rect 19944 7500 21824 7528
rect 19944 7488 19950 7500
rect 21818 7488 21824 7500
rect 21876 7488 21882 7540
rect 22097 7531 22155 7537
rect 22097 7497 22109 7531
rect 22143 7528 22155 7531
rect 22186 7528 22192 7540
rect 22143 7500 22192 7528
rect 22143 7497 22155 7500
rect 22097 7491 22155 7497
rect 22186 7488 22192 7500
rect 22244 7488 22250 7540
rect 22465 7531 22523 7537
rect 22465 7528 22477 7531
rect 22296 7500 22477 7528
rect 2271 7432 11652 7460
rect 11716 7432 17632 7460
rect 18616 7432 19748 7460
rect 2271 7429 2283 7432
rect 2225 7423 2283 7429
rect 1673 7395 1731 7401
rect 1673 7361 1685 7395
rect 1719 7392 1731 7395
rect 11716 7392 11744 7432
rect 1719 7364 11744 7392
rect 1719 7361 1731 7364
rect 1673 7355 1731 7361
rect 12894 7352 12900 7404
rect 12952 7352 12958 7404
rect 17681 7395 17739 7401
rect 17681 7361 17693 7395
rect 17727 7392 17739 7395
rect 18138 7392 18144 7404
rect 17727 7364 18144 7392
rect 17727 7361 17739 7364
rect 17681 7355 17739 7361
rect 18138 7352 18144 7364
rect 18196 7352 18202 7404
rect 18616 7401 18644 7432
rect 20806 7420 20812 7472
rect 20864 7460 20870 7472
rect 22296 7460 22324 7500
rect 22465 7497 22477 7500
rect 22511 7497 22523 7531
rect 22646 7528 22652 7540
rect 22465 7491 22523 7497
rect 22572 7500 22652 7528
rect 20864 7432 22324 7460
rect 20864 7420 20870 7432
rect 22370 7420 22376 7472
rect 22428 7420 22434 7472
rect 18601 7395 18659 7401
rect 18601 7361 18613 7395
rect 18647 7361 18659 7395
rect 18601 7355 18659 7361
rect 19058 7352 19064 7404
rect 19116 7352 19122 7404
rect 19426 7352 19432 7404
rect 19484 7352 19490 7404
rect 19610 7352 19616 7404
rect 19668 7392 19674 7404
rect 19889 7395 19947 7401
rect 19889 7392 19901 7395
rect 19668 7364 19901 7392
rect 19668 7352 19674 7364
rect 19889 7361 19901 7364
rect 19935 7361 19947 7395
rect 19889 7355 19947 7361
rect 21082 7352 21088 7404
rect 21140 7392 21146 7404
rect 21818 7392 21824 7404
rect 21140 7364 21824 7392
rect 21140 7352 21146 7364
rect 21818 7352 21824 7364
rect 21876 7352 21882 7404
rect 21910 7352 21916 7404
rect 21968 7352 21974 7404
rect 22189 7395 22247 7401
rect 22189 7361 22201 7395
rect 22235 7392 22247 7395
rect 22388 7392 22416 7420
rect 22235 7364 22416 7392
rect 22235 7361 22247 7364
rect 22189 7355 22247 7361
rect 4430 7284 4436 7336
rect 4488 7284 4494 7336
rect 6362 7284 6368 7336
rect 6420 7284 6426 7336
rect 11054 7284 11060 7336
rect 11112 7324 11118 7336
rect 12342 7324 12348 7336
rect 11112 7296 12348 7324
rect 11112 7284 11118 7296
rect 12342 7284 12348 7296
rect 12400 7284 12406 7336
rect 12912 7324 12940 7352
rect 12912 7296 21588 7324
rect 4448 7188 4476 7284
rect 6380 7256 6408 7284
rect 21450 7256 21456 7268
rect 6380 7228 21456 7256
rect 21450 7216 21456 7228
rect 21508 7216 21514 7268
rect 21560 7256 21588 7296
rect 21634 7284 21640 7336
rect 21692 7324 21698 7336
rect 22572 7324 22600 7500
rect 22646 7488 22652 7500
rect 22704 7488 22710 7540
rect 22922 7488 22928 7540
rect 22980 7488 22986 7540
rect 23106 7488 23112 7540
rect 23164 7528 23170 7540
rect 24210 7528 24216 7540
rect 23164 7500 24216 7528
rect 23164 7488 23170 7500
rect 24210 7488 24216 7500
rect 24268 7488 24274 7540
rect 24486 7488 24492 7540
rect 24544 7488 24550 7540
rect 27338 7488 27344 7540
rect 27396 7528 27402 7540
rect 30098 7528 30104 7540
rect 27396 7500 30104 7528
rect 27396 7488 27402 7500
rect 30098 7488 30104 7500
rect 30156 7488 30162 7540
rect 30374 7488 30380 7540
rect 30432 7488 30438 7540
rect 30742 7488 30748 7540
rect 30800 7488 30806 7540
rect 43162 7488 43168 7540
rect 43220 7528 43226 7540
rect 43441 7531 43499 7537
rect 43441 7528 43453 7531
rect 43220 7500 43453 7528
rect 43220 7488 43226 7500
rect 43441 7497 43453 7500
rect 43487 7497 43499 7531
rect 43441 7491 43499 7497
rect 44729 7531 44787 7537
rect 44729 7497 44741 7531
rect 44775 7528 44787 7531
rect 45002 7528 45008 7540
rect 44775 7500 45008 7528
rect 44775 7497 44787 7500
rect 44729 7491 44787 7497
rect 45002 7488 45008 7500
rect 45060 7488 45066 7540
rect 45738 7488 45744 7540
rect 45796 7488 45802 7540
rect 22940 7460 22968 7488
rect 24504 7460 24532 7488
rect 22664 7432 22968 7460
rect 23768 7432 24532 7460
rect 22664 7401 22692 7432
rect 22649 7395 22707 7401
rect 22649 7361 22661 7395
rect 22695 7361 22707 7395
rect 22649 7355 22707 7361
rect 22738 7352 22744 7404
rect 22796 7352 22802 7404
rect 22922 7352 22928 7404
rect 22980 7352 22986 7404
rect 23014 7352 23020 7404
rect 23072 7352 23078 7404
rect 23382 7352 23388 7404
rect 23440 7352 23446 7404
rect 23768 7401 23796 7432
rect 25038 7420 25044 7472
rect 25096 7460 25102 7472
rect 30392 7460 30420 7488
rect 25096 7432 30420 7460
rect 25096 7420 25102 7432
rect 23753 7395 23811 7401
rect 23753 7361 23765 7395
rect 23799 7361 23811 7395
rect 23753 7355 23811 7361
rect 24029 7395 24087 7401
rect 24029 7361 24041 7395
rect 24075 7392 24087 7395
rect 30760 7392 30788 7488
rect 44269 7463 44327 7469
rect 44269 7429 44281 7463
rect 44315 7460 44327 7463
rect 45756 7460 45784 7488
rect 44315 7432 45784 7460
rect 44315 7429 44327 7432
rect 44269 7423 44327 7429
rect 24075 7364 30788 7392
rect 31036 7364 31754 7392
rect 24075 7361 24087 7364
rect 24029 7355 24087 7361
rect 21692 7296 22600 7324
rect 22756 7324 22784 7352
rect 31036 7324 31064 7364
rect 22756 7296 31064 7324
rect 21692 7284 21698 7296
rect 31110 7284 31116 7336
rect 31168 7284 31174 7336
rect 26878 7256 26884 7268
rect 21560 7228 26884 7256
rect 26878 7216 26884 7228
rect 26936 7216 26942 7268
rect 14550 7188 14556 7200
rect 4448 7160 14556 7188
rect 14550 7148 14556 7160
rect 14608 7148 14614 7200
rect 15470 7148 15476 7200
rect 15528 7188 15534 7200
rect 21910 7188 21916 7200
rect 15528 7160 21916 7188
rect 15528 7148 15534 7160
rect 21910 7148 21916 7160
rect 21968 7148 21974 7200
rect 22002 7148 22008 7200
rect 22060 7188 22066 7200
rect 22373 7191 22431 7197
rect 22373 7188 22385 7191
rect 22060 7160 22385 7188
rect 22060 7148 22066 7160
rect 22373 7157 22385 7160
rect 22419 7157 22431 7191
rect 22373 7151 22431 7157
rect 22738 7148 22744 7200
rect 22796 7148 22802 7200
rect 23198 7148 23204 7200
rect 23256 7148 23262 7200
rect 23569 7191 23627 7197
rect 23569 7157 23581 7191
rect 23615 7188 23627 7191
rect 23842 7188 23848 7200
rect 23615 7160 23848 7188
rect 23615 7157 23627 7160
rect 23569 7151 23627 7157
rect 23842 7148 23848 7160
rect 23900 7148 23906 7200
rect 23937 7191 23995 7197
rect 23937 7157 23949 7191
rect 23983 7188 23995 7191
rect 24118 7188 24124 7200
rect 23983 7160 24124 7188
rect 23983 7157 23995 7160
rect 23937 7151 23995 7157
rect 24118 7148 24124 7160
rect 24176 7148 24182 7200
rect 24210 7148 24216 7200
rect 24268 7148 24274 7200
rect 24302 7148 24308 7200
rect 24360 7188 24366 7200
rect 31128 7188 31156 7284
rect 24360 7160 31156 7188
rect 31726 7188 31754 7364
rect 43346 7352 43352 7404
rect 43404 7352 43410 7404
rect 43901 7395 43959 7401
rect 43901 7361 43913 7395
rect 43947 7361 43959 7395
rect 43901 7355 43959 7361
rect 43916 7324 43944 7355
rect 44174 7352 44180 7404
rect 44232 7392 44238 7404
rect 44453 7395 44511 7401
rect 44453 7392 44465 7395
rect 44232 7364 44465 7392
rect 44232 7352 44238 7364
rect 44453 7361 44465 7364
rect 44499 7361 44511 7395
rect 44453 7355 44511 7361
rect 45002 7324 45008 7336
rect 43916 7296 45008 7324
rect 45002 7284 45008 7296
rect 45060 7284 45066 7336
rect 37734 7188 37740 7200
rect 31726 7160 37740 7188
rect 24360 7148 24366 7160
rect 37734 7148 37740 7160
rect 37792 7148 37798 7200
rect 1104 7098 45540 7120
rect 1104 7046 6504 7098
rect 6556 7046 6568 7098
rect 6620 7046 6632 7098
rect 6684 7046 6696 7098
rect 6748 7046 6760 7098
rect 6812 7046 17612 7098
rect 17664 7046 17676 7098
rect 17728 7046 17740 7098
rect 17792 7046 17804 7098
rect 17856 7046 17868 7098
rect 17920 7046 28720 7098
rect 28772 7046 28784 7098
rect 28836 7046 28848 7098
rect 28900 7046 28912 7098
rect 28964 7046 28976 7098
rect 29028 7046 39828 7098
rect 39880 7046 39892 7098
rect 39944 7046 39956 7098
rect 40008 7046 40020 7098
rect 40072 7046 40084 7098
rect 40136 7046 45540 7098
rect 1104 7024 45540 7046
rect 9950 6944 9956 6996
rect 10008 6984 10014 6996
rect 10008 6956 12434 6984
rect 10008 6944 10014 6956
rect 12406 6916 12434 6956
rect 14182 6944 14188 6996
rect 14240 6984 14246 6996
rect 22738 6984 22744 6996
rect 14240 6956 22744 6984
rect 14240 6944 14246 6956
rect 22738 6944 22744 6956
rect 22796 6944 22802 6996
rect 17954 6916 17960 6928
rect 12406 6888 17960 6916
rect 17954 6876 17960 6888
rect 18012 6876 18018 6928
rect 21634 6916 21640 6928
rect 18064 6888 21640 6916
rect 1210 6808 1216 6860
rect 1268 6848 1274 6860
rect 1765 6851 1823 6857
rect 1765 6848 1777 6851
rect 1268 6820 1777 6848
rect 1268 6808 1274 6820
rect 1765 6817 1777 6820
rect 1811 6817 1823 6851
rect 1765 6811 1823 6817
rect 16666 6808 16672 6860
rect 16724 6848 16730 6860
rect 18064 6848 18092 6888
rect 21634 6876 21640 6888
rect 21692 6876 21698 6928
rect 22462 6876 22468 6928
rect 22520 6916 22526 6928
rect 27246 6916 27252 6928
rect 22520 6888 27252 6916
rect 22520 6876 22526 6888
rect 27246 6876 27252 6888
rect 27304 6876 27310 6928
rect 16724 6820 18092 6848
rect 16724 6808 16730 6820
rect 19426 6808 19432 6860
rect 19484 6848 19490 6860
rect 26326 6848 26332 6860
rect 19484 6820 26332 6848
rect 19484 6808 19490 6820
rect 26326 6808 26332 6820
rect 26384 6808 26390 6860
rect 44729 6851 44787 6857
rect 44729 6817 44741 6851
rect 44775 6848 44787 6851
rect 45278 6848 45284 6860
rect 44775 6820 45284 6848
rect 44775 6817 44787 6820
rect 44729 6811 44787 6817
rect 45278 6808 45284 6820
rect 45336 6808 45342 6860
rect 46106 6808 46112 6860
rect 46164 6808 46170 6860
rect 14642 6740 14648 6792
rect 14700 6780 14706 6792
rect 20070 6780 20076 6792
rect 14700 6752 20076 6780
rect 14700 6740 14706 6752
rect 20070 6740 20076 6752
rect 20128 6740 20134 6792
rect 20162 6740 20168 6792
rect 20220 6780 20226 6792
rect 24210 6780 24216 6792
rect 20220 6752 24216 6780
rect 20220 6740 20226 6752
rect 24210 6740 24216 6752
rect 24268 6740 24274 6792
rect 44269 6783 44327 6789
rect 44269 6749 44281 6783
rect 44315 6780 44327 6783
rect 46124 6780 46152 6808
rect 44315 6752 46152 6780
rect 44315 6749 44327 6752
rect 44269 6743 44327 6749
rect 1486 6672 1492 6724
rect 1544 6672 1550 6724
rect 12342 6672 12348 6724
rect 12400 6712 12406 6724
rect 12400 6684 17356 6712
rect 12400 6672 12406 6684
rect 3326 6604 3332 6656
rect 3384 6644 3390 6656
rect 17218 6644 17224 6656
rect 3384 6616 17224 6644
rect 3384 6604 3390 6616
rect 17218 6604 17224 6616
rect 17276 6604 17282 6656
rect 17328 6644 17356 6684
rect 43898 6672 43904 6724
rect 43956 6672 43962 6724
rect 44450 6672 44456 6724
rect 44508 6672 44514 6724
rect 23106 6644 23112 6656
rect 17328 6616 23112 6644
rect 23106 6604 23112 6616
rect 23164 6604 23170 6656
rect 1104 6554 45696 6576
rect 1104 6502 12058 6554
rect 12110 6502 12122 6554
rect 12174 6502 12186 6554
rect 12238 6502 12250 6554
rect 12302 6502 12314 6554
rect 12366 6502 23166 6554
rect 23218 6502 23230 6554
rect 23282 6502 23294 6554
rect 23346 6502 23358 6554
rect 23410 6502 23422 6554
rect 23474 6502 34274 6554
rect 34326 6502 34338 6554
rect 34390 6502 34402 6554
rect 34454 6502 34466 6554
rect 34518 6502 34530 6554
rect 34582 6502 45382 6554
rect 45434 6502 45446 6554
rect 45498 6502 45510 6554
rect 45562 6502 45574 6554
rect 45626 6502 45638 6554
rect 45690 6502 45696 6554
rect 1104 6480 45696 6502
rect 1486 6400 1492 6452
rect 1544 6400 1550 6452
rect 14458 6440 14464 6452
rect 6886 6412 14464 6440
rect 1504 6304 1532 6400
rect 2498 6332 2504 6384
rect 2556 6372 2562 6384
rect 6886 6372 6914 6412
rect 14458 6400 14464 6412
rect 14516 6400 14522 6452
rect 14550 6400 14556 6452
rect 14608 6440 14614 6452
rect 14608 6412 17172 6440
rect 14608 6400 14614 6412
rect 2556 6344 6914 6372
rect 17144 6372 17172 6412
rect 17218 6400 17224 6452
rect 17276 6440 17282 6452
rect 25130 6440 25136 6452
rect 17276 6412 25136 6440
rect 17276 6400 17282 6412
rect 25130 6400 25136 6412
rect 25188 6400 25194 6452
rect 44634 6400 44640 6452
rect 44692 6440 44698 6452
rect 44913 6443 44971 6449
rect 44913 6440 44925 6443
rect 44692 6412 44925 6440
rect 44692 6400 44698 6412
rect 44913 6409 44925 6412
rect 44959 6409 44971 6443
rect 44913 6403 44971 6409
rect 22830 6372 22836 6384
rect 17144 6344 22836 6372
rect 2556 6332 2562 6344
rect 22830 6332 22836 6344
rect 22888 6332 22894 6384
rect 24854 6332 24860 6384
rect 24912 6372 24918 6384
rect 32766 6372 32772 6384
rect 24912 6344 32772 6372
rect 24912 6332 24918 6344
rect 32766 6332 32772 6344
rect 32824 6332 32830 6384
rect 18506 6304 18512 6316
rect 1504 6276 18512 6304
rect 18506 6264 18512 6276
rect 18564 6264 18570 6316
rect 24210 6264 24216 6316
rect 24268 6304 24274 6316
rect 35986 6304 35992 6316
rect 24268 6276 35992 6304
rect 24268 6264 24274 6276
rect 35986 6264 35992 6276
rect 36044 6264 36050 6316
rect 44818 6264 44824 6316
rect 44876 6264 44882 6316
rect 2958 6196 2964 6248
rect 3016 6236 3022 6248
rect 3016 6208 9674 6236
rect 3016 6196 3022 6208
rect 9646 6100 9674 6208
rect 14458 6196 14464 6248
rect 14516 6236 14522 6248
rect 25682 6236 25688 6248
rect 14516 6208 25688 6236
rect 14516 6196 14522 6208
rect 25682 6196 25688 6208
rect 25740 6196 25746 6248
rect 27062 6196 27068 6248
rect 27120 6236 27126 6248
rect 42794 6236 42800 6248
rect 27120 6208 42800 6236
rect 27120 6196 27126 6208
rect 42794 6196 42800 6208
rect 42852 6196 42858 6248
rect 25406 6168 25412 6180
rect 19306 6140 25412 6168
rect 19306 6100 19334 6140
rect 25406 6128 25412 6140
rect 25464 6128 25470 6180
rect 25498 6128 25504 6180
rect 25556 6168 25562 6180
rect 42518 6168 42524 6180
rect 25556 6140 42524 6168
rect 25556 6128 25562 6140
rect 42518 6128 42524 6140
rect 42576 6128 42582 6180
rect 9646 6072 19334 6100
rect 1104 6010 45540 6032
rect 1104 5958 6504 6010
rect 6556 5958 6568 6010
rect 6620 5958 6632 6010
rect 6684 5958 6696 6010
rect 6748 5958 6760 6010
rect 6812 5958 17612 6010
rect 17664 5958 17676 6010
rect 17728 5958 17740 6010
rect 17792 5958 17804 6010
rect 17856 5958 17868 6010
rect 17920 5958 28720 6010
rect 28772 5958 28784 6010
rect 28836 5958 28848 6010
rect 28900 5958 28912 6010
rect 28964 5958 28976 6010
rect 29028 5958 39828 6010
rect 39880 5958 39892 6010
rect 39944 5958 39956 6010
rect 40008 5958 40020 6010
rect 40072 5958 40084 6010
rect 40136 5958 45540 6010
rect 1104 5936 45540 5958
rect 1104 5466 45696 5488
rect 1104 5414 12058 5466
rect 12110 5414 12122 5466
rect 12174 5414 12186 5466
rect 12238 5414 12250 5466
rect 12302 5414 12314 5466
rect 12366 5414 23166 5466
rect 23218 5414 23230 5466
rect 23282 5414 23294 5466
rect 23346 5414 23358 5466
rect 23410 5414 23422 5466
rect 23474 5414 34274 5466
rect 34326 5414 34338 5466
rect 34390 5414 34402 5466
rect 34454 5414 34466 5466
rect 34518 5414 34530 5466
rect 34582 5414 45382 5466
rect 45434 5414 45446 5466
rect 45498 5414 45510 5466
rect 45562 5414 45574 5466
rect 45626 5414 45638 5466
rect 45690 5414 45696 5466
rect 1104 5392 45696 5414
rect 23014 5108 23020 5160
rect 23072 5148 23078 5160
rect 33042 5148 33048 5160
rect 23072 5120 33048 5148
rect 23072 5108 23078 5120
rect 33042 5108 33048 5120
rect 33100 5108 33106 5160
rect 22830 5040 22836 5092
rect 22888 5080 22894 5092
rect 35618 5080 35624 5092
rect 22888 5052 35624 5080
rect 22888 5040 22894 5052
rect 35618 5040 35624 5052
rect 35676 5040 35682 5092
rect 20530 4972 20536 5024
rect 20588 5012 20594 5024
rect 33778 5012 33784 5024
rect 20588 4984 33784 5012
rect 20588 4972 20594 4984
rect 33778 4972 33784 4984
rect 33836 4972 33842 5024
rect 1104 4922 45540 4944
rect 1104 4870 6504 4922
rect 6556 4870 6568 4922
rect 6620 4870 6632 4922
rect 6684 4870 6696 4922
rect 6748 4870 6760 4922
rect 6812 4870 17612 4922
rect 17664 4870 17676 4922
rect 17728 4870 17740 4922
rect 17792 4870 17804 4922
rect 17856 4870 17868 4922
rect 17920 4870 28720 4922
rect 28772 4870 28784 4922
rect 28836 4870 28848 4922
rect 28900 4870 28912 4922
rect 28964 4870 28976 4922
rect 29028 4870 39828 4922
rect 39880 4870 39892 4922
rect 39944 4870 39956 4922
rect 40008 4870 40020 4922
rect 40072 4870 40084 4922
rect 40136 4870 45540 4922
rect 1104 4848 45540 4870
rect 29270 4768 29276 4820
rect 29328 4808 29334 4820
rect 43346 4808 43352 4820
rect 29328 4780 43352 4808
rect 29328 4768 29334 4780
rect 43346 4768 43352 4780
rect 43404 4768 43410 4820
rect 1104 4378 45696 4400
rect 1104 4326 12058 4378
rect 12110 4326 12122 4378
rect 12174 4326 12186 4378
rect 12238 4326 12250 4378
rect 12302 4326 12314 4378
rect 12366 4326 23166 4378
rect 23218 4326 23230 4378
rect 23282 4326 23294 4378
rect 23346 4326 23358 4378
rect 23410 4326 23422 4378
rect 23474 4326 34274 4378
rect 34326 4326 34338 4378
rect 34390 4326 34402 4378
rect 34454 4326 34466 4378
rect 34518 4326 34530 4378
rect 34582 4326 45382 4378
rect 45434 4326 45446 4378
rect 45498 4326 45510 4378
rect 45562 4326 45574 4378
rect 45626 4326 45638 4378
rect 45690 4326 45696 4378
rect 1104 4304 45696 4326
rect 1104 3834 45540 3856
rect 1104 3782 6504 3834
rect 6556 3782 6568 3834
rect 6620 3782 6632 3834
rect 6684 3782 6696 3834
rect 6748 3782 6760 3834
rect 6812 3782 17612 3834
rect 17664 3782 17676 3834
rect 17728 3782 17740 3834
rect 17792 3782 17804 3834
rect 17856 3782 17868 3834
rect 17920 3782 28720 3834
rect 28772 3782 28784 3834
rect 28836 3782 28848 3834
rect 28900 3782 28912 3834
rect 28964 3782 28976 3834
rect 29028 3782 39828 3834
rect 39880 3782 39892 3834
rect 39944 3782 39956 3834
rect 40008 3782 40020 3834
rect 40072 3782 40084 3834
rect 40136 3782 45540 3834
rect 1104 3760 45540 3782
rect 23658 3612 23664 3664
rect 23716 3652 23722 3664
rect 33870 3652 33876 3664
rect 23716 3624 33876 3652
rect 23716 3612 23722 3624
rect 33870 3612 33876 3624
rect 33928 3612 33934 3664
rect 22738 3544 22744 3596
rect 22796 3584 22802 3596
rect 35342 3584 35348 3596
rect 22796 3556 35348 3584
rect 22796 3544 22802 3556
rect 35342 3544 35348 3556
rect 35400 3544 35406 3596
rect 23934 3476 23940 3528
rect 23992 3516 23998 3528
rect 37182 3516 37188 3528
rect 23992 3488 37188 3516
rect 23992 3476 23998 3488
rect 37182 3476 37188 3488
rect 37240 3476 37246 3528
rect 20622 3408 20628 3460
rect 20680 3448 20686 3460
rect 38562 3448 38568 3460
rect 20680 3420 38568 3448
rect 20680 3408 20686 3420
rect 38562 3408 38568 3420
rect 38620 3408 38626 3460
rect 1104 3290 45696 3312
rect 1104 3238 12058 3290
rect 12110 3238 12122 3290
rect 12174 3238 12186 3290
rect 12238 3238 12250 3290
rect 12302 3238 12314 3290
rect 12366 3238 23166 3290
rect 23218 3238 23230 3290
rect 23282 3238 23294 3290
rect 23346 3238 23358 3290
rect 23410 3238 23422 3290
rect 23474 3238 34274 3290
rect 34326 3238 34338 3290
rect 34390 3238 34402 3290
rect 34454 3238 34466 3290
rect 34518 3238 34530 3290
rect 34582 3238 45382 3290
rect 45434 3238 45446 3290
rect 45498 3238 45510 3290
rect 45562 3238 45574 3290
rect 45626 3238 45638 3290
rect 45690 3238 45696 3290
rect 1104 3216 45696 3238
rect 1104 2746 45540 2768
rect 1104 2694 6504 2746
rect 6556 2694 6568 2746
rect 6620 2694 6632 2746
rect 6684 2694 6696 2746
rect 6748 2694 6760 2746
rect 6812 2694 17612 2746
rect 17664 2694 17676 2746
rect 17728 2694 17740 2746
rect 17792 2694 17804 2746
rect 17856 2694 17868 2746
rect 17920 2694 28720 2746
rect 28772 2694 28784 2746
rect 28836 2694 28848 2746
rect 28900 2694 28912 2746
rect 28964 2694 28976 2746
rect 29028 2694 39828 2746
rect 39880 2694 39892 2746
rect 39944 2694 39956 2746
rect 40008 2694 40020 2746
rect 40072 2694 40084 2746
rect 40136 2694 45540 2746
rect 1104 2672 45540 2694
rect 20441 2635 20499 2641
rect 20441 2601 20453 2635
rect 20487 2632 20499 2635
rect 20530 2632 20536 2644
rect 20487 2604 20536 2632
rect 20487 2601 20499 2604
rect 20441 2595 20499 2601
rect 20530 2592 20536 2604
rect 20588 2592 20594 2644
rect 22373 2635 22431 2641
rect 22373 2601 22385 2635
rect 22419 2632 22431 2635
rect 22922 2632 22928 2644
rect 22419 2604 22928 2632
rect 22419 2601 22431 2604
rect 22373 2595 22431 2601
rect 22922 2592 22928 2604
rect 22980 2592 22986 2644
rect 23014 2592 23020 2644
rect 23072 2632 23078 2644
rect 23385 2635 23443 2641
rect 23385 2632 23397 2635
rect 23072 2604 23397 2632
rect 23072 2592 23078 2604
rect 23385 2601 23397 2604
rect 23431 2601 23443 2635
rect 23385 2595 23443 2601
rect 23658 2592 23664 2644
rect 23716 2592 23722 2644
rect 23934 2592 23940 2644
rect 23992 2592 23998 2644
rect 24210 2592 24216 2644
rect 24268 2592 24274 2644
rect 24854 2592 24860 2644
rect 24912 2592 24918 2644
rect 27062 2592 27068 2644
rect 27120 2592 27126 2644
rect 29270 2592 29276 2644
rect 29328 2592 29334 2644
rect 43254 2632 43260 2644
rect 31726 2604 43260 2632
rect 22741 2567 22799 2573
rect 22741 2533 22753 2567
rect 22787 2564 22799 2567
rect 31481 2567 31539 2573
rect 22787 2536 26234 2564
rect 22787 2533 22799 2536
rect 22741 2527 22799 2533
rect 22278 2456 22284 2508
rect 22336 2496 22342 2508
rect 22336 2468 23244 2496
rect 22336 2456 22342 2468
rect 22186 2388 22192 2440
rect 22244 2388 22250 2440
rect 22462 2388 22468 2440
rect 22520 2428 22526 2440
rect 23216 2437 23244 2468
rect 23290 2456 23296 2508
rect 23348 2496 23354 2508
rect 25498 2496 25504 2508
rect 23348 2468 25504 2496
rect 23348 2456 23354 2468
rect 25498 2456 25504 2468
rect 25556 2456 25562 2508
rect 22925 2431 22983 2437
rect 22925 2428 22937 2431
rect 22520 2400 22937 2428
rect 22520 2388 22526 2400
rect 22925 2397 22937 2400
rect 22971 2397 22983 2431
rect 22925 2391 22983 2397
rect 23201 2431 23259 2437
rect 23201 2397 23213 2431
rect 23247 2397 23259 2431
rect 23201 2391 23259 2397
rect 23477 2431 23535 2437
rect 23477 2397 23489 2431
rect 23523 2397 23535 2431
rect 23477 2391 23535 2397
rect 20346 2320 20352 2372
rect 20404 2320 20410 2372
rect 21450 2320 21456 2372
rect 21508 2360 21514 2372
rect 22557 2363 22615 2369
rect 22557 2360 22569 2363
rect 21508 2332 22569 2360
rect 21508 2320 21514 2332
rect 22557 2329 22569 2332
rect 22603 2329 22615 2363
rect 22557 2323 22615 2329
rect 22830 2320 22836 2372
rect 22888 2320 22894 2372
rect 23014 2320 23020 2372
rect 23072 2360 23078 2372
rect 23492 2360 23520 2391
rect 23750 2388 23756 2440
rect 23808 2388 23814 2440
rect 23934 2388 23940 2440
rect 23992 2428 23998 2440
rect 24029 2431 24087 2437
rect 24029 2428 24041 2431
rect 23992 2400 24041 2428
rect 23992 2388 23998 2400
rect 24029 2397 24041 2400
rect 24075 2397 24087 2431
rect 24029 2391 24087 2397
rect 24670 2388 24676 2440
rect 24728 2388 24734 2440
rect 23072 2332 23520 2360
rect 26206 2360 26234 2536
rect 31481 2533 31493 2567
rect 31527 2564 31539 2567
rect 31726 2564 31754 2604
rect 43254 2592 43260 2604
rect 43312 2592 43318 2644
rect 43898 2592 43904 2644
rect 43956 2592 43962 2644
rect 44174 2592 44180 2644
rect 44232 2592 44238 2644
rect 44266 2592 44272 2644
rect 44324 2592 44330 2644
rect 44450 2592 44456 2644
rect 44508 2592 44514 2644
rect 45002 2592 45008 2644
rect 45060 2592 45066 2644
rect 31527 2536 31754 2564
rect 33689 2567 33747 2573
rect 31527 2533 31539 2536
rect 31481 2527 31539 2533
rect 33689 2533 33701 2567
rect 33735 2533 33747 2567
rect 33689 2527 33747 2533
rect 35897 2567 35955 2573
rect 35897 2533 35909 2567
rect 35943 2564 35955 2567
rect 39666 2564 39672 2576
rect 35943 2536 39672 2564
rect 35943 2533 35955 2536
rect 35897 2527 35955 2533
rect 33704 2496 33732 2527
rect 39666 2524 39672 2536
rect 39724 2524 39730 2576
rect 44284 2564 44312 2592
rect 41386 2536 44312 2564
rect 41386 2496 41414 2536
rect 33704 2468 41414 2496
rect 41598 2456 41604 2508
rect 41656 2496 41662 2508
rect 41656 2468 44680 2496
rect 41656 2456 41662 2468
rect 26878 2388 26884 2440
rect 26936 2388 26942 2440
rect 29086 2388 29092 2440
rect 29144 2388 29150 2440
rect 31294 2388 31300 2440
rect 31352 2388 31358 2440
rect 33502 2388 33508 2440
rect 33560 2388 33566 2440
rect 35710 2388 35716 2440
rect 35768 2388 35774 2440
rect 37918 2388 37924 2440
rect 37976 2388 37982 2440
rect 44082 2388 44088 2440
rect 44140 2388 44146 2440
rect 44652 2437 44680 2468
rect 44361 2431 44419 2437
rect 44361 2397 44373 2431
rect 44407 2397 44419 2431
rect 44361 2391 44419 2397
rect 44637 2431 44695 2437
rect 44637 2397 44649 2431
rect 44683 2397 44695 2431
rect 44637 2391 44695 2397
rect 36078 2360 36084 2372
rect 26206 2332 36084 2360
rect 23072 2320 23078 2332
rect 36078 2320 36084 2332
rect 36136 2320 36142 2372
rect 43438 2320 43444 2372
rect 43496 2360 43502 2372
rect 44376 2360 44404 2391
rect 44818 2388 44824 2440
rect 44876 2388 44882 2440
rect 45186 2388 45192 2440
rect 45244 2388 45250 2440
rect 43496 2332 44404 2360
rect 43496 2320 43502 2332
rect 22848 2292 22876 2320
rect 23109 2295 23167 2301
rect 23109 2292 23121 2295
rect 22848 2264 23121 2292
rect 23109 2261 23121 2264
rect 23155 2261 23167 2295
rect 23109 2255 23167 2261
rect 38105 2295 38163 2301
rect 38105 2261 38117 2295
rect 38151 2292 38163 2295
rect 44836 2292 44864 2388
rect 38151 2264 44864 2292
rect 38151 2261 38163 2264
rect 38105 2255 38163 2261
rect 1104 2202 45696 2224
rect 1104 2150 12058 2202
rect 12110 2150 12122 2202
rect 12174 2150 12186 2202
rect 12238 2150 12250 2202
rect 12302 2150 12314 2202
rect 12366 2150 23166 2202
rect 23218 2150 23230 2202
rect 23282 2150 23294 2202
rect 23346 2150 23358 2202
rect 23410 2150 23422 2202
rect 23474 2150 34274 2202
rect 34326 2150 34338 2202
rect 34390 2150 34402 2202
rect 34454 2150 34466 2202
rect 34518 2150 34530 2202
rect 34582 2150 45382 2202
rect 45434 2150 45446 2202
rect 45498 2150 45510 2202
rect 45562 2150 45574 2202
rect 45626 2150 45638 2202
rect 45690 2150 45696 2202
rect 1104 2128 45696 2150
rect 19429 2091 19487 2097
rect 19429 2057 19441 2091
rect 19475 2088 19487 2091
rect 20346 2088 20352 2100
rect 19475 2060 20352 2088
rect 19475 2057 19487 2060
rect 19429 2051 19487 2057
rect 20346 2048 20352 2060
rect 20404 2048 20410 2100
rect 20622 2048 20628 2100
rect 20680 2048 20686 2100
rect 21177 2091 21235 2097
rect 21177 2057 21189 2091
rect 21223 2088 21235 2091
rect 22186 2088 22192 2100
rect 21223 2060 22192 2088
rect 21223 2057 21235 2060
rect 21177 2051 21235 2057
rect 22186 2048 22192 2060
rect 22244 2048 22250 2100
rect 22278 2048 22284 2100
rect 22336 2048 22342 2100
rect 22557 2091 22615 2097
rect 22557 2057 22569 2091
rect 22603 2057 22615 2091
rect 22557 2051 22615 2057
rect 20257 2023 20315 2029
rect 6886 1992 20116 2020
rect 1578 1912 1584 1964
rect 1636 1952 1642 1964
rect 6886 1952 6914 1992
rect 1636 1924 6914 1952
rect 1636 1912 1642 1924
rect 19610 1912 19616 1964
rect 19668 1912 19674 1964
rect 20088 1961 20116 1992
rect 20257 1989 20269 2023
rect 20303 2020 20315 2023
rect 20640 2020 20668 2048
rect 20303 1992 20668 2020
rect 22572 2020 22600 2051
rect 23014 2048 23020 2100
rect 23072 2088 23078 2100
rect 23109 2091 23167 2097
rect 23109 2088 23121 2091
rect 23072 2060 23121 2088
rect 23072 2048 23078 2060
rect 23109 2057 23121 2060
rect 23155 2057 23167 2091
rect 23109 2051 23167 2057
rect 23385 2091 23443 2097
rect 23385 2057 23397 2091
rect 23431 2088 23443 2091
rect 23750 2088 23756 2100
rect 23431 2060 23756 2088
rect 23431 2057 23443 2060
rect 23385 2051 23443 2057
rect 23750 2048 23756 2060
rect 23808 2048 23814 2100
rect 23845 2091 23903 2097
rect 23845 2057 23857 2091
rect 23891 2088 23903 2091
rect 24670 2088 24676 2100
rect 23891 2060 24676 2088
rect 23891 2057 23903 2060
rect 23845 2051 23903 2057
rect 24670 2048 24676 2060
rect 24728 2048 24734 2100
rect 26053 2091 26111 2097
rect 26053 2057 26065 2091
rect 26099 2088 26111 2091
rect 26878 2088 26884 2100
rect 26099 2060 26884 2088
rect 26099 2057 26111 2060
rect 26053 2051 26111 2057
rect 26878 2048 26884 2060
rect 26936 2048 26942 2100
rect 28261 2091 28319 2097
rect 28261 2057 28273 2091
rect 28307 2088 28319 2091
rect 29086 2088 29092 2100
rect 28307 2060 29092 2088
rect 28307 2057 28319 2060
rect 28261 2051 28319 2057
rect 29086 2048 29092 2060
rect 29144 2048 29150 2100
rect 30469 2091 30527 2097
rect 30469 2057 30481 2091
rect 30515 2088 30527 2091
rect 31294 2088 31300 2100
rect 30515 2060 31300 2088
rect 30515 2057 30527 2060
rect 30469 2051 30527 2057
rect 31294 2048 31300 2060
rect 31352 2048 31358 2100
rect 32677 2091 32735 2097
rect 32677 2057 32689 2091
rect 32723 2088 32735 2091
rect 33502 2088 33508 2100
rect 32723 2060 33508 2088
rect 32723 2057 32735 2060
rect 32677 2051 32735 2057
rect 33502 2048 33508 2060
rect 33560 2048 33566 2100
rect 34885 2091 34943 2097
rect 34885 2057 34897 2091
rect 34931 2088 34943 2091
rect 35710 2088 35716 2100
rect 34931 2060 35716 2088
rect 34931 2057 34943 2060
rect 34885 2051 34943 2057
rect 35710 2048 35716 2060
rect 35768 2048 35774 2100
rect 37277 2091 37335 2097
rect 37277 2057 37289 2091
rect 37323 2088 37335 2091
rect 37918 2088 37924 2100
rect 37323 2060 37924 2088
rect 37323 2057 37335 2060
rect 37277 2051 37335 2057
rect 37918 2048 37924 2060
rect 37976 2048 37982 2100
rect 41598 2048 41604 2100
rect 41656 2048 41662 2100
rect 43438 2048 43444 2100
rect 43496 2048 43502 2100
rect 43901 2091 43959 2097
rect 43901 2057 43913 2091
rect 43947 2057 43959 2091
rect 43901 2051 43959 2057
rect 23934 2020 23940 2032
rect 22572 1992 23940 2020
rect 20303 1989 20315 1992
rect 20257 1983 20315 1989
rect 23934 1980 23940 1992
rect 23992 1980 23998 2032
rect 43916 2020 43944 2051
rect 44082 2048 44088 2100
rect 44140 2088 44146 2100
rect 44361 2091 44419 2097
rect 44361 2088 44373 2091
rect 44140 2060 44373 2088
rect 44140 2048 44146 2060
rect 44361 2057 44373 2060
rect 44407 2057 44419 2091
rect 44361 2051 44419 2057
rect 45186 2020 45192 2032
rect 43916 1992 45192 2020
rect 45186 1980 45192 1992
rect 45244 1980 45250 2032
rect 20073 1955 20131 1961
rect 20073 1921 20085 1955
rect 20119 1921 20131 1955
rect 20073 1915 20131 1921
rect 20714 1912 20720 1964
rect 20772 1952 20778 1964
rect 21361 1955 21419 1961
rect 21361 1952 21373 1955
rect 20772 1924 21373 1952
rect 20772 1912 20778 1924
rect 21361 1921 21373 1924
rect 21407 1921 21419 1955
rect 21361 1915 21419 1921
rect 21634 1912 21640 1964
rect 21692 1912 21698 1964
rect 22186 1912 22192 1964
rect 22244 1912 22250 1964
rect 22465 1955 22523 1961
rect 22465 1921 22477 1955
rect 22511 1921 22523 1955
rect 22465 1915 22523 1921
rect 22741 1955 22799 1961
rect 22741 1921 22753 1955
rect 22787 1921 22799 1955
rect 22741 1915 22799 1921
rect 20806 1844 20812 1896
rect 20864 1884 20870 1896
rect 22480 1884 22508 1915
rect 22756 1884 22784 1915
rect 22830 1912 22836 1964
rect 22888 1912 22894 1964
rect 23014 1912 23020 1964
rect 23072 1952 23078 1964
rect 23293 1955 23351 1961
rect 23293 1952 23305 1955
rect 23072 1924 23305 1952
rect 23072 1912 23078 1924
rect 23293 1921 23305 1924
rect 23339 1921 23351 1955
rect 23293 1915 23351 1921
rect 23569 1955 23627 1961
rect 23569 1921 23581 1955
rect 23615 1952 23627 1955
rect 23658 1952 23664 1964
rect 23615 1924 23664 1952
rect 23615 1921 23627 1924
rect 23569 1915 23627 1921
rect 23658 1912 23664 1924
rect 23716 1912 23722 1964
rect 24026 1912 24032 1964
rect 24084 1912 24090 1964
rect 26234 1912 26240 1964
rect 26292 1912 26298 1964
rect 28442 1912 28448 1964
rect 28500 1912 28506 1964
rect 30650 1912 30656 1964
rect 30708 1912 30714 1964
rect 32858 1912 32864 1964
rect 32916 1912 32922 1964
rect 35066 1912 35072 1964
rect 35124 1912 35130 1964
rect 37458 1912 37464 1964
rect 37516 1912 37522 1964
rect 41782 1912 41788 1964
rect 41840 1912 41846 1964
rect 43622 1912 43628 1964
rect 43680 1912 43686 1964
rect 44082 1912 44088 1964
rect 44140 1912 44146 1964
rect 44542 1912 44548 1964
rect 44600 1912 44606 1964
rect 20864 1856 22508 1884
rect 22572 1856 22784 1884
rect 20864 1844 20870 1856
rect 22005 1819 22063 1825
rect 22005 1785 22017 1819
rect 22051 1816 22063 1819
rect 22462 1816 22468 1828
rect 22051 1788 22468 1816
rect 22051 1785 22063 1788
rect 22005 1779 22063 1785
rect 22462 1776 22468 1788
rect 22520 1776 22526 1828
rect 21450 1708 21456 1760
rect 21508 1708 21514 1760
rect 21542 1708 21548 1760
rect 21600 1748 21606 1760
rect 22572 1748 22600 1856
rect 21600 1720 22600 1748
rect 21600 1708 21606 1720
rect 22738 1708 22744 1760
rect 22796 1748 22802 1760
rect 23017 1751 23075 1757
rect 23017 1748 23029 1751
rect 22796 1720 23029 1748
rect 22796 1708 22802 1720
rect 23017 1717 23029 1720
rect 23063 1717 23075 1751
rect 23017 1711 23075 1717
rect 1104 1658 45540 1680
rect 1104 1606 6504 1658
rect 6556 1606 6568 1658
rect 6620 1606 6632 1658
rect 6684 1606 6696 1658
rect 6748 1606 6760 1658
rect 6812 1606 17612 1658
rect 17664 1606 17676 1658
rect 17728 1606 17740 1658
rect 17792 1606 17804 1658
rect 17856 1606 17868 1658
rect 17920 1606 28720 1658
rect 28772 1606 28784 1658
rect 28836 1606 28848 1658
rect 28900 1606 28912 1658
rect 28964 1606 28976 1658
rect 29028 1606 39828 1658
rect 39880 1606 39892 1658
rect 39944 1606 39956 1658
rect 40008 1606 40020 1658
rect 40072 1606 40084 1658
rect 40136 1606 45540 1658
rect 1104 1584 45540 1606
rect 1578 1504 1584 1556
rect 1636 1504 1642 1556
rect 19245 1547 19303 1553
rect 19245 1513 19257 1547
rect 19291 1544 19303 1547
rect 19610 1544 19616 1556
rect 19291 1516 19616 1544
rect 19291 1513 19303 1516
rect 19245 1507 19303 1513
rect 19610 1504 19616 1516
rect 19668 1504 19674 1556
rect 21177 1547 21235 1553
rect 21177 1513 21189 1547
rect 21223 1544 21235 1547
rect 21634 1544 21640 1556
rect 21223 1516 21640 1544
rect 21223 1513 21235 1516
rect 21177 1507 21235 1513
rect 21634 1504 21640 1516
rect 21692 1504 21698 1556
rect 22097 1547 22155 1553
rect 22097 1513 22109 1547
rect 22143 1544 22155 1547
rect 22830 1544 22836 1556
rect 22143 1516 22836 1544
rect 22143 1513 22155 1516
rect 22097 1507 22155 1513
rect 22830 1504 22836 1516
rect 22888 1504 22894 1556
rect 23385 1547 23443 1553
rect 23385 1513 23397 1547
rect 23431 1544 23443 1547
rect 24026 1544 24032 1556
rect 23431 1516 24032 1544
rect 23431 1513 23443 1516
rect 23385 1507 23443 1513
rect 24026 1504 24032 1516
rect 24084 1504 24090 1556
rect 27801 1547 27859 1553
rect 27801 1513 27813 1547
rect 27847 1544 27859 1547
rect 28442 1544 28448 1556
rect 27847 1516 28448 1544
rect 27847 1513 27859 1516
rect 27801 1507 27859 1513
rect 28442 1504 28448 1516
rect 28500 1504 28506 1556
rect 32217 1547 32275 1553
rect 32217 1513 32229 1547
rect 32263 1544 32275 1547
rect 32858 1544 32864 1556
rect 32263 1516 32864 1544
rect 32263 1513 32275 1516
rect 32217 1507 32275 1513
rect 32858 1504 32864 1516
rect 32916 1504 32922 1556
rect 34701 1547 34759 1553
rect 34701 1513 34713 1547
rect 34747 1544 34759 1547
rect 35066 1544 35072 1556
rect 34747 1516 35072 1544
rect 34747 1513 34759 1516
rect 34701 1507 34759 1513
rect 35066 1504 35072 1516
rect 35124 1504 35130 1556
rect 43257 1547 43315 1553
rect 43257 1513 43269 1547
rect 43303 1544 43315 1547
rect 44082 1544 44088 1556
rect 43303 1516 44088 1544
rect 43303 1513 43315 1516
rect 43257 1507 43315 1513
rect 44082 1504 44088 1516
rect 44140 1504 44146 1556
rect 44542 1504 44548 1556
rect 44600 1544 44606 1556
rect 45005 1547 45063 1553
rect 45005 1544 45017 1547
rect 44600 1516 45017 1544
rect 44600 1504 44606 1516
rect 45005 1513 45017 1516
rect 45051 1513 45063 1547
rect 45005 1507 45063 1513
rect 14660 1380 14872 1408
rect 1210 1300 1216 1352
rect 1268 1340 1274 1352
rect 1397 1343 1455 1349
rect 1397 1340 1409 1343
rect 1268 1312 1409 1340
rect 1268 1300 1274 1312
rect 1397 1309 1409 1312
rect 1443 1309 1455 1343
rect 1397 1303 1455 1309
rect 3786 1300 3792 1352
rect 3844 1300 3850 1352
rect 5718 1300 5724 1352
rect 5776 1300 5782 1352
rect 7926 1300 7932 1352
rect 7984 1300 7990 1352
rect 10134 1300 10140 1352
rect 10192 1300 10198 1352
rect 12066 1300 12072 1352
rect 12124 1340 12130 1352
rect 12345 1343 12403 1349
rect 12345 1340 12357 1343
rect 12124 1312 12357 1340
rect 12124 1300 12130 1312
rect 12345 1309 12357 1312
rect 12391 1309 12403 1343
rect 14660 1340 14688 1380
rect 12345 1303 12403 1309
rect 12452 1312 14688 1340
rect 12452 1272 12480 1312
rect 14734 1300 14740 1352
rect 14792 1300 14798 1352
rect 14642 1272 14648 1284
rect 6886 1244 12480 1272
rect 12544 1244 14648 1272
rect 3970 1164 3976 1216
rect 4028 1164 4034 1216
rect 5905 1207 5963 1213
rect 5905 1173 5917 1207
rect 5951 1204 5963 1207
rect 6886 1204 6914 1244
rect 5951 1176 6914 1204
rect 5951 1173 5963 1176
rect 5905 1167 5963 1173
rect 8110 1164 8116 1216
rect 8168 1164 8174 1216
rect 10318 1164 10324 1216
rect 10376 1164 10382 1216
rect 12544 1213 12572 1244
rect 14642 1232 14648 1244
rect 14700 1232 14706 1284
rect 14844 1272 14872 1380
rect 16942 1300 16948 1352
rect 17000 1300 17006 1352
rect 19426 1300 19432 1352
rect 19484 1300 19490 1352
rect 19536 1312 20852 1340
rect 19536 1272 19564 1312
rect 14844 1244 19564 1272
rect 20714 1232 20720 1284
rect 20772 1232 20778 1284
rect 20824 1272 20852 1312
rect 21358 1300 21364 1352
rect 21416 1300 21422 1352
rect 22278 1300 22284 1352
rect 22336 1300 22342 1352
rect 23566 1300 23572 1352
rect 23624 1300 23630 1352
rect 25774 1300 25780 1352
rect 25832 1300 25838 1352
rect 27982 1300 27988 1352
rect 28040 1300 28046 1352
rect 30190 1300 30196 1352
rect 30248 1300 30254 1352
rect 30650 1300 30656 1352
rect 30708 1300 30714 1352
rect 32398 1300 32404 1352
rect 32456 1300 32462 1352
rect 34606 1300 34612 1352
rect 34664 1340 34670 1352
rect 34885 1343 34943 1349
rect 34885 1340 34897 1343
rect 34664 1312 34897 1340
rect 34664 1300 34670 1312
rect 34885 1309 34897 1312
rect 34931 1309 34943 1343
rect 34885 1303 34943 1309
rect 36814 1300 36820 1352
rect 36872 1300 36878 1352
rect 37458 1300 37464 1352
rect 37516 1300 37522 1352
rect 39022 1300 39028 1352
rect 39080 1300 39086 1352
rect 41230 1300 41236 1352
rect 41288 1300 41294 1352
rect 43438 1300 43444 1352
rect 43496 1300 43502 1352
rect 45186 1300 45192 1352
rect 45244 1300 45250 1352
rect 22186 1272 22192 1284
rect 20824 1244 22192 1272
rect 22186 1232 22192 1244
rect 22244 1232 22250 1284
rect 12529 1207 12587 1213
rect 12529 1173 12541 1207
rect 12575 1173 12587 1207
rect 12529 1167 12587 1173
rect 14550 1164 14556 1216
rect 14608 1164 14614 1216
rect 16761 1207 16819 1213
rect 16761 1173 16773 1207
rect 16807 1204 16819 1207
rect 20732 1204 20760 1232
rect 16807 1176 20760 1204
rect 25593 1207 25651 1213
rect 16807 1173 16819 1176
rect 16761 1167 16819 1173
rect 25593 1173 25605 1207
rect 25639 1204 25651 1207
rect 26234 1204 26240 1216
rect 25639 1176 26240 1204
rect 25639 1173 25651 1176
rect 25593 1167 25651 1173
rect 26234 1164 26240 1176
rect 26292 1164 26298 1216
rect 30009 1207 30067 1213
rect 30009 1173 30021 1207
rect 30055 1204 30067 1207
rect 30668 1204 30696 1300
rect 30055 1176 30696 1204
rect 36633 1207 36691 1213
rect 30055 1173 30067 1176
rect 30009 1167 30067 1173
rect 36633 1173 36645 1207
rect 36679 1204 36691 1207
rect 37476 1204 37504 1300
rect 43622 1272 43628 1284
rect 38856 1244 43628 1272
rect 38856 1213 38884 1244
rect 43622 1232 43628 1244
rect 43680 1232 43686 1284
rect 36679 1176 37504 1204
rect 38841 1207 38899 1213
rect 36679 1173 36691 1176
rect 36633 1167 36691 1173
rect 38841 1173 38853 1207
rect 38887 1173 38899 1207
rect 38841 1167 38899 1173
rect 41049 1207 41107 1213
rect 41049 1173 41061 1207
rect 41095 1204 41107 1207
rect 41782 1204 41788 1216
rect 41095 1176 41788 1204
rect 41095 1173 41107 1176
rect 41049 1167 41107 1173
rect 41782 1164 41788 1176
rect 41840 1164 41846 1216
rect 1104 1114 45696 1136
rect 1104 1062 12058 1114
rect 12110 1062 12122 1114
rect 12174 1062 12186 1114
rect 12238 1062 12250 1114
rect 12302 1062 12314 1114
rect 12366 1062 23166 1114
rect 23218 1062 23230 1114
rect 23282 1062 23294 1114
rect 23346 1062 23358 1114
rect 23410 1062 23422 1114
rect 23474 1062 34274 1114
rect 34326 1062 34338 1114
rect 34390 1062 34402 1114
rect 34454 1062 34466 1114
rect 34518 1062 34530 1114
rect 34582 1062 45382 1114
rect 45434 1062 45446 1114
rect 45498 1062 45510 1114
rect 45562 1062 45574 1114
rect 45626 1062 45638 1114
rect 45690 1062 45696 1114
rect 1104 1040 45696 1062
rect 3970 960 3976 1012
rect 4028 1000 4034 1012
rect 4028 972 6914 1000
rect 4028 960 4034 972
rect 6886 864 6914 972
rect 14550 960 14556 1012
rect 14608 960 14614 1012
rect 14642 960 14648 1012
rect 14700 1000 14706 1012
rect 20806 1000 20812 1012
rect 14700 972 20812 1000
rect 14700 960 14706 972
rect 20806 960 20812 972
rect 20864 960 20870 1012
rect 22278 960 22284 1012
rect 22336 960 22342 1012
rect 14568 932 14596 960
rect 22296 932 22324 960
rect 14568 904 22324 932
rect 23658 864 23664 876
rect 6886 836 23664 864
rect 23658 824 23664 836
rect 23716 824 23722 876
rect 8110 756 8116 808
rect 8168 756 8174 808
rect 10318 756 10324 808
rect 10376 796 10382 808
rect 23014 796 23020 808
rect 10376 768 23020 796
rect 10376 756 10382 768
rect 23014 756 23020 768
rect 23072 756 23078 808
rect 8128 660 8156 756
rect 21542 660 21548 672
rect 8128 632 21548 660
rect 21542 620 21548 632
rect 21600 620 21606 672
<< via1 >>
rect 13636 9936 13688 9988
rect 14924 9936 14976 9988
rect 18328 9936 18380 9988
rect 18420 9936 18472 9988
rect 19524 9936 19576 9988
rect 20628 9936 20680 9988
rect 35716 9936 35768 9988
rect 8760 9868 8812 9920
rect 14648 9868 14700 9920
rect 16488 9868 16540 9920
rect 19892 9868 19944 9920
rect 9496 9800 9548 9852
rect 14372 9800 14424 9852
rect 17684 9800 17736 9852
rect 28908 9800 28960 9852
rect 5356 9732 5408 9784
rect 8024 9732 8076 9784
rect 14556 9732 14608 9784
rect 16396 9732 16448 9784
rect 20076 9732 20128 9784
rect 22744 9732 22796 9784
rect 7564 9664 7616 9716
rect 17224 9664 17276 9716
rect 17316 9664 17368 9716
rect 24124 9664 24176 9716
rect 5816 9596 5868 9648
rect 14924 9596 14976 9648
rect 15016 9596 15068 9648
rect 19340 9596 19392 9648
rect 19524 9596 19576 9648
rect 28540 9664 28592 9716
rect 32312 9664 32364 9716
rect 4804 9188 4856 9240
rect 19984 9528 20036 9580
rect 7380 9460 7432 9512
rect 22376 9460 22428 9512
rect 17132 9392 17184 9444
rect 17224 9392 17276 9444
rect 24032 9392 24084 9444
rect 36820 9596 36872 9648
rect 27436 9460 27488 9512
rect 38660 9460 38712 9512
rect 34888 9392 34940 9444
rect 36084 9392 36136 9444
rect 26240 9324 26292 9376
rect 26332 9324 26384 9376
rect 33508 9324 33560 9376
rect 33784 9324 33836 9376
rect 13084 9256 13136 9308
rect 13176 9256 13228 9308
rect 16764 9256 16816 9308
rect 8852 9188 8904 9240
rect 9036 9188 9088 9240
rect 16948 9188 17000 9240
rect 17316 9256 17368 9308
rect 19340 9256 19392 9308
rect 19892 9256 19944 9308
rect 28908 9256 28960 9308
rect 35164 9256 35216 9308
rect 35348 9256 35400 9308
rect 41052 9256 41104 9308
rect 10508 9052 10560 9104
rect 18328 9120 18380 9172
rect 22928 9188 22980 9240
rect 27436 9188 27488 9240
rect 27896 9188 27948 9240
rect 17776 9052 17828 9104
rect 5448 8916 5500 8968
rect 13176 8984 13228 9036
rect 22192 8984 22244 9036
rect 23020 9052 23072 9104
rect 32772 9188 32824 9240
rect 34612 9120 34664 9172
rect 43628 9188 43680 9240
rect 34060 9052 34112 9104
rect 42892 9120 42944 9172
rect 20168 8916 20220 8968
rect 22928 8916 22980 8968
rect 27252 8916 27304 8968
rect 33416 8916 33468 8968
rect 33876 8916 33928 8968
rect 14188 8848 14240 8900
rect 16672 8848 16724 8900
rect 16764 8848 16816 8900
rect 20260 8848 20312 8900
rect 23664 8848 23716 8900
rect 31484 8848 31536 8900
rect 35624 8848 35676 8900
rect 39948 8848 40000 8900
rect 43260 8916 43312 8968
rect 3240 8780 3292 8832
rect 8484 8780 8536 8832
rect 11796 8780 11848 8832
rect 13544 8780 13596 8832
rect 17776 8780 17828 8832
rect 19064 8780 19116 8832
rect 22468 8780 22520 8832
rect 23756 8780 23808 8832
rect 32404 8780 32456 8832
rect 35992 8780 36044 8832
rect 40500 8780 40552 8832
rect 40684 8780 40736 8832
rect 12058 8678 12110 8730
rect 12122 8678 12174 8730
rect 12186 8678 12238 8730
rect 12250 8678 12302 8730
rect 12314 8678 12366 8730
rect 23166 8678 23218 8730
rect 23230 8678 23282 8730
rect 23294 8678 23346 8730
rect 23358 8678 23410 8730
rect 23422 8678 23474 8730
rect 34274 8678 34326 8730
rect 34338 8678 34390 8730
rect 34402 8678 34454 8730
rect 34466 8678 34518 8730
rect 34530 8678 34582 8730
rect 45382 8678 45434 8730
rect 45446 8678 45498 8730
rect 45510 8678 45562 8730
rect 45574 8678 45626 8730
rect 45638 8678 45690 8730
rect 2320 8576 2372 8628
rect 756 8508 808 8560
rect 4160 8576 4212 8628
rect 4896 8576 4948 8628
rect 5264 8576 5316 8628
rect 5448 8576 5500 8628
rect 5632 8576 5684 8628
rect 6000 8576 6052 8628
rect 6736 8576 6788 8628
rect 7012 8619 7064 8628
rect 7012 8585 7021 8619
rect 7021 8585 7055 8619
rect 7055 8585 7064 8619
rect 7012 8576 7064 8585
rect 7840 8576 7892 8628
rect 8116 8619 8168 8628
rect 8116 8585 8125 8619
rect 8125 8585 8159 8619
rect 8159 8585 8168 8619
rect 8116 8576 8168 8585
rect 8576 8576 8628 8628
rect 9312 8576 9364 8628
rect 9772 8619 9824 8628
rect 9772 8585 9781 8619
rect 9781 8585 9815 8619
rect 9815 8585 9824 8619
rect 9772 8576 9824 8585
rect 10416 8576 10468 8628
rect 10784 8576 10836 8628
rect 3240 8551 3292 8560
rect 3240 8517 3249 8551
rect 3249 8517 3283 8551
rect 3283 8517 3292 8551
rect 3240 8508 3292 8517
rect 5816 8551 5868 8560
rect 5816 8517 5825 8551
rect 5825 8517 5859 8551
rect 5859 8517 5868 8551
rect 5816 8508 5868 8517
rect 8852 8508 8904 8560
rect 4804 8483 4856 8492
rect 4804 8449 4813 8483
rect 4813 8449 4847 8483
rect 4847 8449 4856 8483
rect 4804 8440 4856 8449
rect 5356 8440 5408 8492
rect 7380 8440 7432 8492
rect 7564 8483 7616 8492
rect 7564 8449 7573 8483
rect 7573 8449 7607 8483
rect 7607 8449 7616 8483
rect 7564 8440 7616 8449
rect 8024 8483 8076 8492
rect 8024 8449 8033 8483
rect 8033 8449 8067 8483
rect 8067 8449 8076 8483
rect 8024 8440 8076 8449
rect 8484 8483 8536 8492
rect 8484 8449 8493 8483
rect 8493 8449 8527 8483
rect 8527 8449 8536 8483
rect 8484 8440 8536 8449
rect 8760 8440 8812 8492
rect 11244 8619 11296 8628
rect 11244 8585 11253 8619
rect 11253 8585 11287 8619
rect 11287 8585 11296 8619
rect 11244 8576 11296 8585
rect 11980 8619 12032 8628
rect 11980 8585 11989 8619
rect 11989 8585 12023 8619
rect 12023 8585 12032 8619
rect 11980 8576 12032 8585
rect 12532 8619 12584 8628
rect 12532 8585 12541 8619
rect 12541 8585 12575 8619
rect 12575 8585 12584 8619
rect 12532 8576 12584 8585
rect 13360 8576 13412 8628
rect 13636 8619 13688 8628
rect 13636 8585 13645 8619
rect 13645 8585 13679 8619
rect 13679 8585 13688 8619
rect 13636 8576 13688 8585
rect 14464 8576 14516 8628
rect 14832 8576 14884 8628
rect 15292 8619 15344 8628
rect 15292 8585 15301 8619
rect 15301 8585 15335 8619
rect 15335 8585 15344 8619
rect 15292 8576 15344 8585
rect 15568 8576 15620 8628
rect 15936 8576 15988 8628
rect 16304 8576 16356 8628
rect 16856 8619 16908 8628
rect 16856 8585 16865 8619
rect 16865 8585 16899 8619
rect 16899 8585 16908 8619
rect 16856 8576 16908 8585
rect 17408 8576 17460 8628
rect 18052 8619 18104 8628
rect 18052 8585 18061 8619
rect 18061 8585 18095 8619
rect 18095 8585 18104 8619
rect 18052 8576 18104 8585
rect 18144 8576 18196 8628
rect 18512 8576 18564 8628
rect 19156 8576 19208 8628
rect 20260 8576 20312 8628
rect 9036 8483 9088 8492
rect 9036 8449 9045 8483
rect 9045 8449 9079 8483
rect 9079 8449 9088 8483
rect 9036 8440 9088 8449
rect 9496 8483 9548 8492
rect 9496 8449 9505 8483
rect 9505 8449 9539 8483
rect 9539 8449 9548 8483
rect 9496 8440 9548 8449
rect 10416 8440 10468 8492
rect 10508 8483 10560 8492
rect 10508 8449 10517 8483
rect 10517 8449 10551 8483
rect 10551 8449 10560 8483
rect 10508 8440 10560 8449
rect 11796 8508 11848 8560
rect 12440 8551 12492 8560
rect 12440 8517 12449 8551
rect 12449 8517 12483 8551
rect 12483 8517 12492 8551
rect 12440 8508 12492 8517
rect 12624 8440 12676 8492
rect 13084 8483 13136 8492
rect 13084 8449 13093 8483
rect 13093 8449 13127 8483
rect 13127 8449 13136 8483
rect 13084 8440 13136 8449
rect 13544 8483 13596 8492
rect 13544 8449 13553 8483
rect 13553 8449 13587 8483
rect 13587 8449 13596 8483
rect 13544 8440 13596 8449
rect 14188 8483 14240 8492
rect 14188 8449 14197 8483
rect 14197 8449 14231 8483
rect 14231 8449 14240 8483
rect 14188 8440 14240 8449
rect 15016 8483 15068 8492
rect 15016 8449 15025 8483
rect 15025 8449 15059 8483
rect 15059 8449 15068 8483
rect 15016 8440 15068 8449
rect 15476 8483 15528 8492
rect 15476 8449 15485 8483
rect 15485 8449 15519 8483
rect 15519 8449 15528 8483
rect 15476 8440 15528 8449
rect 16120 8440 16172 8492
rect 14372 8372 14424 8424
rect 16764 8483 16816 8492
rect 16764 8449 16773 8483
rect 16773 8449 16807 8483
rect 16807 8449 16816 8483
rect 16764 8440 16816 8449
rect 17316 8483 17368 8492
rect 17316 8449 17325 8483
rect 17325 8449 17359 8483
rect 17359 8449 17368 8483
rect 17316 8440 17368 8449
rect 17500 8440 17552 8492
rect 18236 8483 18288 8492
rect 18236 8449 18245 8483
rect 18245 8449 18279 8483
rect 18279 8449 18288 8483
rect 18236 8440 18288 8449
rect 18880 8440 18932 8492
rect 19616 8483 19668 8492
rect 19616 8449 19625 8483
rect 19625 8449 19659 8483
rect 19659 8449 19668 8483
rect 19616 8440 19668 8449
rect 19156 8372 19208 8424
rect 19984 8508 20036 8560
rect 22928 8619 22980 8628
rect 22928 8585 22937 8619
rect 22937 8585 22971 8619
rect 22971 8585 22980 8619
rect 22928 8576 22980 8585
rect 23480 8576 23532 8628
rect 20536 8483 20588 8492
rect 20536 8449 20545 8483
rect 20545 8449 20579 8483
rect 20579 8449 20588 8483
rect 20536 8440 20588 8449
rect 20812 8483 20864 8492
rect 20812 8449 20821 8483
rect 20821 8449 20855 8483
rect 20855 8449 20864 8483
rect 20812 8440 20864 8449
rect 21088 8483 21140 8492
rect 21088 8449 21097 8483
rect 21097 8449 21131 8483
rect 21131 8449 21140 8483
rect 21088 8440 21140 8449
rect 21364 8483 21416 8492
rect 21364 8449 21373 8483
rect 21373 8449 21407 8483
rect 21407 8449 21416 8483
rect 21364 8440 21416 8449
rect 21640 8483 21692 8492
rect 21640 8449 21649 8483
rect 21649 8449 21683 8483
rect 21683 8449 21692 8483
rect 21640 8440 21692 8449
rect 22008 8483 22060 8492
rect 22008 8449 22017 8483
rect 22017 8449 22051 8483
rect 22051 8449 22060 8483
rect 22008 8440 22060 8449
rect 22100 8440 22152 8492
rect 22284 8483 22336 8492
rect 22284 8449 22293 8483
rect 22293 8449 22327 8483
rect 22327 8449 22336 8483
rect 22284 8440 22336 8449
rect 22376 8440 22428 8492
rect 22560 8483 22612 8492
rect 22560 8449 22569 8483
rect 22569 8449 22603 8483
rect 22603 8449 22612 8483
rect 22560 8440 22612 8449
rect 22836 8440 22888 8492
rect 23020 8372 23072 8424
rect 23572 8483 23624 8492
rect 23572 8449 23581 8483
rect 23581 8449 23615 8483
rect 23615 8449 23624 8483
rect 23572 8440 23624 8449
rect 23756 8483 23808 8492
rect 23756 8449 23765 8483
rect 23765 8449 23799 8483
rect 23799 8449 23808 8483
rect 23756 8440 23808 8449
rect 19432 8279 19484 8288
rect 19432 8245 19441 8279
rect 19441 8245 19475 8279
rect 19475 8245 19484 8279
rect 19432 8236 19484 8245
rect 20352 8279 20404 8288
rect 20352 8245 20361 8279
rect 20361 8245 20395 8279
rect 20395 8245 20404 8279
rect 20352 8236 20404 8245
rect 20536 8304 20588 8356
rect 21548 8304 21600 8356
rect 21916 8304 21968 8356
rect 22192 8304 22244 8356
rect 22284 8304 22336 8356
rect 22376 8347 22428 8356
rect 22376 8313 22385 8347
rect 22385 8313 22419 8347
rect 22419 8313 22428 8347
rect 22376 8304 22428 8313
rect 22836 8304 22888 8356
rect 23848 8304 23900 8356
rect 23940 8347 23992 8356
rect 23940 8313 23949 8347
rect 23949 8313 23983 8347
rect 23983 8313 23992 8347
rect 23940 8304 23992 8313
rect 24400 8508 24452 8560
rect 24308 8440 24360 8492
rect 24676 8483 24728 8492
rect 24676 8449 24685 8483
rect 24685 8449 24719 8483
rect 24719 8449 24728 8483
rect 24676 8440 24728 8449
rect 24860 8508 24912 8560
rect 26976 8508 27028 8560
rect 25504 8483 25556 8492
rect 25504 8449 25513 8483
rect 25513 8449 25547 8483
rect 25547 8449 25556 8483
rect 25504 8440 25556 8449
rect 25780 8483 25832 8492
rect 25780 8449 25789 8483
rect 25789 8449 25823 8483
rect 25823 8449 25832 8483
rect 25780 8440 25832 8449
rect 26148 8483 26200 8492
rect 26148 8449 26157 8483
rect 26157 8449 26191 8483
rect 26191 8449 26200 8483
rect 26148 8440 26200 8449
rect 26516 8483 26568 8492
rect 26516 8449 26525 8483
rect 26525 8449 26559 8483
rect 26559 8449 26568 8483
rect 26516 8440 26568 8449
rect 26608 8440 26660 8492
rect 29552 8508 29604 8560
rect 30288 8576 30340 8628
rect 27528 8440 27580 8492
rect 27988 8483 28040 8492
rect 27988 8449 27997 8483
rect 27997 8449 28031 8483
rect 28031 8449 28040 8483
rect 27988 8440 28040 8449
rect 28356 8483 28408 8492
rect 28356 8449 28365 8483
rect 28365 8449 28399 8483
rect 28399 8449 28408 8483
rect 28356 8440 28408 8449
rect 28724 8483 28776 8492
rect 28724 8449 28733 8483
rect 28733 8449 28767 8483
rect 28767 8449 28776 8483
rect 28724 8440 28776 8449
rect 28816 8440 28868 8492
rect 29184 8440 29236 8492
rect 30288 8483 30340 8492
rect 30288 8449 30297 8483
rect 30297 8449 30331 8483
rect 30331 8449 30340 8483
rect 30288 8440 30340 8449
rect 24492 8372 24544 8424
rect 30380 8372 30432 8424
rect 31484 8619 31536 8628
rect 31484 8585 31493 8619
rect 31493 8585 31527 8619
rect 31527 8585 31536 8619
rect 31484 8576 31536 8585
rect 32312 8619 32364 8628
rect 32312 8585 32321 8619
rect 32321 8585 32355 8619
rect 32355 8585 32364 8619
rect 32312 8576 32364 8585
rect 32404 8619 32456 8628
rect 32404 8585 32413 8619
rect 32413 8585 32447 8619
rect 32447 8585 32456 8619
rect 32404 8576 32456 8585
rect 32496 8576 32548 8628
rect 33508 8619 33560 8628
rect 33508 8585 33517 8619
rect 33517 8585 33551 8619
rect 33551 8585 33560 8619
rect 33508 8576 33560 8585
rect 30656 8508 30708 8560
rect 34060 8576 34112 8628
rect 34612 8576 34664 8628
rect 34796 8576 34848 8628
rect 35716 8619 35768 8628
rect 35716 8585 35725 8619
rect 35725 8585 35759 8619
rect 35759 8585 35768 8619
rect 35716 8576 35768 8585
rect 35900 8576 35952 8628
rect 38660 8619 38712 8628
rect 38660 8585 38669 8619
rect 38669 8585 38703 8619
rect 38703 8585 38712 8619
rect 38660 8576 38712 8585
rect 39028 8619 39080 8628
rect 39028 8585 39037 8619
rect 39037 8585 39071 8619
rect 39071 8585 39080 8619
rect 39028 8576 39080 8585
rect 39120 8576 39172 8628
rect 39764 8576 39816 8628
rect 30932 8483 30984 8492
rect 30932 8449 30941 8483
rect 30941 8449 30975 8483
rect 30975 8449 30984 8483
rect 30932 8440 30984 8449
rect 31300 8483 31352 8492
rect 31300 8449 31309 8483
rect 31309 8449 31343 8483
rect 31343 8449 31352 8483
rect 31300 8440 31352 8449
rect 31668 8483 31720 8492
rect 31668 8449 31677 8483
rect 31677 8449 31711 8483
rect 31711 8449 31720 8483
rect 31668 8440 31720 8449
rect 31760 8440 31812 8492
rect 32312 8440 32364 8492
rect 32680 8483 32732 8492
rect 32680 8449 32689 8483
rect 32689 8449 32723 8483
rect 32723 8449 32732 8483
rect 32680 8440 32732 8449
rect 33324 8483 33376 8492
rect 33324 8449 33333 8483
rect 33333 8449 33367 8483
rect 33367 8449 33376 8483
rect 33324 8440 33376 8449
rect 33692 8483 33744 8492
rect 33692 8449 33701 8483
rect 33701 8449 33735 8483
rect 33735 8449 33744 8483
rect 33692 8440 33744 8449
rect 34060 8483 34112 8492
rect 34060 8449 34069 8483
rect 34069 8449 34103 8483
rect 34103 8449 34112 8483
rect 34060 8440 34112 8449
rect 34152 8440 34204 8492
rect 34980 8483 35032 8492
rect 34980 8449 34989 8483
rect 34989 8449 35023 8483
rect 35023 8449 35032 8483
rect 34980 8440 35032 8449
rect 35256 8483 35308 8492
rect 35256 8449 35265 8483
rect 35265 8449 35299 8483
rect 35299 8449 35308 8483
rect 35256 8440 35308 8449
rect 35532 8483 35584 8492
rect 35532 8449 35541 8483
rect 35541 8449 35575 8483
rect 35575 8449 35584 8483
rect 35532 8440 35584 8449
rect 35808 8440 35860 8492
rect 36268 8483 36320 8492
rect 36268 8449 36277 8483
rect 36277 8449 36311 8483
rect 36311 8449 36320 8483
rect 36268 8440 36320 8449
rect 25872 8304 25924 8356
rect 21180 8279 21232 8288
rect 21180 8245 21189 8279
rect 21189 8245 21223 8279
rect 21223 8245 21232 8279
rect 21180 8236 21232 8245
rect 21456 8279 21508 8288
rect 21456 8245 21465 8279
rect 21465 8245 21499 8279
rect 21499 8245 21508 8279
rect 21456 8236 21508 8245
rect 21824 8279 21876 8288
rect 21824 8245 21833 8279
rect 21833 8245 21867 8279
rect 21867 8245 21876 8279
rect 21824 8236 21876 8245
rect 23388 8236 23440 8288
rect 23480 8236 23532 8288
rect 24308 8236 24360 8288
rect 24492 8279 24544 8288
rect 24492 8245 24501 8279
rect 24501 8245 24535 8279
rect 24535 8245 24544 8279
rect 24492 8236 24544 8245
rect 24768 8279 24820 8288
rect 24768 8245 24777 8279
rect 24777 8245 24811 8279
rect 24811 8245 24820 8279
rect 24768 8236 24820 8245
rect 25044 8279 25096 8288
rect 25044 8245 25053 8279
rect 25053 8245 25087 8279
rect 25087 8245 25096 8279
rect 25044 8236 25096 8245
rect 25136 8236 25188 8288
rect 25412 8236 25464 8288
rect 25688 8236 25740 8288
rect 26148 8236 26200 8288
rect 27620 8304 27672 8356
rect 28264 8304 28316 8356
rect 32496 8304 32548 8356
rect 26608 8236 26660 8288
rect 27528 8279 27580 8288
rect 27528 8245 27537 8279
rect 27537 8245 27571 8279
rect 27571 8245 27580 8279
rect 27528 8236 27580 8245
rect 27804 8279 27856 8288
rect 27804 8245 27813 8279
rect 27813 8245 27847 8279
rect 27847 8245 27856 8279
rect 27804 8236 27856 8245
rect 28540 8279 28592 8288
rect 28540 8245 28549 8279
rect 28549 8245 28583 8279
rect 28583 8245 28592 8279
rect 28540 8236 28592 8245
rect 28632 8236 28684 8288
rect 29552 8279 29604 8288
rect 29552 8245 29561 8279
rect 29561 8245 29595 8279
rect 29595 8245 29604 8279
rect 29552 8236 29604 8245
rect 29828 8279 29880 8288
rect 29828 8245 29837 8279
rect 29837 8245 29871 8279
rect 29871 8245 29880 8279
rect 29828 8236 29880 8245
rect 30104 8279 30156 8288
rect 30104 8245 30113 8279
rect 30113 8245 30147 8279
rect 30147 8245 30156 8279
rect 30104 8236 30156 8245
rect 30380 8279 30432 8288
rect 30380 8245 30389 8279
rect 30389 8245 30423 8279
rect 30423 8245 30432 8279
rect 30380 8236 30432 8245
rect 30748 8279 30800 8288
rect 30748 8245 30757 8279
rect 30757 8245 30791 8279
rect 30791 8245 30800 8279
rect 30748 8236 30800 8245
rect 31116 8279 31168 8288
rect 31116 8245 31125 8279
rect 31125 8245 31159 8279
rect 31159 8245 31168 8279
rect 31116 8236 31168 8245
rect 33048 8372 33100 8424
rect 33048 8236 33100 8288
rect 33416 8304 33468 8356
rect 34888 8347 34940 8356
rect 34888 8313 34897 8347
rect 34897 8313 34931 8347
rect 34931 8313 34940 8347
rect 34888 8304 34940 8313
rect 35164 8347 35216 8356
rect 35164 8313 35173 8347
rect 35173 8313 35207 8347
rect 35207 8313 35216 8347
rect 35164 8304 35216 8313
rect 39856 8508 39908 8560
rect 40960 8576 41012 8628
rect 41328 8508 41380 8560
rect 42708 8576 42760 8628
rect 42892 8508 42944 8560
rect 43260 8508 43312 8560
rect 36636 8483 36688 8492
rect 36636 8449 36645 8483
rect 36645 8449 36679 8483
rect 36679 8449 36688 8483
rect 36636 8440 36688 8449
rect 36820 8440 36872 8492
rect 36912 8440 36964 8492
rect 37556 8483 37608 8492
rect 37556 8449 37565 8483
rect 37565 8449 37599 8483
rect 37599 8449 37608 8483
rect 37556 8440 37608 8449
rect 37832 8483 37884 8492
rect 37832 8449 37841 8483
rect 37841 8449 37875 8483
rect 37875 8449 37884 8483
rect 37832 8440 37884 8449
rect 38108 8483 38160 8492
rect 38108 8449 38117 8483
rect 38117 8449 38151 8483
rect 38151 8449 38160 8483
rect 38108 8440 38160 8449
rect 38476 8483 38528 8492
rect 38476 8449 38485 8483
rect 38485 8449 38519 8483
rect 38519 8449 38528 8483
rect 38476 8440 38528 8449
rect 38568 8440 38620 8492
rect 37464 8347 37516 8356
rect 37464 8313 37473 8347
rect 37473 8313 37507 8347
rect 37507 8313 37516 8347
rect 37464 8304 37516 8313
rect 37740 8347 37792 8356
rect 37740 8313 37749 8347
rect 37749 8313 37783 8347
rect 37783 8313 37792 8347
rect 37740 8304 37792 8313
rect 39948 8483 40000 8492
rect 39948 8449 39957 8483
rect 39957 8449 39991 8483
rect 39991 8449 40000 8483
rect 39948 8440 40000 8449
rect 40224 8440 40276 8492
rect 40500 8483 40552 8492
rect 40500 8449 40509 8483
rect 40509 8449 40543 8483
rect 40543 8449 40552 8483
rect 40500 8440 40552 8449
rect 40684 8440 40736 8492
rect 41052 8440 41104 8492
rect 42524 8483 42576 8492
rect 42524 8449 42533 8483
rect 42533 8449 42567 8483
rect 42567 8449 42576 8483
rect 42524 8440 42576 8449
rect 43628 8483 43680 8492
rect 43628 8449 43637 8483
rect 43637 8449 43671 8483
rect 43671 8449 43680 8483
rect 43628 8440 43680 8449
rect 42064 8372 42116 8424
rect 37188 8236 37240 8288
rect 41696 8304 41748 8356
rect 6504 8134 6556 8186
rect 6568 8134 6620 8186
rect 6632 8134 6684 8186
rect 6696 8134 6748 8186
rect 6760 8134 6812 8186
rect 17612 8134 17664 8186
rect 17676 8134 17728 8186
rect 17740 8134 17792 8186
rect 17804 8134 17856 8186
rect 17868 8134 17920 8186
rect 28720 8134 28772 8186
rect 28784 8134 28836 8186
rect 28848 8134 28900 8186
rect 28912 8134 28964 8186
rect 28976 8134 29028 8186
rect 39828 8134 39880 8186
rect 39892 8134 39944 8186
rect 39956 8134 40008 8186
rect 40020 8134 40072 8186
rect 40084 8134 40136 8186
rect 2044 8075 2096 8084
rect 2044 8041 2053 8075
rect 2053 8041 2087 8075
rect 2087 8041 2096 8075
rect 2044 8032 2096 8041
rect 2780 8075 2832 8084
rect 2780 8041 2789 8075
rect 2789 8041 2823 8075
rect 2823 8041 2832 8075
rect 2780 8032 2832 8041
rect 3056 8032 3108 8084
rect 3424 8032 3476 8084
rect 4160 8075 4212 8084
rect 4160 8041 4169 8075
rect 4169 8041 4203 8075
rect 4203 8041 4212 8075
rect 4160 8032 4212 8041
rect 4528 8032 4580 8084
rect 6368 8032 6420 8084
rect 7472 8032 7524 8084
rect 9128 8075 9180 8084
rect 9128 8041 9137 8075
rect 9137 8041 9171 8075
rect 9171 8041 9180 8075
rect 9128 8032 9180 8041
rect 10048 8032 10100 8084
rect 11612 8075 11664 8084
rect 11612 8041 11621 8075
rect 11621 8041 11655 8075
rect 11655 8041 11664 8075
rect 11612 8032 11664 8041
rect 11888 8032 11940 8084
rect 12992 8032 13044 8084
rect 14280 8075 14332 8084
rect 14280 8041 14289 8075
rect 14289 8041 14323 8075
rect 14323 8041 14332 8075
rect 14280 8032 14332 8041
rect 17040 8032 17092 8084
rect 17500 8032 17552 8084
rect 18236 8032 18288 8084
rect 19248 8032 19300 8084
rect 20444 8075 20496 8084
rect 20444 8041 20453 8075
rect 20453 8041 20487 8075
rect 20487 8041 20496 8075
rect 20444 8032 20496 8041
rect 20904 8075 20956 8084
rect 20904 8041 20913 8075
rect 20913 8041 20947 8075
rect 20947 8041 20956 8075
rect 20904 8032 20956 8041
rect 21180 8032 21232 8084
rect 21548 8075 21600 8084
rect 21548 8041 21557 8075
rect 21557 8041 21591 8075
rect 21591 8041 21600 8075
rect 21548 8032 21600 8041
rect 21824 8032 21876 8084
rect 22192 8032 22244 8084
rect 24308 8032 24360 8084
rect 10416 7964 10468 8016
rect 17224 7964 17276 8016
rect 19340 7964 19392 8016
rect 19432 7964 19484 8016
rect 2964 7871 3016 7880
rect 2964 7837 2973 7871
rect 2973 7837 3007 7871
rect 3007 7837 3016 7871
rect 2964 7828 3016 7837
rect 3332 7871 3384 7880
rect 3332 7837 3341 7871
rect 3341 7837 3375 7871
rect 3375 7837 3384 7871
rect 3332 7828 3384 7837
rect 4436 7871 4488 7880
rect 4436 7837 4445 7871
rect 4445 7837 4479 7871
rect 4479 7837 4488 7871
rect 4436 7828 4488 7837
rect 2504 7803 2556 7812
rect 2504 7769 2513 7803
rect 2513 7769 2547 7803
rect 2547 7769 2556 7803
rect 2504 7760 2556 7769
rect 3884 7803 3936 7812
rect 3884 7769 3893 7803
rect 3893 7769 3927 7803
rect 3927 7769 3936 7803
rect 3884 7760 3936 7769
rect 6368 7803 6420 7812
rect 6368 7769 6377 7803
rect 6377 7769 6411 7803
rect 6411 7769 6420 7803
rect 6368 7760 6420 7769
rect 9956 7871 10008 7880
rect 9956 7837 9965 7871
rect 9965 7837 9999 7871
rect 9999 7837 10008 7871
rect 9956 7828 10008 7837
rect 11520 7871 11572 7880
rect 11520 7837 11529 7871
rect 11529 7837 11563 7871
rect 11563 7837 11572 7871
rect 11520 7828 11572 7837
rect 12900 7871 12952 7880
rect 12900 7837 12909 7871
rect 12909 7837 12943 7871
rect 12943 7837 12952 7871
rect 12900 7828 12952 7837
rect 5448 7692 5500 7744
rect 14188 7803 14240 7812
rect 14188 7769 14197 7803
rect 14197 7769 14231 7803
rect 14231 7769 14240 7803
rect 14188 7760 14240 7769
rect 15108 7760 15160 7812
rect 18052 7896 18104 7948
rect 17132 7871 17184 7880
rect 17132 7837 17141 7871
rect 17141 7837 17175 7871
rect 17175 7837 17184 7871
rect 17132 7828 17184 7837
rect 17224 7828 17276 7880
rect 17316 7828 17368 7880
rect 17868 7828 17920 7880
rect 18236 7871 18288 7880
rect 18236 7837 18245 7871
rect 18245 7837 18279 7871
rect 18279 7837 18288 7871
rect 18236 7828 18288 7837
rect 18788 7871 18840 7880
rect 18788 7837 18797 7871
rect 18797 7837 18831 7871
rect 18831 7837 18840 7871
rect 18788 7828 18840 7837
rect 20352 7964 20404 8016
rect 20260 7896 20312 7948
rect 22100 7964 22152 8016
rect 24584 8075 24636 8084
rect 24584 8041 24593 8075
rect 24593 8041 24627 8075
rect 24627 8041 24636 8075
rect 24584 8032 24636 8041
rect 25044 8032 25096 8084
rect 25228 8032 25280 8084
rect 27528 8032 27580 8084
rect 27712 8032 27764 8084
rect 27804 8032 27856 8084
rect 27896 8075 27948 8084
rect 27896 8041 27905 8075
rect 27905 8041 27939 8075
rect 27939 8041 27948 8075
rect 27896 8032 27948 8041
rect 28540 8032 28592 8084
rect 28632 8032 28684 8084
rect 40592 8032 40644 8084
rect 42800 8032 42852 8084
rect 43536 8032 43588 8084
rect 43904 8032 43956 8084
rect 20536 7828 20588 7880
rect 20628 7871 20680 7880
rect 20628 7837 20637 7871
rect 20637 7837 20671 7871
rect 20671 7837 20680 7871
rect 20628 7828 20680 7837
rect 17224 7692 17276 7744
rect 18420 7760 18472 7812
rect 18512 7735 18564 7744
rect 18512 7701 18521 7735
rect 18521 7701 18555 7735
rect 18555 7701 18564 7735
rect 18512 7692 18564 7701
rect 21456 7828 21508 7880
rect 21732 7871 21784 7880
rect 21732 7837 21741 7871
rect 21741 7837 21775 7871
rect 21775 7837 21784 7871
rect 21732 7828 21784 7837
rect 22008 7871 22060 7880
rect 22008 7837 22017 7871
rect 22017 7837 22051 7871
rect 22051 7837 22060 7871
rect 22008 7828 22060 7837
rect 18696 7692 18748 7744
rect 19340 7692 19392 7744
rect 20076 7735 20128 7744
rect 20076 7701 20085 7735
rect 20085 7701 20119 7735
rect 20119 7701 20128 7735
rect 20076 7692 20128 7701
rect 21640 7760 21692 7812
rect 21364 7692 21416 7744
rect 21456 7735 21508 7744
rect 21456 7701 21465 7735
rect 21465 7701 21499 7735
rect 21499 7701 21508 7735
rect 21456 7692 21508 7701
rect 21824 7735 21876 7744
rect 21824 7701 21833 7735
rect 21833 7701 21867 7735
rect 21867 7701 21876 7735
rect 21824 7692 21876 7701
rect 22008 7692 22060 7744
rect 22468 7896 22520 7948
rect 26240 7964 26292 8016
rect 22744 7828 22796 7880
rect 23204 7871 23256 7880
rect 23204 7837 23213 7871
rect 23213 7837 23247 7871
rect 23247 7837 23256 7871
rect 23204 7828 23256 7837
rect 23664 7828 23716 7880
rect 23940 7828 23992 7880
rect 22560 7692 22612 7744
rect 22652 7735 22704 7744
rect 22652 7701 22661 7735
rect 22661 7701 22695 7735
rect 22695 7701 22704 7735
rect 22652 7692 22704 7701
rect 22836 7692 22888 7744
rect 23388 7735 23440 7744
rect 23388 7701 23397 7735
rect 23397 7701 23431 7735
rect 23431 7701 23440 7735
rect 23388 7692 23440 7701
rect 24216 7735 24268 7744
rect 24216 7701 24225 7735
rect 24225 7701 24259 7735
rect 24259 7701 24268 7735
rect 24216 7692 24268 7701
rect 24308 7692 24360 7744
rect 25136 7828 25188 7880
rect 25412 7828 25464 7880
rect 25688 7828 25740 7880
rect 25872 7828 25924 7880
rect 26148 7828 26200 7880
rect 26608 7828 26660 7880
rect 27620 7828 27672 7880
rect 44272 7964 44324 8016
rect 29552 7828 29604 7880
rect 29828 7828 29880 7880
rect 33048 7828 33100 7880
rect 25044 7692 25096 7744
rect 25136 7735 25188 7744
rect 25136 7701 25145 7735
rect 25145 7701 25179 7735
rect 25179 7701 25188 7735
rect 25136 7692 25188 7701
rect 25412 7735 25464 7744
rect 25412 7701 25421 7735
rect 25421 7701 25455 7735
rect 25455 7701 25464 7735
rect 25412 7692 25464 7701
rect 25688 7735 25740 7744
rect 25688 7701 25697 7735
rect 25697 7701 25731 7735
rect 25731 7701 25740 7735
rect 25688 7692 25740 7701
rect 25964 7735 26016 7744
rect 25964 7701 25973 7735
rect 25973 7701 26007 7735
rect 26007 7701 26016 7735
rect 25964 7692 26016 7701
rect 26240 7735 26292 7744
rect 26240 7701 26249 7735
rect 26249 7701 26283 7735
rect 26283 7701 26292 7735
rect 26240 7692 26292 7701
rect 26884 7735 26936 7744
rect 26884 7701 26893 7735
rect 26893 7701 26927 7735
rect 26927 7701 26936 7735
rect 26884 7692 26936 7701
rect 39672 7760 39724 7812
rect 42800 7760 42852 7812
rect 43444 7760 43496 7812
rect 44272 7803 44324 7812
rect 44272 7769 44281 7803
rect 44281 7769 44315 7803
rect 44315 7769 44324 7803
rect 44272 7760 44324 7769
rect 27344 7692 27396 7744
rect 28172 7735 28224 7744
rect 28172 7701 28181 7735
rect 28181 7701 28215 7735
rect 28215 7701 28224 7735
rect 28172 7692 28224 7701
rect 28448 7735 28500 7744
rect 28448 7701 28457 7735
rect 28457 7701 28491 7735
rect 28491 7701 28500 7735
rect 28448 7692 28500 7701
rect 28540 7692 28592 7744
rect 12058 7590 12110 7642
rect 12122 7590 12174 7642
rect 12186 7590 12238 7642
rect 12250 7590 12302 7642
rect 12314 7590 12366 7642
rect 23166 7590 23218 7642
rect 23230 7590 23282 7642
rect 23294 7590 23346 7642
rect 23358 7590 23410 7642
rect 23422 7590 23474 7642
rect 34274 7590 34326 7642
rect 34338 7590 34390 7642
rect 34402 7590 34454 7642
rect 34466 7590 34518 7642
rect 34530 7590 34582 7642
rect 45382 7590 45434 7642
rect 45446 7590 45498 7642
rect 45510 7590 45562 7642
rect 45574 7590 45626 7642
rect 45638 7590 45690 7642
rect 848 7488 900 7540
rect 1584 7420 1636 7472
rect 3884 7488 3936 7540
rect 11060 7488 11112 7540
rect 15108 7488 15160 7540
rect 17132 7488 17184 7540
rect 18696 7488 18748 7540
rect 18788 7531 18840 7540
rect 18788 7497 18797 7531
rect 18797 7497 18831 7531
rect 18831 7497 18840 7531
rect 18788 7488 18840 7497
rect 18880 7531 18932 7540
rect 18880 7497 18889 7531
rect 18889 7497 18923 7531
rect 18923 7497 18932 7531
rect 18880 7488 18932 7497
rect 19156 7488 19208 7540
rect 19892 7488 19944 7540
rect 21824 7488 21876 7540
rect 22192 7488 22244 7540
rect 12900 7352 12952 7404
rect 18144 7352 18196 7404
rect 20812 7420 20864 7472
rect 22376 7420 22428 7472
rect 19064 7395 19116 7404
rect 19064 7361 19073 7395
rect 19073 7361 19107 7395
rect 19107 7361 19116 7395
rect 19064 7352 19116 7361
rect 19432 7395 19484 7404
rect 19432 7361 19441 7395
rect 19441 7361 19475 7395
rect 19475 7361 19484 7395
rect 19432 7352 19484 7361
rect 19616 7352 19668 7404
rect 21088 7352 21140 7404
rect 21824 7352 21876 7404
rect 21916 7395 21968 7404
rect 21916 7361 21925 7395
rect 21925 7361 21959 7395
rect 21959 7361 21968 7395
rect 21916 7352 21968 7361
rect 4436 7284 4488 7336
rect 6368 7284 6420 7336
rect 11060 7284 11112 7336
rect 12348 7284 12400 7336
rect 21456 7216 21508 7268
rect 21640 7284 21692 7336
rect 22652 7488 22704 7540
rect 22928 7488 22980 7540
rect 23112 7488 23164 7540
rect 24216 7488 24268 7540
rect 24492 7488 24544 7540
rect 27344 7488 27396 7540
rect 30104 7488 30156 7540
rect 30380 7488 30432 7540
rect 30748 7488 30800 7540
rect 43168 7488 43220 7540
rect 45008 7488 45060 7540
rect 45744 7488 45796 7540
rect 22744 7352 22796 7404
rect 22928 7395 22980 7404
rect 22928 7361 22937 7395
rect 22937 7361 22971 7395
rect 22971 7361 22980 7395
rect 22928 7352 22980 7361
rect 23020 7395 23072 7404
rect 23020 7361 23029 7395
rect 23029 7361 23063 7395
rect 23063 7361 23072 7395
rect 23020 7352 23072 7361
rect 23388 7395 23440 7404
rect 23388 7361 23397 7395
rect 23397 7361 23431 7395
rect 23431 7361 23440 7395
rect 23388 7352 23440 7361
rect 25044 7420 25096 7472
rect 31116 7284 31168 7336
rect 26884 7216 26936 7268
rect 14556 7148 14608 7200
rect 15476 7148 15528 7200
rect 21916 7148 21968 7200
rect 22008 7148 22060 7200
rect 22744 7191 22796 7200
rect 22744 7157 22753 7191
rect 22753 7157 22787 7191
rect 22787 7157 22796 7191
rect 22744 7148 22796 7157
rect 23204 7191 23256 7200
rect 23204 7157 23213 7191
rect 23213 7157 23247 7191
rect 23247 7157 23256 7191
rect 23204 7148 23256 7157
rect 23848 7148 23900 7200
rect 24124 7148 24176 7200
rect 24216 7191 24268 7200
rect 24216 7157 24225 7191
rect 24225 7157 24259 7191
rect 24259 7157 24268 7191
rect 24216 7148 24268 7157
rect 24308 7148 24360 7200
rect 43352 7395 43404 7404
rect 43352 7361 43361 7395
rect 43361 7361 43395 7395
rect 43395 7361 43404 7395
rect 43352 7352 43404 7361
rect 44180 7352 44232 7404
rect 45008 7284 45060 7336
rect 37740 7148 37792 7200
rect 6504 7046 6556 7098
rect 6568 7046 6620 7098
rect 6632 7046 6684 7098
rect 6696 7046 6748 7098
rect 6760 7046 6812 7098
rect 17612 7046 17664 7098
rect 17676 7046 17728 7098
rect 17740 7046 17792 7098
rect 17804 7046 17856 7098
rect 17868 7046 17920 7098
rect 28720 7046 28772 7098
rect 28784 7046 28836 7098
rect 28848 7046 28900 7098
rect 28912 7046 28964 7098
rect 28976 7046 29028 7098
rect 39828 7046 39880 7098
rect 39892 7046 39944 7098
rect 39956 7046 40008 7098
rect 40020 7046 40072 7098
rect 40084 7046 40136 7098
rect 9956 6944 10008 6996
rect 14188 6944 14240 6996
rect 22744 6944 22796 6996
rect 17960 6876 18012 6928
rect 1216 6808 1268 6860
rect 16672 6808 16724 6860
rect 21640 6876 21692 6928
rect 22468 6876 22520 6928
rect 27252 6876 27304 6928
rect 19432 6808 19484 6860
rect 26332 6808 26384 6860
rect 45284 6808 45336 6860
rect 46112 6808 46164 6860
rect 14648 6740 14700 6792
rect 20076 6740 20128 6792
rect 20168 6740 20220 6792
rect 24216 6740 24268 6792
rect 1492 6715 1544 6724
rect 1492 6681 1501 6715
rect 1501 6681 1535 6715
rect 1535 6681 1544 6715
rect 1492 6672 1544 6681
rect 12348 6672 12400 6724
rect 3332 6604 3384 6656
rect 17224 6604 17276 6656
rect 43904 6715 43956 6724
rect 43904 6681 43913 6715
rect 43913 6681 43947 6715
rect 43947 6681 43956 6715
rect 43904 6672 43956 6681
rect 44456 6715 44508 6724
rect 44456 6681 44465 6715
rect 44465 6681 44499 6715
rect 44499 6681 44508 6715
rect 44456 6672 44508 6681
rect 23112 6604 23164 6656
rect 12058 6502 12110 6554
rect 12122 6502 12174 6554
rect 12186 6502 12238 6554
rect 12250 6502 12302 6554
rect 12314 6502 12366 6554
rect 23166 6502 23218 6554
rect 23230 6502 23282 6554
rect 23294 6502 23346 6554
rect 23358 6502 23410 6554
rect 23422 6502 23474 6554
rect 34274 6502 34326 6554
rect 34338 6502 34390 6554
rect 34402 6502 34454 6554
rect 34466 6502 34518 6554
rect 34530 6502 34582 6554
rect 45382 6502 45434 6554
rect 45446 6502 45498 6554
rect 45510 6502 45562 6554
rect 45574 6502 45626 6554
rect 45638 6502 45690 6554
rect 1492 6400 1544 6452
rect 2504 6332 2556 6384
rect 14464 6400 14516 6452
rect 14556 6400 14608 6452
rect 17224 6400 17276 6452
rect 25136 6400 25188 6452
rect 44640 6400 44692 6452
rect 22836 6332 22888 6384
rect 24860 6332 24912 6384
rect 32772 6332 32824 6384
rect 18512 6264 18564 6316
rect 24216 6264 24268 6316
rect 35992 6264 36044 6316
rect 44824 6307 44876 6316
rect 44824 6273 44833 6307
rect 44833 6273 44867 6307
rect 44867 6273 44876 6307
rect 44824 6264 44876 6273
rect 2964 6196 3016 6248
rect 14464 6196 14516 6248
rect 25688 6196 25740 6248
rect 27068 6196 27120 6248
rect 42800 6196 42852 6248
rect 25412 6128 25464 6180
rect 25504 6128 25556 6180
rect 42524 6128 42576 6180
rect 6504 5958 6556 6010
rect 6568 5958 6620 6010
rect 6632 5958 6684 6010
rect 6696 5958 6748 6010
rect 6760 5958 6812 6010
rect 17612 5958 17664 6010
rect 17676 5958 17728 6010
rect 17740 5958 17792 6010
rect 17804 5958 17856 6010
rect 17868 5958 17920 6010
rect 28720 5958 28772 6010
rect 28784 5958 28836 6010
rect 28848 5958 28900 6010
rect 28912 5958 28964 6010
rect 28976 5958 29028 6010
rect 39828 5958 39880 6010
rect 39892 5958 39944 6010
rect 39956 5958 40008 6010
rect 40020 5958 40072 6010
rect 40084 5958 40136 6010
rect 12058 5414 12110 5466
rect 12122 5414 12174 5466
rect 12186 5414 12238 5466
rect 12250 5414 12302 5466
rect 12314 5414 12366 5466
rect 23166 5414 23218 5466
rect 23230 5414 23282 5466
rect 23294 5414 23346 5466
rect 23358 5414 23410 5466
rect 23422 5414 23474 5466
rect 34274 5414 34326 5466
rect 34338 5414 34390 5466
rect 34402 5414 34454 5466
rect 34466 5414 34518 5466
rect 34530 5414 34582 5466
rect 45382 5414 45434 5466
rect 45446 5414 45498 5466
rect 45510 5414 45562 5466
rect 45574 5414 45626 5466
rect 45638 5414 45690 5466
rect 23020 5108 23072 5160
rect 33048 5108 33100 5160
rect 22836 5040 22888 5092
rect 35624 5040 35676 5092
rect 20536 4972 20588 5024
rect 33784 4972 33836 5024
rect 6504 4870 6556 4922
rect 6568 4870 6620 4922
rect 6632 4870 6684 4922
rect 6696 4870 6748 4922
rect 6760 4870 6812 4922
rect 17612 4870 17664 4922
rect 17676 4870 17728 4922
rect 17740 4870 17792 4922
rect 17804 4870 17856 4922
rect 17868 4870 17920 4922
rect 28720 4870 28772 4922
rect 28784 4870 28836 4922
rect 28848 4870 28900 4922
rect 28912 4870 28964 4922
rect 28976 4870 29028 4922
rect 39828 4870 39880 4922
rect 39892 4870 39944 4922
rect 39956 4870 40008 4922
rect 40020 4870 40072 4922
rect 40084 4870 40136 4922
rect 29276 4768 29328 4820
rect 43352 4768 43404 4820
rect 12058 4326 12110 4378
rect 12122 4326 12174 4378
rect 12186 4326 12238 4378
rect 12250 4326 12302 4378
rect 12314 4326 12366 4378
rect 23166 4326 23218 4378
rect 23230 4326 23282 4378
rect 23294 4326 23346 4378
rect 23358 4326 23410 4378
rect 23422 4326 23474 4378
rect 34274 4326 34326 4378
rect 34338 4326 34390 4378
rect 34402 4326 34454 4378
rect 34466 4326 34518 4378
rect 34530 4326 34582 4378
rect 45382 4326 45434 4378
rect 45446 4326 45498 4378
rect 45510 4326 45562 4378
rect 45574 4326 45626 4378
rect 45638 4326 45690 4378
rect 6504 3782 6556 3834
rect 6568 3782 6620 3834
rect 6632 3782 6684 3834
rect 6696 3782 6748 3834
rect 6760 3782 6812 3834
rect 17612 3782 17664 3834
rect 17676 3782 17728 3834
rect 17740 3782 17792 3834
rect 17804 3782 17856 3834
rect 17868 3782 17920 3834
rect 28720 3782 28772 3834
rect 28784 3782 28836 3834
rect 28848 3782 28900 3834
rect 28912 3782 28964 3834
rect 28976 3782 29028 3834
rect 39828 3782 39880 3834
rect 39892 3782 39944 3834
rect 39956 3782 40008 3834
rect 40020 3782 40072 3834
rect 40084 3782 40136 3834
rect 23664 3612 23716 3664
rect 33876 3612 33928 3664
rect 22744 3544 22796 3596
rect 35348 3544 35400 3596
rect 23940 3476 23992 3528
rect 37188 3476 37240 3528
rect 20628 3408 20680 3460
rect 38568 3408 38620 3460
rect 12058 3238 12110 3290
rect 12122 3238 12174 3290
rect 12186 3238 12238 3290
rect 12250 3238 12302 3290
rect 12314 3238 12366 3290
rect 23166 3238 23218 3290
rect 23230 3238 23282 3290
rect 23294 3238 23346 3290
rect 23358 3238 23410 3290
rect 23422 3238 23474 3290
rect 34274 3238 34326 3290
rect 34338 3238 34390 3290
rect 34402 3238 34454 3290
rect 34466 3238 34518 3290
rect 34530 3238 34582 3290
rect 45382 3238 45434 3290
rect 45446 3238 45498 3290
rect 45510 3238 45562 3290
rect 45574 3238 45626 3290
rect 45638 3238 45690 3290
rect 6504 2694 6556 2746
rect 6568 2694 6620 2746
rect 6632 2694 6684 2746
rect 6696 2694 6748 2746
rect 6760 2694 6812 2746
rect 17612 2694 17664 2746
rect 17676 2694 17728 2746
rect 17740 2694 17792 2746
rect 17804 2694 17856 2746
rect 17868 2694 17920 2746
rect 28720 2694 28772 2746
rect 28784 2694 28836 2746
rect 28848 2694 28900 2746
rect 28912 2694 28964 2746
rect 28976 2694 29028 2746
rect 39828 2694 39880 2746
rect 39892 2694 39944 2746
rect 39956 2694 40008 2746
rect 40020 2694 40072 2746
rect 40084 2694 40136 2746
rect 20536 2592 20588 2644
rect 22928 2592 22980 2644
rect 23020 2592 23072 2644
rect 23664 2635 23716 2644
rect 23664 2601 23673 2635
rect 23673 2601 23707 2635
rect 23707 2601 23716 2635
rect 23664 2592 23716 2601
rect 23940 2635 23992 2644
rect 23940 2601 23949 2635
rect 23949 2601 23983 2635
rect 23983 2601 23992 2635
rect 23940 2592 23992 2601
rect 24216 2635 24268 2644
rect 24216 2601 24225 2635
rect 24225 2601 24259 2635
rect 24259 2601 24268 2635
rect 24216 2592 24268 2601
rect 24860 2635 24912 2644
rect 24860 2601 24869 2635
rect 24869 2601 24903 2635
rect 24903 2601 24912 2635
rect 24860 2592 24912 2601
rect 27068 2635 27120 2644
rect 27068 2601 27077 2635
rect 27077 2601 27111 2635
rect 27111 2601 27120 2635
rect 27068 2592 27120 2601
rect 29276 2635 29328 2644
rect 29276 2601 29285 2635
rect 29285 2601 29319 2635
rect 29319 2601 29328 2635
rect 29276 2592 29328 2601
rect 22284 2456 22336 2508
rect 22192 2431 22244 2440
rect 22192 2397 22201 2431
rect 22201 2397 22235 2431
rect 22235 2397 22244 2431
rect 22192 2388 22244 2397
rect 22468 2388 22520 2440
rect 23296 2456 23348 2508
rect 25504 2456 25556 2508
rect 20352 2363 20404 2372
rect 20352 2329 20361 2363
rect 20361 2329 20395 2363
rect 20395 2329 20404 2363
rect 20352 2320 20404 2329
rect 21456 2320 21508 2372
rect 22836 2320 22888 2372
rect 23020 2320 23072 2372
rect 23756 2431 23808 2440
rect 23756 2397 23765 2431
rect 23765 2397 23799 2431
rect 23799 2397 23808 2431
rect 23756 2388 23808 2397
rect 23940 2388 23992 2440
rect 24676 2431 24728 2440
rect 24676 2397 24685 2431
rect 24685 2397 24719 2431
rect 24719 2397 24728 2431
rect 24676 2388 24728 2397
rect 43260 2592 43312 2644
rect 43904 2635 43956 2644
rect 43904 2601 43913 2635
rect 43913 2601 43947 2635
rect 43947 2601 43956 2635
rect 43904 2592 43956 2601
rect 44180 2635 44232 2644
rect 44180 2601 44189 2635
rect 44189 2601 44223 2635
rect 44223 2601 44232 2635
rect 44180 2592 44232 2601
rect 44272 2592 44324 2644
rect 44456 2635 44508 2644
rect 44456 2601 44465 2635
rect 44465 2601 44499 2635
rect 44499 2601 44508 2635
rect 44456 2592 44508 2601
rect 45008 2635 45060 2644
rect 45008 2601 45017 2635
rect 45017 2601 45051 2635
rect 45051 2601 45060 2635
rect 45008 2592 45060 2601
rect 39672 2524 39724 2576
rect 41604 2456 41656 2508
rect 26884 2431 26936 2440
rect 26884 2397 26893 2431
rect 26893 2397 26927 2431
rect 26927 2397 26936 2431
rect 26884 2388 26936 2397
rect 29092 2431 29144 2440
rect 29092 2397 29101 2431
rect 29101 2397 29135 2431
rect 29135 2397 29144 2431
rect 29092 2388 29144 2397
rect 31300 2431 31352 2440
rect 31300 2397 31309 2431
rect 31309 2397 31343 2431
rect 31343 2397 31352 2431
rect 31300 2388 31352 2397
rect 33508 2431 33560 2440
rect 33508 2397 33517 2431
rect 33517 2397 33551 2431
rect 33551 2397 33560 2431
rect 33508 2388 33560 2397
rect 35716 2431 35768 2440
rect 35716 2397 35725 2431
rect 35725 2397 35759 2431
rect 35759 2397 35768 2431
rect 35716 2388 35768 2397
rect 37924 2431 37976 2440
rect 37924 2397 37933 2431
rect 37933 2397 37967 2431
rect 37967 2397 37976 2431
rect 37924 2388 37976 2397
rect 44088 2431 44140 2440
rect 44088 2397 44097 2431
rect 44097 2397 44131 2431
rect 44131 2397 44140 2431
rect 44088 2388 44140 2397
rect 36084 2320 36136 2372
rect 43444 2320 43496 2372
rect 44824 2388 44876 2440
rect 45192 2431 45244 2440
rect 45192 2397 45201 2431
rect 45201 2397 45235 2431
rect 45235 2397 45244 2431
rect 45192 2388 45244 2397
rect 12058 2150 12110 2202
rect 12122 2150 12174 2202
rect 12186 2150 12238 2202
rect 12250 2150 12302 2202
rect 12314 2150 12366 2202
rect 23166 2150 23218 2202
rect 23230 2150 23282 2202
rect 23294 2150 23346 2202
rect 23358 2150 23410 2202
rect 23422 2150 23474 2202
rect 34274 2150 34326 2202
rect 34338 2150 34390 2202
rect 34402 2150 34454 2202
rect 34466 2150 34518 2202
rect 34530 2150 34582 2202
rect 45382 2150 45434 2202
rect 45446 2150 45498 2202
rect 45510 2150 45562 2202
rect 45574 2150 45626 2202
rect 45638 2150 45690 2202
rect 20352 2048 20404 2100
rect 20628 2048 20680 2100
rect 22192 2048 22244 2100
rect 22284 2091 22336 2100
rect 22284 2057 22293 2091
rect 22293 2057 22327 2091
rect 22327 2057 22336 2091
rect 22284 2048 22336 2057
rect 1584 1912 1636 1964
rect 19616 1955 19668 1964
rect 19616 1921 19625 1955
rect 19625 1921 19659 1955
rect 19659 1921 19668 1955
rect 19616 1912 19668 1921
rect 23020 2048 23072 2100
rect 23756 2048 23808 2100
rect 24676 2048 24728 2100
rect 26884 2048 26936 2100
rect 29092 2048 29144 2100
rect 31300 2048 31352 2100
rect 33508 2048 33560 2100
rect 35716 2048 35768 2100
rect 37924 2048 37976 2100
rect 41604 2091 41656 2100
rect 41604 2057 41613 2091
rect 41613 2057 41647 2091
rect 41647 2057 41656 2091
rect 41604 2048 41656 2057
rect 43444 2091 43496 2100
rect 43444 2057 43453 2091
rect 43453 2057 43487 2091
rect 43487 2057 43496 2091
rect 43444 2048 43496 2057
rect 23940 1980 23992 2032
rect 44088 2048 44140 2100
rect 45192 1980 45244 2032
rect 20720 1912 20772 1964
rect 21640 1955 21692 1964
rect 21640 1921 21649 1955
rect 21649 1921 21683 1955
rect 21683 1921 21692 1955
rect 21640 1912 21692 1921
rect 22192 1955 22244 1964
rect 22192 1921 22201 1955
rect 22201 1921 22235 1955
rect 22235 1921 22244 1955
rect 22192 1912 22244 1921
rect 20812 1844 20864 1896
rect 22836 1955 22888 1964
rect 22836 1921 22845 1955
rect 22845 1921 22879 1955
rect 22879 1921 22888 1955
rect 22836 1912 22888 1921
rect 23020 1912 23072 1964
rect 23664 1912 23716 1964
rect 24032 1955 24084 1964
rect 24032 1921 24041 1955
rect 24041 1921 24075 1955
rect 24075 1921 24084 1955
rect 24032 1912 24084 1921
rect 26240 1955 26292 1964
rect 26240 1921 26249 1955
rect 26249 1921 26283 1955
rect 26283 1921 26292 1955
rect 26240 1912 26292 1921
rect 28448 1955 28500 1964
rect 28448 1921 28457 1955
rect 28457 1921 28491 1955
rect 28491 1921 28500 1955
rect 28448 1912 28500 1921
rect 30656 1955 30708 1964
rect 30656 1921 30665 1955
rect 30665 1921 30699 1955
rect 30699 1921 30708 1955
rect 30656 1912 30708 1921
rect 32864 1955 32916 1964
rect 32864 1921 32873 1955
rect 32873 1921 32907 1955
rect 32907 1921 32916 1955
rect 32864 1912 32916 1921
rect 35072 1955 35124 1964
rect 35072 1921 35081 1955
rect 35081 1921 35115 1955
rect 35115 1921 35124 1955
rect 35072 1912 35124 1921
rect 37464 1955 37516 1964
rect 37464 1921 37473 1955
rect 37473 1921 37507 1955
rect 37507 1921 37516 1955
rect 37464 1912 37516 1921
rect 41788 1955 41840 1964
rect 41788 1921 41797 1955
rect 41797 1921 41831 1955
rect 41831 1921 41840 1955
rect 41788 1912 41840 1921
rect 43628 1955 43680 1964
rect 43628 1921 43637 1955
rect 43637 1921 43671 1955
rect 43671 1921 43680 1955
rect 43628 1912 43680 1921
rect 44088 1955 44140 1964
rect 44088 1921 44097 1955
rect 44097 1921 44131 1955
rect 44131 1921 44140 1955
rect 44088 1912 44140 1921
rect 44548 1955 44600 1964
rect 44548 1921 44557 1955
rect 44557 1921 44591 1955
rect 44591 1921 44600 1955
rect 44548 1912 44600 1921
rect 22468 1776 22520 1828
rect 21456 1751 21508 1760
rect 21456 1717 21465 1751
rect 21465 1717 21499 1751
rect 21499 1717 21508 1751
rect 21456 1708 21508 1717
rect 21548 1708 21600 1760
rect 22744 1708 22796 1760
rect 6504 1606 6556 1658
rect 6568 1606 6620 1658
rect 6632 1606 6684 1658
rect 6696 1606 6748 1658
rect 6760 1606 6812 1658
rect 17612 1606 17664 1658
rect 17676 1606 17728 1658
rect 17740 1606 17792 1658
rect 17804 1606 17856 1658
rect 17868 1606 17920 1658
rect 28720 1606 28772 1658
rect 28784 1606 28836 1658
rect 28848 1606 28900 1658
rect 28912 1606 28964 1658
rect 28976 1606 29028 1658
rect 39828 1606 39880 1658
rect 39892 1606 39944 1658
rect 39956 1606 40008 1658
rect 40020 1606 40072 1658
rect 40084 1606 40136 1658
rect 1584 1547 1636 1556
rect 1584 1513 1593 1547
rect 1593 1513 1627 1547
rect 1627 1513 1636 1547
rect 1584 1504 1636 1513
rect 19616 1504 19668 1556
rect 21640 1504 21692 1556
rect 22836 1504 22888 1556
rect 24032 1504 24084 1556
rect 28448 1504 28500 1556
rect 32864 1504 32916 1556
rect 35072 1504 35124 1556
rect 44088 1504 44140 1556
rect 44548 1504 44600 1556
rect 1216 1300 1268 1352
rect 3792 1343 3844 1352
rect 3792 1309 3801 1343
rect 3801 1309 3835 1343
rect 3835 1309 3844 1343
rect 3792 1300 3844 1309
rect 5724 1343 5776 1352
rect 5724 1309 5733 1343
rect 5733 1309 5767 1343
rect 5767 1309 5776 1343
rect 5724 1300 5776 1309
rect 7932 1343 7984 1352
rect 7932 1309 7941 1343
rect 7941 1309 7975 1343
rect 7975 1309 7984 1343
rect 7932 1300 7984 1309
rect 10140 1343 10192 1352
rect 10140 1309 10149 1343
rect 10149 1309 10183 1343
rect 10183 1309 10192 1343
rect 10140 1300 10192 1309
rect 12072 1300 12124 1352
rect 14740 1343 14792 1352
rect 14740 1309 14749 1343
rect 14749 1309 14783 1343
rect 14783 1309 14792 1343
rect 14740 1300 14792 1309
rect 3976 1207 4028 1216
rect 3976 1173 3985 1207
rect 3985 1173 4019 1207
rect 4019 1173 4028 1207
rect 3976 1164 4028 1173
rect 8116 1207 8168 1216
rect 8116 1173 8125 1207
rect 8125 1173 8159 1207
rect 8159 1173 8168 1207
rect 8116 1164 8168 1173
rect 10324 1207 10376 1216
rect 10324 1173 10333 1207
rect 10333 1173 10367 1207
rect 10367 1173 10376 1207
rect 10324 1164 10376 1173
rect 14648 1232 14700 1284
rect 16948 1343 17000 1352
rect 16948 1309 16957 1343
rect 16957 1309 16991 1343
rect 16991 1309 17000 1343
rect 16948 1300 17000 1309
rect 19432 1343 19484 1352
rect 19432 1309 19441 1343
rect 19441 1309 19475 1343
rect 19475 1309 19484 1343
rect 19432 1300 19484 1309
rect 20720 1232 20772 1284
rect 21364 1343 21416 1352
rect 21364 1309 21373 1343
rect 21373 1309 21407 1343
rect 21407 1309 21416 1343
rect 21364 1300 21416 1309
rect 22284 1343 22336 1352
rect 22284 1309 22293 1343
rect 22293 1309 22327 1343
rect 22327 1309 22336 1343
rect 22284 1300 22336 1309
rect 23572 1343 23624 1352
rect 23572 1309 23581 1343
rect 23581 1309 23615 1343
rect 23615 1309 23624 1343
rect 23572 1300 23624 1309
rect 25780 1343 25832 1352
rect 25780 1309 25789 1343
rect 25789 1309 25823 1343
rect 25823 1309 25832 1343
rect 25780 1300 25832 1309
rect 27988 1343 28040 1352
rect 27988 1309 27997 1343
rect 27997 1309 28031 1343
rect 28031 1309 28040 1343
rect 27988 1300 28040 1309
rect 30196 1343 30248 1352
rect 30196 1309 30205 1343
rect 30205 1309 30239 1343
rect 30239 1309 30248 1343
rect 30196 1300 30248 1309
rect 30656 1300 30708 1352
rect 32404 1343 32456 1352
rect 32404 1309 32413 1343
rect 32413 1309 32447 1343
rect 32447 1309 32456 1343
rect 32404 1300 32456 1309
rect 34612 1300 34664 1352
rect 36820 1343 36872 1352
rect 36820 1309 36829 1343
rect 36829 1309 36863 1343
rect 36863 1309 36872 1343
rect 36820 1300 36872 1309
rect 37464 1300 37516 1352
rect 39028 1343 39080 1352
rect 39028 1309 39037 1343
rect 39037 1309 39071 1343
rect 39071 1309 39080 1343
rect 39028 1300 39080 1309
rect 41236 1343 41288 1352
rect 41236 1309 41245 1343
rect 41245 1309 41279 1343
rect 41279 1309 41288 1343
rect 41236 1300 41288 1309
rect 43444 1343 43496 1352
rect 43444 1309 43453 1343
rect 43453 1309 43487 1343
rect 43487 1309 43496 1343
rect 43444 1300 43496 1309
rect 45192 1343 45244 1352
rect 45192 1309 45201 1343
rect 45201 1309 45235 1343
rect 45235 1309 45244 1343
rect 45192 1300 45244 1309
rect 22192 1232 22244 1284
rect 14556 1207 14608 1216
rect 14556 1173 14565 1207
rect 14565 1173 14599 1207
rect 14599 1173 14608 1207
rect 14556 1164 14608 1173
rect 26240 1164 26292 1216
rect 43628 1232 43680 1284
rect 41788 1164 41840 1216
rect 12058 1062 12110 1114
rect 12122 1062 12174 1114
rect 12186 1062 12238 1114
rect 12250 1062 12302 1114
rect 12314 1062 12366 1114
rect 23166 1062 23218 1114
rect 23230 1062 23282 1114
rect 23294 1062 23346 1114
rect 23358 1062 23410 1114
rect 23422 1062 23474 1114
rect 34274 1062 34326 1114
rect 34338 1062 34390 1114
rect 34402 1062 34454 1114
rect 34466 1062 34518 1114
rect 34530 1062 34582 1114
rect 45382 1062 45434 1114
rect 45446 1062 45498 1114
rect 45510 1062 45562 1114
rect 45574 1062 45626 1114
rect 45638 1062 45690 1114
rect 3976 960 4028 1012
rect 14556 960 14608 1012
rect 14648 960 14700 1012
rect 20812 960 20864 1012
rect 22284 960 22336 1012
rect 23664 824 23716 876
rect 8116 756 8168 808
rect 10324 756 10376 808
rect 23020 756 23072 808
rect 21548 620 21600 672
<< metal2 >>
rect 478 9840 534 10300
rect 584 9846 796 9874
rect 492 9738 520 9840
rect 584 9738 612 9846
rect 492 9710 612 9738
rect 768 8566 796 9846
rect 846 9840 902 10300
rect 1214 9840 1270 10300
rect 1582 9840 1638 10300
rect 1950 9840 2006 10300
rect 2318 9840 2374 10300
rect 2686 9840 2742 10300
rect 3054 9840 3110 10300
rect 3422 9840 3478 10300
rect 3790 9840 3846 10300
rect 3896 9846 4108 9874
rect 756 8560 808 8566
rect 756 8502 808 8508
rect 860 7546 888 9840
rect 848 7540 900 7546
rect 848 7482 900 7488
rect 1228 6866 1256 9840
rect 1596 7478 1624 9840
rect 1964 8786 1992 9840
rect 1964 8758 2084 8786
rect 2056 8090 2084 8758
rect 2332 8634 2360 9840
rect 2320 8628 2372 8634
rect 2320 8570 2372 8576
rect 2700 8242 2728 9840
rect 2700 8214 2820 8242
rect 2792 8090 2820 8214
rect 3068 8090 3096 9840
rect 3240 8832 3292 8838
rect 3240 8774 3292 8780
rect 3252 8566 3280 8774
rect 3240 8560 3292 8566
rect 3240 8502 3292 8508
rect 3436 8090 3464 9840
rect 3804 9738 3832 9840
rect 3896 9738 3924 9846
rect 3804 9710 3924 9738
rect 4080 8242 4108 9846
rect 4158 9840 4214 10300
rect 4526 9840 4582 10300
rect 4894 9840 4950 10300
rect 5262 9840 5318 10300
rect 5630 9840 5686 10300
rect 5998 9840 6054 10300
rect 6366 9840 6422 10300
rect 6734 9840 6790 10300
rect 7102 9840 7158 10300
rect 7470 9840 7526 10300
rect 7838 9840 7894 10300
rect 8206 9840 8262 10300
rect 8574 9840 8630 10300
rect 8760 9920 8812 9926
rect 8760 9862 8812 9868
rect 4172 8634 4200 9840
rect 4160 8628 4212 8634
rect 4160 8570 4212 8576
rect 4080 8214 4200 8242
rect 4172 8090 4200 8214
rect 4540 8090 4568 9840
rect 4804 9240 4856 9246
rect 4804 9182 4856 9188
rect 4816 8498 4844 9182
rect 4908 8634 4936 9840
rect 5276 8634 5304 9840
rect 5356 9784 5408 9790
rect 5356 9726 5408 9732
rect 4896 8628 4948 8634
rect 4896 8570 4948 8576
rect 5264 8628 5316 8634
rect 5264 8570 5316 8576
rect 5368 8498 5396 9726
rect 5448 8968 5500 8974
rect 5448 8910 5500 8916
rect 5460 8634 5488 8910
rect 5644 8634 5672 9840
rect 5816 9648 5868 9654
rect 5816 9590 5868 9596
rect 5448 8628 5500 8634
rect 5448 8570 5500 8576
rect 5632 8628 5684 8634
rect 5632 8570 5684 8576
rect 5828 8566 5856 9590
rect 6012 8634 6040 9840
rect 6000 8628 6052 8634
rect 6000 8570 6052 8576
rect 5816 8560 5868 8566
rect 5816 8502 5868 8508
rect 4804 8492 4856 8498
rect 4804 8434 4856 8440
rect 5356 8492 5408 8498
rect 5356 8434 5408 8440
rect 6380 8090 6408 9840
rect 6748 8634 6776 9840
rect 6736 8628 6788 8634
rect 6736 8570 6788 8576
rect 7012 8628 7064 8634
rect 7116 8616 7144 9840
rect 7380 9512 7432 9518
rect 7380 9454 7432 9460
rect 7064 8588 7144 8616
rect 7012 8570 7064 8576
rect 7392 8498 7420 9454
rect 7380 8492 7432 8498
rect 7380 8434 7432 8440
rect 6504 8188 6812 8197
rect 6504 8186 6510 8188
rect 6566 8186 6590 8188
rect 6646 8186 6670 8188
rect 6726 8186 6750 8188
rect 6806 8186 6812 8188
rect 6566 8134 6568 8186
rect 6748 8134 6750 8186
rect 6504 8132 6510 8134
rect 6566 8132 6590 8134
rect 6646 8132 6670 8134
rect 6726 8132 6750 8134
rect 6806 8132 6812 8134
rect 6504 8123 6812 8132
rect 7484 8090 7512 9840
rect 7564 9716 7616 9722
rect 7564 9658 7616 9664
rect 7576 8498 7604 9658
rect 7852 8634 7880 9840
rect 8024 9784 8076 9790
rect 8024 9726 8076 9732
rect 7840 8628 7892 8634
rect 7840 8570 7892 8576
rect 8036 8498 8064 9726
rect 8116 8628 8168 8634
rect 8220 8616 8248 9840
rect 8484 8832 8536 8838
rect 8484 8774 8536 8780
rect 8168 8588 8248 8616
rect 8116 8570 8168 8576
rect 8496 8498 8524 8774
rect 8588 8634 8616 9840
rect 8576 8628 8628 8634
rect 8576 8570 8628 8576
rect 8772 8498 8800 9862
rect 8942 9840 8998 10300
rect 9048 9846 9168 9874
rect 9048 9840 9076 9846
rect 8956 9812 9076 9840
rect 8852 9240 8904 9246
rect 8852 9182 8904 9188
rect 9036 9240 9088 9246
rect 9036 9182 9088 9188
rect 8864 8566 8892 9182
rect 8852 8560 8904 8566
rect 8852 8502 8904 8508
rect 9048 8498 9076 9182
rect 7564 8492 7616 8498
rect 7564 8434 7616 8440
rect 8024 8492 8076 8498
rect 8024 8434 8076 8440
rect 8484 8492 8536 8498
rect 8484 8434 8536 8440
rect 8760 8492 8812 8498
rect 8760 8434 8812 8440
rect 9036 8492 9088 8498
rect 9036 8434 9088 8440
rect 9140 8090 9168 9846
rect 9310 9840 9366 10300
rect 9496 9852 9548 9858
rect 9324 8634 9352 9840
rect 9678 9840 9734 10300
rect 10046 9840 10102 10300
rect 10414 9840 10470 10300
rect 10782 9840 10838 10300
rect 11150 9840 11206 10300
rect 11518 9840 11574 10300
rect 11886 9840 11942 10300
rect 11992 9846 12204 9874
rect 9496 9794 9548 9800
rect 9312 8628 9364 8634
rect 9312 8570 9364 8576
rect 9508 8498 9536 9794
rect 9692 8616 9720 9840
rect 9772 8628 9824 8634
rect 9692 8588 9772 8616
rect 9772 8570 9824 8576
rect 9496 8492 9548 8498
rect 9496 8434 9548 8440
rect 10060 8090 10088 9840
rect 10428 8634 10456 9840
rect 10508 9104 10560 9110
rect 10508 9046 10560 9052
rect 10416 8628 10468 8634
rect 10416 8570 10468 8576
rect 10520 8498 10548 9046
rect 10796 8634 10824 9840
rect 10784 8628 10836 8634
rect 11164 8616 11192 9840
rect 11532 8786 11560 9840
rect 11796 8832 11848 8838
rect 11532 8758 11652 8786
rect 11796 8774 11848 8780
rect 11244 8628 11296 8634
rect 11164 8588 11244 8616
rect 10784 8570 10836 8576
rect 11244 8570 11296 8576
rect 10416 8492 10468 8498
rect 10416 8434 10468 8440
rect 10508 8492 10560 8498
rect 10508 8434 10560 8440
rect 2044 8084 2096 8090
rect 2044 8026 2096 8032
rect 2780 8084 2832 8090
rect 2780 8026 2832 8032
rect 3056 8084 3108 8090
rect 3056 8026 3108 8032
rect 3424 8084 3476 8090
rect 3424 8026 3476 8032
rect 4160 8084 4212 8090
rect 4160 8026 4212 8032
rect 4528 8084 4580 8090
rect 4528 8026 4580 8032
rect 6368 8084 6420 8090
rect 6368 8026 6420 8032
rect 7472 8084 7524 8090
rect 7472 8026 7524 8032
rect 9128 8084 9180 8090
rect 9128 8026 9180 8032
rect 10048 8084 10100 8090
rect 10048 8026 10100 8032
rect 10428 8022 10456 8434
rect 11624 8090 11652 8758
rect 11808 8566 11836 8774
rect 11796 8560 11848 8566
rect 11796 8502 11848 8508
rect 11900 8090 11928 9840
rect 11992 8634 12020 9846
rect 12176 9840 12204 9846
rect 12254 9840 12310 10300
rect 12622 9840 12678 10300
rect 12990 9840 13046 10300
rect 13358 9840 13414 10300
rect 13636 9988 13688 9994
rect 13636 9930 13688 9936
rect 12176 9812 12296 9840
rect 12438 8936 12494 8945
rect 12438 8871 12494 8880
rect 12058 8732 12366 8741
rect 12058 8730 12064 8732
rect 12120 8730 12144 8732
rect 12200 8730 12224 8732
rect 12280 8730 12304 8732
rect 12360 8730 12366 8732
rect 12120 8678 12122 8730
rect 12302 8678 12304 8730
rect 12058 8676 12064 8678
rect 12120 8676 12144 8678
rect 12200 8676 12224 8678
rect 12280 8676 12304 8678
rect 12360 8676 12366 8678
rect 12058 8667 12366 8676
rect 11980 8628 12032 8634
rect 11980 8570 12032 8576
rect 12452 8566 12480 8871
rect 12532 8628 12584 8634
rect 12636 8616 12664 9840
rect 12584 8588 12664 8616
rect 12532 8570 12584 8576
rect 12440 8560 12492 8566
rect 12440 8502 12492 8508
rect 12624 8492 12676 8498
rect 12624 8434 12676 8440
rect 11612 8084 11664 8090
rect 11612 8026 11664 8032
rect 11888 8084 11940 8090
rect 11888 8026 11940 8032
rect 10416 8016 10468 8022
rect 10416 7958 10468 7964
rect 2964 7880 3016 7886
rect 2964 7822 3016 7828
rect 3332 7880 3384 7886
rect 3332 7822 3384 7828
rect 4436 7880 4488 7886
rect 4436 7822 4488 7828
rect 9956 7880 10008 7886
rect 9956 7822 10008 7828
rect 11520 7880 11572 7886
rect 11520 7822 11572 7828
rect 2504 7812 2556 7818
rect 2504 7754 2556 7760
rect 1584 7472 1636 7478
rect 1584 7414 1636 7420
rect 1216 6860 1268 6866
rect 1216 6802 1268 6808
rect 1492 6724 1544 6730
rect 1492 6666 1544 6672
rect 1504 6458 1532 6666
rect 1492 6452 1544 6458
rect 1492 6394 1544 6400
rect 2516 6390 2544 7754
rect 2504 6384 2556 6390
rect 2504 6326 2556 6332
rect 2976 6254 3004 7822
rect 3344 6662 3372 7822
rect 3884 7812 3936 7818
rect 3884 7754 3936 7760
rect 3896 7546 3924 7754
rect 3884 7540 3936 7546
rect 3884 7482 3936 7488
rect 4448 7342 4476 7822
rect 6368 7812 6420 7818
rect 6368 7754 6420 7760
rect 5448 7744 5500 7750
rect 5448 7686 5500 7692
rect 4436 7336 4488 7342
rect 4436 7278 4488 7284
rect 5460 6905 5488 7686
rect 6380 7342 6408 7754
rect 6368 7336 6420 7342
rect 6368 7278 6420 7284
rect 6504 7100 6812 7109
rect 6504 7098 6510 7100
rect 6566 7098 6590 7100
rect 6646 7098 6670 7100
rect 6726 7098 6750 7100
rect 6806 7098 6812 7100
rect 6566 7046 6568 7098
rect 6748 7046 6750 7098
rect 6504 7044 6510 7046
rect 6566 7044 6590 7046
rect 6646 7044 6670 7046
rect 6726 7044 6750 7046
rect 6806 7044 6812 7046
rect 6504 7035 6812 7044
rect 9968 7002 9996 7822
rect 11060 7540 11112 7546
rect 11060 7482 11112 7488
rect 11072 7342 11100 7482
rect 11532 7449 11560 7822
rect 12058 7644 12366 7653
rect 12058 7642 12064 7644
rect 12120 7642 12144 7644
rect 12200 7642 12224 7644
rect 12280 7642 12304 7644
rect 12360 7642 12366 7644
rect 12120 7590 12122 7642
rect 12302 7590 12304 7642
rect 12058 7588 12064 7590
rect 12120 7588 12144 7590
rect 12200 7588 12224 7590
rect 12280 7588 12304 7590
rect 12360 7588 12366 7590
rect 12058 7579 12366 7588
rect 11518 7440 11574 7449
rect 11518 7375 11574 7384
rect 11060 7336 11112 7342
rect 11060 7278 11112 7284
rect 12348 7336 12400 7342
rect 12348 7278 12400 7284
rect 9956 6996 10008 7002
rect 9956 6938 10008 6944
rect 5446 6896 5502 6905
rect 5446 6831 5502 6840
rect 12360 6730 12388 7278
rect 12636 6769 12664 8434
rect 13004 8090 13032 9840
rect 13084 9308 13136 9314
rect 13084 9250 13136 9256
rect 13176 9308 13228 9314
rect 13176 9250 13228 9256
rect 13096 8498 13124 9250
rect 13188 9042 13216 9250
rect 13176 9036 13228 9042
rect 13176 8978 13228 8984
rect 13372 8634 13400 9840
rect 13648 9625 13676 9930
rect 13726 9840 13782 10300
rect 14094 9840 14150 10300
rect 14370 9888 14426 9897
rect 14200 9846 14320 9874
rect 14200 9840 14228 9846
rect 13634 9616 13690 9625
rect 13634 9551 13690 9560
rect 13544 8832 13596 8838
rect 13544 8774 13596 8780
rect 13360 8628 13412 8634
rect 13360 8570 13412 8576
rect 13556 8498 13584 8774
rect 13636 8628 13688 8634
rect 13740 8616 13768 9840
rect 14108 9812 14228 9840
rect 14188 8900 14240 8906
rect 14188 8842 14240 8848
rect 13688 8588 13768 8616
rect 13636 8570 13688 8576
rect 14200 8498 14228 8842
rect 13084 8492 13136 8498
rect 13084 8434 13136 8440
rect 13544 8492 13596 8498
rect 13544 8434 13596 8440
rect 14188 8492 14240 8498
rect 14188 8434 14240 8440
rect 14292 8090 14320 9846
rect 14462 9840 14518 10300
rect 14648 9920 14700 9926
rect 14648 9862 14700 9868
rect 14370 9823 14372 9832
rect 14424 9823 14426 9832
rect 14372 9794 14424 9800
rect 14370 9208 14426 9217
rect 14370 9143 14426 9152
rect 14384 8430 14412 9143
rect 14476 8634 14504 9840
rect 14556 9784 14608 9790
rect 14554 9752 14556 9761
rect 14608 9752 14610 9761
rect 14554 9687 14610 9696
rect 14464 8628 14516 8634
rect 14464 8570 14516 8576
rect 14372 8424 14424 8430
rect 14372 8366 14424 8372
rect 12992 8084 13044 8090
rect 12992 8026 13044 8032
rect 14280 8084 14332 8090
rect 14280 8026 14332 8032
rect 12900 7880 12952 7886
rect 12900 7822 12952 7828
rect 12912 7410 12940 7822
rect 14188 7812 14240 7818
rect 14188 7754 14240 7760
rect 12900 7404 12952 7410
rect 12900 7346 12952 7352
rect 14200 7002 14228 7754
rect 14556 7200 14608 7206
rect 14556 7142 14608 7148
rect 14188 6996 14240 7002
rect 14188 6938 14240 6944
rect 12622 6760 12678 6769
rect 12348 6724 12400 6730
rect 12622 6695 12678 6704
rect 12348 6666 12400 6672
rect 3332 6656 3384 6662
rect 3332 6598 3384 6604
rect 12058 6556 12366 6565
rect 12058 6554 12064 6556
rect 12120 6554 12144 6556
rect 12200 6554 12224 6556
rect 12280 6554 12304 6556
rect 12360 6554 12366 6556
rect 12120 6502 12122 6554
rect 12302 6502 12304 6554
rect 12058 6500 12064 6502
rect 12120 6500 12144 6502
rect 12200 6500 12224 6502
rect 12280 6500 12304 6502
rect 12360 6500 12366 6502
rect 12058 6491 12366 6500
rect 14568 6458 14596 7142
rect 14660 6798 14688 9862
rect 14830 9840 14886 10300
rect 14924 9988 14976 9994
rect 14924 9930 14976 9936
rect 14844 8634 14872 9840
rect 14936 9654 14964 9930
rect 15198 9840 15254 10300
rect 15566 9840 15622 10300
rect 15934 9840 15990 10300
rect 16302 9840 16358 10300
rect 16488 9920 16540 9926
rect 16394 9888 16450 9897
rect 14924 9648 14976 9654
rect 14924 9590 14976 9596
rect 15016 9648 15068 9654
rect 15016 9590 15068 9596
rect 14832 8628 14884 8634
rect 14832 8570 14884 8576
rect 15028 8498 15056 9590
rect 15212 8616 15240 9840
rect 15580 8634 15608 9840
rect 15948 8634 15976 9840
rect 16316 8634 16344 9840
rect 16488 9862 16540 9868
rect 16394 9823 16450 9832
rect 16408 9790 16436 9823
rect 16396 9784 16448 9790
rect 16500 9761 16528 9862
rect 16670 9840 16726 10300
rect 16776 9846 16896 9874
rect 16776 9840 16804 9846
rect 16684 9812 16804 9840
rect 16396 9726 16448 9732
rect 16486 9752 16542 9761
rect 16486 9687 16542 9696
rect 16762 9480 16818 9489
rect 16762 9415 16818 9424
rect 16776 9314 16804 9415
rect 16764 9308 16816 9314
rect 16764 9250 16816 9256
rect 16672 8900 16724 8906
rect 16672 8842 16724 8848
rect 16764 8900 16816 8906
rect 16764 8842 16816 8848
rect 15292 8628 15344 8634
rect 15212 8588 15292 8616
rect 15292 8570 15344 8576
rect 15568 8628 15620 8634
rect 15568 8570 15620 8576
rect 15936 8628 15988 8634
rect 15936 8570 15988 8576
rect 16304 8628 16356 8634
rect 16304 8570 16356 8576
rect 15016 8492 15068 8498
rect 15016 8434 15068 8440
rect 15476 8492 15528 8498
rect 15476 8434 15528 8440
rect 16120 8492 16172 8498
rect 16120 8434 16172 8440
rect 15106 7848 15162 7857
rect 15106 7783 15108 7792
rect 15160 7783 15162 7792
rect 15108 7754 15160 7760
rect 15106 7576 15162 7585
rect 15106 7511 15108 7520
rect 15160 7511 15162 7520
rect 15108 7482 15160 7488
rect 15488 7206 15516 8434
rect 16132 8401 16160 8434
rect 16118 8392 16174 8401
rect 16118 8327 16174 8336
rect 15476 7200 15528 7206
rect 15476 7142 15528 7148
rect 16684 6866 16712 8842
rect 16776 8498 16804 8842
rect 16868 8634 16896 9846
rect 17038 9840 17094 10300
rect 17406 9840 17462 10300
rect 17684 9852 17736 9858
rect 16948 9240 17000 9246
rect 16948 9182 17000 9188
rect 16856 8628 16908 8634
rect 16856 8570 16908 8576
rect 16764 8492 16816 8498
rect 16764 8434 16816 8440
rect 16960 7449 16988 9182
rect 17052 8090 17080 9840
rect 17224 9716 17276 9722
rect 17224 9658 17276 9664
rect 17316 9716 17368 9722
rect 17316 9658 17368 9664
rect 17236 9450 17264 9658
rect 17132 9444 17184 9450
rect 17132 9386 17184 9392
rect 17224 9444 17276 9450
rect 17224 9386 17276 9392
rect 17144 9353 17172 9386
rect 17130 9344 17186 9353
rect 17328 9314 17356 9658
rect 17130 9279 17186 9288
rect 17316 9308 17368 9314
rect 17316 9250 17368 9256
rect 17420 8634 17448 9840
rect 17774 9840 17830 10300
rect 17880 9846 18092 9874
rect 17880 9840 17908 9846
rect 17788 9812 17908 9840
rect 17684 9794 17736 9800
rect 17408 8628 17460 8634
rect 17408 8570 17460 8576
rect 17316 8492 17368 8498
rect 17316 8434 17368 8440
rect 17500 8492 17552 8498
rect 17500 8434 17552 8440
rect 17040 8084 17092 8090
rect 17040 8026 17092 8032
rect 17224 8016 17276 8022
rect 17224 7958 17276 7964
rect 17236 7886 17264 7958
rect 17328 7886 17356 8434
rect 17512 8090 17540 8434
rect 17696 8276 17724 9794
rect 17776 9104 17828 9110
rect 17776 9046 17828 9052
rect 17958 9072 18014 9081
rect 17788 8838 17816 9046
rect 17958 9007 18014 9016
rect 17776 8832 17828 8838
rect 17776 8774 17828 8780
rect 17972 8514 18000 9007
rect 18064 8634 18092 9846
rect 18142 9840 18198 10300
rect 18328 9988 18380 9994
rect 18328 9930 18380 9936
rect 18420 9988 18472 9994
rect 18420 9930 18472 9936
rect 18156 8634 18184 9840
rect 18340 9761 18368 9930
rect 18326 9752 18382 9761
rect 18326 9687 18382 9696
rect 18328 9172 18380 9178
rect 18328 9114 18380 9120
rect 18052 8628 18104 8634
rect 18052 8570 18104 8576
rect 18144 8628 18196 8634
rect 18144 8570 18196 8576
rect 17972 8486 18184 8514
rect 17696 8248 18000 8276
rect 17612 8188 17920 8197
rect 17612 8186 17618 8188
rect 17674 8186 17698 8188
rect 17754 8186 17778 8188
rect 17834 8186 17858 8188
rect 17914 8186 17920 8188
rect 17674 8134 17676 8186
rect 17856 8134 17858 8186
rect 17612 8132 17618 8134
rect 17674 8132 17698 8134
rect 17754 8132 17778 8134
rect 17834 8132 17858 8134
rect 17914 8132 17920 8134
rect 17612 8123 17920 8132
rect 17500 8084 17552 8090
rect 17972 8072 18000 8248
rect 17500 8026 17552 8032
rect 17880 8044 18000 8072
rect 18050 8120 18106 8129
rect 18050 8055 18106 8064
rect 17880 7886 17908 8044
rect 17958 7984 18014 7993
rect 18064 7954 18092 8055
rect 17958 7919 18014 7928
rect 18052 7948 18104 7954
rect 17132 7880 17184 7886
rect 17132 7822 17184 7828
rect 17224 7880 17276 7886
rect 17224 7822 17276 7828
rect 17316 7880 17368 7886
rect 17316 7822 17368 7828
rect 17868 7880 17920 7886
rect 17868 7822 17920 7828
rect 17144 7546 17172 7822
rect 17224 7744 17276 7750
rect 17222 7712 17224 7721
rect 17276 7712 17278 7721
rect 17222 7647 17278 7656
rect 17132 7540 17184 7546
rect 17132 7482 17184 7488
rect 16946 7440 17002 7449
rect 16946 7375 17002 7384
rect 17612 7100 17920 7109
rect 17612 7098 17618 7100
rect 17674 7098 17698 7100
rect 17754 7098 17778 7100
rect 17834 7098 17858 7100
rect 17914 7098 17920 7100
rect 17674 7046 17676 7098
rect 17856 7046 17858 7098
rect 17612 7044 17618 7046
rect 17674 7044 17698 7046
rect 17754 7044 17778 7046
rect 17834 7044 17858 7046
rect 17914 7044 17920 7046
rect 17612 7035 17920 7044
rect 17972 6934 18000 7919
rect 18052 7890 18104 7896
rect 18156 7410 18184 8486
rect 18236 8492 18288 8498
rect 18236 8434 18288 8440
rect 18248 8090 18276 8434
rect 18236 8084 18288 8090
rect 18236 8026 18288 8032
rect 18236 7880 18288 7886
rect 18340 7868 18368 9114
rect 18288 7840 18368 7868
rect 18236 7822 18288 7828
rect 18432 7818 18460 9930
rect 18510 9840 18566 10300
rect 18878 9840 18934 10300
rect 18984 9846 19196 9874
rect 18984 9840 19012 9846
rect 18524 8634 18552 9840
rect 18892 9812 19012 9840
rect 19064 8832 19116 8838
rect 19064 8774 19116 8780
rect 18512 8628 18564 8634
rect 18512 8570 18564 8576
rect 18880 8492 18932 8498
rect 18880 8434 18932 8440
rect 18786 8256 18842 8265
rect 18786 8191 18842 8200
rect 18800 7886 18828 8191
rect 18788 7880 18840 7886
rect 18788 7822 18840 7828
rect 18420 7812 18472 7818
rect 18420 7754 18472 7760
rect 18512 7744 18564 7750
rect 18512 7686 18564 7692
rect 18696 7744 18748 7750
rect 18696 7686 18748 7692
rect 18144 7404 18196 7410
rect 18144 7346 18196 7352
rect 17960 6928 18012 6934
rect 17960 6870 18012 6876
rect 16672 6860 16724 6866
rect 16672 6802 16724 6808
rect 14648 6792 14700 6798
rect 14648 6734 14700 6740
rect 17224 6656 17276 6662
rect 17224 6598 17276 6604
rect 17236 6458 17264 6598
rect 14464 6452 14516 6458
rect 14464 6394 14516 6400
rect 14556 6452 14608 6458
rect 14556 6394 14608 6400
rect 17224 6452 17276 6458
rect 17224 6394 17276 6400
rect 14476 6254 14504 6394
rect 18524 6322 18552 7686
rect 18708 7546 18736 7686
rect 18786 7576 18842 7585
rect 18696 7540 18748 7546
rect 18892 7546 18920 8434
rect 18786 7511 18788 7520
rect 18696 7482 18748 7488
rect 18840 7511 18842 7520
rect 18880 7540 18932 7546
rect 18788 7482 18840 7488
rect 18880 7482 18932 7488
rect 19076 7410 19104 8774
rect 19168 8634 19196 9846
rect 19246 9840 19302 10300
rect 19524 9988 19576 9994
rect 19524 9930 19576 9936
rect 19156 8628 19208 8634
rect 19156 8570 19208 8576
rect 19156 8424 19208 8430
rect 19156 8366 19208 8372
rect 19168 7546 19196 8366
rect 19260 8090 19288 9840
rect 19536 9654 19564 9930
rect 19614 9840 19670 10300
rect 19892 9920 19944 9926
rect 19890 9888 19892 9897
rect 19944 9888 19946 9897
rect 19340 9648 19392 9654
rect 19340 9590 19392 9596
rect 19524 9648 19576 9654
rect 19524 9590 19576 9596
rect 19352 9314 19380 9590
rect 19340 9308 19392 9314
rect 19340 9250 19392 9256
rect 19628 8650 19656 9840
rect 19982 9840 20038 10300
rect 20350 9840 20406 10300
rect 20628 9988 20680 9994
rect 20628 9930 20680 9936
rect 20456 9846 20576 9874
rect 20456 9840 20484 9846
rect 19890 9823 19946 9832
rect 19996 9738 20024 9840
rect 20364 9812 20484 9840
rect 19536 8622 19656 8650
rect 19720 9710 20024 9738
rect 20076 9784 20128 9790
rect 20076 9726 20128 9732
rect 19432 8288 19484 8294
rect 19432 8230 19484 8236
rect 19248 8084 19300 8090
rect 19248 8026 19300 8032
rect 19444 8022 19472 8230
rect 19340 8016 19392 8022
rect 19340 7958 19392 7964
rect 19432 8016 19484 8022
rect 19432 7958 19484 7964
rect 19352 7750 19380 7958
rect 19340 7744 19392 7750
rect 19340 7686 19392 7692
rect 19156 7540 19208 7546
rect 19156 7482 19208 7488
rect 19064 7404 19116 7410
rect 19064 7346 19116 7352
rect 19432 7404 19484 7410
rect 19536 7392 19564 8622
rect 19616 8492 19668 8498
rect 19720 8480 19748 9710
rect 19984 9580 20036 9586
rect 19984 9522 20036 9528
rect 19892 9308 19944 9314
rect 19892 9250 19944 9256
rect 19668 8452 19748 8480
rect 19616 8434 19668 8440
rect 19904 7546 19932 9250
rect 19996 8566 20024 9522
rect 19984 8560 20036 8566
rect 19984 8502 20036 8508
rect 20088 7834 20116 9726
rect 20166 9480 20222 9489
rect 20166 9415 20222 9424
rect 20180 8974 20208 9415
rect 20168 8968 20220 8974
rect 20168 8910 20220 8916
rect 20260 8900 20312 8906
rect 20312 8860 20484 8888
rect 20260 8842 20312 8848
rect 20260 8628 20312 8634
rect 20260 8570 20312 8576
rect 20272 7954 20300 8570
rect 20352 8288 20404 8294
rect 20352 8230 20404 8236
rect 20364 8022 20392 8230
rect 20456 8090 20484 8860
rect 20548 8498 20576 9846
rect 20536 8492 20588 8498
rect 20536 8434 20588 8440
rect 20640 8378 20668 9930
rect 20718 9840 20774 10300
rect 21086 9840 21142 10300
rect 21454 9840 21510 10300
rect 21652 9846 21772 9874
rect 20732 8480 20760 9840
rect 20810 9344 20866 9353
rect 20866 9302 20944 9330
rect 20810 9279 20866 9288
rect 20812 8492 20864 8498
rect 20732 8452 20812 8480
rect 20812 8434 20864 8440
rect 20810 8392 20866 8401
rect 20536 8356 20588 8362
rect 20640 8350 20760 8378
rect 20536 8298 20588 8304
rect 20444 8084 20496 8090
rect 20444 8026 20496 8032
rect 20352 8016 20404 8022
rect 20352 7958 20404 7964
rect 20260 7948 20312 7954
rect 20260 7890 20312 7896
rect 20548 7886 20576 8298
rect 20732 7970 20760 8350
rect 20810 8327 20866 8336
rect 20640 7942 20760 7970
rect 20640 7886 20668 7942
rect 20536 7880 20588 7886
rect 20088 7806 20208 7834
rect 20536 7822 20588 7828
rect 20628 7880 20680 7886
rect 20628 7822 20680 7828
rect 20076 7744 20128 7750
rect 20076 7686 20128 7692
rect 19892 7540 19944 7546
rect 19892 7482 19944 7488
rect 19616 7404 19668 7410
rect 19536 7364 19616 7392
rect 19432 7346 19484 7352
rect 19616 7346 19668 7352
rect 19444 6866 19472 7346
rect 19432 6860 19484 6866
rect 19432 6802 19484 6808
rect 20088 6798 20116 7686
rect 20180 6798 20208 7806
rect 20824 7478 20852 8327
rect 20916 8090 20944 9302
rect 21100 8498 21128 9840
rect 21178 9752 21234 9761
rect 21234 9710 21312 9738
rect 21178 9687 21234 9696
rect 21178 9616 21234 9625
rect 21178 9551 21234 9560
rect 21088 8492 21140 8498
rect 21088 8434 21140 8440
rect 21192 8378 21220 9551
rect 21100 8350 21220 8378
rect 20904 8084 20956 8090
rect 20904 8026 20956 8032
rect 20812 7472 20864 7478
rect 20812 7414 20864 7420
rect 21100 7410 21128 8350
rect 21284 8344 21312 9710
rect 21364 8492 21416 8498
rect 21468 8480 21496 9840
rect 21652 8498 21680 9846
rect 21744 9840 21772 9846
rect 21822 9840 21878 10300
rect 21928 9846 22140 9874
rect 21744 9812 21864 9840
rect 21416 8452 21496 8480
rect 21640 8492 21692 8498
rect 21364 8434 21416 8440
rect 21928 8480 21956 9846
rect 22112 9840 22140 9846
rect 22190 9840 22246 10300
rect 22296 9846 22508 9874
rect 22112 9812 22232 9840
rect 22192 9036 22244 9042
rect 22192 8978 22244 8984
rect 22008 8492 22060 8498
rect 21928 8452 22008 8480
rect 21640 8434 21692 8440
rect 22008 8434 22060 8440
rect 22100 8492 22152 8498
rect 22100 8434 22152 8440
rect 21548 8356 21600 8362
rect 21284 8316 21404 8344
rect 21180 8288 21232 8294
rect 21180 8230 21232 8236
rect 21270 8256 21326 8265
rect 21192 8090 21220 8230
rect 21270 8191 21326 8200
rect 21180 8084 21232 8090
rect 21180 8026 21232 8032
rect 21284 7993 21312 8191
rect 21270 7984 21326 7993
rect 21270 7919 21326 7928
rect 21376 7750 21404 8316
rect 21548 8298 21600 8304
rect 21916 8356 21968 8362
rect 21916 8298 21968 8304
rect 21456 8288 21508 8294
rect 21456 8230 21508 8236
rect 21468 7886 21496 8230
rect 21560 8090 21588 8298
rect 21824 8288 21876 8294
rect 21824 8230 21876 8236
rect 21836 8090 21864 8230
rect 21548 8084 21600 8090
rect 21548 8026 21600 8032
rect 21824 8084 21876 8090
rect 21824 8026 21876 8032
rect 21456 7880 21508 7886
rect 21456 7822 21508 7828
rect 21732 7880 21784 7886
rect 21732 7822 21784 7828
rect 21640 7812 21692 7818
rect 21640 7754 21692 7760
rect 21364 7744 21416 7750
rect 21364 7686 21416 7692
rect 21456 7744 21508 7750
rect 21652 7721 21680 7754
rect 21456 7686 21508 7692
rect 21638 7712 21694 7721
rect 21088 7404 21140 7410
rect 21088 7346 21140 7352
rect 21468 7274 21496 7686
rect 21638 7647 21694 7656
rect 21640 7336 21692 7342
rect 21744 7313 21772 7822
rect 21824 7744 21876 7750
rect 21824 7686 21876 7692
rect 21836 7546 21864 7686
rect 21824 7540 21876 7546
rect 21824 7482 21876 7488
rect 21928 7410 21956 8298
rect 22112 8106 22140 8434
rect 22204 8362 22232 8978
rect 22296 8498 22324 9846
rect 22480 9840 22508 9846
rect 22558 9840 22614 10300
rect 22664 9846 22876 9874
rect 22480 9812 22600 9840
rect 22376 9512 22428 9518
rect 22376 9454 22428 9460
rect 22388 8498 22416 9454
rect 22468 8832 22520 8838
rect 22468 8774 22520 8780
rect 22480 8537 22508 8774
rect 22466 8528 22522 8537
rect 22284 8492 22336 8498
rect 22284 8434 22336 8440
rect 22376 8492 22428 8498
rect 22466 8463 22522 8472
rect 22560 8492 22612 8498
rect 22376 8434 22428 8440
rect 22664 8480 22692 9846
rect 22848 9840 22876 9846
rect 22926 9840 22982 10300
rect 23294 9840 23350 10300
rect 23400 9846 23612 9874
rect 23400 9840 23428 9846
rect 22848 9812 22968 9840
rect 23308 9812 23428 9840
rect 22744 9784 22796 9790
rect 22744 9726 22796 9732
rect 22612 8452 22692 8480
rect 22560 8434 22612 8440
rect 22756 8378 22784 9726
rect 22928 9240 22980 9246
rect 22848 9188 22928 9194
rect 22848 9182 22980 9188
rect 22848 9166 22968 9182
rect 22848 8498 22876 9166
rect 23020 9104 23072 9110
rect 23020 9046 23072 9052
rect 22928 8968 22980 8974
rect 22928 8910 22980 8916
rect 22940 8634 22968 8910
rect 22928 8628 22980 8634
rect 22928 8570 22980 8576
rect 23032 8514 23060 9046
rect 23166 8732 23474 8741
rect 23166 8730 23172 8732
rect 23228 8730 23252 8732
rect 23308 8730 23332 8732
rect 23388 8730 23412 8732
rect 23468 8730 23474 8732
rect 23228 8678 23230 8730
rect 23410 8678 23412 8730
rect 23166 8676 23172 8678
rect 23228 8676 23252 8678
rect 23308 8676 23332 8678
rect 23388 8676 23412 8678
rect 23468 8676 23474 8678
rect 23166 8667 23474 8676
rect 23480 8628 23532 8634
rect 23480 8570 23532 8576
rect 22836 8492 22888 8498
rect 22836 8434 22888 8440
rect 22940 8486 23060 8514
rect 22192 8356 22244 8362
rect 22192 8298 22244 8304
rect 22284 8356 22336 8362
rect 22284 8298 22336 8304
rect 22376 8356 22428 8362
rect 22376 8298 22428 8304
rect 22572 8350 22784 8378
rect 22834 8392 22890 8401
rect 22112 8090 22232 8106
rect 22112 8084 22244 8090
rect 22112 8078 22192 8084
rect 22192 8026 22244 8032
rect 22100 8016 22152 8022
rect 22006 7984 22062 7993
rect 22100 7958 22152 7964
rect 22006 7919 22062 7928
rect 22020 7886 22048 7919
rect 22008 7880 22060 7886
rect 22008 7822 22060 7828
rect 22008 7744 22060 7750
rect 22008 7686 22060 7692
rect 21824 7404 21876 7410
rect 21824 7346 21876 7352
rect 21916 7404 21968 7410
rect 21916 7346 21968 7352
rect 21640 7278 21692 7284
rect 21730 7304 21786 7313
rect 21456 7268 21508 7274
rect 21456 7210 21508 7216
rect 21652 6934 21680 7278
rect 21730 7239 21786 7248
rect 21836 7018 21864 7346
rect 22020 7290 22048 7686
rect 22112 7449 22140 7958
rect 22192 7540 22244 7546
rect 22296 7528 22324 8298
rect 22244 7500 22324 7528
rect 22192 7482 22244 7488
rect 22388 7478 22416 8298
rect 22468 7948 22520 7954
rect 22468 7890 22520 7896
rect 22376 7472 22428 7478
rect 22098 7440 22154 7449
rect 22376 7414 22428 7420
rect 22098 7375 22154 7384
rect 21928 7262 22048 7290
rect 21928 7206 21956 7262
rect 21916 7200 21968 7206
rect 21916 7142 21968 7148
rect 22008 7200 22060 7206
rect 22008 7142 22060 7148
rect 22020 7018 22048 7142
rect 21836 6990 22048 7018
rect 22480 6934 22508 7890
rect 22572 7750 22600 8350
rect 22834 8327 22836 8336
rect 22888 8327 22890 8336
rect 22836 8298 22888 8304
rect 22744 7880 22796 7886
rect 22744 7822 22796 7828
rect 22560 7744 22612 7750
rect 22560 7686 22612 7692
rect 22652 7744 22704 7750
rect 22652 7686 22704 7692
rect 22664 7546 22692 7686
rect 22652 7540 22704 7546
rect 22652 7482 22704 7488
rect 22756 7410 22784 7822
rect 22836 7744 22888 7750
rect 22836 7686 22888 7692
rect 22744 7404 22796 7410
rect 22744 7346 22796 7352
rect 22744 7200 22796 7206
rect 22744 7142 22796 7148
rect 22756 7002 22784 7142
rect 22744 6996 22796 7002
rect 22744 6938 22796 6944
rect 21640 6928 21692 6934
rect 21640 6870 21692 6876
rect 22468 6928 22520 6934
rect 22468 6870 22520 6876
rect 20076 6792 20128 6798
rect 20076 6734 20128 6740
rect 20168 6792 20220 6798
rect 20168 6734 20220 6740
rect 22848 6390 22876 7686
rect 22940 7546 22968 8486
rect 23020 8424 23072 8430
rect 23020 8366 23072 8372
rect 23202 8392 23258 8401
rect 22928 7540 22980 7546
rect 22928 7482 22980 7488
rect 22926 7440 22982 7449
rect 23032 7410 23060 8366
rect 23492 8378 23520 8570
rect 23584 8498 23612 9846
rect 23662 9840 23718 10300
rect 23938 9888 23994 9897
rect 23676 9353 23704 9840
rect 24030 9840 24086 10300
rect 24136 9846 24348 9874
rect 24136 9840 24164 9846
rect 23938 9823 23994 9832
rect 23662 9344 23718 9353
rect 23662 9279 23718 9288
rect 23664 8900 23716 8906
rect 23664 8842 23716 8848
rect 23572 8492 23624 8498
rect 23572 8434 23624 8440
rect 23492 8350 23612 8378
rect 23202 8327 23258 8336
rect 23216 7886 23244 8327
rect 23388 8288 23440 8294
rect 23388 8230 23440 8236
rect 23480 8288 23532 8294
rect 23480 8230 23532 8236
rect 23204 7880 23256 7886
rect 23204 7822 23256 7828
rect 23400 7750 23428 8230
rect 23492 8129 23520 8230
rect 23478 8120 23534 8129
rect 23478 8055 23534 8064
rect 23388 7744 23440 7750
rect 23388 7686 23440 7692
rect 23166 7644 23474 7653
rect 23166 7642 23172 7644
rect 23228 7642 23252 7644
rect 23308 7642 23332 7644
rect 23388 7642 23412 7644
rect 23468 7642 23474 7644
rect 23228 7590 23230 7642
rect 23410 7590 23412 7642
rect 23166 7588 23172 7590
rect 23228 7588 23252 7590
rect 23308 7588 23332 7590
rect 23388 7588 23412 7590
rect 23468 7588 23474 7590
rect 23166 7579 23474 7588
rect 23112 7540 23164 7546
rect 23584 7528 23612 8350
rect 23676 7886 23704 8842
rect 23756 8832 23808 8838
rect 23756 8774 23808 8780
rect 23768 8498 23796 8774
rect 23846 8664 23902 8673
rect 23846 8599 23902 8608
rect 23756 8492 23808 8498
rect 23756 8434 23808 8440
rect 23860 8362 23888 8599
rect 23952 8362 23980 9823
rect 24044 9812 24164 9840
rect 24124 9716 24176 9722
rect 24124 9658 24176 9664
rect 24032 9444 24084 9450
rect 24032 9386 24084 9392
rect 23848 8356 23900 8362
rect 23848 8298 23900 8304
rect 23940 8356 23992 8362
rect 23940 8298 23992 8304
rect 23938 8120 23994 8129
rect 23938 8055 23994 8064
rect 23952 7886 23980 8055
rect 23664 7880 23716 7886
rect 23664 7822 23716 7828
rect 23940 7880 23992 7886
rect 23940 7822 23992 7828
rect 23112 7482 23164 7488
rect 23400 7500 23612 7528
rect 22926 7375 22928 7384
rect 22980 7375 22982 7384
rect 23020 7404 23072 7410
rect 22928 7346 22980 7352
rect 23020 7346 23072 7352
rect 23124 6662 23152 7482
rect 23400 7410 23428 7500
rect 23388 7404 23440 7410
rect 23388 7346 23440 7352
rect 23204 7200 23256 7206
rect 23202 7168 23204 7177
rect 23848 7200 23900 7206
rect 23256 7168 23258 7177
rect 24044 7188 24072 9386
rect 24136 7206 24164 9658
rect 24320 9466 24348 9846
rect 24398 9840 24454 10300
rect 24504 9846 24716 9874
rect 24504 9840 24532 9846
rect 24412 9812 24532 9840
rect 24320 9438 24440 9466
rect 24306 9344 24362 9353
rect 24306 9279 24362 9288
rect 24320 8498 24348 9279
rect 24412 8566 24440 9438
rect 24400 8560 24452 8566
rect 24400 8502 24452 8508
rect 24490 8528 24546 8537
rect 24308 8492 24360 8498
rect 24688 8498 24716 9846
rect 24766 9840 24822 10300
rect 25134 9840 25190 10300
rect 25240 9846 25452 9874
rect 25240 9840 25268 9846
rect 24780 9194 24808 9840
rect 25148 9812 25268 9840
rect 24780 9166 24900 9194
rect 24872 8566 24900 9166
rect 25226 8936 25282 8945
rect 25226 8871 25282 8880
rect 24860 8560 24912 8566
rect 24860 8502 24912 8508
rect 24490 8463 24546 8472
rect 24676 8492 24728 8498
rect 24308 8434 24360 8440
rect 24504 8430 24532 8463
rect 24676 8434 24728 8440
rect 24492 8424 24544 8430
rect 24492 8366 24544 8372
rect 24308 8288 24360 8294
rect 24308 8230 24360 8236
rect 24492 8288 24544 8294
rect 24768 8288 24820 8294
rect 24492 8230 24544 8236
rect 24582 8256 24638 8265
rect 24320 8090 24348 8230
rect 24308 8084 24360 8090
rect 24308 8026 24360 8032
rect 24216 7744 24268 7750
rect 24216 7686 24268 7692
rect 24308 7744 24360 7750
rect 24308 7686 24360 7692
rect 24228 7546 24256 7686
rect 24216 7540 24268 7546
rect 24216 7482 24268 7488
rect 24320 7206 24348 7686
rect 24504 7546 24532 8230
rect 24768 8230 24820 8236
rect 25044 8288 25096 8294
rect 25044 8230 25096 8236
rect 25136 8288 25188 8294
rect 25136 8230 25188 8236
rect 24582 8191 24638 8200
rect 24596 8090 24624 8191
rect 24780 8129 24808 8230
rect 24766 8120 24822 8129
rect 24584 8084 24636 8090
rect 25056 8090 25084 8230
rect 24766 8055 24822 8064
rect 25044 8084 25096 8090
rect 24584 8026 24636 8032
rect 25044 8026 25096 8032
rect 25148 7886 25176 8230
rect 25240 8090 25268 8871
rect 25424 8480 25452 9846
rect 25502 9840 25558 10300
rect 25608 9846 25820 9874
rect 25608 9840 25636 9846
rect 25516 9812 25636 9840
rect 25792 8498 25820 9846
rect 25870 9840 25926 10300
rect 25976 9846 26188 9874
rect 25976 9840 26004 9846
rect 25884 9812 26004 9840
rect 26160 8498 26188 9846
rect 26238 9840 26294 10300
rect 26344 9846 26556 9874
rect 26344 9840 26372 9846
rect 26252 9812 26372 9840
rect 26240 9376 26292 9382
rect 26240 9318 26292 9324
rect 26332 9376 26384 9382
rect 26332 9318 26384 9324
rect 25504 8492 25556 8498
rect 25424 8452 25504 8480
rect 25504 8434 25556 8440
rect 25780 8492 25832 8498
rect 25780 8434 25832 8440
rect 26148 8492 26200 8498
rect 26148 8434 26200 8440
rect 25872 8356 25924 8362
rect 25872 8298 25924 8304
rect 25412 8288 25464 8294
rect 25412 8230 25464 8236
rect 25688 8288 25740 8294
rect 25688 8230 25740 8236
rect 25228 8084 25280 8090
rect 25228 8026 25280 8032
rect 25424 7886 25452 8230
rect 25700 7886 25728 8230
rect 25884 7886 25912 8298
rect 26148 8288 26200 8294
rect 26148 8230 26200 8236
rect 26160 7886 26188 8230
rect 26252 8022 26280 9318
rect 26240 8016 26292 8022
rect 26240 7958 26292 7964
rect 25136 7880 25188 7886
rect 25136 7822 25188 7828
rect 25412 7880 25464 7886
rect 25412 7822 25464 7828
rect 25688 7880 25740 7886
rect 25688 7822 25740 7828
rect 25872 7880 25924 7886
rect 25872 7822 25924 7828
rect 26148 7880 26200 7886
rect 26148 7822 26200 7828
rect 25044 7744 25096 7750
rect 25044 7686 25096 7692
rect 25136 7744 25188 7750
rect 25136 7686 25188 7692
rect 25412 7744 25464 7750
rect 25412 7686 25464 7692
rect 25688 7744 25740 7750
rect 25688 7686 25740 7692
rect 25964 7744 26016 7750
rect 25964 7686 26016 7692
rect 26240 7744 26292 7750
rect 26240 7686 26292 7692
rect 24492 7540 24544 7546
rect 24492 7482 24544 7488
rect 25056 7478 25084 7686
rect 25044 7472 25096 7478
rect 25044 7414 25096 7420
rect 23900 7160 24072 7188
rect 24124 7200 24176 7206
rect 23848 7142 23900 7148
rect 24124 7142 24176 7148
rect 24216 7200 24268 7206
rect 24216 7142 24268 7148
rect 24308 7200 24360 7206
rect 24308 7142 24360 7148
rect 23202 7103 23258 7112
rect 24228 6798 24256 7142
rect 24216 6792 24268 6798
rect 24216 6734 24268 6740
rect 23112 6656 23164 6662
rect 23112 6598 23164 6604
rect 23166 6556 23474 6565
rect 23166 6554 23172 6556
rect 23228 6554 23252 6556
rect 23308 6554 23332 6556
rect 23388 6554 23412 6556
rect 23468 6554 23474 6556
rect 23228 6502 23230 6554
rect 23410 6502 23412 6554
rect 23166 6500 23172 6502
rect 23228 6500 23252 6502
rect 23308 6500 23332 6502
rect 23388 6500 23412 6502
rect 23468 6500 23474 6502
rect 23166 6491 23474 6500
rect 25148 6458 25176 7686
rect 25136 6452 25188 6458
rect 25136 6394 25188 6400
rect 22836 6384 22888 6390
rect 22836 6326 22888 6332
rect 24860 6384 24912 6390
rect 24860 6326 24912 6332
rect 18512 6316 18564 6322
rect 18512 6258 18564 6264
rect 24216 6316 24268 6322
rect 24216 6258 24268 6264
rect 2964 6248 3016 6254
rect 2964 6190 3016 6196
rect 14464 6248 14516 6254
rect 14464 6190 14516 6196
rect 6504 6012 6812 6021
rect 6504 6010 6510 6012
rect 6566 6010 6590 6012
rect 6646 6010 6670 6012
rect 6726 6010 6750 6012
rect 6806 6010 6812 6012
rect 6566 5958 6568 6010
rect 6748 5958 6750 6010
rect 6504 5956 6510 5958
rect 6566 5956 6590 5958
rect 6646 5956 6670 5958
rect 6726 5956 6750 5958
rect 6806 5956 6812 5958
rect 6504 5947 6812 5956
rect 17612 6012 17920 6021
rect 17612 6010 17618 6012
rect 17674 6010 17698 6012
rect 17754 6010 17778 6012
rect 17834 6010 17858 6012
rect 17914 6010 17920 6012
rect 17674 5958 17676 6010
rect 17856 5958 17858 6010
rect 17612 5956 17618 5958
rect 17674 5956 17698 5958
rect 17754 5956 17778 5958
rect 17834 5956 17858 5958
rect 17914 5956 17920 5958
rect 17612 5947 17920 5956
rect 12058 5468 12366 5477
rect 12058 5466 12064 5468
rect 12120 5466 12144 5468
rect 12200 5466 12224 5468
rect 12280 5466 12304 5468
rect 12360 5466 12366 5468
rect 12120 5414 12122 5466
rect 12302 5414 12304 5466
rect 12058 5412 12064 5414
rect 12120 5412 12144 5414
rect 12200 5412 12224 5414
rect 12280 5412 12304 5414
rect 12360 5412 12366 5414
rect 12058 5403 12366 5412
rect 23166 5468 23474 5477
rect 23166 5466 23172 5468
rect 23228 5466 23252 5468
rect 23308 5466 23332 5468
rect 23388 5466 23412 5468
rect 23468 5466 23474 5468
rect 23228 5414 23230 5466
rect 23410 5414 23412 5466
rect 23166 5412 23172 5414
rect 23228 5412 23252 5414
rect 23308 5412 23332 5414
rect 23388 5412 23412 5414
rect 23468 5412 23474 5414
rect 23166 5403 23474 5412
rect 23020 5160 23072 5166
rect 23020 5102 23072 5108
rect 22836 5092 22888 5098
rect 22836 5034 22888 5040
rect 20536 5024 20588 5030
rect 20536 4966 20588 4972
rect 6504 4924 6812 4933
rect 6504 4922 6510 4924
rect 6566 4922 6590 4924
rect 6646 4922 6670 4924
rect 6726 4922 6750 4924
rect 6806 4922 6812 4924
rect 6566 4870 6568 4922
rect 6748 4870 6750 4922
rect 6504 4868 6510 4870
rect 6566 4868 6590 4870
rect 6646 4868 6670 4870
rect 6726 4868 6750 4870
rect 6806 4868 6812 4870
rect 6504 4859 6812 4868
rect 17612 4924 17920 4933
rect 17612 4922 17618 4924
rect 17674 4922 17698 4924
rect 17754 4922 17778 4924
rect 17834 4922 17858 4924
rect 17914 4922 17920 4924
rect 17674 4870 17676 4922
rect 17856 4870 17858 4922
rect 17612 4868 17618 4870
rect 17674 4868 17698 4870
rect 17754 4868 17778 4870
rect 17834 4868 17858 4870
rect 17914 4868 17920 4870
rect 17612 4859 17920 4868
rect 12058 4380 12366 4389
rect 12058 4378 12064 4380
rect 12120 4378 12144 4380
rect 12200 4378 12224 4380
rect 12280 4378 12304 4380
rect 12360 4378 12366 4380
rect 12120 4326 12122 4378
rect 12302 4326 12304 4378
rect 12058 4324 12064 4326
rect 12120 4324 12144 4326
rect 12200 4324 12224 4326
rect 12280 4324 12304 4326
rect 12360 4324 12366 4326
rect 12058 4315 12366 4324
rect 6504 3836 6812 3845
rect 6504 3834 6510 3836
rect 6566 3834 6590 3836
rect 6646 3834 6670 3836
rect 6726 3834 6750 3836
rect 6806 3834 6812 3836
rect 6566 3782 6568 3834
rect 6748 3782 6750 3834
rect 6504 3780 6510 3782
rect 6566 3780 6590 3782
rect 6646 3780 6670 3782
rect 6726 3780 6750 3782
rect 6806 3780 6812 3782
rect 6504 3771 6812 3780
rect 17612 3836 17920 3845
rect 17612 3834 17618 3836
rect 17674 3834 17698 3836
rect 17754 3834 17778 3836
rect 17834 3834 17858 3836
rect 17914 3834 17920 3836
rect 17674 3782 17676 3834
rect 17856 3782 17858 3834
rect 17612 3780 17618 3782
rect 17674 3780 17698 3782
rect 17754 3780 17778 3782
rect 17834 3780 17858 3782
rect 17914 3780 17920 3782
rect 17612 3771 17920 3780
rect 12058 3292 12366 3301
rect 12058 3290 12064 3292
rect 12120 3290 12144 3292
rect 12200 3290 12224 3292
rect 12280 3290 12304 3292
rect 12360 3290 12366 3292
rect 12120 3238 12122 3290
rect 12302 3238 12304 3290
rect 12058 3236 12064 3238
rect 12120 3236 12144 3238
rect 12200 3236 12224 3238
rect 12280 3236 12304 3238
rect 12360 3236 12366 3238
rect 12058 3227 12366 3236
rect 6504 2748 6812 2757
rect 6504 2746 6510 2748
rect 6566 2746 6590 2748
rect 6646 2746 6670 2748
rect 6726 2746 6750 2748
rect 6806 2746 6812 2748
rect 6566 2694 6568 2746
rect 6748 2694 6750 2746
rect 6504 2692 6510 2694
rect 6566 2692 6590 2694
rect 6646 2692 6670 2694
rect 6726 2692 6750 2694
rect 6806 2692 6812 2694
rect 6504 2683 6812 2692
rect 17612 2748 17920 2757
rect 17612 2746 17618 2748
rect 17674 2746 17698 2748
rect 17754 2746 17778 2748
rect 17834 2746 17858 2748
rect 17914 2746 17920 2748
rect 17674 2694 17676 2746
rect 17856 2694 17858 2746
rect 17612 2692 17618 2694
rect 17674 2692 17698 2694
rect 17754 2692 17778 2694
rect 17834 2692 17858 2694
rect 17914 2692 17920 2694
rect 17612 2683 17920 2692
rect 20548 2650 20576 4966
rect 22744 3596 22796 3602
rect 22744 3538 22796 3544
rect 20628 3460 20680 3466
rect 20628 3402 20680 3408
rect 20536 2644 20588 2650
rect 20536 2586 20588 2592
rect 20352 2372 20404 2378
rect 20352 2314 20404 2320
rect 12058 2204 12366 2213
rect 12058 2202 12064 2204
rect 12120 2202 12144 2204
rect 12200 2202 12224 2204
rect 12280 2202 12304 2204
rect 12360 2202 12366 2204
rect 12120 2150 12122 2202
rect 12302 2150 12304 2202
rect 12058 2148 12064 2150
rect 12120 2148 12144 2150
rect 12200 2148 12224 2150
rect 12280 2148 12304 2150
rect 12360 2148 12366 2150
rect 12058 2139 12366 2148
rect 20364 2106 20392 2314
rect 20640 2106 20668 3402
rect 22284 2508 22336 2514
rect 22284 2450 22336 2456
rect 22192 2440 22244 2446
rect 22192 2382 22244 2388
rect 21456 2372 21508 2378
rect 21456 2314 21508 2320
rect 20352 2100 20404 2106
rect 20352 2042 20404 2048
rect 20628 2100 20680 2106
rect 20628 2042 20680 2048
rect 1584 1964 1636 1970
rect 1584 1906 1636 1912
rect 19616 1964 19668 1970
rect 19616 1906 19668 1912
rect 20720 1964 20772 1970
rect 20720 1906 20772 1912
rect 1596 1562 1624 1906
rect 6504 1660 6812 1669
rect 6504 1658 6510 1660
rect 6566 1658 6590 1660
rect 6646 1658 6670 1660
rect 6726 1658 6750 1660
rect 6806 1658 6812 1660
rect 6566 1606 6568 1658
rect 6748 1606 6750 1658
rect 6504 1604 6510 1606
rect 6566 1604 6590 1606
rect 6646 1604 6670 1606
rect 6726 1604 6750 1606
rect 6806 1604 6812 1606
rect 6504 1595 6812 1604
rect 17612 1660 17920 1669
rect 17612 1658 17618 1660
rect 17674 1658 17698 1660
rect 17754 1658 17778 1660
rect 17834 1658 17858 1660
rect 17914 1658 17920 1660
rect 17674 1606 17676 1658
rect 17856 1606 17858 1658
rect 17612 1604 17618 1606
rect 17674 1604 17698 1606
rect 17754 1604 17778 1606
rect 17834 1604 17858 1606
rect 17914 1604 17920 1606
rect 17612 1595 17920 1604
rect 19628 1562 19656 1906
rect 1584 1556 1636 1562
rect 1584 1498 1636 1504
rect 19616 1556 19668 1562
rect 19616 1498 19668 1504
rect 1216 1352 1268 1358
rect 1216 1294 1268 1300
rect 3792 1352 3844 1358
rect 3792 1294 3844 1300
rect 5724 1352 5776 1358
rect 5724 1294 5776 1300
rect 7932 1352 7984 1358
rect 7932 1294 7984 1300
rect 10140 1352 10192 1358
rect 12072 1352 12124 1358
rect 10140 1294 10192 1300
rect 11992 1312 12072 1340
rect 1228 160 1256 1294
rect 1214 -300 1270 160
rect 3422 82 3478 160
rect 3804 82 3832 1294
rect 3976 1216 4028 1222
rect 3976 1158 4028 1164
rect 3988 1018 4016 1158
rect 3976 1012 4028 1018
rect 3976 954 4028 960
rect 3422 54 3832 82
rect 5630 82 5686 160
rect 5736 82 5764 1294
rect 5630 54 5764 82
rect 7838 82 7894 160
rect 7944 82 7972 1294
rect 8116 1216 8168 1222
rect 8116 1158 8168 1164
rect 8128 814 8156 1158
rect 8116 808 8168 814
rect 8116 750 8168 756
rect 7838 54 7972 82
rect 10046 82 10102 160
rect 10152 82 10180 1294
rect 10324 1216 10376 1222
rect 10324 1158 10376 1164
rect 10336 814 10364 1158
rect 10324 808 10376 814
rect 10324 750 10376 756
rect 10046 54 10180 82
rect 11992 82 12020 1312
rect 12072 1294 12124 1300
rect 14740 1352 14792 1358
rect 14740 1294 14792 1300
rect 16948 1352 17000 1358
rect 19432 1352 19484 1358
rect 16948 1294 17000 1300
rect 19352 1312 19432 1340
rect 14648 1284 14700 1290
rect 14648 1226 14700 1232
rect 14556 1216 14608 1222
rect 14556 1158 14608 1164
rect 12058 1116 12366 1125
rect 12058 1114 12064 1116
rect 12120 1114 12144 1116
rect 12200 1114 12224 1116
rect 12280 1114 12304 1116
rect 12360 1114 12366 1116
rect 12120 1062 12122 1114
rect 12302 1062 12304 1114
rect 12058 1060 12064 1062
rect 12120 1060 12144 1062
rect 12200 1060 12224 1062
rect 12280 1060 12304 1062
rect 12360 1060 12366 1062
rect 12058 1051 12366 1060
rect 14568 1018 14596 1158
rect 14660 1018 14688 1226
rect 14556 1012 14608 1018
rect 14556 954 14608 960
rect 14648 1012 14700 1018
rect 14648 954 14700 960
rect 12254 82 12310 160
rect 11992 54 12310 82
rect 3422 -300 3478 54
rect 5630 -300 5686 54
rect 7838 -300 7894 54
rect 10046 -300 10102 54
rect 12254 -300 12310 54
rect 14462 82 14518 160
rect 14752 82 14780 1294
rect 14462 54 14780 82
rect 16670 82 16726 160
rect 16960 82 16988 1294
rect 16670 54 16988 82
rect 18878 82 18934 160
rect 19352 82 19380 1312
rect 19432 1294 19484 1300
rect 20732 1290 20760 1906
rect 20812 1896 20864 1902
rect 20812 1838 20864 1844
rect 20720 1284 20772 1290
rect 20720 1226 20772 1232
rect 20824 1018 20852 1838
rect 21468 1766 21496 2314
rect 22204 2106 22232 2382
rect 22296 2106 22324 2450
rect 22468 2440 22520 2446
rect 22468 2382 22520 2388
rect 22192 2100 22244 2106
rect 22192 2042 22244 2048
rect 22284 2100 22336 2106
rect 22284 2042 22336 2048
rect 21640 1964 21692 1970
rect 21640 1906 21692 1912
rect 22192 1964 22244 1970
rect 22192 1906 22244 1912
rect 21456 1760 21508 1766
rect 21456 1702 21508 1708
rect 21548 1760 21600 1766
rect 21548 1702 21600 1708
rect 21364 1352 21416 1358
rect 21364 1294 21416 1300
rect 20812 1012 20864 1018
rect 20812 954 20864 960
rect 18878 54 19380 82
rect 21086 82 21142 160
rect 21376 82 21404 1294
rect 21560 678 21588 1702
rect 21652 1562 21680 1906
rect 21640 1556 21692 1562
rect 21640 1498 21692 1504
rect 22204 1290 22232 1906
rect 22480 1834 22508 2382
rect 22468 1828 22520 1834
rect 22468 1770 22520 1776
rect 22756 1766 22784 3538
rect 22848 2378 22876 5034
rect 23032 2650 23060 5102
rect 23166 4380 23474 4389
rect 23166 4378 23172 4380
rect 23228 4378 23252 4380
rect 23308 4378 23332 4380
rect 23388 4378 23412 4380
rect 23468 4378 23474 4380
rect 23228 4326 23230 4378
rect 23410 4326 23412 4378
rect 23166 4324 23172 4326
rect 23228 4324 23252 4326
rect 23308 4324 23332 4326
rect 23388 4324 23412 4326
rect 23468 4324 23474 4326
rect 23166 4315 23474 4324
rect 23664 3664 23716 3670
rect 23664 3606 23716 3612
rect 23166 3292 23474 3301
rect 23166 3290 23172 3292
rect 23228 3290 23252 3292
rect 23308 3290 23332 3292
rect 23388 3290 23412 3292
rect 23468 3290 23474 3292
rect 23228 3238 23230 3290
rect 23410 3238 23412 3290
rect 23166 3236 23172 3238
rect 23228 3236 23252 3238
rect 23308 3236 23332 3238
rect 23388 3236 23412 3238
rect 23468 3236 23474 3238
rect 23166 3227 23474 3236
rect 23676 2650 23704 3606
rect 23940 3528 23992 3534
rect 23940 3470 23992 3476
rect 23952 2650 23980 3470
rect 24228 2650 24256 6258
rect 24872 2650 24900 6326
rect 25424 6186 25452 7686
rect 25700 6254 25728 7686
rect 25976 6769 26004 7686
rect 26252 6905 26280 7686
rect 26238 6896 26294 6905
rect 26344 6866 26372 9318
rect 26528 8498 26556 9846
rect 26606 9840 26662 10300
rect 26974 9840 27030 10300
rect 27342 9840 27398 10300
rect 27448 9846 27568 9874
rect 27448 9840 27476 9846
rect 26620 8498 26648 9840
rect 26988 8566 27016 9840
rect 27356 9812 27476 9840
rect 27436 9512 27488 9518
rect 27436 9454 27488 9460
rect 27448 9246 27476 9454
rect 27436 9240 27488 9246
rect 27436 9182 27488 9188
rect 27252 8968 27304 8974
rect 27252 8910 27304 8916
rect 26976 8560 27028 8566
rect 26976 8502 27028 8508
rect 26516 8492 26568 8498
rect 26516 8434 26568 8440
rect 26608 8492 26660 8498
rect 26608 8434 26660 8440
rect 26608 8288 26660 8294
rect 26608 8230 26660 8236
rect 26620 7886 26648 8230
rect 26608 7880 26660 7886
rect 26608 7822 26660 7828
rect 26884 7744 26936 7750
rect 26884 7686 26936 7692
rect 26896 7274 26924 7686
rect 26884 7268 26936 7274
rect 26884 7210 26936 7216
rect 27264 6934 27292 8910
rect 27540 8498 27568 9846
rect 27710 9840 27766 10300
rect 27816 9846 28028 9874
rect 27816 9840 27844 9846
rect 27724 9812 27844 9840
rect 27618 9480 27674 9489
rect 27674 9438 27752 9466
rect 27618 9415 27674 9424
rect 27528 8492 27580 8498
rect 27528 8434 27580 8440
rect 27620 8356 27672 8362
rect 27620 8298 27672 8304
rect 27528 8288 27580 8294
rect 27528 8230 27580 8236
rect 27540 8090 27568 8230
rect 27528 8084 27580 8090
rect 27528 8026 27580 8032
rect 27632 7886 27660 8298
rect 27724 8090 27752 9438
rect 27896 9240 27948 9246
rect 27896 9182 27948 9188
rect 27804 8288 27856 8294
rect 27804 8230 27856 8236
rect 27816 8090 27844 8230
rect 27908 8090 27936 9182
rect 28000 8498 28028 9846
rect 28078 9840 28134 10300
rect 28184 9846 28396 9874
rect 28184 9840 28212 9846
rect 28092 9812 28212 9840
rect 28262 8664 28318 8673
rect 28262 8599 28318 8608
rect 27988 8492 28040 8498
rect 27988 8434 28040 8440
rect 28276 8362 28304 8599
rect 28368 8498 28396 9846
rect 28446 9840 28502 10300
rect 28552 9846 28764 9874
rect 28552 9840 28580 9846
rect 28460 9812 28580 9840
rect 28540 9716 28592 9722
rect 28540 9658 28592 9664
rect 28446 9208 28502 9217
rect 28446 9143 28502 9152
rect 28356 8492 28408 8498
rect 28356 8434 28408 8440
rect 28264 8356 28316 8362
rect 28264 8298 28316 8304
rect 27712 8084 27764 8090
rect 27712 8026 27764 8032
rect 27804 8084 27856 8090
rect 27804 8026 27856 8032
rect 27896 8084 27948 8090
rect 27896 8026 27948 8032
rect 27620 7880 27672 7886
rect 27620 7822 27672 7828
rect 28170 7848 28226 7857
rect 28460 7834 28488 9143
rect 28552 8401 28580 9658
rect 28736 8498 28764 9846
rect 28814 9840 28870 10300
rect 28908 9852 28960 9858
rect 28828 8498 28856 9840
rect 29182 9840 29238 10300
rect 29550 9840 29606 10300
rect 29918 9840 29974 10300
rect 30024 9846 30236 9874
rect 30024 9840 30052 9846
rect 28908 9794 28960 9800
rect 28920 9314 28948 9794
rect 28908 9308 28960 9314
rect 28908 9250 28960 9256
rect 29196 8498 29224 9840
rect 29564 8566 29592 9840
rect 29932 9812 30052 9840
rect 29552 8560 29604 8566
rect 29552 8502 29604 8508
rect 28724 8492 28776 8498
rect 28724 8434 28776 8440
rect 28816 8492 28868 8498
rect 28816 8434 28868 8440
rect 29184 8492 29236 8498
rect 30208 8480 30236 9846
rect 30286 9840 30342 10300
rect 30654 9840 30710 10300
rect 30760 9846 30972 9874
rect 30760 9840 30788 9846
rect 30300 8634 30328 9840
rect 30668 9812 30788 9840
rect 30288 8628 30340 8634
rect 30288 8570 30340 8576
rect 30656 8560 30708 8566
rect 30392 8520 30656 8548
rect 30288 8492 30340 8498
rect 30208 8452 30288 8480
rect 29184 8434 29236 8440
rect 30288 8434 30340 8440
rect 30392 8430 30420 8520
rect 30656 8502 30708 8508
rect 30944 8498 30972 9846
rect 31022 9840 31078 10300
rect 31128 9846 31340 9874
rect 31128 9840 31156 9846
rect 31036 9812 31156 9840
rect 31312 8498 31340 9846
rect 31390 9840 31446 10300
rect 31496 9846 31708 9874
rect 31496 9840 31524 9846
rect 31404 9812 31524 9840
rect 31484 8900 31536 8906
rect 31484 8842 31536 8848
rect 31496 8634 31524 8842
rect 31484 8628 31536 8634
rect 31484 8570 31536 8576
rect 31680 8498 31708 9846
rect 31758 9840 31814 10300
rect 32126 9840 32182 10300
rect 32494 9840 32550 10300
rect 32600 9846 32720 9874
rect 32600 9840 32628 9846
rect 31772 8498 31800 9840
rect 30932 8492 30984 8498
rect 30932 8434 30984 8440
rect 31300 8492 31352 8498
rect 31300 8434 31352 8440
rect 31668 8492 31720 8498
rect 31668 8434 31720 8440
rect 31760 8492 31812 8498
rect 32140 8480 32168 9840
rect 32508 9812 32628 9840
rect 32312 9716 32364 9722
rect 32312 9658 32364 9664
rect 32324 8634 32352 9658
rect 32404 8832 32456 8838
rect 32404 8774 32456 8780
rect 32416 8634 32444 8774
rect 32312 8628 32364 8634
rect 32312 8570 32364 8576
rect 32404 8628 32456 8634
rect 32404 8570 32456 8576
rect 32496 8628 32548 8634
rect 32496 8570 32548 8576
rect 32312 8492 32364 8498
rect 32140 8452 32312 8480
rect 31760 8434 31812 8440
rect 32312 8434 32364 8440
rect 30380 8424 30432 8430
rect 28538 8392 28594 8401
rect 30380 8366 30432 8372
rect 32508 8362 32536 8570
rect 32692 8498 32720 9846
rect 32862 9840 32918 10300
rect 32968 9846 33088 9874
rect 32968 9840 32996 9846
rect 32876 9812 32996 9840
rect 32772 9240 32824 9246
rect 32772 9182 32824 9188
rect 32680 8492 32732 8498
rect 32680 8434 32732 8440
rect 28538 8327 28594 8336
rect 32496 8356 32548 8362
rect 32496 8298 32548 8304
rect 28540 8288 28592 8294
rect 28540 8230 28592 8236
rect 28632 8288 28684 8294
rect 28632 8230 28684 8236
rect 29552 8288 29604 8294
rect 29552 8230 29604 8236
rect 29828 8288 29880 8294
rect 29828 8230 29880 8236
rect 30104 8288 30156 8294
rect 30104 8230 30156 8236
rect 30380 8288 30432 8294
rect 30380 8230 30432 8236
rect 30748 8288 30800 8294
rect 30748 8230 30800 8236
rect 31116 8288 31168 8294
rect 31116 8230 31168 8236
rect 28552 8090 28580 8230
rect 28644 8090 28672 8230
rect 28720 8188 29028 8197
rect 28720 8186 28726 8188
rect 28782 8186 28806 8188
rect 28862 8186 28886 8188
rect 28942 8186 28966 8188
rect 29022 8186 29028 8188
rect 28782 8134 28784 8186
rect 28964 8134 28966 8186
rect 28720 8132 28726 8134
rect 28782 8132 28806 8134
rect 28862 8132 28886 8134
rect 28942 8132 28966 8134
rect 29022 8132 29028 8134
rect 28720 8123 29028 8132
rect 28540 8084 28592 8090
rect 28540 8026 28592 8032
rect 28632 8084 28684 8090
rect 28632 8026 28684 8032
rect 29564 7886 29592 8230
rect 29840 7886 29868 8230
rect 29552 7880 29604 7886
rect 28460 7806 28580 7834
rect 29552 7822 29604 7828
rect 29828 7880 29880 7886
rect 29828 7822 29880 7828
rect 28170 7783 28226 7792
rect 28184 7750 28212 7783
rect 28552 7750 28580 7806
rect 27344 7744 27396 7750
rect 27344 7686 27396 7692
rect 28172 7744 28224 7750
rect 28172 7686 28224 7692
rect 28448 7744 28500 7750
rect 28448 7686 28500 7692
rect 28540 7744 28592 7750
rect 28540 7686 28592 7692
rect 27356 7546 27384 7686
rect 27344 7540 27396 7546
rect 27344 7482 27396 7488
rect 28460 7041 28488 7686
rect 30116 7546 30144 8230
rect 30392 7546 30420 8230
rect 30760 7546 30788 8230
rect 30104 7540 30156 7546
rect 30104 7482 30156 7488
rect 30380 7540 30432 7546
rect 30380 7482 30432 7488
rect 30748 7540 30800 7546
rect 30748 7482 30800 7488
rect 31128 7342 31156 8230
rect 31116 7336 31168 7342
rect 31116 7278 31168 7284
rect 28720 7100 29028 7109
rect 28720 7098 28726 7100
rect 28782 7098 28806 7100
rect 28862 7098 28886 7100
rect 28942 7098 28966 7100
rect 29022 7098 29028 7100
rect 28782 7046 28784 7098
rect 28964 7046 28966 7098
rect 28720 7044 28726 7046
rect 28782 7044 28806 7046
rect 28862 7044 28886 7046
rect 28942 7044 28966 7046
rect 29022 7044 29028 7046
rect 28446 7032 28502 7041
rect 28720 7035 29028 7044
rect 28446 6967 28502 6976
rect 27252 6928 27304 6934
rect 27252 6870 27304 6876
rect 26238 6831 26294 6840
rect 26332 6860 26384 6866
rect 26332 6802 26384 6808
rect 25962 6760 26018 6769
rect 25962 6695 26018 6704
rect 32784 6390 32812 9182
rect 33060 8430 33088 9846
rect 33230 9840 33286 10300
rect 33598 9840 33654 10300
rect 33966 9840 34022 10300
rect 34164 9846 34284 9874
rect 33244 8480 33272 9840
rect 33508 9376 33560 9382
rect 33508 9318 33560 9324
rect 33416 8968 33468 8974
rect 33416 8910 33468 8916
rect 33324 8492 33376 8498
rect 33244 8452 33324 8480
rect 33324 8434 33376 8440
rect 33048 8424 33100 8430
rect 33048 8366 33100 8372
rect 33428 8362 33456 8910
rect 33520 8634 33548 9318
rect 33508 8628 33560 8634
rect 33508 8570 33560 8576
rect 33612 8480 33640 9840
rect 33784 9376 33836 9382
rect 33784 9318 33836 9324
rect 33692 8492 33744 8498
rect 33612 8452 33692 8480
rect 33692 8434 33744 8440
rect 33416 8356 33468 8362
rect 33416 8298 33468 8304
rect 33048 8288 33100 8294
rect 33048 8230 33100 8236
rect 33060 7970 33088 8230
rect 32968 7942 33088 7970
rect 32968 7313 32996 7942
rect 33048 7880 33100 7886
rect 33048 7822 33100 7828
rect 32954 7304 33010 7313
rect 32954 7239 33010 7248
rect 32772 6384 32824 6390
rect 32772 6326 32824 6332
rect 25688 6248 25740 6254
rect 25688 6190 25740 6196
rect 27068 6248 27120 6254
rect 27068 6190 27120 6196
rect 25412 6180 25464 6186
rect 25412 6122 25464 6128
rect 25504 6180 25556 6186
rect 25504 6122 25556 6128
rect 22928 2644 22980 2650
rect 22928 2586 22980 2592
rect 23020 2644 23072 2650
rect 23020 2586 23072 2592
rect 23664 2644 23716 2650
rect 23664 2586 23716 2592
rect 23940 2644 23992 2650
rect 23940 2586 23992 2592
rect 24216 2644 24268 2650
rect 24216 2586 24268 2592
rect 24860 2644 24912 2650
rect 24860 2586 24912 2592
rect 22940 2530 22968 2586
rect 22940 2514 23336 2530
rect 25516 2514 25544 6122
rect 27080 2650 27108 6190
rect 28720 6012 29028 6021
rect 28720 6010 28726 6012
rect 28782 6010 28806 6012
rect 28862 6010 28886 6012
rect 28942 6010 28966 6012
rect 29022 6010 29028 6012
rect 28782 5958 28784 6010
rect 28964 5958 28966 6010
rect 28720 5956 28726 5958
rect 28782 5956 28806 5958
rect 28862 5956 28886 5958
rect 28942 5956 28966 5958
rect 29022 5956 29028 5958
rect 28720 5947 29028 5956
rect 33060 5166 33088 7822
rect 33048 5160 33100 5166
rect 33048 5102 33100 5108
rect 33796 5030 33824 9318
rect 33876 8968 33928 8974
rect 33876 8910 33928 8916
rect 33784 5024 33836 5030
rect 33784 4966 33836 4972
rect 28720 4924 29028 4933
rect 28720 4922 28726 4924
rect 28782 4922 28806 4924
rect 28862 4922 28886 4924
rect 28942 4922 28966 4924
rect 29022 4922 29028 4924
rect 28782 4870 28784 4922
rect 28964 4870 28966 4922
rect 28720 4868 28726 4870
rect 28782 4868 28806 4870
rect 28862 4868 28886 4870
rect 28942 4868 28966 4870
rect 29022 4868 29028 4870
rect 28720 4859 29028 4868
rect 29276 4820 29328 4826
rect 29276 4762 29328 4768
rect 28720 3836 29028 3845
rect 28720 3834 28726 3836
rect 28782 3834 28806 3836
rect 28862 3834 28886 3836
rect 28942 3834 28966 3836
rect 29022 3834 29028 3836
rect 28782 3782 28784 3834
rect 28964 3782 28966 3834
rect 28720 3780 28726 3782
rect 28782 3780 28806 3782
rect 28862 3780 28886 3782
rect 28942 3780 28966 3782
rect 29022 3780 29028 3782
rect 28720 3771 29028 3780
rect 28720 2748 29028 2757
rect 28720 2746 28726 2748
rect 28782 2746 28806 2748
rect 28862 2746 28886 2748
rect 28942 2746 28966 2748
rect 29022 2746 29028 2748
rect 28782 2694 28784 2746
rect 28964 2694 28966 2746
rect 28720 2692 28726 2694
rect 28782 2692 28806 2694
rect 28862 2692 28886 2694
rect 28942 2692 28966 2694
rect 29022 2692 29028 2694
rect 28720 2683 29028 2692
rect 29288 2650 29316 4762
rect 33888 3670 33916 8910
rect 33980 8480 34008 9840
rect 34060 9104 34112 9110
rect 34060 9046 34112 9052
rect 34072 8634 34100 9046
rect 34060 8628 34112 8634
rect 34060 8570 34112 8576
rect 34164 8498 34192 9846
rect 34256 9840 34284 9846
rect 34334 9840 34390 10300
rect 34702 9840 34758 10300
rect 34808 9846 35020 9874
rect 34808 9840 34836 9846
rect 34256 9812 34376 9840
rect 34716 9812 34836 9840
rect 34888 9444 34940 9450
rect 34888 9386 34940 9392
rect 34612 9172 34664 9178
rect 34612 9114 34664 9120
rect 34274 8732 34582 8741
rect 34274 8730 34280 8732
rect 34336 8730 34360 8732
rect 34416 8730 34440 8732
rect 34496 8730 34520 8732
rect 34576 8730 34582 8732
rect 34336 8678 34338 8730
rect 34518 8678 34520 8730
rect 34274 8676 34280 8678
rect 34336 8676 34360 8678
rect 34416 8676 34440 8678
rect 34496 8676 34520 8678
rect 34576 8676 34582 8678
rect 34274 8667 34582 8676
rect 34624 8634 34652 9114
rect 34794 9072 34850 9081
rect 34794 9007 34850 9016
rect 34808 8634 34836 9007
rect 34612 8628 34664 8634
rect 34612 8570 34664 8576
rect 34796 8628 34848 8634
rect 34796 8570 34848 8576
rect 34060 8492 34112 8498
rect 33980 8452 34060 8480
rect 34060 8434 34112 8440
rect 34152 8492 34204 8498
rect 34152 8434 34204 8440
rect 34900 8362 34928 9386
rect 34992 8498 35020 9846
rect 35070 9840 35126 10300
rect 35176 9846 35296 9874
rect 35176 9840 35204 9846
rect 35084 9812 35204 9840
rect 35164 9308 35216 9314
rect 35164 9250 35216 9256
rect 34980 8492 35032 8498
rect 34980 8434 35032 8440
rect 35176 8362 35204 9250
rect 35268 8498 35296 9846
rect 35438 9840 35494 10300
rect 35716 9988 35768 9994
rect 35716 9930 35768 9936
rect 35348 9308 35400 9314
rect 35348 9250 35400 9256
rect 35256 8492 35308 8498
rect 35256 8434 35308 8440
rect 34888 8356 34940 8362
rect 34888 8298 34940 8304
rect 35164 8356 35216 8362
rect 35164 8298 35216 8304
rect 34274 7644 34582 7653
rect 34274 7642 34280 7644
rect 34336 7642 34360 7644
rect 34416 7642 34440 7644
rect 34496 7642 34520 7644
rect 34576 7642 34582 7644
rect 34336 7590 34338 7642
rect 34518 7590 34520 7642
rect 34274 7588 34280 7590
rect 34336 7588 34360 7590
rect 34416 7588 34440 7590
rect 34496 7588 34520 7590
rect 34576 7588 34582 7590
rect 34274 7579 34582 7588
rect 34274 6556 34582 6565
rect 34274 6554 34280 6556
rect 34336 6554 34360 6556
rect 34416 6554 34440 6556
rect 34496 6554 34520 6556
rect 34576 6554 34582 6556
rect 34336 6502 34338 6554
rect 34518 6502 34520 6554
rect 34274 6500 34280 6502
rect 34336 6500 34360 6502
rect 34416 6500 34440 6502
rect 34496 6500 34520 6502
rect 34576 6500 34582 6502
rect 34274 6491 34582 6500
rect 34274 5468 34582 5477
rect 34274 5466 34280 5468
rect 34336 5466 34360 5468
rect 34416 5466 34440 5468
rect 34496 5466 34520 5468
rect 34576 5466 34582 5468
rect 34336 5414 34338 5466
rect 34518 5414 34520 5466
rect 34274 5412 34280 5414
rect 34336 5412 34360 5414
rect 34416 5412 34440 5414
rect 34496 5412 34520 5414
rect 34576 5412 34582 5414
rect 34274 5403 34582 5412
rect 34274 4380 34582 4389
rect 34274 4378 34280 4380
rect 34336 4378 34360 4380
rect 34416 4378 34440 4380
rect 34496 4378 34520 4380
rect 34576 4378 34582 4380
rect 34336 4326 34338 4378
rect 34518 4326 34520 4378
rect 34274 4324 34280 4326
rect 34336 4324 34360 4326
rect 34416 4324 34440 4326
rect 34496 4324 34520 4326
rect 34576 4324 34582 4326
rect 34274 4315 34582 4324
rect 33876 3664 33928 3670
rect 33876 3606 33928 3612
rect 35360 3602 35388 9250
rect 35452 8480 35480 9840
rect 35624 8900 35676 8906
rect 35624 8842 35676 8848
rect 35532 8492 35584 8498
rect 35452 8452 35532 8480
rect 35532 8434 35584 8440
rect 35636 5098 35664 8842
rect 35728 8634 35756 9930
rect 35806 9840 35862 10300
rect 36174 9840 36230 10300
rect 36542 9840 36598 10300
rect 36910 9840 36966 10300
rect 37278 9840 37334 10300
rect 37384 9846 37596 9874
rect 37384 9840 37412 9846
rect 35716 8628 35768 8634
rect 35716 8570 35768 8576
rect 35820 8498 35848 9840
rect 36084 9444 36136 9450
rect 36084 9386 36136 9392
rect 35992 8832 36044 8838
rect 35992 8774 36044 8780
rect 35900 8628 35952 8634
rect 35900 8570 35952 8576
rect 35808 8492 35860 8498
rect 35808 8434 35860 8440
rect 35912 7449 35940 8570
rect 35898 7440 35954 7449
rect 35898 7375 35954 7384
rect 36004 6322 36032 8774
rect 35992 6316 36044 6322
rect 35992 6258 36044 6264
rect 35624 5092 35676 5098
rect 35624 5034 35676 5040
rect 35348 3596 35400 3602
rect 35348 3538 35400 3544
rect 34274 3292 34582 3301
rect 34274 3290 34280 3292
rect 34336 3290 34360 3292
rect 34416 3290 34440 3292
rect 34496 3290 34520 3292
rect 34576 3290 34582 3292
rect 34336 3238 34338 3290
rect 34518 3238 34520 3290
rect 34274 3236 34280 3238
rect 34336 3236 34360 3238
rect 34416 3236 34440 3238
rect 34496 3236 34520 3238
rect 34576 3236 34582 3238
rect 34274 3227 34582 3236
rect 27068 2644 27120 2650
rect 27068 2586 27120 2592
rect 29276 2644 29328 2650
rect 29276 2586 29328 2592
rect 22940 2508 23348 2514
rect 22940 2502 23296 2508
rect 23296 2450 23348 2456
rect 25504 2508 25556 2514
rect 25504 2450 25556 2456
rect 23756 2440 23808 2446
rect 23756 2382 23808 2388
rect 23940 2440 23992 2446
rect 23940 2382 23992 2388
rect 24676 2440 24728 2446
rect 24676 2382 24728 2388
rect 26884 2440 26936 2446
rect 26884 2382 26936 2388
rect 29092 2440 29144 2446
rect 29092 2382 29144 2388
rect 31300 2440 31352 2446
rect 31300 2382 31352 2388
rect 33508 2440 33560 2446
rect 33508 2382 33560 2388
rect 35716 2440 35768 2446
rect 35716 2382 35768 2388
rect 22836 2372 22888 2378
rect 22836 2314 22888 2320
rect 23020 2372 23072 2378
rect 23020 2314 23072 2320
rect 23032 2106 23060 2314
rect 23166 2204 23474 2213
rect 23166 2202 23172 2204
rect 23228 2202 23252 2204
rect 23308 2202 23332 2204
rect 23388 2202 23412 2204
rect 23468 2202 23474 2204
rect 23228 2150 23230 2202
rect 23410 2150 23412 2202
rect 23166 2148 23172 2150
rect 23228 2148 23252 2150
rect 23308 2148 23332 2150
rect 23388 2148 23412 2150
rect 23468 2148 23474 2150
rect 23166 2139 23474 2148
rect 23768 2106 23796 2382
rect 23020 2100 23072 2106
rect 23020 2042 23072 2048
rect 23756 2100 23808 2106
rect 23756 2042 23808 2048
rect 23952 2038 23980 2382
rect 24688 2106 24716 2382
rect 26896 2106 26924 2382
rect 29104 2106 29132 2382
rect 31312 2106 31340 2382
rect 33520 2106 33548 2382
rect 34274 2204 34582 2213
rect 34274 2202 34280 2204
rect 34336 2202 34360 2204
rect 34416 2202 34440 2204
rect 34496 2202 34520 2204
rect 34576 2202 34582 2204
rect 34336 2150 34338 2202
rect 34518 2150 34520 2202
rect 34274 2148 34280 2150
rect 34336 2148 34360 2150
rect 34416 2148 34440 2150
rect 34496 2148 34520 2150
rect 34576 2148 34582 2150
rect 34274 2139 34582 2148
rect 35728 2106 35756 2382
rect 36096 2378 36124 9386
rect 36188 8480 36216 9840
rect 36268 8492 36320 8498
rect 36188 8452 36268 8480
rect 36556 8480 36584 9840
rect 36820 9648 36872 9654
rect 36820 9590 36872 9596
rect 36832 8498 36860 9590
rect 36924 8498 36952 9840
rect 37292 9812 37412 9840
rect 37568 8498 37596 9846
rect 37646 9840 37702 10300
rect 37752 9846 37872 9874
rect 37752 9840 37780 9846
rect 37660 9812 37780 9840
rect 37844 8498 37872 9846
rect 38014 9840 38070 10300
rect 38382 9840 38438 10300
rect 38750 9840 38806 10300
rect 38856 9846 39068 9874
rect 38856 9840 38884 9846
rect 36636 8492 36688 8498
rect 36556 8452 36636 8480
rect 36268 8434 36320 8440
rect 36636 8434 36688 8440
rect 36820 8492 36872 8498
rect 36820 8434 36872 8440
rect 36912 8492 36964 8498
rect 36912 8434 36964 8440
rect 37556 8492 37608 8498
rect 37556 8434 37608 8440
rect 37832 8492 37884 8498
rect 38028 8480 38056 9840
rect 38108 8492 38160 8498
rect 38028 8452 38108 8480
rect 37832 8434 37884 8440
rect 38396 8480 38424 9840
rect 38764 9812 38884 9840
rect 38660 9512 38712 9518
rect 38660 9454 38712 9460
rect 38672 8634 38700 9454
rect 39040 8634 39068 9846
rect 39118 9840 39174 10300
rect 39486 9840 39542 10300
rect 39592 9846 39804 9874
rect 39592 9840 39620 9846
rect 39132 8634 39160 9840
rect 39500 9812 39620 9840
rect 39776 8634 39804 9846
rect 39854 9840 39910 10300
rect 40222 9840 40278 10300
rect 40590 9840 40646 10300
rect 40958 9840 41014 10300
rect 41326 9840 41382 10300
rect 41694 9840 41750 10300
rect 42062 9840 42118 10300
rect 42430 9840 42486 10300
rect 42536 9846 42748 9874
rect 38660 8628 38712 8634
rect 38660 8570 38712 8576
rect 39028 8628 39080 8634
rect 39028 8570 39080 8576
rect 39120 8628 39172 8634
rect 39120 8570 39172 8576
rect 39764 8628 39816 8634
rect 39764 8570 39816 8576
rect 39868 8566 39896 9840
rect 39948 8900 40000 8906
rect 39948 8842 40000 8848
rect 39856 8560 39908 8566
rect 39856 8502 39908 8508
rect 39960 8498 39988 8842
rect 40236 8498 40264 9840
rect 40500 8832 40552 8838
rect 40500 8774 40552 8780
rect 40512 8498 40540 8774
rect 38476 8492 38528 8498
rect 38396 8452 38476 8480
rect 38108 8434 38160 8440
rect 38476 8434 38528 8440
rect 38568 8492 38620 8498
rect 38568 8434 38620 8440
rect 39948 8492 40000 8498
rect 39948 8434 40000 8440
rect 40224 8492 40276 8498
rect 40224 8434 40276 8440
rect 40500 8492 40552 8498
rect 40500 8434 40552 8440
rect 37464 8356 37516 8362
rect 37464 8298 37516 8304
rect 37740 8356 37792 8362
rect 37740 8298 37792 8304
rect 37188 8288 37240 8294
rect 37188 8230 37240 8236
rect 37200 3534 37228 8230
rect 37476 7993 37504 8298
rect 37462 7984 37518 7993
rect 37462 7919 37518 7928
rect 37752 7206 37780 8298
rect 37740 7200 37792 7206
rect 37740 7142 37792 7148
rect 37188 3528 37240 3534
rect 37188 3470 37240 3476
rect 38580 3466 38608 8434
rect 39828 8188 40136 8197
rect 39828 8186 39834 8188
rect 39890 8186 39914 8188
rect 39970 8186 39994 8188
rect 40050 8186 40074 8188
rect 40130 8186 40136 8188
rect 39890 8134 39892 8186
rect 40072 8134 40074 8186
rect 39828 8132 39834 8134
rect 39890 8132 39914 8134
rect 39970 8132 39994 8134
rect 40050 8132 40074 8134
rect 40130 8132 40136 8134
rect 39828 8123 40136 8132
rect 40604 8090 40632 9840
rect 40684 8832 40736 8838
rect 40684 8774 40736 8780
rect 40696 8498 40724 8774
rect 40972 8634 41000 9840
rect 41052 9308 41104 9314
rect 41052 9250 41104 9256
rect 40960 8628 41012 8634
rect 40960 8570 41012 8576
rect 41064 8498 41092 9250
rect 41340 8566 41368 9840
rect 41328 8560 41380 8566
rect 41328 8502 41380 8508
rect 40684 8492 40736 8498
rect 40684 8434 40736 8440
rect 41052 8492 41104 8498
rect 41052 8434 41104 8440
rect 41708 8362 41736 9840
rect 42076 8430 42104 9840
rect 42444 9738 42472 9840
rect 42536 9738 42564 9846
rect 42444 9710 42564 9738
rect 42720 8634 42748 9846
rect 42798 9840 42854 10300
rect 43166 9840 43222 10300
rect 43534 9840 43590 10300
rect 43902 9840 43958 10300
rect 44270 9840 44326 10300
rect 44638 9840 44694 10300
rect 45006 9840 45062 10300
rect 45374 9840 45430 10300
rect 45742 9840 45798 10300
rect 46110 9840 46166 10300
rect 42708 8628 42760 8634
rect 42708 8570 42760 8576
rect 42524 8492 42576 8498
rect 42524 8434 42576 8440
rect 42064 8424 42116 8430
rect 42064 8366 42116 8372
rect 41696 8356 41748 8362
rect 41696 8298 41748 8304
rect 40592 8084 40644 8090
rect 40592 8026 40644 8032
rect 39672 7812 39724 7818
rect 39672 7754 39724 7760
rect 38568 3460 38620 3466
rect 38568 3402 38620 3408
rect 39684 2582 39712 7754
rect 39828 7100 40136 7109
rect 39828 7098 39834 7100
rect 39890 7098 39914 7100
rect 39970 7098 39994 7100
rect 40050 7098 40074 7100
rect 40130 7098 40136 7100
rect 39890 7046 39892 7098
rect 40072 7046 40074 7098
rect 39828 7044 39834 7046
rect 39890 7044 39914 7046
rect 39970 7044 39994 7046
rect 40050 7044 40074 7046
rect 40130 7044 40136 7046
rect 39828 7035 40136 7044
rect 42536 6186 42564 8434
rect 42812 8090 42840 9840
rect 42892 9172 42944 9178
rect 42892 9114 42944 9120
rect 42904 8566 42932 9114
rect 42892 8560 42944 8566
rect 42892 8502 42944 8508
rect 42800 8084 42852 8090
rect 42800 8026 42852 8032
rect 42800 7812 42852 7818
rect 42800 7754 42852 7760
rect 42812 6254 42840 7754
rect 43180 7546 43208 9840
rect 43260 8968 43312 8974
rect 43260 8910 43312 8916
rect 43272 8566 43300 8910
rect 43260 8560 43312 8566
rect 43260 8502 43312 8508
rect 43548 8090 43576 9840
rect 43628 9240 43680 9246
rect 43628 9182 43680 9188
rect 43640 8498 43668 9182
rect 43628 8492 43680 8498
rect 43628 8434 43680 8440
rect 43916 8090 43944 9840
rect 43536 8084 43588 8090
rect 43536 8026 43588 8032
rect 43904 8084 43956 8090
rect 43904 8026 43956 8032
rect 44284 8022 44312 9840
rect 44272 8016 44324 8022
rect 44272 7958 44324 7964
rect 43444 7812 43496 7818
rect 43444 7754 43496 7760
rect 44272 7812 44324 7818
rect 44272 7754 44324 7760
rect 43456 7562 43484 7754
rect 43168 7540 43220 7546
rect 43168 7482 43220 7488
rect 43272 7534 43484 7562
rect 42800 6248 42852 6254
rect 42800 6190 42852 6196
rect 42524 6180 42576 6186
rect 42524 6122 42576 6128
rect 39828 6012 40136 6021
rect 39828 6010 39834 6012
rect 39890 6010 39914 6012
rect 39970 6010 39994 6012
rect 40050 6010 40074 6012
rect 40130 6010 40136 6012
rect 39890 5958 39892 6010
rect 40072 5958 40074 6010
rect 39828 5956 39834 5958
rect 39890 5956 39914 5958
rect 39970 5956 39994 5958
rect 40050 5956 40074 5958
rect 40130 5956 40136 5958
rect 39828 5947 40136 5956
rect 39828 4924 40136 4933
rect 39828 4922 39834 4924
rect 39890 4922 39914 4924
rect 39970 4922 39994 4924
rect 40050 4922 40074 4924
rect 40130 4922 40136 4924
rect 39890 4870 39892 4922
rect 40072 4870 40074 4922
rect 39828 4868 39834 4870
rect 39890 4868 39914 4870
rect 39970 4868 39994 4870
rect 40050 4868 40074 4870
rect 40130 4868 40136 4870
rect 39828 4859 40136 4868
rect 39828 3836 40136 3845
rect 39828 3834 39834 3836
rect 39890 3834 39914 3836
rect 39970 3834 39994 3836
rect 40050 3834 40074 3836
rect 40130 3834 40136 3836
rect 39890 3782 39892 3834
rect 40072 3782 40074 3834
rect 39828 3780 39834 3782
rect 39890 3780 39914 3782
rect 39970 3780 39994 3782
rect 40050 3780 40074 3782
rect 40130 3780 40136 3782
rect 39828 3771 40136 3780
rect 39828 2748 40136 2757
rect 39828 2746 39834 2748
rect 39890 2746 39914 2748
rect 39970 2746 39994 2748
rect 40050 2746 40074 2748
rect 40130 2746 40136 2748
rect 39890 2694 39892 2746
rect 40072 2694 40074 2746
rect 39828 2692 39834 2694
rect 39890 2692 39914 2694
rect 39970 2692 39994 2694
rect 40050 2692 40074 2694
rect 40130 2692 40136 2694
rect 39828 2683 40136 2692
rect 43272 2650 43300 7534
rect 43352 7404 43404 7410
rect 43352 7346 43404 7352
rect 44180 7404 44232 7410
rect 44180 7346 44232 7352
rect 43364 4826 43392 7346
rect 43904 6724 43956 6730
rect 43904 6666 43956 6672
rect 43352 4820 43404 4826
rect 43352 4762 43404 4768
rect 43916 2650 43944 6666
rect 44192 2650 44220 7346
rect 44284 2650 44312 7754
rect 44456 6724 44508 6730
rect 44456 6666 44508 6672
rect 44468 2650 44496 6666
rect 44652 6458 44680 9840
rect 45020 7546 45048 9840
rect 45388 8922 45416 9840
rect 45296 8894 45416 8922
rect 45008 7540 45060 7546
rect 45008 7482 45060 7488
rect 45008 7336 45060 7342
rect 45008 7278 45060 7284
rect 44640 6452 44692 6458
rect 44640 6394 44692 6400
rect 44824 6316 44876 6322
rect 44824 6258 44876 6264
rect 43260 2644 43312 2650
rect 43260 2586 43312 2592
rect 43904 2644 43956 2650
rect 43904 2586 43956 2592
rect 44180 2644 44232 2650
rect 44180 2586 44232 2592
rect 44272 2644 44324 2650
rect 44272 2586 44324 2592
rect 44456 2644 44508 2650
rect 44456 2586 44508 2592
rect 39672 2576 39724 2582
rect 39672 2518 39724 2524
rect 41604 2508 41656 2514
rect 41604 2450 41656 2456
rect 37924 2440 37976 2446
rect 37924 2382 37976 2388
rect 36084 2372 36136 2378
rect 36084 2314 36136 2320
rect 37936 2106 37964 2382
rect 41616 2106 41644 2450
rect 44836 2446 44864 6258
rect 45020 2650 45048 7278
rect 45296 6866 45324 8894
rect 45382 8732 45690 8741
rect 45382 8730 45388 8732
rect 45444 8730 45468 8732
rect 45524 8730 45548 8732
rect 45604 8730 45628 8732
rect 45684 8730 45690 8732
rect 45444 8678 45446 8730
rect 45626 8678 45628 8730
rect 45382 8676 45388 8678
rect 45444 8676 45468 8678
rect 45524 8676 45548 8678
rect 45604 8676 45628 8678
rect 45684 8676 45690 8678
rect 45382 8667 45690 8676
rect 45382 7644 45690 7653
rect 45382 7642 45388 7644
rect 45444 7642 45468 7644
rect 45524 7642 45548 7644
rect 45604 7642 45628 7644
rect 45684 7642 45690 7644
rect 45444 7590 45446 7642
rect 45626 7590 45628 7642
rect 45382 7588 45388 7590
rect 45444 7588 45468 7590
rect 45524 7588 45548 7590
rect 45604 7588 45628 7590
rect 45684 7588 45690 7590
rect 45382 7579 45690 7588
rect 45756 7546 45784 9840
rect 45744 7540 45796 7546
rect 45744 7482 45796 7488
rect 46124 6866 46152 9840
rect 45284 6860 45336 6866
rect 45284 6802 45336 6808
rect 46112 6860 46164 6866
rect 46112 6802 46164 6808
rect 45382 6556 45690 6565
rect 45382 6554 45388 6556
rect 45444 6554 45468 6556
rect 45524 6554 45548 6556
rect 45604 6554 45628 6556
rect 45684 6554 45690 6556
rect 45444 6502 45446 6554
rect 45626 6502 45628 6554
rect 45382 6500 45388 6502
rect 45444 6500 45468 6502
rect 45524 6500 45548 6502
rect 45604 6500 45628 6502
rect 45684 6500 45690 6502
rect 45382 6491 45690 6500
rect 45382 5468 45690 5477
rect 45382 5466 45388 5468
rect 45444 5466 45468 5468
rect 45524 5466 45548 5468
rect 45604 5466 45628 5468
rect 45684 5466 45690 5468
rect 45444 5414 45446 5466
rect 45626 5414 45628 5466
rect 45382 5412 45388 5414
rect 45444 5412 45468 5414
rect 45524 5412 45548 5414
rect 45604 5412 45628 5414
rect 45684 5412 45690 5414
rect 45382 5403 45690 5412
rect 45382 4380 45690 4389
rect 45382 4378 45388 4380
rect 45444 4378 45468 4380
rect 45524 4378 45548 4380
rect 45604 4378 45628 4380
rect 45684 4378 45690 4380
rect 45444 4326 45446 4378
rect 45626 4326 45628 4378
rect 45382 4324 45388 4326
rect 45444 4324 45468 4326
rect 45524 4324 45548 4326
rect 45604 4324 45628 4326
rect 45684 4324 45690 4326
rect 45382 4315 45690 4324
rect 45382 3292 45690 3301
rect 45382 3290 45388 3292
rect 45444 3290 45468 3292
rect 45524 3290 45548 3292
rect 45604 3290 45628 3292
rect 45684 3290 45690 3292
rect 45444 3238 45446 3290
rect 45626 3238 45628 3290
rect 45382 3236 45388 3238
rect 45444 3236 45468 3238
rect 45524 3236 45548 3238
rect 45604 3236 45628 3238
rect 45684 3236 45690 3238
rect 45382 3227 45690 3236
rect 45008 2644 45060 2650
rect 45008 2586 45060 2592
rect 44088 2440 44140 2446
rect 44088 2382 44140 2388
rect 44824 2440 44876 2446
rect 44824 2382 44876 2388
rect 45192 2440 45244 2446
rect 45192 2382 45244 2388
rect 43444 2372 43496 2378
rect 43444 2314 43496 2320
rect 43456 2106 43484 2314
rect 44100 2106 44128 2382
rect 24676 2100 24728 2106
rect 24676 2042 24728 2048
rect 26884 2100 26936 2106
rect 26884 2042 26936 2048
rect 29092 2100 29144 2106
rect 29092 2042 29144 2048
rect 31300 2100 31352 2106
rect 31300 2042 31352 2048
rect 33508 2100 33560 2106
rect 33508 2042 33560 2048
rect 35716 2100 35768 2106
rect 35716 2042 35768 2048
rect 37924 2100 37976 2106
rect 37924 2042 37976 2048
rect 41604 2100 41656 2106
rect 41604 2042 41656 2048
rect 43444 2100 43496 2106
rect 43444 2042 43496 2048
rect 44088 2100 44140 2106
rect 44088 2042 44140 2048
rect 45204 2038 45232 2382
rect 45382 2204 45690 2213
rect 45382 2202 45388 2204
rect 45444 2202 45468 2204
rect 45524 2202 45548 2204
rect 45604 2202 45628 2204
rect 45684 2202 45690 2204
rect 45444 2150 45446 2202
rect 45626 2150 45628 2202
rect 45382 2148 45388 2150
rect 45444 2148 45468 2150
rect 45524 2148 45548 2150
rect 45604 2148 45628 2150
rect 45684 2148 45690 2150
rect 45382 2139 45690 2148
rect 23940 2032 23992 2038
rect 23940 1974 23992 1980
rect 45192 2032 45244 2038
rect 45192 1974 45244 1980
rect 22836 1964 22888 1970
rect 22836 1906 22888 1912
rect 23020 1964 23072 1970
rect 23020 1906 23072 1912
rect 23664 1964 23716 1970
rect 23664 1906 23716 1912
rect 24032 1964 24084 1970
rect 24032 1906 24084 1912
rect 26240 1964 26292 1970
rect 26240 1906 26292 1912
rect 28448 1964 28500 1970
rect 28448 1906 28500 1912
rect 30656 1964 30708 1970
rect 30656 1906 30708 1912
rect 32864 1964 32916 1970
rect 32864 1906 32916 1912
rect 35072 1964 35124 1970
rect 35072 1906 35124 1912
rect 37464 1964 37516 1970
rect 37464 1906 37516 1912
rect 41788 1964 41840 1970
rect 41788 1906 41840 1912
rect 43628 1964 43680 1970
rect 43628 1906 43680 1912
rect 44088 1964 44140 1970
rect 44088 1906 44140 1912
rect 44548 1964 44600 1970
rect 44548 1906 44600 1912
rect 22744 1760 22796 1766
rect 22744 1702 22796 1708
rect 22848 1562 22876 1906
rect 22836 1556 22888 1562
rect 22836 1498 22888 1504
rect 22284 1352 22336 1358
rect 22284 1294 22336 1300
rect 22192 1284 22244 1290
rect 22192 1226 22244 1232
rect 22296 1018 22324 1294
rect 22284 1012 22336 1018
rect 22284 954 22336 960
rect 23032 814 23060 1906
rect 23572 1352 23624 1358
rect 23572 1294 23624 1300
rect 23166 1116 23474 1125
rect 23166 1114 23172 1116
rect 23228 1114 23252 1116
rect 23308 1114 23332 1116
rect 23388 1114 23412 1116
rect 23468 1114 23474 1116
rect 23228 1062 23230 1114
rect 23410 1062 23412 1114
rect 23166 1060 23172 1062
rect 23228 1060 23252 1062
rect 23308 1060 23332 1062
rect 23388 1060 23412 1062
rect 23468 1060 23474 1062
rect 23166 1051 23474 1060
rect 23020 808 23072 814
rect 23020 750 23072 756
rect 21548 672 21600 678
rect 21548 614 21600 620
rect 23308 190 23428 218
rect 23308 160 23336 190
rect 21086 54 21404 82
rect 14462 -300 14518 54
rect 16670 -300 16726 54
rect 18878 -300 18934 54
rect 21086 -300 21142 54
rect 23294 -300 23350 160
rect 23400 82 23428 190
rect 23584 82 23612 1294
rect 23676 882 23704 1906
rect 24044 1562 24072 1906
rect 24032 1556 24084 1562
rect 24032 1498 24084 1504
rect 25780 1352 25832 1358
rect 25780 1294 25832 1300
rect 23664 876 23716 882
rect 23664 818 23716 824
rect 23400 54 23612 82
rect 25502 82 25558 160
rect 25792 82 25820 1294
rect 26252 1222 26280 1906
rect 28460 1562 28488 1906
rect 28720 1660 29028 1669
rect 28720 1658 28726 1660
rect 28782 1658 28806 1660
rect 28862 1658 28886 1660
rect 28942 1658 28966 1660
rect 29022 1658 29028 1660
rect 28782 1606 28784 1658
rect 28964 1606 28966 1658
rect 28720 1604 28726 1606
rect 28782 1604 28806 1606
rect 28862 1604 28886 1606
rect 28942 1604 28966 1606
rect 29022 1604 29028 1606
rect 28720 1595 29028 1604
rect 28448 1556 28500 1562
rect 28448 1498 28500 1504
rect 30668 1358 30696 1906
rect 32876 1562 32904 1906
rect 35084 1562 35112 1906
rect 32864 1556 32916 1562
rect 32864 1498 32916 1504
rect 35072 1556 35124 1562
rect 35072 1498 35124 1504
rect 37476 1358 37504 1906
rect 39828 1660 40136 1669
rect 39828 1658 39834 1660
rect 39890 1658 39914 1660
rect 39970 1658 39994 1660
rect 40050 1658 40074 1660
rect 40130 1658 40136 1660
rect 39890 1606 39892 1658
rect 40072 1606 40074 1658
rect 39828 1604 39834 1606
rect 39890 1604 39914 1606
rect 39970 1604 39994 1606
rect 40050 1604 40074 1606
rect 40130 1604 40136 1606
rect 39828 1595 40136 1604
rect 27988 1352 28040 1358
rect 27988 1294 28040 1300
rect 30196 1352 30248 1358
rect 30196 1294 30248 1300
rect 30656 1352 30708 1358
rect 30656 1294 30708 1300
rect 32404 1352 32456 1358
rect 32404 1294 32456 1300
rect 34612 1352 34664 1358
rect 34612 1294 34664 1300
rect 36820 1352 36872 1358
rect 36820 1294 36872 1300
rect 37464 1352 37516 1358
rect 37464 1294 37516 1300
rect 39028 1352 39080 1358
rect 39028 1294 39080 1300
rect 41236 1352 41288 1358
rect 41236 1294 41288 1300
rect 26240 1216 26292 1222
rect 26240 1158 26292 1164
rect 25502 54 25820 82
rect 27710 82 27766 160
rect 28000 82 28028 1294
rect 27710 54 28028 82
rect 29918 82 29974 160
rect 30208 82 30236 1294
rect 29918 54 30236 82
rect 32126 82 32182 160
rect 32416 82 32444 1294
rect 34274 1116 34582 1125
rect 34274 1114 34280 1116
rect 34336 1114 34360 1116
rect 34416 1114 34440 1116
rect 34496 1114 34520 1116
rect 34576 1114 34582 1116
rect 34336 1062 34338 1114
rect 34518 1062 34520 1114
rect 34274 1060 34280 1062
rect 34336 1060 34360 1062
rect 34416 1060 34440 1062
rect 34496 1060 34520 1062
rect 34576 1060 34582 1062
rect 34274 1051 34582 1060
rect 32126 54 32444 82
rect 34334 82 34390 160
rect 34624 82 34652 1294
rect 34334 54 34652 82
rect 36542 82 36598 160
rect 36832 82 36860 1294
rect 36542 54 36860 82
rect 38750 82 38806 160
rect 39040 82 39068 1294
rect 38750 54 39068 82
rect 40958 82 41014 160
rect 41248 82 41276 1294
rect 41800 1222 41828 1906
rect 43444 1352 43496 1358
rect 43444 1294 43496 1300
rect 41788 1216 41840 1222
rect 41788 1158 41840 1164
rect 40958 54 41276 82
rect 43166 82 43222 160
rect 43456 82 43484 1294
rect 43640 1290 43668 1906
rect 44100 1562 44128 1906
rect 44560 1562 44588 1906
rect 44088 1556 44140 1562
rect 44088 1498 44140 1504
rect 44548 1556 44600 1562
rect 44548 1498 44600 1504
rect 45192 1352 45244 1358
rect 45192 1294 45244 1300
rect 43628 1284 43680 1290
rect 43628 1226 43680 1232
rect 43166 54 43484 82
rect 45204 82 45232 1294
rect 45382 1116 45690 1125
rect 45382 1114 45388 1116
rect 45444 1114 45468 1116
rect 45524 1114 45548 1116
rect 45604 1114 45628 1116
rect 45684 1114 45690 1116
rect 45444 1062 45446 1114
rect 45626 1062 45628 1114
rect 45382 1060 45388 1062
rect 45444 1060 45468 1062
rect 45524 1060 45548 1062
rect 45604 1060 45628 1062
rect 45684 1060 45690 1062
rect 45382 1051 45690 1060
rect 45374 82 45430 160
rect 45204 54 45430 82
rect 25502 -300 25558 54
rect 27710 -300 27766 54
rect 29918 -300 29974 54
rect 32126 -300 32182 54
rect 34334 -300 34390 54
rect 36542 -300 36598 54
rect 38750 -300 38806 54
rect 40958 -300 41014 54
rect 43166 -300 43222 54
rect 45374 -300 45430 54
<< via2 >>
rect 6510 8186 6566 8188
rect 6590 8186 6646 8188
rect 6670 8186 6726 8188
rect 6750 8186 6806 8188
rect 6510 8134 6556 8186
rect 6556 8134 6566 8186
rect 6590 8134 6620 8186
rect 6620 8134 6632 8186
rect 6632 8134 6646 8186
rect 6670 8134 6684 8186
rect 6684 8134 6696 8186
rect 6696 8134 6726 8186
rect 6750 8134 6760 8186
rect 6760 8134 6806 8186
rect 6510 8132 6566 8134
rect 6590 8132 6646 8134
rect 6670 8132 6726 8134
rect 6750 8132 6806 8134
rect 12438 8880 12494 8936
rect 12064 8730 12120 8732
rect 12144 8730 12200 8732
rect 12224 8730 12280 8732
rect 12304 8730 12360 8732
rect 12064 8678 12110 8730
rect 12110 8678 12120 8730
rect 12144 8678 12174 8730
rect 12174 8678 12186 8730
rect 12186 8678 12200 8730
rect 12224 8678 12238 8730
rect 12238 8678 12250 8730
rect 12250 8678 12280 8730
rect 12304 8678 12314 8730
rect 12314 8678 12360 8730
rect 12064 8676 12120 8678
rect 12144 8676 12200 8678
rect 12224 8676 12280 8678
rect 12304 8676 12360 8678
rect 6510 7098 6566 7100
rect 6590 7098 6646 7100
rect 6670 7098 6726 7100
rect 6750 7098 6806 7100
rect 6510 7046 6556 7098
rect 6556 7046 6566 7098
rect 6590 7046 6620 7098
rect 6620 7046 6632 7098
rect 6632 7046 6646 7098
rect 6670 7046 6684 7098
rect 6684 7046 6696 7098
rect 6696 7046 6726 7098
rect 6750 7046 6760 7098
rect 6760 7046 6806 7098
rect 6510 7044 6566 7046
rect 6590 7044 6646 7046
rect 6670 7044 6726 7046
rect 6750 7044 6806 7046
rect 12064 7642 12120 7644
rect 12144 7642 12200 7644
rect 12224 7642 12280 7644
rect 12304 7642 12360 7644
rect 12064 7590 12110 7642
rect 12110 7590 12120 7642
rect 12144 7590 12174 7642
rect 12174 7590 12186 7642
rect 12186 7590 12200 7642
rect 12224 7590 12238 7642
rect 12238 7590 12250 7642
rect 12250 7590 12280 7642
rect 12304 7590 12314 7642
rect 12314 7590 12360 7642
rect 12064 7588 12120 7590
rect 12144 7588 12200 7590
rect 12224 7588 12280 7590
rect 12304 7588 12360 7590
rect 11518 7384 11574 7440
rect 5446 6840 5502 6896
rect 13634 9560 13690 9616
rect 14370 9852 14426 9888
rect 14370 9832 14372 9852
rect 14372 9832 14424 9852
rect 14424 9832 14426 9852
rect 14370 9152 14426 9208
rect 14554 9732 14556 9752
rect 14556 9732 14608 9752
rect 14608 9732 14610 9752
rect 14554 9696 14610 9732
rect 12622 6704 12678 6760
rect 12064 6554 12120 6556
rect 12144 6554 12200 6556
rect 12224 6554 12280 6556
rect 12304 6554 12360 6556
rect 12064 6502 12110 6554
rect 12110 6502 12120 6554
rect 12144 6502 12174 6554
rect 12174 6502 12186 6554
rect 12186 6502 12200 6554
rect 12224 6502 12238 6554
rect 12238 6502 12250 6554
rect 12250 6502 12280 6554
rect 12304 6502 12314 6554
rect 12314 6502 12360 6554
rect 12064 6500 12120 6502
rect 12144 6500 12200 6502
rect 12224 6500 12280 6502
rect 12304 6500 12360 6502
rect 16394 9832 16450 9888
rect 16486 9696 16542 9752
rect 16762 9424 16818 9480
rect 15106 7812 15162 7848
rect 15106 7792 15108 7812
rect 15108 7792 15160 7812
rect 15160 7792 15162 7812
rect 15106 7540 15162 7576
rect 15106 7520 15108 7540
rect 15108 7520 15160 7540
rect 15160 7520 15162 7540
rect 16118 8336 16174 8392
rect 17130 9288 17186 9344
rect 17958 9016 18014 9072
rect 18326 9696 18382 9752
rect 17618 8186 17674 8188
rect 17698 8186 17754 8188
rect 17778 8186 17834 8188
rect 17858 8186 17914 8188
rect 17618 8134 17664 8186
rect 17664 8134 17674 8186
rect 17698 8134 17728 8186
rect 17728 8134 17740 8186
rect 17740 8134 17754 8186
rect 17778 8134 17792 8186
rect 17792 8134 17804 8186
rect 17804 8134 17834 8186
rect 17858 8134 17868 8186
rect 17868 8134 17914 8186
rect 17618 8132 17674 8134
rect 17698 8132 17754 8134
rect 17778 8132 17834 8134
rect 17858 8132 17914 8134
rect 18050 8064 18106 8120
rect 17958 7928 18014 7984
rect 17222 7692 17224 7712
rect 17224 7692 17276 7712
rect 17276 7692 17278 7712
rect 17222 7656 17278 7692
rect 16946 7384 17002 7440
rect 17618 7098 17674 7100
rect 17698 7098 17754 7100
rect 17778 7098 17834 7100
rect 17858 7098 17914 7100
rect 17618 7046 17664 7098
rect 17664 7046 17674 7098
rect 17698 7046 17728 7098
rect 17728 7046 17740 7098
rect 17740 7046 17754 7098
rect 17778 7046 17792 7098
rect 17792 7046 17804 7098
rect 17804 7046 17834 7098
rect 17858 7046 17868 7098
rect 17868 7046 17914 7098
rect 17618 7044 17674 7046
rect 17698 7044 17754 7046
rect 17778 7044 17834 7046
rect 17858 7044 17914 7046
rect 18786 8200 18842 8256
rect 18786 7540 18842 7576
rect 18786 7520 18788 7540
rect 18788 7520 18840 7540
rect 18840 7520 18842 7540
rect 19890 9868 19892 9888
rect 19892 9868 19944 9888
rect 19944 9868 19946 9888
rect 19890 9832 19946 9868
rect 20166 9424 20222 9480
rect 20810 9288 20866 9344
rect 20810 8336 20866 8392
rect 21178 9696 21234 9752
rect 21178 9560 21234 9616
rect 21270 8200 21326 8256
rect 21270 7928 21326 7984
rect 21638 7656 21694 7712
rect 22466 8472 22522 8528
rect 23172 8730 23228 8732
rect 23252 8730 23308 8732
rect 23332 8730 23388 8732
rect 23412 8730 23468 8732
rect 23172 8678 23218 8730
rect 23218 8678 23228 8730
rect 23252 8678 23282 8730
rect 23282 8678 23294 8730
rect 23294 8678 23308 8730
rect 23332 8678 23346 8730
rect 23346 8678 23358 8730
rect 23358 8678 23388 8730
rect 23412 8678 23422 8730
rect 23422 8678 23468 8730
rect 23172 8676 23228 8678
rect 23252 8676 23308 8678
rect 23332 8676 23388 8678
rect 23412 8676 23468 8678
rect 22834 8356 22890 8392
rect 22006 7928 22062 7984
rect 21730 7248 21786 7304
rect 22098 7384 22154 7440
rect 22834 8336 22836 8356
rect 22836 8336 22888 8356
rect 22888 8336 22890 8356
rect 22926 7404 22982 7440
rect 23202 8336 23258 8392
rect 23938 9832 23994 9888
rect 23662 9288 23718 9344
rect 23478 8064 23534 8120
rect 23172 7642 23228 7644
rect 23252 7642 23308 7644
rect 23332 7642 23388 7644
rect 23412 7642 23468 7644
rect 23172 7590 23218 7642
rect 23218 7590 23228 7642
rect 23252 7590 23282 7642
rect 23282 7590 23294 7642
rect 23294 7590 23308 7642
rect 23332 7590 23346 7642
rect 23346 7590 23358 7642
rect 23358 7590 23388 7642
rect 23412 7590 23422 7642
rect 23422 7590 23468 7642
rect 23172 7588 23228 7590
rect 23252 7588 23308 7590
rect 23332 7588 23388 7590
rect 23412 7588 23468 7590
rect 23846 8608 23902 8664
rect 23938 8064 23994 8120
rect 22926 7384 22928 7404
rect 22928 7384 22980 7404
rect 22980 7384 22982 7404
rect 23202 7148 23204 7168
rect 23204 7148 23256 7168
rect 23256 7148 23258 7168
rect 23202 7112 23258 7148
rect 24306 9288 24362 9344
rect 24490 8472 24546 8528
rect 25226 8880 25282 8936
rect 24582 8200 24638 8256
rect 24766 8064 24822 8120
rect 23172 6554 23228 6556
rect 23252 6554 23308 6556
rect 23332 6554 23388 6556
rect 23412 6554 23468 6556
rect 23172 6502 23218 6554
rect 23218 6502 23228 6554
rect 23252 6502 23282 6554
rect 23282 6502 23294 6554
rect 23294 6502 23308 6554
rect 23332 6502 23346 6554
rect 23346 6502 23358 6554
rect 23358 6502 23388 6554
rect 23412 6502 23422 6554
rect 23422 6502 23468 6554
rect 23172 6500 23228 6502
rect 23252 6500 23308 6502
rect 23332 6500 23388 6502
rect 23412 6500 23468 6502
rect 6510 6010 6566 6012
rect 6590 6010 6646 6012
rect 6670 6010 6726 6012
rect 6750 6010 6806 6012
rect 6510 5958 6556 6010
rect 6556 5958 6566 6010
rect 6590 5958 6620 6010
rect 6620 5958 6632 6010
rect 6632 5958 6646 6010
rect 6670 5958 6684 6010
rect 6684 5958 6696 6010
rect 6696 5958 6726 6010
rect 6750 5958 6760 6010
rect 6760 5958 6806 6010
rect 6510 5956 6566 5958
rect 6590 5956 6646 5958
rect 6670 5956 6726 5958
rect 6750 5956 6806 5958
rect 17618 6010 17674 6012
rect 17698 6010 17754 6012
rect 17778 6010 17834 6012
rect 17858 6010 17914 6012
rect 17618 5958 17664 6010
rect 17664 5958 17674 6010
rect 17698 5958 17728 6010
rect 17728 5958 17740 6010
rect 17740 5958 17754 6010
rect 17778 5958 17792 6010
rect 17792 5958 17804 6010
rect 17804 5958 17834 6010
rect 17858 5958 17868 6010
rect 17868 5958 17914 6010
rect 17618 5956 17674 5958
rect 17698 5956 17754 5958
rect 17778 5956 17834 5958
rect 17858 5956 17914 5958
rect 12064 5466 12120 5468
rect 12144 5466 12200 5468
rect 12224 5466 12280 5468
rect 12304 5466 12360 5468
rect 12064 5414 12110 5466
rect 12110 5414 12120 5466
rect 12144 5414 12174 5466
rect 12174 5414 12186 5466
rect 12186 5414 12200 5466
rect 12224 5414 12238 5466
rect 12238 5414 12250 5466
rect 12250 5414 12280 5466
rect 12304 5414 12314 5466
rect 12314 5414 12360 5466
rect 12064 5412 12120 5414
rect 12144 5412 12200 5414
rect 12224 5412 12280 5414
rect 12304 5412 12360 5414
rect 23172 5466 23228 5468
rect 23252 5466 23308 5468
rect 23332 5466 23388 5468
rect 23412 5466 23468 5468
rect 23172 5414 23218 5466
rect 23218 5414 23228 5466
rect 23252 5414 23282 5466
rect 23282 5414 23294 5466
rect 23294 5414 23308 5466
rect 23332 5414 23346 5466
rect 23346 5414 23358 5466
rect 23358 5414 23388 5466
rect 23412 5414 23422 5466
rect 23422 5414 23468 5466
rect 23172 5412 23228 5414
rect 23252 5412 23308 5414
rect 23332 5412 23388 5414
rect 23412 5412 23468 5414
rect 6510 4922 6566 4924
rect 6590 4922 6646 4924
rect 6670 4922 6726 4924
rect 6750 4922 6806 4924
rect 6510 4870 6556 4922
rect 6556 4870 6566 4922
rect 6590 4870 6620 4922
rect 6620 4870 6632 4922
rect 6632 4870 6646 4922
rect 6670 4870 6684 4922
rect 6684 4870 6696 4922
rect 6696 4870 6726 4922
rect 6750 4870 6760 4922
rect 6760 4870 6806 4922
rect 6510 4868 6566 4870
rect 6590 4868 6646 4870
rect 6670 4868 6726 4870
rect 6750 4868 6806 4870
rect 17618 4922 17674 4924
rect 17698 4922 17754 4924
rect 17778 4922 17834 4924
rect 17858 4922 17914 4924
rect 17618 4870 17664 4922
rect 17664 4870 17674 4922
rect 17698 4870 17728 4922
rect 17728 4870 17740 4922
rect 17740 4870 17754 4922
rect 17778 4870 17792 4922
rect 17792 4870 17804 4922
rect 17804 4870 17834 4922
rect 17858 4870 17868 4922
rect 17868 4870 17914 4922
rect 17618 4868 17674 4870
rect 17698 4868 17754 4870
rect 17778 4868 17834 4870
rect 17858 4868 17914 4870
rect 12064 4378 12120 4380
rect 12144 4378 12200 4380
rect 12224 4378 12280 4380
rect 12304 4378 12360 4380
rect 12064 4326 12110 4378
rect 12110 4326 12120 4378
rect 12144 4326 12174 4378
rect 12174 4326 12186 4378
rect 12186 4326 12200 4378
rect 12224 4326 12238 4378
rect 12238 4326 12250 4378
rect 12250 4326 12280 4378
rect 12304 4326 12314 4378
rect 12314 4326 12360 4378
rect 12064 4324 12120 4326
rect 12144 4324 12200 4326
rect 12224 4324 12280 4326
rect 12304 4324 12360 4326
rect 6510 3834 6566 3836
rect 6590 3834 6646 3836
rect 6670 3834 6726 3836
rect 6750 3834 6806 3836
rect 6510 3782 6556 3834
rect 6556 3782 6566 3834
rect 6590 3782 6620 3834
rect 6620 3782 6632 3834
rect 6632 3782 6646 3834
rect 6670 3782 6684 3834
rect 6684 3782 6696 3834
rect 6696 3782 6726 3834
rect 6750 3782 6760 3834
rect 6760 3782 6806 3834
rect 6510 3780 6566 3782
rect 6590 3780 6646 3782
rect 6670 3780 6726 3782
rect 6750 3780 6806 3782
rect 17618 3834 17674 3836
rect 17698 3834 17754 3836
rect 17778 3834 17834 3836
rect 17858 3834 17914 3836
rect 17618 3782 17664 3834
rect 17664 3782 17674 3834
rect 17698 3782 17728 3834
rect 17728 3782 17740 3834
rect 17740 3782 17754 3834
rect 17778 3782 17792 3834
rect 17792 3782 17804 3834
rect 17804 3782 17834 3834
rect 17858 3782 17868 3834
rect 17868 3782 17914 3834
rect 17618 3780 17674 3782
rect 17698 3780 17754 3782
rect 17778 3780 17834 3782
rect 17858 3780 17914 3782
rect 12064 3290 12120 3292
rect 12144 3290 12200 3292
rect 12224 3290 12280 3292
rect 12304 3290 12360 3292
rect 12064 3238 12110 3290
rect 12110 3238 12120 3290
rect 12144 3238 12174 3290
rect 12174 3238 12186 3290
rect 12186 3238 12200 3290
rect 12224 3238 12238 3290
rect 12238 3238 12250 3290
rect 12250 3238 12280 3290
rect 12304 3238 12314 3290
rect 12314 3238 12360 3290
rect 12064 3236 12120 3238
rect 12144 3236 12200 3238
rect 12224 3236 12280 3238
rect 12304 3236 12360 3238
rect 6510 2746 6566 2748
rect 6590 2746 6646 2748
rect 6670 2746 6726 2748
rect 6750 2746 6806 2748
rect 6510 2694 6556 2746
rect 6556 2694 6566 2746
rect 6590 2694 6620 2746
rect 6620 2694 6632 2746
rect 6632 2694 6646 2746
rect 6670 2694 6684 2746
rect 6684 2694 6696 2746
rect 6696 2694 6726 2746
rect 6750 2694 6760 2746
rect 6760 2694 6806 2746
rect 6510 2692 6566 2694
rect 6590 2692 6646 2694
rect 6670 2692 6726 2694
rect 6750 2692 6806 2694
rect 17618 2746 17674 2748
rect 17698 2746 17754 2748
rect 17778 2746 17834 2748
rect 17858 2746 17914 2748
rect 17618 2694 17664 2746
rect 17664 2694 17674 2746
rect 17698 2694 17728 2746
rect 17728 2694 17740 2746
rect 17740 2694 17754 2746
rect 17778 2694 17792 2746
rect 17792 2694 17804 2746
rect 17804 2694 17834 2746
rect 17858 2694 17868 2746
rect 17868 2694 17914 2746
rect 17618 2692 17674 2694
rect 17698 2692 17754 2694
rect 17778 2692 17834 2694
rect 17858 2692 17914 2694
rect 12064 2202 12120 2204
rect 12144 2202 12200 2204
rect 12224 2202 12280 2204
rect 12304 2202 12360 2204
rect 12064 2150 12110 2202
rect 12110 2150 12120 2202
rect 12144 2150 12174 2202
rect 12174 2150 12186 2202
rect 12186 2150 12200 2202
rect 12224 2150 12238 2202
rect 12238 2150 12250 2202
rect 12250 2150 12280 2202
rect 12304 2150 12314 2202
rect 12314 2150 12360 2202
rect 12064 2148 12120 2150
rect 12144 2148 12200 2150
rect 12224 2148 12280 2150
rect 12304 2148 12360 2150
rect 6510 1658 6566 1660
rect 6590 1658 6646 1660
rect 6670 1658 6726 1660
rect 6750 1658 6806 1660
rect 6510 1606 6556 1658
rect 6556 1606 6566 1658
rect 6590 1606 6620 1658
rect 6620 1606 6632 1658
rect 6632 1606 6646 1658
rect 6670 1606 6684 1658
rect 6684 1606 6696 1658
rect 6696 1606 6726 1658
rect 6750 1606 6760 1658
rect 6760 1606 6806 1658
rect 6510 1604 6566 1606
rect 6590 1604 6646 1606
rect 6670 1604 6726 1606
rect 6750 1604 6806 1606
rect 17618 1658 17674 1660
rect 17698 1658 17754 1660
rect 17778 1658 17834 1660
rect 17858 1658 17914 1660
rect 17618 1606 17664 1658
rect 17664 1606 17674 1658
rect 17698 1606 17728 1658
rect 17728 1606 17740 1658
rect 17740 1606 17754 1658
rect 17778 1606 17792 1658
rect 17792 1606 17804 1658
rect 17804 1606 17834 1658
rect 17858 1606 17868 1658
rect 17868 1606 17914 1658
rect 17618 1604 17674 1606
rect 17698 1604 17754 1606
rect 17778 1604 17834 1606
rect 17858 1604 17914 1606
rect 12064 1114 12120 1116
rect 12144 1114 12200 1116
rect 12224 1114 12280 1116
rect 12304 1114 12360 1116
rect 12064 1062 12110 1114
rect 12110 1062 12120 1114
rect 12144 1062 12174 1114
rect 12174 1062 12186 1114
rect 12186 1062 12200 1114
rect 12224 1062 12238 1114
rect 12238 1062 12250 1114
rect 12250 1062 12280 1114
rect 12304 1062 12314 1114
rect 12314 1062 12360 1114
rect 12064 1060 12120 1062
rect 12144 1060 12200 1062
rect 12224 1060 12280 1062
rect 12304 1060 12360 1062
rect 23172 4378 23228 4380
rect 23252 4378 23308 4380
rect 23332 4378 23388 4380
rect 23412 4378 23468 4380
rect 23172 4326 23218 4378
rect 23218 4326 23228 4378
rect 23252 4326 23282 4378
rect 23282 4326 23294 4378
rect 23294 4326 23308 4378
rect 23332 4326 23346 4378
rect 23346 4326 23358 4378
rect 23358 4326 23388 4378
rect 23412 4326 23422 4378
rect 23422 4326 23468 4378
rect 23172 4324 23228 4326
rect 23252 4324 23308 4326
rect 23332 4324 23388 4326
rect 23412 4324 23468 4326
rect 23172 3290 23228 3292
rect 23252 3290 23308 3292
rect 23332 3290 23388 3292
rect 23412 3290 23468 3292
rect 23172 3238 23218 3290
rect 23218 3238 23228 3290
rect 23252 3238 23282 3290
rect 23282 3238 23294 3290
rect 23294 3238 23308 3290
rect 23332 3238 23346 3290
rect 23346 3238 23358 3290
rect 23358 3238 23388 3290
rect 23412 3238 23422 3290
rect 23422 3238 23468 3290
rect 23172 3236 23228 3238
rect 23252 3236 23308 3238
rect 23332 3236 23388 3238
rect 23412 3236 23468 3238
rect 26238 6840 26294 6896
rect 27618 9424 27674 9480
rect 28262 8608 28318 8664
rect 28446 9152 28502 9208
rect 28170 7792 28226 7848
rect 28538 8336 28594 8392
rect 28726 8186 28782 8188
rect 28806 8186 28862 8188
rect 28886 8186 28942 8188
rect 28966 8186 29022 8188
rect 28726 8134 28772 8186
rect 28772 8134 28782 8186
rect 28806 8134 28836 8186
rect 28836 8134 28848 8186
rect 28848 8134 28862 8186
rect 28886 8134 28900 8186
rect 28900 8134 28912 8186
rect 28912 8134 28942 8186
rect 28966 8134 28976 8186
rect 28976 8134 29022 8186
rect 28726 8132 28782 8134
rect 28806 8132 28862 8134
rect 28886 8132 28942 8134
rect 28966 8132 29022 8134
rect 28726 7098 28782 7100
rect 28806 7098 28862 7100
rect 28886 7098 28942 7100
rect 28966 7098 29022 7100
rect 28726 7046 28772 7098
rect 28772 7046 28782 7098
rect 28806 7046 28836 7098
rect 28836 7046 28848 7098
rect 28848 7046 28862 7098
rect 28886 7046 28900 7098
rect 28900 7046 28912 7098
rect 28912 7046 28942 7098
rect 28966 7046 28976 7098
rect 28976 7046 29022 7098
rect 28726 7044 28782 7046
rect 28806 7044 28862 7046
rect 28886 7044 28942 7046
rect 28966 7044 29022 7046
rect 28446 6976 28502 7032
rect 25962 6704 26018 6760
rect 32954 7248 33010 7304
rect 28726 6010 28782 6012
rect 28806 6010 28862 6012
rect 28886 6010 28942 6012
rect 28966 6010 29022 6012
rect 28726 5958 28772 6010
rect 28772 5958 28782 6010
rect 28806 5958 28836 6010
rect 28836 5958 28848 6010
rect 28848 5958 28862 6010
rect 28886 5958 28900 6010
rect 28900 5958 28912 6010
rect 28912 5958 28942 6010
rect 28966 5958 28976 6010
rect 28976 5958 29022 6010
rect 28726 5956 28782 5958
rect 28806 5956 28862 5958
rect 28886 5956 28942 5958
rect 28966 5956 29022 5958
rect 28726 4922 28782 4924
rect 28806 4922 28862 4924
rect 28886 4922 28942 4924
rect 28966 4922 29022 4924
rect 28726 4870 28772 4922
rect 28772 4870 28782 4922
rect 28806 4870 28836 4922
rect 28836 4870 28848 4922
rect 28848 4870 28862 4922
rect 28886 4870 28900 4922
rect 28900 4870 28912 4922
rect 28912 4870 28942 4922
rect 28966 4870 28976 4922
rect 28976 4870 29022 4922
rect 28726 4868 28782 4870
rect 28806 4868 28862 4870
rect 28886 4868 28942 4870
rect 28966 4868 29022 4870
rect 28726 3834 28782 3836
rect 28806 3834 28862 3836
rect 28886 3834 28942 3836
rect 28966 3834 29022 3836
rect 28726 3782 28772 3834
rect 28772 3782 28782 3834
rect 28806 3782 28836 3834
rect 28836 3782 28848 3834
rect 28848 3782 28862 3834
rect 28886 3782 28900 3834
rect 28900 3782 28912 3834
rect 28912 3782 28942 3834
rect 28966 3782 28976 3834
rect 28976 3782 29022 3834
rect 28726 3780 28782 3782
rect 28806 3780 28862 3782
rect 28886 3780 28942 3782
rect 28966 3780 29022 3782
rect 28726 2746 28782 2748
rect 28806 2746 28862 2748
rect 28886 2746 28942 2748
rect 28966 2746 29022 2748
rect 28726 2694 28772 2746
rect 28772 2694 28782 2746
rect 28806 2694 28836 2746
rect 28836 2694 28848 2746
rect 28848 2694 28862 2746
rect 28886 2694 28900 2746
rect 28900 2694 28912 2746
rect 28912 2694 28942 2746
rect 28966 2694 28976 2746
rect 28976 2694 29022 2746
rect 28726 2692 28782 2694
rect 28806 2692 28862 2694
rect 28886 2692 28942 2694
rect 28966 2692 29022 2694
rect 34280 8730 34336 8732
rect 34360 8730 34416 8732
rect 34440 8730 34496 8732
rect 34520 8730 34576 8732
rect 34280 8678 34326 8730
rect 34326 8678 34336 8730
rect 34360 8678 34390 8730
rect 34390 8678 34402 8730
rect 34402 8678 34416 8730
rect 34440 8678 34454 8730
rect 34454 8678 34466 8730
rect 34466 8678 34496 8730
rect 34520 8678 34530 8730
rect 34530 8678 34576 8730
rect 34280 8676 34336 8678
rect 34360 8676 34416 8678
rect 34440 8676 34496 8678
rect 34520 8676 34576 8678
rect 34794 9016 34850 9072
rect 34280 7642 34336 7644
rect 34360 7642 34416 7644
rect 34440 7642 34496 7644
rect 34520 7642 34576 7644
rect 34280 7590 34326 7642
rect 34326 7590 34336 7642
rect 34360 7590 34390 7642
rect 34390 7590 34402 7642
rect 34402 7590 34416 7642
rect 34440 7590 34454 7642
rect 34454 7590 34466 7642
rect 34466 7590 34496 7642
rect 34520 7590 34530 7642
rect 34530 7590 34576 7642
rect 34280 7588 34336 7590
rect 34360 7588 34416 7590
rect 34440 7588 34496 7590
rect 34520 7588 34576 7590
rect 34280 6554 34336 6556
rect 34360 6554 34416 6556
rect 34440 6554 34496 6556
rect 34520 6554 34576 6556
rect 34280 6502 34326 6554
rect 34326 6502 34336 6554
rect 34360 6502 34390 6554
rect 34390 6502 34402 6554
rect 34402 6502 34416 6554
rect 34440 6502 34454 6554
rect 34454 6502 34466 6554
rect 34466 6502 34496 6554
rect 34520 6502 34530 6554
rect 34530 6502 34576 6554
rect 34280 6500 34336 6502
rect 34360 6500 34416 6502
rect 34440 6500 34496 6502
rect 34520 6500 34576 6502
rect 34280 5466 34336 5468
rect 34360 5466 34416 5468
rect 34440 5466 34496 5468
rect 34520 5466 34576 5468
rect 34280 5414 34326 5466
rect 34326 5414 34336 5466
rect 34360 5414 34390 5466
rect 34390 5414 34402 5466
rect 34402 5414 34416 5466
rect 34440 5414 34454 5466
rect 34454 5414 34466 5466
rect 34466 5414 34496 5466
rect 34520 5414 34530 5466
rect 34530 5414 34576 5466
rect 34280 5412 34336 5414
rect 34360 5412 34416 5414
rect 34440 5412 34496 5414
rect 34520 5412 34576 5414
rect 34280 4378 34336 4380
rect 34360 4378 34416 4380
rect 34440 4378 34496 4380
rect 34520 4378 34576 4380
rect 34280 4326 34326 4378
rect 34326 4326 34336 4378
rect 34360 4326 34390 4378
rect 34390 4326 34402 4378
rect 34402 4326 34416 4378
rect 34440 4326 34454 4378
rect 34454 4326 34466 4378
rect 34466 4326 34496 4378
rect 34520 4326 34530 4378
rect 34530 4326 34576 4378
rect 34280 4324 34336 4326
rect 34360 4324 34416 4326
rect 34440 4324 34496 4326
rect 34520 4324 34576 4326
rect 35898 7384 35954 7440
rect 34280 3290 34336 3292
rect 34360 3290 34416 3292
rect 34440 3290 34496 3292
rect 34520 3290 34576 3292
rect 34280 3238 34326 3290
rect 34326 3238 34336 3290
rect 34360 3238 34390 3290
rect 34390 3238 34402 3290
rect 34402 3238 34416 3290
rect 34440 3238 34454 3290
rect 34454 3238 34466 3290
rect 34466 3238 34496 3290
rect 34520 3238 34530 3290
rect 34530 3238 34576 3290
rect 34280 3236 34336 3238
rect 34360 3236 34416 3238
rect 34440 3236 34496 3238
rect 34520 3236 34576 3238
rect 23172 2202 23228 2204
rect 23252 2202 23308 2204
rect 23332 2202 23388 2204
rect 23412 2202 23468 2204
rect 23172 2150 23218 2202
rect 23218 2150 23228 2202
rect 23252 2150 23282 2202
rect 23282 2150 23294 2202
rect 23294 2150 23308 2202
rect 23332 2150 23346 2202
rect 23346 2150 23358 2202
rect 23358 2150 23388 2202
rect 23412 2150 23422 2202
rect 23422 2150 23468 2202
rect 23172 2148 23228 2150
rect 23252 2148 23308 2150
rect 23332 2148 23388 2150
rect 23412 2148 23468 2150
rect 34280 2202 34336 2204
rect 34360 2202 34416 2204
rect 34440 2202 34496 2204
rect 34520 2202 34576 2204
rect 34280 2150 34326 2202
rect 34326 2150 34336 2202
rect 34360 2150 34390 2202
rect 34390 2150 34402 2202
rect 34402 2150 34416 2202
rect 34440 2150 34454 2202
rect 34454 2150 34466 2202
rect 34466 2150 34496 2202
rect 34520 2150 34530 2202
rect 34530 2150 34576 2202
rect 34280 2148 34336 2150
rect 34360 2148 34416 2150
rect 34440 2148 34496 2150
rect 34520 2148 34576 2150
rect 37462 7928 37518 7984
rect 39834 8186 39890 8188
rect 39914 8186 39970 8188
rect 39994 8186 40050 8188
rect 40074 8186 40130 8188
rect 39834 8134 39880 8186
rect 39880 8134 39890 8186
rect 39914 8134 39944 8186
rect 39944 8134 39956 8186
rect 39956 8134 39970 8186
rect 39994 8134 40008 8186
rect 40008 8134 40020 8186
rect 40020 8134 40050 8186
rect 40074 8134 40084 8186
rect 40084 8134 40130 8186
rect 39834 8132 39890 8134
rect 39914 8132 39970 8134
rect 39994 8132 40050 8134
rect 40074 8132 40130 8134
rect 39834 7098 39890 7100
rect 39914 7098 39970 7100
rect 39994 7098 40050 7100
rect 40074 7098 40130 7100
rect 39834 7046 39880 7098
rect 39880 7046 39890 7098
rect 39914 7046 39944 7098
rect 39944 7046 39956 7098
rect 39956 7046 39970 7098
rect 39994 7046 40008 7098
rect 40008 7046 40020 7098
rect 40020 7046 40050 7098
rect 40074 7046 40084 7098
rect 40084 7046 40130 7098
rect 39834 7044 39890 7046
rect 39914 7044 39970 7046
rect 39994 7044 40050 7046
rect 40074 7044 40130 7046
rect 39834 6010 39890 6012
rect 39914 6010 39970 6012
rect 39994 6010 40050 6012
rect 40074 6010 40130 6012
rect 39834 5958 39880 6010
rect 39880 5958 39890 6010
rect 39914 5958 39944 6010
rect 39944 5958 39956 6010
rect 39956 5958 39970 6010
rect 39994 5958 40008 6010
rect 40008 5958 40020 6010
rect 40020 5958 40050 6010
rect 40074 5958 40084 6010
rect 40084 5958 40130 6010
rect 39834 5956 39890 5958
rect 39914 5956 39970 5958
rect 39994 5956 40050 5958
rect 40074 5956 40130 5958
rect 39834 4922 39890 4924
rect 39914 4922 39970 4924
rect 39994 4922 40050 4924
rect 40074 4922 40130 4924
rect 39834 4870 39880 4922
rect 39880 4870 39890 4922
rect 39914 4870 39944 4922
rect 39944 4870 39956 4922
rect 39956 4870 39970 4922
rect 39994 4870 40008 4922
rect 40008 4870 40020 4922
rect 40020 4870 40050 4922
rect 40074 4870 40084 4922
rect 40084 4870 40130 4922
rect 39834 4868 39890 4870
rect 39914 4868 39970 4870
rect 39994 4868 40050 4870
rect 40074 4868 40130 4870
rect 39834 3834 39890 3836
rect 39914 3834 39970 3836
rect 39994 3834 40050 3836
rect 40074 3834 40130 3836
rect 39834 3782 39880 3834
rect 39880 3782 39890 3834
rect 39914 3782 39944 3834
rect 39944 3782 39956 3834
rect 39956 3782 39970 3834
rect 39994 3782 40008 3834
rect 40008 3782 40020 3834
rect 40020 3782 40050 3834
rect 40074 3782 40084 3834
rect 40084 3782 40130 3834
rect 39834 3780 39890 3782
rect 39914 3780 39970 3782
rect 39994 3780 40050 3782
rect 40074 3780 40130 3782
rect 39834 2746 39890 2748
rect 39914 2746 39970 2748
rect 39994 2746 40050 2748
rect 40074 2746 40130 2748
rect 39834 2694 39880 2746
rect 39880 2694 39890 2746
rect 39914 2694 39944 2746
rect 39944 2694 39956 2746
rect 39956 2694 39970 2746
rect 39994 2694 40008 2746
rect 40008 2694 40020 2746
rect 40020 2694 40050 2746
rect 40074 2694 40084 2746
rect 40084 2694 40130 2746
rect 39834 2692 39890 2694
rect 39914 2692 39970 2694
rect 39994 2692 40050 2694
rect 40074 2692 40130 2694
rect 45388 8730 45444 8732
rect 45468 8730 45524 8732
rect 45548 8730 45604 8732
rect 45628 8730 45684 8732
rect 45388 8678 45434 8730
rect 45434 8678 45444 8730
rect 45468 8678 45498 8730
rect 45498 8678 45510 8730
rect 45510 8678 45524 8730
rect 45548 8678 45562 8730
rect 45562 8678 45574 8730
rect 45574 8678 45604 8730
rect 45628 8678 45638 8730
rect 45638 8678 45684 8730
rect 45388 8676 45444 8678
rect 45468 8676 45524 8678
rect 45548 8676 45604 8678
rect 45628 8676 45684 8678
rect 45388 7642 45444 7644
rect 45468 7642 45524 7644
rect 45548 7642 45604 7644
rect 45628 7642 45684 7644
rect 45388 7590 45434 7642
rect 45434 7590 45444 7642
rect 45468 7590 45498 7642
rect 45498 7590 45510 7642
rect 45510 7590 45524 7642
rect 45548 7590 45562 7642
rect 45562 7590 45574 7642
rect 45574 7590 45604 7642
rect 45628 7590 45638 7642
rect 45638 7590 45684 7642
rect 45388 7588 45444 7590
rect 45468 7588 45524 7590
rect 45548 7588 45604 7590
rect 45628 7588 45684 7590
rect 45388 6554 45444 6556
rect 45468 6554 45524 6556
rect 45548 6554 45604 6556
rect 45628 6554 45684 6556
rect 45388 6502 45434 6554
rect 45434 6502 45444 6554
rect 45468 6502 45498 6554
rect 45498 6502 45510 6554
rect 45510 6502 45524 6554
rect 45548 6502 45562 6554
rect 45562 6502 45574 6554
rect 45574 6502 45604 6554
rect 45628 6502 45638 6554
rect 45638 6502 45684 6554
rect 45388 6500 45444 6502
rect 45468 6500 45524 6502
rect 45548 6500 45604 6502
rect 45628 6500 45684 6502
rect 45388 5466 45444 5468
rect 45468 5466 45524 5468
rect 45548 5466 45604 5468
rect 45628 5466 45684 5468
rect 45388 5414 45434 5466
rect 45434 5414 45444 5466
rect 45468 5414 45498 5466
rect 45498 5414 45510 5466
rect 45510 5414 45524 5466
rect 45548 5414 45562 5466
rect 45562 5414 45574 5466
rect 45574 5414 45604 5466
rect 45628 5414 45638 5466
rect 45638 5414 45684 5466
rect 45388 5412 45444 5414
rect 45468 5412 45524 5414
rect 45548 5412 45604 5414
rect 45628 5412 45684 5414
rect 45388 4378 45444 4380
rect 45468 4378 45524 4380
rect 45548 4378 45604 4380
rect 45628 4378 45684 4380
rect 45388 4326 45434 4378
rect 45434 4326 45444 4378
rect 45468 4326 45498 4378
rect 45498 4326 45510 4378
rect 45510 4326 45524 4378
rect 45548 4326 45562 4378
rect 45562 4326 45574 4378
rect 45574 4326 45604 4378
rect 45628 4326 45638 4378
rect 45638 4326 45684 4378
rect 45388 4324 45444 4326
rect 45468 4324 45524 4326
rect 45548 4324 45604 4326
rect 45628 4324 45684 4326
rect 45388 3290 45444 3292
rect 45468 3290 45524 3292
rect 45548 3290 45604 3292
rect 45628 3290 45684 3292
rect 45388 3238 45434 3290
rect 45434 3238 45444 3290
rect 45468 3238 45498 3290
rect 45498 3238 45510 3290
rect 45510 3238 45524 3290
rect 45548 3238 45562 3290
rect 45562 3238 45574 3290
rect 45574 3238 45604 3290
rect 45628 3238 45638 3290
rect 45638 3238 45684 3290
rect 45388 3236 45444 3238
rect 45468 3236 45524 3238
rect 45548 3236 45604 3238
rect 45628 3236 45684 3238
rect 45388 2202 45444 2204
rect 45468 2202 45524 2204
rect 45548 2202 45604 2204
rect 45628 2202 45684 2204
rect 45388 2150 45434 2202
rect 45434 2150 45444 2202
rect 45468 2150 45498 2202
rect 45498 2150 45510 2202
rect 45510 2150 45524 2202
rect 45548 2150 45562 2202
rect 45562 2150 45574 2202
rect 45574 2150 45604 2202
rect 45628 2150 45638 2202
rect 45638 2150 45684 2202
rect 45388 2148 45444 2150
rect 45468 2148 45524 2150
rect 45548 2148 45604 2150
rect 45628 2148 45684 2150
rect 23172 1114 23228 1116
rect 23252 1114 23308 1116
rect 23332 1114 23388 1116
rect 23412 1114 23468 1116
rect 23172 1062 23218 1114
rect 23218 1062 23228 1114
rect 23252 1062 23282 1114
rect 23282 1062 23294 1114
rect 23294 1062 23308 1114
rect 23332 1062 23346 1114
rect 23346 1062 23358 1114
rect 23358 1062 23388 1114
rect 23412 1062 23422 1114
rect 23422 1062 23468 1114
rect 23172 1060 23228 1062
rect 23252 1060 23308 1062
rect 23332 1060 23388 1062
rect 23412 1060 23468 1062
rect 28726 1658 28782 1660
rect 28806 1658 28862 1660
rect 28886 1658 28942 1660
rect 28966 1658 29022 1660
rect 28726 1606 28772 1658
rect 28772 1606 28782 1658
rect 28806 1606 28836 1658
rect 28836 1606 28848 1658
rect 28848 1606 28862 1658
rect 28886 1606 28900 1658
rect 28900 1606 28912 1658
rect 28912 1606 28942 1658
rect 28966 1606 28976 1658
rect 28976 1606 29022 1658
rect 28726 1604 28782 1606
rect 28806 1604 28862 1606
rect 28886 1604 28942 1606
rect 28966 1604 29022 1606
rect 39834 1658 39890 1660
rect 39914 1658 39970 1660
rect 39994 1658 40050 1660
rect 40074 1658 40130 1660
rect 39834 1606 39880 1658
rect 39880 1606 39890 1658
rect 39914 1606 39944 1658
rect 39944 1606 39956 1658
rect 39956 1606 39970 1658
rect 39994 1606 40008 1658
rect 40008 1606 40020 1658
rect 40020 1606 40050 1658
rect 40074 1606 40084 1658
rect 40084 1606 40130 1658
rect 39834 1604 39890 1606
rect 39914 1604 39970 1606
rect 39994 1604 40050 1606
rect 40074 1604 40130 1606
rect 34280 1114 34336 1116
rect 34360 1114 34416 1116
rect 34440 1114 34496 1116
rect 34520 1114 34576 1116
rect 34280 1062 34326 1114
rect 34326 1062 34336 1114
rect 34360 1062 34390 1114
rect 34390 1062 34402 1114
rect 34402 1062 34416 1114
rect 34440 1062 34454 1114
rect 34454 1062 34466 1114
rect 34466 1062 34496 1114
rect 34520 1062 34530 1114
rect 34530 1062 34576 1114
rect 34280 1060 34336 1062
rect 34360 1060 34416 1062
rect 34440 1060 34496 1062
rect 34520 1060 34576 1062
rect 45388 1114 45444 1116
rect 45468 1114 45524 1116
rect 45548 1114 45604 1116
rect 45628 1114 45684 1116
rect 45388 1062 45434 1114
rect 45434 1062 45444 1114
rect 45468 1062 45498 1114
rect 45498 1062 45510 1114
rect 45510 1062 45524 1114
rect 45548 1062 45562 1114
rect 45562 1062 45574 1114
rect 45574 1062 45604 1114
rect 45628 1062 45638 1114
rect 45638 1062 45684 1114
rect 45388 1060 45444 1062
rect 45468 1060 45524 1062
rect 45548 1060 45604 1062
rect 45628 1060 45684 1062
<< metal3 >>
rect 14365 9890 14431 9893
rect 16389 9890 16455 9893
rect 14365 9888 16455 9890
rect 14365 9832 14370 9888
rect 14426 9832 16394 9888
rect 16450 9832 16455 9888
rect 14365 9830 16455 9832
rect 14365 9827 14431 9830
rect 16389 9827 16455 9830
rect 19885 9890 19951 9893
rect 23933 9890 23999 9893
rect 19885 9888 23999 9890
rect 19885 9832 19890 9888
rect 19946 9832 23938 9888
rect 23994 9832 23999 9888
rect 19885 9830 23999 9832
rect 19885 9827 19951 9830
rect 23933 9827 23999 9830
rect 14549 9754 14615 9757
rect 16481 9754 16547 9757
rect 14549 9752 16547 9754
rect 14549 9696 14554 9752
rect 14610 9696 16486 9752
rect 16542 9696 16547 9752
rect 14549 9694 16547 9696
rect 14549 9691 14615 9694
rect 16481 9691 16547 9694
rect 18321 9754 18387 9757
rect 21173 9754 21239 9757
rect 18321 9752 21239 9754
rect 18321 9696 18326 9752
rect 18382 9696 21178 9752
rect 21234 9696 21239 9752
rect 18321 9694 21239 9696
rect 18321 9691 18387 9694
rect 21173 9691 21239 9694
rect 13629 9618 13695 9621
rect 21173 9618 21239 9621
rect 13629 9616 21239 9618
rect 13629 9560 13634 9616
rect 13690 9560 21178 9616
rect 21234 9560 21239 9616
rect 13629 9558 21239 9560
rect 13629 9555 13695 9558
rect 21173 9555 21239 9558
rect 16757 9482 16823 9485
rect 19374 9482 19380 9484
rect 16757 9480 19380 9482
rect 16757 9424 16762 9480
rect 16818 9424 19380 9480
rect 16757 9422 19380 9424
rect 16757 9419 16823 9422
rect 19374 9420 19380 9422
rect 19444 9420 19450 9484
rect 20161 9482 20227 9485
rect 27613 9482 27679 9485
rect 20161 9480 27679 9482
rect 20161 9424 20166 9480
rect 20222 9424 27618 9480
rect 27674 9424 27679 9480
rect 20161 9422 27679 9424
rect 20161 9419 20227 9422
rect 27613 9419 27679 9422
rect 17125 9346 17191 9349
rect 20805 9346 20871 9349
rect 17125 9344 20871 9346
rect 17125 9288 17130 9344
rect 17186 9288 20810 9344
rect 20866 9288 20871 9344
rect 17125 9286 20871 9288
rect 17125 9283 17191 9286
rect 20805 9283 20871 9286
rect 23657 9346 23723 9349
rect 24301 9346 24367 9349
rect 23657 9344 24367 9346
rect 23657 9288 23662 9344
rect 23718 9288 24306 9344
rect 24362 9288 24367 9344
rect 23657 9286 24367 9288
rect 23657 9283 23723 9286
rect 24301 9283 24367 9286
rect 14365 9210 14431 9213
rect 28441 9210 28507 9213
rect 14365 9208 28507 9210
rect 14365 9152 14370 9208
rect 14426 9152 28446 9208
rect 28502 9152 28507 9208
rect 14365 9150 28507 9152
rect 14365 9147 14431 9150
rect 28441 9147 28507 9150
rect 17953 9074 18019 9077
rect 34789 9074 34855 9077
rect 17953 9072 34855 9074
rect 17953 9016 17958 9072
rect 18014 9016 34794 9072
rect 34850 9016 34855 9072
rect 17953 9014 34855 9016
rect 17953 9011 18019 9014
rect 34789 9011 34855 9014
rect 12433 8938 12499 8941
rect 25221 8938 25287 8941
rect 12433 8936 25287 8938
rect 12433 8880 12438 8936
rect 12494 8880 25226 8936
rect 25282 8880 25287 8936
rect 12433 8878 25287 8880
rect 12433 8875 12499 8878
rect 25221 8875 25287 8878
rect 12054 8736 12370 8737
rect 12054 8672 12060 8736
rect 12124 8672 12140 8736
rect 12204 8672 12220 8736
rect 12284 8672 12300 8736
rect 12364 8672 12370 8736
rect 12054 8671 12370 8672
rect 23162 8736 23478 8737
rect 23162 8672 23168 8736
rect 23232 8672 23248 8736
rect 23312 8672 23328 8736
rect 23392 8672 23408 8736
rect 23472 8672 23478 8736
rect 23162 8671 23478 8672
rect 34270 8736 34586 8737
rect 34270 8672 34276 8736
rect 34340 8672 34356 8736
rect 34420 8672 34436 8736
rect 34500 8672 34516 8736
rect 34580 8672 34586 8736
rect 34270 8671 34586 8672
rect 45378 8736 45694 8737
rect 45378 8672 45384 8736
rect 45448 8672 45464 8736
rect 45528 8672 45544 8736
rect 45608 8672 45624 8736
rect 45688 8672 45694 8736
rect 45378 8671 45694 8672
rect 23841 8666 23907 8669
rect 28257 8666 28323 8669
rect 23841 8664 28323 8666
rect 23841 8608 23846 8664
rect 23902 8608 28262 8664
rect 28318 8608 28323 8664
rect 23841 8606 28323 8608
rect 23841 8603 23907 8606
rect 28257 8603 28323 8606
rect 22461 8530 22527 8533
rect 24485 8530 24551 8533
rect 22461 8528 24551 8530
rect 22461 8472 22466 8528
rect 22522 8472 24490 8528
rect 24546 8472 24551 8528
rect 22461 8470 24551 8472
rect 22461 8467 22527 8470
rect 24485 8467 24551 8470
rect 16113 8394 16179 8397
rect 20805 8394 20871 8397
rect 22829 8394 22895 8397
rect 16113 8392 20871 8394
rect 16113 8336 16118 8392
rect 16174 8336 20810 8392
rect 20866 8336 20871 8392
rect 16113 8334 20871 8336
rect 16113 8331 16179 8334
rect 20805 8331 20871 8334
rect 21038 8392 22895 8394
rect 21038 8336 22834 8392
rect 22890 8336 22895 8392
rect 21038 8334 22895 8336
rect 18781 8258 18847 8261
rect 21038 8258 21098 8334
rect 22829 8331 22895 8334
rect 23197 8394 23263 8397
rect 28533 8394 28599 8397
rect 23197 8392 28599 8394
rect 23197 8336 23202 8392
rect 23258 8336 28538 8392
rect 28594 8336 28599 8392
rect 23197 8334 28599 8336
rect 23197 8331 23263 8334
rect 28533 8331 28599 8334
rect 18781 8256 21098 8258
rect 18781 8200 18786 8256
rect 18842 8200 21098 8256
rect 18781 8198 21098 8200
rect 21265 8258 21331 8261
rect 24577 8258 24643 8261
rect 21265 8256 24643 8258
rect 21265 8200 21270 8256
rect 21326 8200 24582 8256
rect 24638 8200 24643 8256
rect 21265 8198 24643 8200
rect 18781 8195 18847 8198
rect 21265 8195 21331 8198
rect 24577 8195 24643 8198
rect 6500 8192 6816 8193
rect 6500 8128 6506 8192
rect 6570 8128 6586 8192
rect 6650 8128 6666 8192
rect 6730 8128 6746 8192
rect 6810 8128 6816 8192
rect 6500 8127 6816 8128
rect 17608 8192 17924 8193
rect 17608 8128 17614 8192
rect 17678 8128 17694 8192
rect 17758 8128 17774 8192
rect 17838 8128 17854 8192
rect 17918 8128 17924 8192
rect 17608 8127 17924 8128
rect 28716 8192 29032 8193
rect 28716 8128 28722 8192
rect 28786 8128 28802 8192
rect 28866 8128 28882 8192
rect 28946 8128 28962 8192
rect 29026 8128 29032 8192
rect 28716 8127 29032 8128
rect 39824 8192 40140 8193
rect 39824 8128 39830 8192
rect 39894 8128 39910 8192
rect 39974 8128 39990 8192
rect 40054 8128 40070 8192
rect 40134 8128 40140 8192
rect 39824 8127 40140 8128
rect 18045 8122 18111 8125
rect 23473 8122 23539 8125
rect 18045 8120 23539 8122
rect 18045 8064 18050 8120
rect 18106 8064 23478 8120
rect 23534 8064 23539 8120
rect 18045 8062 23539 8064
rect 18045 8059 18111 8062
rect 23473 8059 23539 8062
rect 23933 8122 23999 8125
rect 24761 8122 24827 8125
rect 23933 8120 24827 8122
rect 23933 8064 23938 8120
rect 23994 8064 24766 8120
rect 24822 8064 24827 8120
rect 23933 8062 24827 8064
rect 23933 8059 23999 8062
rect 24761 8059 24827 8062
rect 17953 7986 18019 7989
rect 21265 7986 21331 7989
rect 17953 7984 21331 7986
rect 17953 7928 17958 7984
rect 18014 7928 21270 7984
rect 21326 7928 21331 7984
rect 17953 7926 21331 7928
rect 17953 7923 18019 7926
rect 21265 7923 21331 7926
rect 22001 7986 22067 7989
rect 37457 7986 37523 7989
rect 22001 7984 37523 7986
rect 22001 7928 22006 7984
rect 22062 7928 37462 7984
rect 37518 7928 37523 7984
rect 22001 7926 37523 7928
rect 22001 7923 22067 7926
rect 37457 7923 37523 7926
rect 15101 7850 15167 7853
rect 28165 7850 28231 7853
rect 15101 7848 28231 7850
rect 15101 7792 15106 7848
rect 15162 7792 28170 7848
rect 28226 7792 28231 7848
rect 15101 7790 28231 7792
rect 15101 7787 15167 7790
rect 28165 7787 28231 7790
rect 17217 7714 17283 7717
rect 21633 7714 21699 7717
rect 17217 7712 21699 7714
rect 17217 7656 17222 7712
rect 17278 7656 21638 7712
rect 21694 7656 21699 7712
rect 17217 7654 21699 7656
rect 17217 7651 17283 7654
rect 21633 7651 21699 7654
rect 12054 7648 12370 7649
rect 12054 7584 12060 7648
rect 12124 7584 12140 7648
rect 12204 7584 12220 7648
rect 12284 7584 12300 7648
rect 12364 7584 12370 7648
rect 12054 7583 12370 7584
rect 23162 7648 23478 7649
rect 23162 7584 23168 7648
rect 23232 7584 23248 7648
rect 23312 7584 23328 7648
rect 23392 7584 23408 7648
rect 23472 7584 23478 7648
rect 23162 7583 23478 7584
rect 34270 7648 34586 7649
rect 34270 7584 34276 7648
rect 34340 7584 34356 7648
rect 34420 7584 34436 7648
rect 34500 7584 34516 7648
rect 34580 7584 34586 7648
rect 34270 7583 34586 7584
rect 45378 7648 45694 7649
rect 45378 7584 45384 7648
rect 45448 7584 45464 7648
rect 45528 7584 45544 7648
rect 45608 7584 45624 7648
rect 45688 7584 45694 7648
rect 45378 7583 45694 7584
rect 15101 7578 15167 7581
rect 18781 7578 18847 7581
rect 15101 7576 18847 7578
rect 15101 7520 15106 7576
rect 15162 7520 18786 7576
rect 18842 7520 18847 7576
rect 15101 7518 18847 7520
rect 15101 7515 15167 7518
rect 18781 7515 18847 7518
rect 11513 7442 11579 7445
rect 16941 7442 17007 7445
rect 22093 7442 22159 7445
rect 11513 7440 16866 7442
rect 11513 7384 11518 7440
rect 11574 7384 16866 7440
rect 11513 7382 16866 7384
rect 11513 7379 11579 7382
rect 16806 7306 16866 7382
rect 16941 7440 22159 7442
rect 16941 7384 16946 7440
rect 17002 7384 22098 7440
rect 22154 7384 22159 7440
rect 16941 7382 22159 7384
rect 16941 7379 17007 7382
rect 22093 7379 22159 7382
rect 22921 7442 22987 7445
rect 35893 7442 35959 7445
rect 22921 7440 35959 7442
rect 22921 7384 22926 7440
rect 22982 7384 35898 7440
rect 35954 7384 35959 7440
rect 22921 7382 35959 7384
rect 22921 7379 22987 7382
rect 35893 7379 35959 7382
rect 21725 7306 21791 7309
rect 32949 7306 33015 7309
rect 16806 7246 18108 7306
rect 6500 7104 6816 7105
rect 6500 7040 6506 7104
rect 6570 7040 6586 7104
rect 6650 7040 6666 7104
rect 6730 7040 6746 7104
rect 6810 7040 6816 7104
rect 6500 7039 6816 7040
rect 17608 7104 17924 7105
rect 17608 7040 17614 7104
rect 17678 7040 17694 7104
rect 17758 7040 17774 7104
rect 17838 7040 17854 7104
rect 17918 7040 17924 7104
rect 17608 7039 17924 7040
rect 18048 7034 18108 7246
rect 21725 7304 33015 7306
rect 21725 7248 21730 7304
rect 21786 7248 32954 7304
rect 33010 7248 33015 7304
rect 21725 7246 33015 7248
rect 21725 7243 21791 7246
rect 32949 7243 33015 7246
rect 19374 7108 19380 7172
rect 19444 7170 19450 7172
rect 23197 7170 23263 7173
rect 19444 7168 23263 7170
rect 19444 7112 23202 7168
rect 23258 7112 23263 7168
rect 19444 7110 23263 7112
rect 19444 7108 19450 7110
rect 23197 7107 23263 7110
rect 28716 7104 29032 7105
rect 28716 7040 28722 7104
rect 28786 7040 28802 7104
rect 28866 7040 28882 7104
rect 28946 7040 28962 7104
rect 29026 7040 29032 7104
rect 28716 7039 29032 7040
rect 39824 7104 40140 7105
rect 39824 7040 39830 7104
rect 39894 7040 39910 7104
rect 39974 7040 39990 7104
rect 40054 7040 40070 7104
rect 40134 7040 40140 7104
rect 39824 7039 40140 7040
rect 28441 7034 28507 7037
rect 18048 7032 28507 7034
rect 18048 6976 28446 7032
rect 28502 6976 28507 7032
rect 18048 6974 28507 6976
rect 28441 6971 28507 6974
rect 5441 6898 5507 6901
rect 26233 6898 26299 6901
rect 5441 6896 26299 6898
rect 5441 6840 5446 6896
rect 5502 6840 26238 6896
rect 26294 6840 26299 6896
rect 5441 6838 26299 6840
rect 5441 6835 5507 6838
rect 26233 6835 26299 6838
rect 12617 6762 12683 6765
rect 25957 6762 26023 6765
rect 12617 6760 26023 6762
rect 12617 6704 12622 6760
rect 12678 6704 25962 6760
rect 26018 6704 26023 6760
rect 12617 6702 26023 6704
rect 12617 6699 12683 6702
rect 25957 6699 26023 6702
rect 12054 6560 12370 6561
rect 12054 6496 12060 6560
rect 12124 6496 12140 6560
rect 12204 6496 12220 6560
rect 12284 6496 12300 6560
rect 12364 6496 12370 6560
rect 12054 6495 12370 6496
rect 23162 6560 23478 6561
rect 23162 6496 23168 6560
rect 23232 6496 23248 6560
rect 23312 6496 23328 6560
rect 23392 6496 23408 6560
rect 23472 6496 23478 6560
rect 23162 6495 23478 6496
rect 34270 6560 34586 6561
rect 34270 6496 34276 6560
rect 34340 6496 34356 6560
rect 34420 6496 34436 6560
rect 34500 6496 34516 6560
rect 34580 6496 34586 6560
rect 34270 6495 34586 6496
rect 45378 6560 45694 6561
rect 45378 6496 45384 6560
rect 45448 6496 45464 6560
rect 45528 6496 45544 6560
rect 45608 6496 45624 6560
rect 45688 6496 45694 6560
rect 45378 6495 45694 6496
rect 6500 6016 6816 6017
rect 6500 5952 6506 6016
rect 6570 5952 6586 6016
rect 6650 5952 6666 6016
rect 6730 5952 6746 6016
rect 6810 5952 6816 6016
rect 6500 5951 6816 5952
rect 17608 6016 17924 6017
rect 17608 5952 17614 6016
rect 17678 5952 17694 6016
rect 17758 5952 17774 6016
rect 17838 5952 17854 6016
rect 17918 5952 17924 6016
rect 17608 5951 17924 5952
rect 28716 6016 29032 6017
rect 28716 5952 28722 6016
rect 28786 5952 28802 6016
rect 28866 5952 28882 6016
rect 28946 5952 28962 6016
rect 29026 5952 29032 6016
rect 28716 5951 29032 5952
rect 39824 6016 40140 6017
rect 39824 5952 39830 6016
rect 39894 5952 39910 6016
rect 39974 5952 39990 6016
rect 40054 5952 40070 6016
rect 40134 5952 40140 6016
rect 39824 5951 40140 5952
rect 12054 5472 12370 5473
rect 12054 5408 12060 5472
rect 12124 5408 12140 5472
rect 12204 5408 12220 5472
rect 12284 5408 12300 5472
rect 12364 5408 12370 5472
rect 12054 5407 12370 5408
rect 23162 5472 23478 5473
rect 23162 5408 23168 5472
rect 23232 5408 23248 5472
rect 23312 5408 23328 5472
rect 23392 5408 23408 5472
rect 23472 5408 23478 5472
rect 23162 5407 23478 5408
rect 34270 5472 34586 5473
rect 34270 5408 34276 5472
rect 34340 5408 34356 5472
rect 34420 5408 34436 5472
rect 34500 5408 34516 5472
rect 34580 5408 34586 5472
rect 34270 5407 34586 5408
rect 45378 5472 45694 5473
rect 45378 5408 45384 5472
rect 45448 5408 45464 5472
rect 45528 5408 45544 5472
rect 45608 5408 45624 5472
rect 45688 5408 45694 5472
rect 45378 5407 45694 5408
rect 6500 4928 6816 4929
rect 6500 4864 6506 4928
rect 6570 4864 6586 4928
rect 6650 4864 6666 4928
rect 6730 4864 6746 4928
rect 6810 4864 6816 4928
rect 6500 4863 6816 4864
rect 17608 4928 17924 4929
rect 17608 4864 17614 4928
rect 17678 4864 17694 4928
rect 17758 4864 17774 4928
rect 17838 4864 17854 4928
rect 17918 4864 17924 4928
rect 17608 4863 17924 4864
rect 28716 4928 29032 4929
rect 28716 4864 28722 4928
rect 28786 4864 28802 4928
rect 28866 4864 28882 4928
rect 28946 4864 28962 4928
rect 29026 4864 29032 4928
rect 28716 4863 29032 4864
rect 39824 4928 40140 4929
rect 39824 4864 39830 4928
rect 39894 4864 39910 4928
rect 39974 4864 39990 4928
rect 40054 4864 40070 4928
rect 40134 4864 40140 4928
rect 39824 4863 40140 4864
rect 12054 4384 12370 4385
rect 12054 4320 12060 4384
rect 12124 4320 12140 4384
rect 12204 4320 12220 4384
rect 12284 4320 12300 4384
rect 12364 4320 12370 4384
rect 12054 4319 12370 4320
rect 23162 4384 23478 4385
rect 23162 4320 23168 4384
rect 23232 4320 23248 4384
rect 23312 4320 23328 4384
rect 23392 4320 23408 4384
rect 23472 4320 23478 4384
rect 23162 4319 23478 4320
rect 34270 4384 34586 4385
rect 34270 4320 34276 4384
rect 34340 4320 34356 4384
rect 34420 4320 34436 4384
rect 34500 4320 34516 4384
rect 34580 4320 34586 4384
rect 34270 4319 34586 4320
rect 45378 4384 45694 4385
rect 45378 4320 45384 4384
rect 45448 4320 45464 4384
rect 45528 4320 45544 4384
rect 45608 4320 45624 4384
rect 45688 4320 45694 4384
rect 45378 4319 45694 4320
rect 6500 3840 6816 3841
rect 6500 3776 6506 3840
rect 6570 3776 6586 3840
rect 6650 3776 6666 3840
rect 6730 3776 6746 3840
rect 6810 3776 6816 3840
rect 6500 3775 6816 3776
rect 17608 3840 17924 3841
rect 17608 3776 17614 3840
rect 17678 3776 17694 3840
rect 17758 3776 17774 3840
rect 17838 3776 17854 3840
rect 17918 3776 17924 3840
rect 17608 3775 17924 3776
rect 28716 3840 29032 3841
rect 28716 3776 28722 3840
rect 28786 3776 28802 3840
rect 28866 3776 28882 3840
rect 28946 3776 28962 3840
rect 29026 3776 29032 3840
rect 28716 3775 29032 3776
rect 39824 3840 40140 3841
rect 39824 3776 39830 3840
rect 39894 3776 39910 3840
rect 39974 3776 39990 3840
rect 40054 3776 40070 3840
rect 40134 3776 40140 3840
rect 39824 3775 40140 3776
rect 12054 3296 12370 3297
rect 12054 3232 12060 3296
rect 12124 3232 12140 3296
rect 12204 3232 12220 3296
rect 12284 3232 12300 3296
rect 12364 3232 12370 3296
rect 12054 3231 12370 3232
rect 23162 3296 23478 3297
rect 23162 3232 23168 3296
rect 23232 3232 23248 3296
rect 23312 3232 23328 3296
rect 23392 3232 23408 3296
rect 23472 3232 23478 3296
rect 23162 3231 23478 3232
rect 34270 3296 34586 3297
rect 34270 3232 34276 3296
rect 34340 3232 34356 3296
rect 34420 3232 34436 3296
rect 34500 3232 34516 3296
rect 34580 3232 34586 3296
rect 34270 3231 34586 3232
rect 45378 3296 45694 3297
rect 45378 3232 45384 3296
rect 45448 3232 45464 3296
rect 45528 3232 45544 3296
rect 45608 3232 45624 3296
rect 45688 3232 45694 3296
rect 45378 3231 45694 3232
rect 6500 2752 6816 2753
rect 6500 2688 6506 2752
rect 6570 2688 6586 2752
rect 6650 2688 6666 2752
rect 6730 2688 6746 2752
rect 6810 2688 6816 2752
rect 6500 2687 6816 2688
rect 17608 2752 17924 2753
rect 17608 2688 17614 2752
rect 17678 2688 17694 2752
rect 17758 2688 17774 2752
rect 17838 2688 17854 2752
rect 17918 2688 17924 2752
rect 17608 2687 17924 2688
rect 28716 2752 29032 2753
rect 28716 2688 28722 2752
rect 28786 2688 28802 2752
rect 28866 2688 28882 2752
rect 28946 2688 28962 2752
rect 29026 2688 29032 2752
rect 28716 2687 29032 2688
rect 39824 2752 40140 2753
rect 39824 2688 39830 2752
rect 39894 2688 39910 2752
rect 39974 2688 39990 2752
rect 40054 2688 40070 2752
rect 40134 2688 40140 2752
rect 39824 2687 40140 2688
rect 12054 2208 12370 2209
rect 12054 2144 12060 2208
rect 12124 2144 12140 2208
rect 12204 2144 12220 2208
rect 12284 2144 12300 2208
rect 12364 2144 12370 2208
rect 12054 2143 12370 2144
rect 23162 2208 23478 2209
rect 23162 2144 23168 2208
rect 23232 2144 23248 2208
rect 23312 2144 23328 2208
rect 23392 2144 23408 2208
rect 23472 2144 23478 2208
rect 23162 2143 23478 2144
rect 34270 2208 34586 2209
rect 34270 2144 34276 2208
rect 34340 2144 34356 2208
rect 34420 2144 34436 2208
rect 34500 2144 34516 2208
rect 34580 2144 34586 2208
rect 34270 2143 34586 2144
rect 45378 2208 45694 2209
rect 45378 2144 45384 2208
rect 45448 2144 45464 2208
rect 45528 2144 45544 2208
rect 45608 2144 45624 2208
rect 45688 2144 45694 2208
rect 45378 2143 45694 2144
rect 6500 1664 6816 1665
rect 6500 1600 6506 1664
rect 6570 1600 6586 1664
rect 6650 1600 6666 1664
rect 6730 1600 6746 1664
rect 6810 1600 6816 1664
rect 6500 1599 6816 1600
rect 17608 1664 17924 1665
rect 17608 1600 17614 1664
rect 17678 1600 17694 1664
rect 17758 1600 17774 1664
rect 17838 1600 17854 1664
rect 17918 1600 17924 1664
rect 17608 1599 17924 1600
rect 28716 1664 29032 1665
rect 28716 1600 28722 1664
rect 28786 1600 28802 1664
rect 28866 1600 28882 1664
rect 28946 1600 28962 1664
rect 29026 1600 29032 1664
rect 28716 1599 29032 1600
rect 39824 1664 40140 1665
rect 39824 1600 39830 1664
rect 39894 1600 39910 1664
rect 39974 1600 39990 1664
rect 40054 1600 40070 1664
rect 40134 1600 40140 1664
rect 39824 1599 40140 1600
rect 12054 1120 12370 1121
rect 12054 1056 12060 1120
rect 12124 1056 12140 1120
rect 12204 1056 12220 1120
rect 12284 1056 12300 1120
rect 12364 1056 12370 1120
rect 12054 1055 12370 1056
rect 23162 1120 23478 1121
rect 23162 1056 23168 1120
rect 23232 1056 23248 1120
rect 23312 1056 23328 1120
rect 23392 1056 23408 1120
rect 23472 1056 23478 1120
rect 23162 1055 23478 1056
rect 34270 1120 34586 1121
rect 34270 1056 34276 1120
rect 34340 1056 34356 1120
rect 34420 1056 34436 1120
rect 34500 1056 34516 1120
rect 34580 1056 34586 1120
rect 34270 1055 34586 1056
rect 45378 1120 45694 1121
rect 45378 1056 45384 1120
rect 45448 1056 45464 1120
rect 45528 1056 45544 1120
rect 45608 1056 45624 1120
rect 45688 1056 45694 1120
rect 45378 1055 45694 1056
<< via3 >>
rect 19380 9420 19444 9484
rect 12060 8732 12124 8736
rect 12060 8676 12064 8732
rect 12064 8676 12120 8732
rect 12120 8676 12124 8732
rect 12060 8672 12124 8676
rect 12140 8732 12204 8736
rect 12140 8676 12144 8732
rect 12144 8676 12200 8732
rect 12200 8676 12204 8732
rect 12140 8672 12204 8676
rect 12220 8732 12284 8736
rect 12220 8676 12224 8732
rect 12224 8676 12280 8732
rect 12280 8676 12284 8732
rect 12220 8672 12284 8676
rect 12300 8732 12364 8736
rect 12300 8676 12304 8732
rect 12304 8676 12360 8732
rect 12360 8676 12364 8732
rect 12300 8672 12364 8676
rect 23168 8732 23232 8736
rect 23168 8676 23172 8732
rect 23172 8676 23228 8732
rect 23228 8676 23232 8732
rect 23168 8672 23232 8676
rect 23248 8732 23312 8736
rect 23248 8676 23252 8732
rect 23252 8676 23308 8732
rect 23308 8676 23312 8732
rect 23248 8672 23312 8676
rect 23328 8732 23392 8736
rect 23328 8676 23332 8732
rect 23332 8676 23388 8732
rect 23388 8676 23392 8732
rect 23328 8672 23392 8676
rect 23408 8732 23472 8736
rect 23408 8676 23412 8732
rect 23412 8676 23468 8732
rect 23468 8676 23472 8732
rect 23408 8672 23472 8676
rect 34276 8732 34340 8736
rect 34276 8676 34280 8732
rect 34280 8676 34336 8732
rect 34336 8676 34340 8732
rect 34276 8672 34340 8676
rect 34356 8732 34420 8736
rect 34356 8676 34360 8732
rect 34360 8676 34416 8732
rect 34416 8676 34420 8732
rect 34356 8672 34420 8676
rect 34436 8732 34500 8736
rect 34436 8676 34440 8732
rect 34440 8676 34496 8732
rect 34496 8676 34500 8732
rect 34436 8672 34500 8676
rect 34516 8732 34580 8736
rect 34516 8676 34520 8732
rect 34520 8676 34576 8732
rect 34576 8676 34580 8732
rect 34516 8672 34580 8676
rect 45384 8732 45448 8736
rect 45384 8676 45388 8732
rect 45388 8676 45444 8732
rect 45444 8676 45448 8732
rect 45384 8672 45448 8676
rect 45464 8732 45528 8736
rect 45464 8676 45468 8732
rect 45468 8676 45524 8732
rect 45524 8676 45528 8732
rect 45464 8672 45528 8676
rect 45544 8732 45608 8736
rect 45544 8676 45548 8732
rect 45548 8676 45604 8732
rect 45604 8676 45608 8732
rect 45544 8672 45608 8676
rect 45624 8732 45688 8736
rect 45624 8676 45628 8732
rect 45628 8676 45684 8732
rect 45684 8676 45688 8732
rect 45624 8672 45688 8676
rect 6506 8188 6570 8192
rect 6506 8132 6510 8188
rect 6510 8132 6566 8188
rect 6566 8132 6570 8188
rect 6506 8128 6570 8132
rect 6586 8188 6650 8192
rect 6586 8132 6590 8188
rect 6590 8132 6646 8188
rect 6646 8132 6650 8188
rect 6586 8128 6650 8132
rect 6666 8188 6730 8192
rect 6666 8132 6670 8188
rect 6670 8132 6726 8188
rect 6726 8132 6730 8188
rect 6666 8128 6730 8132
rect 6746 8188 6810 8192
rect 6746 8132 6750 8188
rect 6750 8132 6806 8188
rect 6806 8132 6810 8188
rect 6746 8128 6810 8132
rect 17614 8188 17678 8192
rect 17614 8132 17618 8188
rect 17618 8132 17674 8188
rect 17674 8132 17678 8188
rect 17614 8128 17678 8132
rect 17694 8188 17758 8192
rect 17694 8132 17698 8188
rect 17698 8132 17754 8188
rect 17754 8132 17758 8188
rect 17694 8128 17758 8132
rect 17774 8188 17838 8192
rect 17774 8132 17778 8188
rect 17778 8132 17834 8188
rect 17834 8132 17838 8188
rect 17774 8128 17838 8132
rect 17854 8188 17918 8192
rect 17854 8132 17858 8188
rect 17858 8132 17914 8188
rect 17914 8132 17918 8188
rect 17854 8128 17918 8132
rect 28722 8188 28786 8192
rect 28722 8132 28726 8188
rect 28726 8132 28782 8188
rect 28782 8132 28786 8188
rect 28722 8128 28786 8132
rect 28802 8188 28866 8192
rect 28802 8132 28806 8188
rect 28806 8132 28862 8188
rect 28862 8132 28866 8188
rect 28802 8128 28866 8132
rect 28882 8188 28946 8192
rect 28882 8132 28886 8188
rect 28886 8132 28942 8188
rect 28942 8132 28946 8188
rect 28882 8128 28946 8132
rect 28962 8188 29026 8192
rect 28962 8132 28966 8188
rect 28966 8132 29022 8188
rect 29022 8132 29026 8188
rect 28962 8128 29026 8132
rect 39830 8188 39894 8192
rect 39830 8132 39834 8188
rect 39834 8132 39890 8188
rect 39890 8132 39894 8188
rect 39830 8128 39894 8132
rect 39910 8188 39974 8192
rect 39910 8132 39914 8188
rect 39914 8132 39970 8188
rect 39970 8132 39974 8188
rect 39910 8128 39974 8132
rect 39990 8188 40054 8192
rect 39990 8132 39994 8188
rect 39994 8132 40050 8188
rect 40050 8132 40054 8188
rect 39990 8128 40054 8132
rect 40070 8188 40134 8192
rect 40070 8132 40074 8188
rect 40074 8132 40130 8188
rect 40130 8132 40134 8188
rect 40070 8128 40134 8132
rect 12060 7644 12124 7648
rect 12060 7588 12064 7644
rect 12064 7588 12120 7644
rect 12120 7588 12124 7644
rect 12060 7584 12124 7588
rect 12140 7644 12204 7648
rect 12140 7588 12144 7644
rect 12144 7588 12200 7644
rect 12200 7588 12204 7644
rect 12140 7584 12204 7588
rect 12220 7644 12284 7648
rect 12220 7588 12224 7644
rect 12224 7588 12280 7644
rect 12280 7588 12284 7644
rect 12220 7584 12284 7588
rect 12300 7644 12364 7648
rect 12300 7588 12304 7644
rect 12304 7588 12360 7644
rect 12360 7588 12364 7644
rect 12300 7584 12364 7588
rect 23168 7644 23232 7648
rect 23168 7588 23172 7644
rect 23172 7588 23228 7644
rect 23228 7588 23232 7644
rect 23168 7584 23232 7588
rect 23248 7644 23312 7648
rect 23248 7588 23252 7644
rect 23252 7588 23308 7644
rect 23308 7588 23312 7644
rect 23248 7584 23312 7588
rect 23328 7644 23392 7648
rect 23328 7588 23332 7644
rect 23332 7588 23388 7644
rect 23388 7588 23392 7644
rect 23328 7584 23392 7588
rect 23408 7644 23472 7648
rect 23408 7588 23412 7644
rect 23412 7588 23468 7644
rect 23468 7588 23472 7644
rect 23408 7584 23472 7588
rect 34276 7644 34340 7648
rect 34276 7588 34280 7644
rect 34280 7588 34336 7644
rect 34336 7588 34340 7644
rect 34276 7584 34340 7588
rect 34356 7644 34420 7648
rect 34356 7588 34360 7644
rect 34360 7588 34416 7644
rect 34416 7588 34420 7644
rect 34356 7584 34420 7588
rect 34436 7644 34500 7648
rect 34436 7588 34440 7644
rect 34440 7588 34496 7644
rect 34496 7588 34500 7644
rect 34436 7584 34500 7588
rect 34516 7644 34580 7648
rect 34516 7588 34520 7644
rect 34520 7588 34576 7644
rect 34576 7588 34580 7644
rect 34516 7584 34580 7588
rect 45384 7644 45448 7648
rect 45384 7588 45388 7644
rect 45388 7588 45444 7644
rect 45444 7588 45448 7644
rect 45384 7584 45448 7588
rect 45464 7644 45528 7648
rect 45464 7588 45468 7644
rect 45468 7588 45524 7644
rect 45524 7588 45528 7644
rect 45464 7584 45528 7588
rect 45544 7644 45608 7648
rect 45544 7588 45548 7644
rect 45548 7588 45604 7644
rect 45604 7588 45608 7644
rect 45544 7584 45608 7588
rect 45624 7644 45688 7648
rect 45624 7588 45628 7644
rect 45628 7588 45684 7644
rect 45684 7588 45688 7644
rect 45624 7584 45688 7588
rect 6506 7100 6570 7104
rect 6506 7044 6510 7100
rect 6510 7044 6566 7100
rect 6566 7044 6570 7100
rect 6506 7040 6570 7044
rect 6586 7100 6650 7104
rect 6586 7044 6590 7100
rect 6590 7044 6646 7100
rect 6646 7044 6650 7100
rect 6586 7040 6650 7044
rect 6666 7100 6730 7104
rect 6666 7044 6670 7100
rect 6670 7044 6726 7100
rect 6726 7044 6730 7100
rect 6666 7040 6730 7044
rect 6746 7100 6810 7104
rect 6746 7044 6750 7100
rect 6750 7044 6806 7100
rect 6806 7044 6810 7100
rect 6746 7040 6810 7044
rect 17614 7100 17678 7104
rect 17614 7044 17618 7100
rect 17618 7044 17674 7100
rect 17674 7044 17678 7100
rect 17614 7040 17678 7044
rect 17694 7100 17758 7104
rect 17694 7044 17698 7100
rect 17698 7044 17754 7100
rect 17754 7044 17758 7100
rect 17694 7040 17758 7044
rect 17774 7100 17838 7104
rect 17774 7044 17778 7100
rect 17778 7044 17834 7100
rect 17834 7044 17838 7100
rect 17774 7040 17838 7044
rect 17854 7100 17918 7104
rect 17854 7044 17858 7100
rect 17858 7044 17914 7100
rect 17914 7044 17918 7100
rect 17854 7040 17918 7044
rect 19380 7108 19444 7172
rect 28722 7100 28786 7104
rect 28722 7044 28726 7100
rect 28726 7044 28782 7100
rect 28782 7044 28786 7100
rect 28722 7040 28786 7044
rect 28802 7100 28866 7104
rect 28802 7044 28806 7100
rect 28806 7044 28862 7100
rect 28862 7044 28866 7100
rect 28802 7040 28866 7044
rect 28882 7100 28946 7104
rect 28882 7044 28886 7100
rect 28886 7044 28942 7100
rect 28942 7044 28946 7100
rect 28882 7040 28946 7044
rect 28962 7100 29026 7104
rect 28962 7044 28966 7100
rect 28966 7044 29022 7100
rect 29022 7044 29026 7100
rect 28962 7040 29026 7044
rect 39830 7100 39894 7104
rect 39830 7044 39834 7100
rect 39834 7044 39890 7100
rect 39890 7044 39894 7100
rect 39830 7040 39894 7044
rect 39910 7100 39974 7104
rect 39910 7044 39914 7100
rect 39914 7044 39970 7100
rect 39970 7044 39974 7100
rect 39910 7040 39974 7044
rect 39990 7100 40054 7104
rect 39990 7044 39994 7100
rect 39994 7044 40050 7100
rect 40050 7044 40054 7100
rect 39990 7040 40054 7044
rect 40070 7100 40134 7104
rect 40070 7044 40074 7100
rect 40074 7044 40130 7100
rect 40130 7044 40134 7100
rect 40070 7040 40134 7044
rect 12060 6556 12124 6560
rect 12060 6500 12064 6556
rect 12064 6500 12120 6556
rect 12120 6500 12124 6556
rect 12060 6496 12124 6500
rect 12140 6556 12204 6560
rect 12140 6500 12144 6556
rect 12144 6500 12200 6556
rect 12200 6500 12204 6556
rect 12140 6496 12204 6500
rect 12220 6556 12284 6560
rect 12220 6500 12224 6556
rect 12224 6500 12280 6556
rect 12280 6500 12284 6556
rect 12220 6496 12284 6500
rect 12300 6556 12364 6560
rect 12300 6500 12304 6556
rect 12304 6500 12360 6556
rect 12360 6500 12364 6556
rect 12300 6496 12364 6500
rect 23168 6556 23232 6560
rect 23168 6500 23172 6556
rect 23172 6500 23228 6556
rect 23228 6500 23232 6556
rect 23168 6496 23232 6500
rect 23248 6556 23312 6560
rect 23248 6500 23252 6556
rect 23252 6500 23308 6556
rect 23308 6500 23312 6556
rect 23248 6496 23312 6500
rect 23328 6556 23392 6560
rect 23328 6500 23332 6556
rect 23332 6500 23388 6556
rect 23388 6500 23392 6556
rect 23328 6496 23392 6500
rect 23408 6556 23472 6560
rect 23408 6500 23412 6556
rect 23412 6500 23468 6556
rect 23468 6500 23472 6556
rect 23408 6496 23472 6500
rect 34276 6556 34340 6560
rect 34276 6500 34280 6556
rect 34280 6500 34336 6556
rect 34336 6500 34340 6556
rect 34276 6496 34340 6500
rect 34356 6556 34420 6560
rect 34356 6500 34360 6556
rect 34360 6500 34416 6556
rect 34416 6500 34420 6556
rect 34356 6496 34420 6500
rect 34436 6556 34500 6560
rect 34436 6500 34440 6556
rect 34440 6500 34496 6556
rect 34496 6500 34500 6556
rect 34436 6496 34500 6500
rect 34516 6556 34580 6560
rect 34516 6500 34520 6556
rect 34520 6500 34576 6556
rect 34576 6500 34580 6556
rect 34516 6496 34580 6500
rect 45384 6556 45448 6560
rect 45384 6500 45388 6556
rect 45388 6500 45444 6556
rect 45444 6500 45448 6556
rect 45384 6496 45448 6500
rect 45464 6556 45528 6560
rect 45464 6500 45468 6556
rect 45468 6500 45524 6556
rect 45524 6500 45528 6556
rect 45464 6496 45528 6500
rect 45544 6556 45608 6560
rect 45544 6500 45548 6556
rect 45548 6500 45604 6556
rect 45604 6500 45608 6556
rect 45544 6496 45608 6500
rect 45624 6556 45688 6560
rect 45624 6500 45628 6556
rect 45628 6500 45684 6556
rect 45684 6500 45688 6556
rect 45624 6496 45688 6500
rect 6506 6012 6570 6016
rect 6506 5956 6510 6012
rect 6510 5956 6566 6012
rect 6566 5956 6570 6012
rect 6506 5952 6570 5956
rect 6586 6012 6650 6016
rect 6586 5956 6590 6012
rect 6590 5956 6646 6012
rect 6646 5956 6650 6012
rect 6586 5952 6650 5956
rect 6666 6012 6730 6016
rect 6666 5956 6670 6012
rect 6670 5956 6726 6012
rect 6726 5956 6730 6012
rect 6666 5952 6730 5956
rect 6746 6012 6810 6016
rect 6746 5956 6750 6012
rect 6750 5956 6806 6012
rect 6806 5956 6810 6012
rect 6746 5952 6810 5956
rect 17614 6012 17678 6016
rect 17614 5956 17618 6012
rect 17618 5956 17674 6012
rect 17674 5956 17678 6012
rect 17614 5952 17678 5956
rect 17694 6012 17758 6016
rect 17694 5956 17698 6012
rect 17698 5956 17754 6012
rect 17754 5956 17758 6012
rect 17694 5952 17758 5956
rect 17774 6012 17838 6016
rect 17774 5956 17778 6012
rect 17778 5956 17834 6012
rect 17834 5956 17838 6012
rect 17774 5952 17838 5956
rect 17854 6012 17918 6016
rect 17854 5956 17858 6012
rect 17858 5956 17914 6012
rect 17914 5956 17918 6012
rect 17854 5952 17918 5956
rect 28722 6012 28786 6016
rect 28722 5956 28726 6012
rect 28726 5956 28782 6012
rect 28782 5956 28786 6012
rect 28722 5952 28786 5956
rect 28802 6012 28866 6016
rect 28802 5956 28806 6012
rect 28806 5956 28862 6012
rect 28862 5956 28866 6012
rect 28802 5952 28866 5956
rect 28882 6012 28946 6016
rect 28882 5956 28886 6012
rect 28886 5956 28942 6012
rect 28942 5956 28946 6012
rect 28882 5952 28946 5956
rect 28962 6012 29026 6016
rect 28962 5956 28966 6012
rect 28966 5956 29022 6012
rect 29022 5956 29026 6012
rect 28962 5952 29026 5956
rect 39830 6012 39894 6016
rect 39830 5956 39834 6012
rect 39834 5956 39890 6012
rect 39890 5956 39894 6012
rect 39830 5952 39894 5956
rect 39910 6012 39974 6016
rect 39910 5956 39914 6012
rect 39914 5956 39970 6012
rect 39970 5956 39974 6012
rect 39910 5952 39974 5956
rect 39990 6012 40054 6016
rect 39990 5956 39994 6012
rect 39994 5956 40050 6012
rect 40050 5956 40054 6012
rect 39990 5952 40054 5956
rect 40070 6012 40134 6016
rect 40070 5956 40074 6012
rect 40074 5956 40130 6012
rect 40130 5956 40134 6012
rect 40070 5952 40134 5956
rect 12060 5468 12124 5472
rect 12060 5412 12064 5468
rect 12064 5412 12120 5468
rect 12120 5412 12124 5468
rect 12060 5408 12124 5412
rect 12140 5468 12204 5472
rect 12140 5412 12144 5468
rect 12144 5412 12200 5468
rect 12200 5412 12204 5468
rect 12140 5408 12204 5412
rect 12220 5468 12284 5472
rect 12220 5412 12224 5468
rect 12224 5412 12280 5468
rect 12280 5412 12284 5468
rect 12220 5408 12284 5412
rect 12300 5468 12364 5472
rect 12300 5412 12304 5468
rect 12304 5412 12360 5468
rect 12360 5412 12364 5468
rect 12300 5408 12364 5412
rect 23168 5468 23232 5472
rect 23168 5412 23172 5468
rect 23172 5412 23228 5468
rect 23228 5412 23232 5468
rect 23168 5408 23232 5412
rect 23248 5468 23312 5472
rect 23248 5412 23252 5468
rect 23252 5412 23308 5468
rect 23308 5412 23312 5468
rect 23248 5408 23312 5412
rect 23328 5468 23392 5472
rect 23328 5412 23332 5468
rect 23332 5412 23388 5468
rect 23388 5412 23392 5468
rect 23328 5408 23392 5412
rect 23408 5468 23472 5472
rect 23408 5412 23412 5468
rect 23412 5412 23468 5468
rect 23468 5412 23472 5468
rect 23408 5408 23472 5412
rect 34276 5468 34340 5472
rect 34276 5412 34280 5468
rect 34280 5412 34336 5468
rect 34336 5412 34340 5468
rect 34276 5408 34340 5412
rect 34356 5468 34420 5472
rect 34356 5412 34360 5468
rect 34360 5412 34416 5468
rect 34416 5412 34420 5468
rect 34356 5408 34420 5412
rect 34436 5468 34500 5472
rect 34436 5412 34440 5468
rect 34440 5412 34496 5468
rect 34496 5412 34500 5468
rect 34436 5408 34500 5412
rect 34516 5468 34580 5472
rect 34516 5412 34520 5468
rect 34520 5412 34576 5468
rect 34576 5412 34580 5468
rect 34516 5408 34580 5412
rect 45384 5468 45448 5472
rect 45384 5412 45388 5468
rect 45388 5412 45444 5468
rect 45444 5412 45448 5468
rect 45384 5408 45448 5412
rect 45464 5468 45528 5472
rect 45464 5412 45468 5468
rect 45468 5412 45524 5468
rect 45524 5412 45528 5468
rect 45464 5408 45528 5412
rect 45544 5468 45608 5472
rect 45544 5412 45548 5468
rect 45548 5412 45604 5468
rect 45604 5412 45608 5468
rect 45544 5408 45608 5412
rect 45624 5468 45688 5472
rect 45624 5412 45628 5468
rect 45628 5412 45684 5468
rect 45684 5412 45688 5468
rect 45624 5408 45688 5412
rect 6506 4924 6570 4928
rect 6506 4868 6510 4924
rect 6510 4868 6566 4924
rect 6566 4868 6570 4924
rect 6506 4864 6570 4868
rect 6586 4924 6650 4928
rect 6586 4868 6590 4924
rect 6590 4868 6646 4924
rect 6646 4868 6650 4924
rect 6586 4864 6650 4868
rect 6666 4924 6730 4928
rect 6666 4868 6670 4924
rect 6670 4868 6726 4924
rect 6726 4868 6730 4924
rect 6666 4864 6730 4868
rect 6746 4924 6810 4928
rect 6746 4868 6750 4924
rect 6750 4868 6806 4924
rect 6806 4868 6810 4924
rect 6746 4864 6810 4868
rect 17614 4924 17678 4928
rect 17614 4868 17618 4924
rect 17618 4868 17674 4924
rect 17674 4868 17678 4924
rect 17614 4864 17678 4868
rect 17694 4924 17758 4928
rect 17694 4868 17698 4924
rect 17698 4868 17754 4924
rect 17754 4868 17758 4924
rect 17694 4864 17758 4868
rect 17774 4924 17838 4928
rect 17774 4868 17778 4924
rect 17778 4868 17834 4924
rect 17834 4868 17838 4924
rect 17774 4864 17838 4868
rect 17854 4924 17918 4928
rect 17854 4868 17858 4924
rect 17858 4868 17914 4924
rect 17914 4868 17918 4924
rect 17854 4864 17918 4868
rect 28722 4924 28786 4928
rect 28722 4868 28726 4924
rect 28726 4868 28782 4924
rect 28782 4868 28786 4924
rect 28722 4864 28786 4868
rect 28802 4924 28866 4928
rect 28802 4868 28806 4924
rect 28806 4868 28862 4924
rect 28862 4868 28866 4924
rect 28802 4864 28866 4868
rect 28882 4924 28946 4928
rect 28882 4868 28886 4924
rect 28886 4868 28942 4924
rect 28942 4868 28946 4924
rect 28882 4864 28946 4868
rect 28962 4924 29026 4928
rect 28962 4868 28966 4924
rect 28966 4868 29022 4924
rect 29022 4868 29026 4924
rect 28962 4864 29026 4868
rect 39830 4924 39894 4928
rect 39830 4868 39834 4924
rect 39834 4868 39890 4924
rect 39890 4868 39894 4924
rect 39830 4864 39894 4868
rect 39910 4924 39974 4928
rect 39910 4868 39914 4924
rect 39914 4868 39970 4924
rect 39970 4868 39974 4924
rect 39910 4864 39974 4868
rect 39990 4924 40054 4928
rect 39990 4868 39994 4924
rect 39994 4868 40050 4924
rect 40050 4868 40054 4924
rect 39990 4864 40054 4868
rect 40070 4924 40134 4928
rect 40070 4868 40074 4924
rect 40074 4868 40130 4924
rect 40130 4868 40134 4924
rect 40070 4864 40134 4868
rect 12060 4380 12124 4384
rect 12060 4324 12064 4380
rect 12064 4324 12120 4380
rect 12120 4324 12124 4380
rect 12060 4320 12124 4324
rect 12140 4380 12204 4384
rect 12140 4324 12144 4380
rect 12144 4324 12200 4380
rect 12200 4324 12204 4380
rect 12140 4320 12204 4324
rect 12220 4380 12284 4384
rect 12220 4324 12224 4380
rect 12224 4324 12280 4380
rect 12280 4324 12284 4380
rect 12220 4320 12284 4324
rect 12300 4380 12364 4384
rect 12300 4324 12304 4380
rect 12304 4324 12360 4380
rect 12360 4324 12364 4380
rect 12300 4320 12364 4324
rect 23168 4380 23232 4384
rect 23168 4324 23172 4380
rect 23172 4324 23228 4380
rect 23228 4324 23232 4380
rect 23168 4320 23232 4324
rect 23248 4380 23312 4384
rect 23248 4324 23252 4380
rect 23252 4324 23308 4380
rect 23308 4324 23312 4380
rect 23248 4320 23312 4324
rect 23328 4380 23392 4384
rect 23328 4324 23332 4380
rect 23332 4324 23388 4380
rect 23388 4324 23392 4380
rect 23328 4320 23392 4324
rect 23408 4380 23472 4384
rect 23408 4324 23412 4380
rect 23412 4324 23468 4380
rect 23468 4324 23472 4380
rect 23408 4320 23472 4324
rect 34276 4380 34340 4384
rect 34276 4324 34280 4380
rect 34280 4324 34336 4380
rect 34336 4324 34340 4380
rect 34276 4320 34340 4324
rect 34356 4380 34420 4384
rect 34356 4324 34360 4380
rect 34360 4324 34416 4380
rect 34416 4324 34420 4380
rect 34356 4320 34420 4324
rect 34436 4380 34500 4384
rect 34436 4324 34440 4380
rect 34440 4324 34496 4380
rect 34496 4324 34500 4380
rect 34436 4320 34500 4324
rect 34516 4380 34580 4384
rect 34516 4324 34520 4380
rect 34520 4324 34576 4380
rect 34576 4324 34580 4380
rect 34516 4320 34580 4324
rect 45384 4380 45448 4384
rect 45384 4324 45388 4380
rect 45388 4324 45444 4380
rect 45444 4324 45448 4380
rect 45384 4320 45448 4324
rect 45464 4380 45528 4384
rect 45464 4324 45468 4380
rect 45468 4324 45524 4380
rect 45524 4324 45528 4380
rect 45464 4320 45528 4324
rect 45544 4380 45608 4384
rect 45544 4324 45548 4380
rect 45548 4324 45604 4380
rect 45604 4324 45608 4380
rect 45544 4320 45608 4324
rect 45624 4380 45688 4384
rect 45624 4324 45628 4380
rect 45628 4324 45684 4380
rect 45684 4324 45688 4380
rect 45624 4320 45688 4324
rect 6506 3836 6570 3840
rect 6506 3780 6510 3836
rect 6510 3780 6566 3836
rect 6566 3780 6570 3836
rect 6506 3776 6570 3780
rect 6586 3836 6650 3840
rect 6586 3780 6590 3836
rect 6590 3780 6646 3836
rect 6646 3780 6650 3836
rect 6586 3776 6650 3780
rect 6666 3836 6730 3840
rect 6666 3780 6670 3836
rect 6670 3780 6726 3836
rect 6726 3780 6730 3836
rect 6666 3776 6730 3780
rect 6746 3836 6810 3840
rect 6746 3780 6750 3836
rect 6750 3780 6806 3836
rect 6806 3780 6810 3836
rect 6746 3776 6810 3780
rect 17614 3836 17678 3840
rect 17614 3780 17618 3836
rect 17618 3780 17674 3836
rect 17674 3780 17678 3836
rect 17614 3776 17678 3780
rect 17694 3836 17758 3840
rect 17694 3780 17698 3836
rect 17698 3780 17754 3836
rect 17754 3780 17758 3836
rect 17694 3776 17758 3780
rect 17774 3836 17838 3840
rect 17774 3780 17778 3836
rect 17778 3780 17834 3836
rect 17834 3780 17838 3836
rect 17774 3776 17838 3780
rect 17854 3836 17918 3840
rect 17854 3780 17858 3836
rect 17858 3780 17914 3836
rect 17914 3780 17918 3836
rect 17854 3776 17918 3780
rect 28722 3836 28786 3840
rect 28722 3780 28726 3836
rect 28726 3780 28782 3836
rect 28782 3780 28786 3836
rect 28722 3776 28786 3780
rect 28802 3836 28866 3840
rect 28802 3780 28806 3836
rect 28806 3780 28862 3836
rect 28862 3780 28866 3836
rect 28802 3776 28866 3780
rect 28882 3836 28946 3840
rect 28882 3780 28886 3836
rect 28886 3780 28942 3836
rect 28942 3780 28946 3836
rect 28882 3776 28946 3780
rect 28962 3836 29026 3840
rect 28962 3780 28966 3836
rect 28966 3780 29022 3836
rect 29022 3780 29026 3836
rect 28962 3776 29026 3780
rect 39830 3836 39894 3840
rect 39830 3780 39834 3836
rect 39834 3780 39890 3836
rect 39890 3780 39894 3836
rect 39830 3776 39894 3780
rect 39910 3836 39974 3840
rect 39910 3780 39914 3836
rect 39914 3780 39970 3836
rect 39970 3780 39974 3836
rect 39910 3776 39974 3780
rect 39990 3836 40054 3840
rect 39990 3780 39994 3836
rect 39994 3780 40050 3836
rect 40050 3780 40054 3836
rect 39990 3776 40054 3780
rect 40070 3836 40134 3840
rect 40070 3780 40074 3836
rect 40074 3780 40130 3836
rect 40130 3780 40134 3836
rect 40070 3776 40134 3780
rect 12060 3292 12124 3296
rect 12060 3236 12064 3292
rect 12064 3236 12120 3292
rect 12120 3236 12124 3292
rect 12060 3232 12124 3236
rect 12140 3292 12204 3296
rect 12140 3236 12144 3292
rect 12144 3236 12200 3292
rect 12200 3236 12204 3292
rect 12140 3232 12204 3236
rect 12220 3292 12284 3296
rect 12220 3236 12224 3292
rect 12224 3236 12280 3292
rect 12280 3236 12284 3292
rect 12220 3232 12284 3236
rect 12300 3292 12364 3296
rect 12300 3236 12304 3292
rect 12304 3236 12360 3292
rect 12360 3236 12364 3292
rect 12300 3232 12364 3236
rect 23168 3292 23232 3296
rect 23168 3236 23172 3292
rect 23172 3236 23228 3292
rect 23228 3236 23232 3292
rect 23168 3232 23232 3236
rect 23248 3292 23312 3296
rect 23248 3236 23252 3292
rect 23252 3236 23308 3292
rect 23308 3236 23312 3292
rect 23248 3232 23312 3236
rect 23328 3292 23392 3296
rect 23328 3236 23332 3292
rect 23332 3236 23388 3292
rect 23388 3236 23392 3292
rect 23328 3232 23392 3236
rect 23408 3292 23472 3296
rect 23408 3236 23412 3292
rect 23412 3236 23468 3292
rect 23468 3236 23472 3292
rect 23408 3232 23472 3236
rect 34276 3292 34340 3296
rect 34276 3236 34280 3292
rect 34280 3236 34336 3292
rect 34336 3236 34340 3292
rect 34276 3232 34340 3236
rect 34356 3292 34420 3296
rect 34356 3236 34360 3292
rect 34360 3236 34416 3292
rect 34416 3236 34420 3292
rect 34356 3232 34420 3236
rect 34436 3292 34500 3296
rect 34436 3236 34440 3292
rect 34440 3236 34496 3292
rect 34496 3236 34500 3292
rect 34436 3232 34500 3236
rect 34516 3292 34580 3296
rect 34516 3236 34520 3292
rect 34520 3236 34576 3292
rect 34576 3236 34580 3292
rect 34516 3232 34580 3236
rect 45384 3292 45448 3296
rect 45384 3236 45388 3292
rect 45388 3236 45444 3292
rect 45444 3236 45448 3292
rect 45384 3232 45448 3236
rect 45464 3292 45528 3296
rect 45464 3236 45468 3292
rect 45468 3236 45524 3292
rect 45524 3236 45528 3292
rect 45464 3232 45528 3236
rect 45544 3292 45608 3296
rect 45544 3236 45548 3292
rect 45548 3236 45604 3292
rect 45604 3236 45608 3292
rect 45544 3232 45608 3236
rect 45624 3292 45688 3296
rect 45624 3236 45628 3292
rect 45628 3236 45684 3292
rect 45684 3236 45688 3292
rect 45624 3232 45688 3236
rect 6506 2748 6570 2752
rect 6506 2692 6510 2748
rect 6510 2692 6566 2748
rect 6566 2692 6570 2748
rect 6506 2688 6570 2692
rect 6586 2748 6650 2752
rect 6586 2692 6590 2748
rect 6590 2692 6646 2748
rect 6646 2692 6650 2748
rect 6586 2688 6650 2692
rect 6666 2748 6730 2752
rect 6666 2692 6670 2748
rect 6670 2692 6726 2748
rect 6726 2692 6730 2748
rect 6666 2688 6730 2692
rect 6746 2748 6810 2752
rect 6746 2692 6750 2748
rect 6750 2692 6806 2748
rect 6806 2692 6810 2748
rect 6746 2688 6810 2692
rect 17614 2748 17678 2752
rect 17614 2692 17618 2748
rect 17618 2692 17674 2748
rect 17674 2692 17678 2748
rect 17614 2688 17678 2692
rect 17694 2748 17758 2752
rect 17694 2692 17698 2748
rect 17698 2692 17754 2748
rect 17754 2692 17758 2748
rect 17694 2688 17758 2692
rect 17774 2748 17838 2752
rect 17774 2692 17778 2748
rect 17778 2692 17834 2748
rect 17834 2692 17838 2748
rect 17774 2688 17838 2692
rect 17854 2748 17918 2752
rect 17854 2692 17858 2748
rect 17858 2692 17914 2748
rect 17914 2692 17918 2748
rect 17854 2688 17918 2692
rect 28722 2748 28786 2752
rect 28722 2692 28726 2748
rect 28726 2692 28782 2748
rect 28782 2692 28786 2748
rect 28722 2688 28786 2692
rect 28802 2748 28866 2752
rect 28802 2692 28806 2748
rect 28806 2692 28862 2748
rect 28862 2692 28866 2748
rect 28802 2688 28866 2692
rect 28882 2748 28946 2752
rect 28882 2692 28886 2748
rect 28886 2692 28942 2748
rect 28942 2692 28946 2748
rect 28882 2688 28946 2692
rect 28962 2748 29026 2752
rect 28962 2692 28966 2748
rect 28966 2692 29022 2748
rect 29022 2692 29026 2748
rect 28962 2688 29026 2692
rect 39830 2748 39894 2752
rect 39830 2692 39834 2748
rect 39834 2692 39890 2748
rect 39890 2692 39894 2748
rect 39830 2688 39894 2692
rect 39910 2748 39974 2752
rect 39910 2692 39914 2748
rect 39914 2692 39970 2748
rect 39970 2692 39974 2748
rect 39910 2688 39974 2692
rect 39990 2748 40054 2752
rect 39990 2692 39994 2748
rect 39994 2692 40050 2748
rect 40050 2692 40054 2748
rect 39990 2688 40054 2692
rect 40070 2748 40134 2752
rect 40070 2692 40074 2748
rect 40074 2692 40130 2748
rect 40130 2692 40134 2748
rect 40070 2688 40134 2692
rect 12060 2204 12124 2208
rect 12060 2148 12064 2204
rect 12064 2148 12120 2204
rect 12120 2148 12124 2204
rect 12060 2144 12124 2148
rect 12140 2204 12204 2208
rect 12140 2148 12144 2204
rect 12144 2148 12200 2204
rect 12200 2148 12204 2204
rect 12140 2144 12204 2148
rect 12220 2204 12284 2208
rect 12220 2148 12224 2204
rect 12224 2148 12280 2204
rect 12280 2148 12284 2204
rect 12220 2144 12284 2148
rect 12300 2204 12364 2208
rect 12300 2148 12304 2204
rect 12304 2148 12360 2204
rect 12360 2148 12364 2204
rect 12300 2144 12364 2148
rect 23168 2204 23232 2208
rect 23168 2148 23172 2204
rect 23172 2148 23228 2204
rect 23228 2148 23232 2204
rect 23168 2144 23232 2148
rect 23248 2204 23312 2208
rect 23248 2148 23252 2204
rect 23252 2148 23308 2204
rect 23308 2148 23312 2204
rect 23248 2144 23312 2148
rect 23328 2204 23392 2208
rect 23328 2148 23332 2204
rect 23332 2148 23388 2204
rect 23388 2148 23392 2204
rect 23328 2144 23392 2148
rect 23408 2204 23472 2208
rect 23408 2148 23412 2204
rect 23412 2148 23468 2204
rect 23468 2148 23472 2204
rect 23408 2144 23472 2148
rect 34276 2204 34340 2208
rect 34276 2148 34280 2204
rect 34280 2148 34336 2204
rect 34336 2148 34340 2204
rect 34276 2144 34340 2148
rect 34356 2204 34420 2208
rect 34356 2148 34360 2204
rect 34360 2148 34416 2204
rect 34416 2148 34420 2204
rect 34356 2144 34420 2148
rect 34436 2204 34500 2208
rect 34436 2148 34440 2204
rect 34440 2148 34496 2204
rect 34496 2148 34500 2204
rect 34436 2144 34500 2148
rect 34516 2204 34580 2208
rect 34516 2148 34520 2204
rect 34520 2148 34576 2204
rect 34576 2148 34580 2204
rect 34516 2144 34580 2148
rect 45384 2204 45448 2208
rect 45384 2148 45388 2204
rect 45388 2148 45444 2204
rect 45444 2148 45448 2204
rect 45384 2144 45448 2148
rect 45464 2204 45528 2208
rect 45464 2148 45468 2204
rect 45468 2148 45524 2204
rect 45524 2148 45528 2204
rect 45464 2144 45528 2148
rect 45544 2204 45608 2208
rect 45544 2148 45548 2204
rect 45548 2148 45604 2204
rect 45604 2148 45608 2204
rect 45544 2144 45608 2148
rect 45624 2204 45688 2208
rect 45624 2148 45628 2204
rect 45628 2148 45684 2204
rect 45684 2148 45688 2204
rect 45624 2144 45688 2148
rect 6506 1660 6570 1664
rect 6506 1604 6510 1660
rect 6510 1604 6566 1660
rect 6566 1604 6570 1660
rect 6506 1600 6570 1604
rect 6586 1660 6650 1664
rect 6586 1604 6590 1660
rect 6590 1604 6646 1660
rect 6646 1604 6650 1660
rect 6586 1600 6650 1604
rect 6666 1660 6730 1664
rect 6666 1604 6670 1660
rect 6670 1604 6726 1660
rect 6726 1604 6730 1660
rect 6666 1600 6730 1604
rect 6746 1660 6810 1664
rect 6746 1604 6750 1660
rect 6750 1604 6806 1660
rect 6806 1604 6810 1660
rect 6746 1600 6810 1604
rect 17614 1660 17678 1664
rect 17614 1604 17618 1660
rect 17618 1604 17674 1660
rect 17674 1604 17678 1660
rect 17614 1600 17678 1604
rect 17694 1660 17758 1664
rect 17694 1604 17698 1660
rect 17698 1604 17754 1660
rect 17754 1604 17758 1660
rect 17694 1600 17758 1604
rect 17774 1660 17838 1664
rect 17774 1604 17778 1660
rect 17778 1604 17834 1660
rect 17834 1604 17838 1660
rect 17774 1600 17838 1604
rect 17854 1660 17918 1664
rect 17854 1604 17858 1660
rect 17858 1604 17914 1660
rect 17914 1604 17918 1660
rect 17854 1600 17918 1604
rect 28722 1660 28786 1664
rect 28722 1604 28726 1660
rect 28726 1604 28782 1660
rect 28782 1604 28786 1660
rect 28722 1600 28786 1604
rect 28802 1660 28866 1664
rect 28802 1604 28806 1660
rect 28806 1604 28862 1660
rect 28862 1604 28866 1660
rect 28802 1600 28866 1604
rect 28882 1660 28946 1664
rect 28882 1604 28886 1660
rect 28886 1604 28942 1660
rect 28942 1604 28946 1660
rect 28882 1600 28946 1604
rect 28962 1660 29026 1664
rect 28962 1604 28966 1660
rect 28966 1604 29022 1660
rect 29022 1604 29026 1660
rect 28962 1600 29026 1604
rect 39830 1660 39894 1664
rect 39830 1604 39834 1660
rect 39834 1604 39890 1660
rect 39890 1604 39894 1660
rect 39830 1600 39894 1604
rect 39910 1660 39974 1664
rect 39910 1604 39914 1660
rect 39914 1604 39970 1660
rect 39970 1604 39974 1660
rect 39910 1600 39974 1604
rect 39990 1660 40054 1664
rect 39990 1604 39994 1660
rect 39994 1604 40050 1660
rect 40050 1604 40054 1660
rect 39990 1600 40054 1604
rect 40070 1660 40134 1664
rect 40070 1604 40074 1660
rect 40074 1604 40130 1660
rect 40130 1604 40134 1660
rect 40070 1600 40134 1604
rect 12060 1116 12124 1120
rect 12060 1060 12064 1116
rect 12064 1060 12120 1116
rect 12120 1060 12124 1116
rect 12060 1056 12124 1060
rect 12140 1116 12204 1120
rect 12140 1060 12144 1116
rect 12144 1060 12200 1116
rect 12200 1060 12204 1116
rect 12140 1056 12204 1060
rect 12220 1116 12284 1120
rect 12220 1060 12224 1116
rect 12224 1060 12280 1116
rect 12280 1060 12284 1116
rect 12220 1056 12284 1060
rect 12300 1116 12364 1120
rect 12300 1060 12304 1116
rect 12304 1060 12360 1116
rect 12360 1060 12364 1116
rect 12300 1056 12364 1060
rect 23168 1116 23232 1120
rect 23168 1060 23172 1116
rect 23172 1060 23228 1116
rect 23228 1060 23232 1116
rect 23168 1056 23232 1060
rect 23248 1116 23312 1120
rect 23248 1060 23252 1116
rect 23252 1060 23308 1116
rect 23308 1060 23312 1116
rect 23248 1056 23312 1060
rect 23328 1116 23392 1120
rect 23328 1060 23332 1116
rect 23332 1060 23388 1116
rect 23388 1060 23392 1116
rect 23328 1056 23392 1060
rect 23408 1116 23472 1120
rect 23408 1060 23412 1116
rect 23412 1060 23468 1116
rect 23468 1060 23472 1116
rect 23408 1056 23472 1060
rect 34276 1116 34340 1120
rect 34276 1060 34280 1116
rect 34280 1060 34336 1116
rect 34336 1060 34340 1116
rect 34276 1056 34340 1060
rect 34356 1116 34420 1120
rect 34356 1060 34360 1116
rect 34360 1060 34416 1116
rect 34416 1060 34420 1116
rect 34356 1056 34420 1060
rect 34436 1116 34500 1120
rect 34436 1060 34440 1116
rect 34440 1060 34496 1116
rect 34496 1060 34500 1116
rect 34436 1056 34500 1060
rect 34516 1116 34580 1120
rect 34516 1060 34520 1116
rect 34520 1060 34576 1116
rect 34576 1060 34580 1116
rect 34516 1056 34580 1060
rect 45384 1116 45448 1120
rect 45384 1060 45388 1116
rect 45388 1060 45444 1116
rect 45444 1060 45448 1116
rect 45384 1056 45448 1060
rect 45464 1116 45528 1120
rect 45464 1060 45468 1116
rect 45468 1060 45524 1116
rect 45524 1060 45528 1116
rect 45464 1056 45528 1060
rect 45544 1116 45608 1120
rect 45544 1060 45548 1116
rect 45548 1060 45604 1116
rect 45604 1060 45608 1116
rect 45544 1056 45608 1060
rect 45624 1116 45688 1120
rect 45624 1060 45628 1116
rect 45628 1060 45684 1116
rect 45684 1060 45688 1116
rect 45624 1056 45688 1060
<< metal4 >>
rect 19379 9484 19445 9485
rect 19379 9420 19380 9484
rect 19444 9420 19445 9484
rect 19379 9419 19445 9420
rect 6498 8192 6818 8752
rect 6498 8128 6506 8192
rect 6570 8128 6586 8192
rect 6650 8128 6666 8192
rect 6730 8128 6746 8192
rect 6810 8128 6818 8192
rect 6498 7104 6818 8128
rect 6498 7040 6506 7104
rect 6570 7040 6586 7104
rect 6650 7040 6666 7104
rect 6730 7040 6746 7104
rect 6810 7040 6818 7104
rect 6498 6016 6818 7040
rect 6498 5952 6506 6016
rect 6570 5952 6586 6016
rect 6650 5952 6666 6016
rect 6730 5952 6746 6016
rect 6810 5952 6818 6016
rect 6498 4928 6818 5952
rect 6498 4864 6506 4928
rect 6570 4864 6586 4928
rect 6650 4864 6666 4928
rect 6730 4864 6746 4928
rect 6810 4864 6818 4928
rect 6498 3840 6818 4864
rect 6498 3776 6506 3840
rect 6570 3776 6586 3840
rect 6650 3776 6666 3840
rect 6730 3776 6746 3840
rect 6810 3776 6818 3840
rect 6498 2752 6818 3776
rect 6498 2688 6506 2752
rect 6570 2688 6586 2752
rect 6650 2688 6666 2752
rect 6730 2688 6746 2752
rect 6810 2688 6818 2752
rect 6498 1664 6818 2688
rect 6498 1600 6506 1664
rect 6570 1600 6586 1664
rect 6650 1600 6666 1664
rect 6730 1600 6746 1664
rect 6810 1600 6818 1664
rect 6498 1040 6818 1600
rect 12052 8736 12372 8752
rect 12052 8672 12060 8736
rect 12124 8672 12140 8736
rect 12204 8672 12220 8736
rect 12284 8672 12300 8736
rect 12364 8672 12372 8736
rect 12052 7648 12372 8672
rect 12052 7584 12060 7648
rect 12124 7584 12140 7648
rect 12204 7584 12220 7648
rect 12284 7584 12300 7648
rect 12364 7584 12372 7648
rect 12052 6560 12372 7584
rect 12052 6496 12060 6560
rect 12124 6496 12140 6560
rect 12204 6496 12220 6560
rect 12284 6496 12300 6560
rect 12364 6496 12372 6560
rect 12052 5472 12372 6496
rect 12052 5408 12060 5472
rect 12124 5408 12140 5472
rect 12204 5408 12220 5472
rect 12284 5408 12300 5472
rect 12364 5408 12372 5472
rect 12052 4384 12372 5408
rect 12052 4320 12060 4384
rect 12124 4320 12140 4384
rect 12204 4320 12220 4384
rect 12284 4320 12300 4384
rect 12364 4320 12372 4384
rect 12052 3296 12372 4320
rect 12052 3232 12060 3296
rect 12124 3232 12140 3296
rect 12204 3232 12220 3296
rect 12284 3232 12300 3296
rect 12364 3232 12372 3296
rect 12052 2208 12372 3232
rect 12052 2144 12060 2208
rect 12124 2144 12140 2208
rect 12204 2144 12220 2208
rect 12284 2144 12300 2208
rect 12364 2144 12372 2208
rect 12052 1120 12372 2144
rect 12052 1056 12060 1120
rect 12124 1056 12140 1120
rect 12204 1056 12220 1120
rect 12284 1056 12300 1120
rect 12364 1056 12372 1120
rect 12052 1040 12372 1056
rect 17606 8192 17926 8752
rect 17606 8128 17614 8192
rect 17678 8128 17694 8192
rect 17758 8128 17774 8192
rect 17838 8128 17854 8192
rect 17918 8128 17926 8192
rect 17606 7104 17926 8128
rect 19382 7173 19442 9419
rect 23160 8736 23480 8752
rect 23160 8672 23168 8736
rect 23232 8672 23248 8736
rect 23312 8672 23328 8736
rect 23392 8672 23408 8736
rect 23472 8672 23480 8736
rect 23160 7648 23480 8672
rect 23160 7584 23168 7648
rect 23232 7584 23248 7648
rect 23312 7584 23328 7648
rect 23392 7584 23408 7648
rect 23472 7584 23480 7648
rect 19379 7172 19445 7173
rect 19379 7108 19380 7172
rect 19444 7108 19445 7172
rect 19379 7107 19445 7108
rect 17606 7040 17614 7104
rect 17678 7040 17694 7104
rect 17758 7040 17774 7104
rect 17838 7040 17854 7104
rect 17918 7040 17926 7104
rect 17606 6016 17926 7040
rect 17606 5952 17614 6016
rect 17678 5952 17694 6016
rect 17758 5952 17774 6016
rect 17838 5952 17854 6016
rect 17918 5952 17926 6016
rect 17606 4928 17926 5952
rect 17606 4864 17614 4928
rect 17678 4864 17694 4928
rect 17758 4864 17774 4928
rect 17838 4864 17854 4928
rect 17918 4864 17926 4928
rect 17606 3840 17926 4864
rect 17606 3776 17614 3840
rect 17678 3776 17694 3840
rect 17758 3776 17774 3840
rect 17838 3776 17854 3840
rect 17918 3776 17926 3840
rect 17606 2752 17926 3776
rect 17606 2688 17614 2752
rect 17678 2688 17694 2752
rect 17758 2688 17774 2752
rect 17838 2688 17854 2752
rect 17918 2688 17926 2752
rect 17606 1664 17926 2688
rect 17606 1600 17614 1664
rect 17678 1600 17694 1664
rect 17758 1600 17774 1664
rect 17838 1600 17854 1664
rect 17918 1600 17926 1664
rect 17606 1040 17926 1600
rect 23160 6560 23480 7584
rect 23160 6496 23168 6560
rect 23232 6496 23248 6560
rect 23312 6496 23328 6560
rect 23392 6496 23408 6560
rect 23472 6496 23480 6560
rect 23160 5472 23480 6496
rect 23160 5408 23168 5472
rect 23232 5408 23248 5472
rect 23312 5408 23328 5472
rect 23392 5408 23408 5472
rect 23472 5408 23480 5472
rect 23160 4384 23480 5408
rect 23160 4320 23168 4384
rect 23232 4320 23248 4384
rect 23312 4320 23328 4384
rect 23392 4320 23408 4384
rect 23472 4320 23480 4384
rect 23160 3296 23480 4320
rect 23160 3232 23168 3296
rect 23232 3232 23248 3296
rect 23312 3232 23328 3296
rect 23392 3232 23408 3296
rect 23472 3232 23480 3296
rect 23160 2208 23480 3232
rect 23160 2144 23168 2208
rect 23232 2144 23248 2208
rect 23312 2144 23328 2208
rect 23392 2144 23408 2208
rect 23472 2144 23480 2208
rect 23160 1120 23480 2144
rect 23160 1056 23168 1120
rect 23232 1056 23248 1120
rect 23312 1056 23328 1120
rect 23392 1056 23408 1120
rect 23472 1056 23480 1120
rect 23160 1040 23480 1056
rect 28714 8192 29034 8752
rect 28714 8128 28722 8192
rect 28786 8128 28802 8192
rect 28866 8128 28882 8192
rect 28946 8128 28962 8192
rect 29026 8128 29034 8192
rect 28714 7104 29034 8128
rect 28714 7040 28722 7104
rect 28786 7040 28802 7104
rect 28866 7040 28882 7104
rect 28946 7040 28962 7104
rect 29026 7040 29034 7104
rect 28714 6016 29034 7040
rect 28714 5952 28722 6016
rect 28786 5952 28802 6016
rect 28866 5952 28882 6016
rect 28946 5952 28962 6016
rect 29026 5952 29034 6016
rect 28714 4928 29034 5952
rect 28714 4864 28722 4928
rect 28786 4864 28802 4928
rect 28866 4864 28882 4928
rect 28946 4864 28962 4928
rect 29026 4864 29034 4928
rect 28714 3840 29034 4864
rect 28714 3776 28722 3840
rect 28786 3776 28802 3840
rect 28866 3776 28882 3840
rect 28946 3776 28962 3840
rect 29026 3776 29034 3840
rect 28714 2752 29034 3776
rect 28714 2688 28722 2752
rect 28786 2688 28802 2752
rect 28866 2688 28882 2752
rect 28946 2688 28962 2752
rect 29026 2688 29034 2752
rect 28714 1664 29034 2688
rect 28714 1600 28722 1664
rect 28786 1600 28802 1664
rect 28866 1600 28882 1664
rect 28946 1600 28962 1664
rect 29026 1600 29034 1664
rect 28714 1040 29034 1600
rect 34268 8736 34588 8752
rect 34268 8672 34276 8736
rect 34340 8672 34356 8736
rect 34420 8672 34436 8736
rect 34500 8672 34516 8736
rect 34580 8672 34588 8736
rect 34268 7648 34588 8672
rect 34268 7584 34276 7648
rect 34340 7584 34356 7648
rect 34420 7584 34436 7648
rect 34500 7584 34516 7648
rect 34580 7584 34588 7648
rect 34268 6560 34588 7584
rect 34268 6496 34276 6560
rect 34340 6496 34356 6560
rect 34420 6496 34436 6560
rect 34500 6496 34516 6560
rect 34580 6496 34588 6560
rect 34268 5472 34588 6496
rect 34268 5408 34276 5472
rect 34340 5408 34356 5472
rect 34420 5408 34436 5472
rect 34500 5408 34516 5472
rect 34580 5408 34588 5472
rect 34268 4384 34588 5408
rect 34268 4320 34276 4384
rect 34340 4320 34356 4384
rect 34420 4320 34436 4384
rect 34500 4320 34516 4384
rect 34580 4320 34588 4384
rect 34268 3296 34588 4320
rect 34268 3232 34276 3296
rect 34340 3232 34356 3296
rect 34420 3232 34436 3296
rect 34500 3232 34516 3296
rect 34580 3232 34588 3296
rect 34268 2208 34588 3232
rect 34268 2144 34276 2208
rect 34340 2144 34356 2208
rect 34420 2144 34436 2208
rect 34500 2144 34516 2208
rect 34580 2144 34588 2208
rect 34268 1120 34588 2144
rect 34268 1056 34276 1120
rect 34340 1056 34356 1120
rect 34420 1056 34436 1120
rect 34500 1056 34516 1120
rect 34580 1056 34588 1120
rect 34268 1040 34588 1056
rect 39822 8192 40142 8752
rect 39822 8128 39830 8192
rect 39894 8128 39910 8192
rect 39974 8128 39990 8192
rect 40054 8128 40070 8192
rect 40134 8128 40142 8192
rect 39822 7104 40142 8128
rect 39822 7040 39830 7104
rect 39894 7040 39910 7104
rect 39974 7040 39990 7104
rect 40054 7040 40070 7104
rect 40134 7040 40142 7104
rect 39822 6016 40142 7040
rect 39822 5952 39830 6016
rect 39894 5952 39910 6016
rect 39974 5952 39990 6016
rect 40054 5952 40070 6016
rect 40134 5952 40142 6016
rect 39822 4928 40142 5952
rect 39822 4864 39830 4928
rect 39894 4864 39910 4928
rect 39974 4864 39990 4928
rect 40054 4864 40070 4928
rect 40134 4864 40142 4928
rect 39822 3840 40142 4864
rect 39822 3776 39830 3840
rect 39894 3776 39910 3840
rect 39974 3776 39990 3840
rect 40054 3776 40070 3840
rect 40134 3776 40142 3840
rect 39822 2752 40142 3776
rect 39822 2688 39830 2752
rect 39894 2688 39910 2752
rect 39974 2688 39990 2752
rect 40054 2688 40070 2752
rect 40134 2688 40142 2752
rect 39822 1664 40142 2688
rect 39822 1600 39830 1664
rect 39894 1600 39910 1664
rect 39974 1600 39990 1664
rect 40054 1600 40070 1664
rect 40134 1600 40142 1664
rect 39822 1040 40142 1600
rect 45376 8736 45696 8752
rect 45376 8672 45384 8736
rect 45448 8672 45464 8736
rect 45528 8672 45544 8736
rect 45608 8672 45624 8736
rect 45688 8672 45696 8736
rect 45376 7648 45696 8672
rect 45376 7584 45384 7648
rect 45448 7584 45464 7648
rect 45528 7584 45544 7648
rect 45608 7584 45624 7648
rect 45688 7584 45696 7648
rect 45376 6560 45696 7584
rect 45376 6496 45384 6560
rect 45448 6496 45464 6560
rect 45528 6496 45544 6560
rect 45608 6496 45624 6560
rect 45688 6496 45696 6560
rect 45376 5472 45696 6496
rect 45376 5408 45384 5472
rect 45448 5408 45464 5472
rect 45528 5408 45544 5472
rect 45608 5408 45624 5472
rect 45688 5408 45696 5472
rect 45376 4384 45696 5408
rect 45376 4320 45384 4384
rect 45448 4320 45464 4384
rect 45528 4320 45544 4384
rect 45608 4320 45624 4384
rect 45688 4320 45696 4384
rect 45376 3296 45696 4320
rect 45376 3232 45384 3296
rect 45448 3232 45464 3296
rect 45528 3232 45544 3296
rect 45608 3232 45624 3296
rect 45688 3232 45696 3296
rect 45376 2208 45696 3232
rect 45376 2144 45384 2208
rect 45448 2144 45464 2208
rect 45528 2144 45544 2208
rect 45608 2144 45624 2208
rect 45688 2144 45696 2208
rect 45376 1120 45696 2144
rect 45376 1056 45384 1120
rect 45448 1056 45464 1120
rect 45528 1056 45544 1120
rect 45608 1056 45624 1120
rect 45688 1056 45696 1120
rect 45376 1040 45696 1056
use sky130_fd_sc_hd__diode_2  ANTENNA_1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 1840 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1688980957
transform -1 0 4232 0 -1 8704
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_6 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1656 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_18 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2760 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_26 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3496 0 1 1088
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_32
timestamp 1688980957
transform 1 0 4048 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_44 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5152 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_53 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5980 0 1 1088
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_57
timestamp 1688980957
transform 1 0 6348 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_69 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 7452 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_73 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 7820 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_77
timestamp 1688980957
transform 1 0 8188 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_83
timestamp 1688980957
transform 1 0 8740 0 1 1088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_85
timestamp 1688980957
transform 1 0 8924 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_97
timestamp 1688980957
transform 1 0 10028 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_101
timestamp 1688980957
transform 1 0 10396 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_109
timestamp 1688980957
transform 1 0 11132 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_113
timestamp 1688980957
transform 1 0 11500 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_121
timestamp 1688980957
transform 1 0 12236 0 1 1088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_125
timestamp 1688980957
transform 1 0 12604 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_137
timestamp 1688980957
transform 1 0 13708 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_141
timestamp 1688980957
transform 1 0 14076 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_145
timestamp 1688980957
transform 1 0 14444 0 1 1088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_149
timestamp 1688980957
transform 1 0 14812 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_161
timestamp 1688980957
transform 1 0 15916 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_167
timestamp 1688980957
transform 1 0 16468 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_169
timestamp 1688980957
transform 1 0 16652 0 1 1088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_173
timestamp 1688980957
transform 1 0 17020 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_185
timestamp 1688980957
transform 1 0 18124 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_193
timestamp 1688980957
transform 1 0 18860 0 1 1088
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_200
timestamp 1688980957
transform 1 0 19504 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_212
timestamp 1688980957
transform 1 0 20608 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_221
timestamp 1688980957
transform 1 0 21436 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_225
timestamp 1688980957
transform 1 0 21804 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_231
timestamp 1688980957
transform 1 0 22356 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_239
timestamp 1688980957
transform 1 0 23092 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_245
timestamp 1688980957
transform 1 0 23644 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_251
timestamp 1688980957
transform 1 0 24196 0 1 1088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_253
timestamp 1688980957
transform 1 0 24380 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_265
timestamp 1688980957
transform 1 0 25484 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_269
timestamp 1688980957
transform 1 0 25852 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_277
timestamp 1688980957
transform 1 0 26588 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_281
timestamp 1688980957
transform 1 0 26956 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_289
timestamp 1688980957
transform 1 0 27692 0 1 1088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_293
timestamp 1688980957
transform 1 0 28060 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_305
timestamp 1688980957
transform 1 0 29164 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_309
timestamp 1688980957
transform 1 0 29532 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_313
timestamp 1688980957
transform 1 0 29900 0 1 1088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_317
timestamp 1688980957
transform 1 0 30268 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_329
timestamp 1688980957
transform 1 0 31372 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_335
timestamp 1688980957
transform 1 0 31924 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_337
timestamp 1688980957
transform 1 0 32108 0 1 1088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_341
timestamp 1688980957
transform 1 0 32476 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_353
timestamp 1688980957
transform 1 0 33580 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_361
timestamp 1688980957
transform 1 0 34316 0 1 1088
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_368
timestamp 1688980957
transform 1 0 34960 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_380
timestamp 1688980957
transform 1 0 36064 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_389
timestamp 1688980957
transform 1 0 36892 0 1 1088
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_393
timestamp 1688980957
transform 1 0 37260 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_405
timestamp 1688980957
transform 1 0 38364 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_409
timestamp 1688980957
transform 1 0 38732 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_413
timestamp 1688980957
transform 1 0 39100 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_419
timestamp 1688980957
transform 1 0 39652 0 1 1088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_421
timestamp 1688980957
transform 1 0 39836 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_433
timestamp 1688980957
transform 1 0 40940 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_437
timestamp 1688980957
transform 1 0 41308 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_445
timestamp 1688980957
transform 1 0 42044 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_449
timestamp 1688980957
transform 1 0 42412 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_457
timestamp 1688980957
transform 1 0 43148 0 1 1088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_461
timestamp 1688980957
transform 1 0 43516 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_473
timestamp 1688980957
transform 1 0 44620 0 1 1088
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 1688980957
transform 1 0 1380 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 1688980957
transform 1 0 2484 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_27
timestamp 1688980957
transform 1 0 3588 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_39
timestamp 1688980957
transform 1 0 4692 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_51
timestamp 1688980957
transform 1 0 5796 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 1688980957
transform 1 0 6164 0 -1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_57
timestamp 1688980957
transform 1 0 6348 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_69
timestamp 1688980957
transform 1 0 7452 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_81
timestamp 1688980957
transform 1 0 8556 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_93
timestamp 1688980957
transform 1 0 9660 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_105
timestamp 1688980957
transform 1 0 10764 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_111
timestamp 1688980957
transform 1 0 11316 0 -1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_113
timestamp 1688980957
transform 1 0 11500 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_125
timestamp 1688980957
transform 1 0 12604 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_137
timestamp 1688980957
transform 1 0 13708 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_149
timestamp 1688980957
transform 1 0 14812 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_161
timestamp 1688980957
transform 1 0 15916 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_167
timestamp 1688980957
transform 1 0 16468 0 -1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_169
timestamp 1688980957
transform 1 0 16652 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_181
timestamp 1688980957
transform 1 0 17756 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_193
timestamp 1688980957
transform 1 0 18860 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_202
timestamp 1688980957
transform 1 0 19688 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_209
timestamp 1688980957
transform 1 0 20332 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_217
timestamp 1688980957
transform 1 0 21068 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_225
timestamp 1688980957
transform 1 0 21804 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_245
timestamp 1688980957
transform 1 0 23644 0 -1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_250
timestamp 1688980957
transform 1 0 24104 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_262
timestamp 1688980957
transform 1 0 25208 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_270
timestamp 1688980957
transform 1 0 25944 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_274
timestamp 1688980957
transform 1 0 26312 0 -1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_281
timestamp 1688980957
transform 1 0 26956 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_293
timestamp 1688980957
transform 1 0 28060 0 -1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_298
timestamp 1688980957
transform 1 0 28520 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_310
timestamp 1688980957
transform 1 0 29624 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_318
timestamp 1688980957
transform 1 0 30360 0 -1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_322
timestamp 1688980957
transform 1 0 30728 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_334
timestamp 1688980957
transform 1 0 31832 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_337
timestamp 1688980957
transform 1 0 32108 0 -1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_346
timestamp 1688980957
transform 1 0 32936 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_358
timestamp 1688980957
transform 1 0 34040 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_366
timestamp 1688980957
transform 1 0 34776 0 -1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_370
timestamp 1688980957
transform 1 0 35144 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_382
timestamp 1688980957
transform 1 0 36248 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_390
timestamp 1688980957
transform 1 0 36984 0 -1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_396
timestamp 1688980957
transform 1 0 37536 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_408
timestamp 1688980957
transform 1 0 38640 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_420
timestamp 1688980957
transform 1 0 39744 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_432
timestamp 1688980957
transform 1 0 40848 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_443
timestamp 1688980957
transform 1 0 41860 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_447
timestamp 1688980957
transform 1 0 42228 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_449
timestamp 1688980957
transform 1 0 42412 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_457
timestamp 1688980957
transform 1 0 43148 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_463
timestamp 1688980957
transform 1 0 43700 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_468
timestamp 1688980957
transform 1 0 44160 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_473
timestamp 1688980957
transform 1 0 44620 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_479
timestamp 1688980957
transform 1 0 45172 0 -1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1688980957
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 1688980957
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1688980957
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 1688980957
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 1688980957
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_53
timestamp 1688980957
transform 1 0 5980 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_65
timestamp 1688980957
transform 1 0 7084 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_77
timestamp 1688980957
transform 1 0 8188 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 1688980957
transform 1 0 8740 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_85
timestamp 1688980957
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_97
timestamp 1688980957
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_109
timestamp 1688980957
transform 1 0 11132 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_121
timestamp 1688980957
transform 1 0 12236 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_133
timestamp 1688980957
transform 1 0 13340 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_139
timestamp 1688980957
transform 1 0 13892 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_141
timestamp 1688980957
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_153
timestamp 1688980957
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_165
timestamp 1688980957
transform 1 0 16284 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_177
timestamp 1688980957
transform 1 0 17388 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_189
timestamp 1688980957
transform 1 0 18492 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_195
timestamp 1688980957
transform 1 0 19044 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_197
timestamp 1688980957
transform 1 0 19228 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_205
timestamp 1688980957
transform 1 0 19964 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_212
timestamp 1688980957
transform 1 0 20608 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_224
timestamp 1688980957
transform 1 0 21712 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_228
timestamp 1688980957
transform 1 0 22080 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_236
timestamp 1688980957
transform 1 0 22816 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_253
timestamp 1688980957
transform 1 0 24380 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_259
timestamp 1688980957
transform 1 0 24932 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_271
timestamp 1688980957
transform 1 0 26036 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_279
timestamp 1688980957
transform 1 0 26772 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_283
timestamp 1688980957
transform 1 0 27140 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_295
timestamp 1688980957
transform 1 0 28244 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_303
timestamp 1688980957
transform 1 0 28980 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_307
timestamp 1688980957
transform 1 0 29348 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_309
timestamp 1688980957
transform 1 0 29532 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_321
timestamp 1688980957
transform 1 0 30636 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_327
timestamp 1688980957
transform 1 0 31188 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_331
timestamp 1688980957
transform 1 0 31556 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_343
timestamp 1688980957
transform 1 0 32660 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_351
timestamp 1688980957
transform 1 0 33396 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_355
timestamp 1688980957
transform 1 0 33764 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_363
timestamp 1688980957
transform 1 0 34500 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_365
timestamp 1688980957
transform 1 0 34684 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_373
timestamp 1688980957
transform 1 0 35420 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_379
timestamp 1688980957
transform 1 0 35972 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_391
timestamp 1688980957
transform 1 0 37076 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_399
timestamp 1688980957
transform 1 0 37812 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_403
timestamp 1688980957
transform 1 0 38180 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_415
timestamp 1688980957
transform 1 0 39284 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_419
timestamp 1688980957
transform 1 0 39652 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_421
timestamp 1688980957
transform 1 0 39836 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_433
timestamp 1688980957
transform 1 0 40940 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_445
timestamp 1688980957
transform 1 0 42044 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_457
timestamp 1688980957
transform 1 0 43148 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_474
timestamp 1688980957
transform 1 0 44712 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1688980957
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1688980957
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 1688980957
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 1688980957
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 1688980957
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1688980957
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 1688980957
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_69
timestamp 1688980957
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_81
timestamp 1688980957
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_93
timestamp 1688980957
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_105
timestamp 1688980957
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_111
timestamp 1688980957
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_113
timestamp 1688980957
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_125
timestamp 1688980957
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_137
timestamp 1688980957
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_149
timestamp 1688980957
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_161
timestamp 1688980957
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_167
timestamp 1688980957
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_169
timestamp 1688980957
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_181
timestamp 1688980957
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_193
timestamp 1688980957
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_205
timestamp 1688980957
transform 1 0 19964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_217
timestamp 1688980957
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_223
timestamp 1688980957
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_225
timestamp 1688980957
transform 1 0 21804 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_237
timestamp 1688980957
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_249
timestamp 1688980957
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_261
timestamp 1688980957
transform 1 0 25116 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_273
timestamp 1688980957
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_279
timestamp 1688980957
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_281
timestamp 1688980957
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_293
timestamp 1688980957
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_305
timestamp 1688980957
transform 1 0 29164 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_317
timestamp 1688980957
transform 1 0 30268 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_329
timestamp 1688980957
transform 1 0 31372 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_335
timestamp 1688980957
transform 1 0 31924 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_337
timestamp 1688980957
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_349
timestamp 1688980957
transform 1 0 33212 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_361
timestamp 1688980957
transform 1 0 34316 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_373
timestamp 1688980957
transform 1 0 35420 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_385
timestamp 1688980957
transform 1 0 36524 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_391
timestamp 1688980957
transform 1 0 37076 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_393
timestamp 1688980957
transform 1 0 37260 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_405
timestamp 1688980957
transform 1 0 38364 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_417
timestamp 1688980957
transform 1 0 39468 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_429
timestamp 1688980957
transform 1 0 40572 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_441
timestamp 1688980957
transform 1 0 41676 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_447
timestamp 1688980957
transform 1 0 42228 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_449
timestamp 1688980957
transform 1 0 42412 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_461
timestamp 1688980957
transform 1 0 43516 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_473
timestamp 1688980957
transform 1 0 44620 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_479
timestamp 1688980957
transform 1 0 45172 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1688980957
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 1688980957
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1688980957
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 1688980957
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 1688980957
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_53
timestamp 1688980957
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_65
timestamp 1688980957
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_77
timestamp 1688980957
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp 1688980957
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_85
timestamp 1688980957
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_97
timestamp 1688980957
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_109
timestamp 1688980957
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_121
timestamp 1688980957
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_133
timestamp 1688980957
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_139
timestamp 1688980957
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_141
timestamp 1688980957
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_153
timestamp 1688980957
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_165
timestamp 1688980957
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_177
timestamp 1688980957
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_189
timestamp 1688980957
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_195
timestamp 1688980957
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_197
timestamp 1688980957
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_209
timestamp 1688980957
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_221
timestamp 1688980957
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_233
timestamp 1688980957
transform 1 0 22540 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_245
timestamp 1688980957
transform 1 0 23644 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_251
timestamp 1688980957
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_253
timestamp 1688980957
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_265
timestamp 1688980957
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_277
timestamp 1688980957
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_289
timestamp 1688980957
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_301
timestamp 1688980957
transform 1 0 28796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_307
timestamp 1688980957
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_309
timestamp 1688980957
transform 1 0 29532 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_321
timestamp 1688980957
transform 1 0 30636 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_333
timestamp 1688980957
transform 1 0 31740 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_345
timestamp 1688980957
transform 1 0 32844 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_357
timestamp 1688980957
transform 1 0 33948 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_363
timestamp 1688980957
transform 1 0 34500 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_365
timestamp 1688980957
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_377
timestamp 1688980957
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_389
timestamp 1688980957
transform 1 0 36892 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_401
timestamp 1688980957
transform 1 0 37996 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_413
timestamp 1688980957
transform 1 0 39100 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_419
timestamp 1688980957
transform 1 0 39652 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_421
timestamp 1688980957
transform 1 0 39836 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_433
timestamp 1688980957
transform 1 0 40940 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_445
timestamp 1688980957
transform 1 0 42044 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_457
timestamp 1688980957
transform 1 0 43148 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_469
timestamp 1688980957
transform 1 0 44252 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_475
timestamp 1688980957
transform 1 0 44804 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_477
timestamp 1688980957
transform 1 0 44988 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 1688980957
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 1688980957
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_27
timestamp 1688980957
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_39
timestamp 1688980957
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_51
timestamp 1688980957
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 1688980957
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_57
timestamp 1688980957
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_69
timestamp 1688980957
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_81
timestamp 1688980957
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_93
timestamp 1688980957
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_105
timestamp 1688980957
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_111
timestamp 1688980957
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_113
timestamp 1688980957
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_125
timestamp 1688980957
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_137
timestamp 1688980957
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_149
timestamp 1688980957
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_161
timestamp 1688980957
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_167
timestamp 1688980957
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_169
timestamp 1688980957
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_181
timestamp 1688980957
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_193
timestamp 1688980957
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_205
timestamp 1688980957
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_217
timestamp 1688980957
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_223
timestamp 1688980957
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_225
timestamp 1688980957
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_237
timestamp 1688980957
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_249
timestamp 1688980957
transform 1 0 24012 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_261
timestamp 1688980957
transform 1 0 25116 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_273
timestamp 1688980957
transform 1 0 26220 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_279
timestamp 1688980957
transform 1 0 26772 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_281
timestamp 1688980957
transform 1 0 26956 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_293
timestamp 1688980957
transform 1 0 28060 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_305
timestamp 1688980957
transform 1 0 29164 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_317
timestamp 1688980957
transform 1 0 30268 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_329
timestamp 1688980957
transform 1 0 31372 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_335
timestamp 1688980957
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_337
timestamp 1688980957
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_349
timestamp 1688980957
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_361
timestamp 1688980957
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_373
timestamp 1688980957
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_385
timestamp 1688980957
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_391
timestamp 1688980957
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_393
timestamp 1688980957
transform 1 0 37260 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_405
timestamp 1688980957
transform 1 0 38364 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_417
timestamp 1688980957
transform 1 0 39468 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_429
timestamp 1688980957
transform 1 0 40572 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_441
timestamp 1688980957
transform 1 0 41676 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_447
timestamp 1688980957
transform 1 0 42228 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_449
timestamp 1688980957
transform 1 0 42412 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_461
timestamp 1688980957
transform 1 0 43516 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_473
timestamp 1688980957
transform 1 0 44620 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_479
timestamp 1688980957
transform 1 0 45172 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 1688980957
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_15
timestamp 1688980957
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1688980957
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 1688980957
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_41
timestamp 1688980957
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_53
timestamp 1688980957
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_65
timestamp 1688980957
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_77
timestamp 1688980957
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_83
timestamp 1688980957
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_85
timestamp 1688980957
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_97
timestamp 1688980957
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_109
timestamp 1688980957
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_121
timestamp 1688980957
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_133
timestamp 1688980957
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_139
timestamp 1688980957
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_141
timestamp 1688980957
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_153
timestamp 1688980957
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_165
timestamp 1688980957
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_177
timestamp 1688980957
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_189
timestamp 1688980957
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_195
timestamp 1688980957
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_197
timestamp 1688980957
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_209
timestamp 1688980957
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_221
timestamp 1688980957
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_233
timestamp 1688980957
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_245
timestamp 1688980957
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_251
timestamp 1688980957
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_253
timestamp 1688980957
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_265
timestamp 1688980957
transform 1 0 25484 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_277
timestamp 1688980957
transform 1 0 26588 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_289
timestamp 1688980957
transform 1 0 27692 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_301
timestamp 1688980957
transform 1 0 28796 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_307
timestamp 1688980957
transform 1 0 29348 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_309
timestamp 1688980957
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_321
timestamp 1688980957
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_333
timestamp 1688980957
transform 1 0 31740 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_345
timestamp 1688980957
transform 1 0 32844 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_357
timestamp 1688980957
transform 1 0 33948 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_363
timestamp 1688980957
transform 1 0 34500 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_365
timestamp 1688980957
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_377
timestamp 1688980957
transform 1 0 35788 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_389
timestamp 1688980957
transform 1 0 36892 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_401
timestamp 1688980957
transform 1 0 37996 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_413
timestamp 1688980957
transform 1 0 39100 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_419
timestamp 1688980957
transform 1 0 39652 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_421
timestamp 1688980957
transform 1 0 39836 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_433
timestamp 1688980957
transform 1 0 40940 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_445
timestamp 1688980957
transform 1 0 42044 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_457
timestamp 1688980957
transform 1 0 43148 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_469
timestamp 1688980957
transform 1 0 44252 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_475
timestamp 1688980957
transform 1 0 44804 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_477
timestamp 1688980957
transform 1 0 44988 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 1688980957
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 1688980957
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_27
timestamp 1688980957
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_39
timestamp 1688980957
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_51
timestamp 1688980957
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 1688980957
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_57
timestamp 1688980957
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_69
timestamp 1688980957
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_81
timestamp 1688980957
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_93
timestamp 1688980957
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_105
timestamp 1688980957
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_111
timestamp 1688980957
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_113
timestamp 1688980957
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_125
timestamp 1688980957
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_137
timestamp 1688980957
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_149
timestamp 1688980957
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_161
timestamp 1688980957
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_167
timestamp 1688980957
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_169
timestamp 1688980957
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_181
timestamp 1688980957
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_193
timestamp 1688980957
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_205
timestamp 1688980957
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_217
timestamp 1688980957
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_223
timestamp 1688980957
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_225
timestamp 1688980957
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_237
timestamp 1688980957
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_249
timestamp 1688980957
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_261
timestamp 1688980957
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_273
timestamp 1688980957
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_279
timestamp 1688980957
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_281
timestamp 1688980957
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_293
timestamp 1688980957
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_305
timestamp 1688980957
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_317
timestamp 1688980957
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_329
timestamp 1688980957
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_335
timestamp 1688980957
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_337
timestamp 1688980957
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_349
timestamp 1688980957
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_361
timestamp 1688980957
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_373
timestamp 1688980957
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_385
timestamp 1688980957
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_391
timestamp 1688980957
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_393
timestamp 1688980957
transform 1 0 37260 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_405
timestamp 1688980957
transform 1 0 38364 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_417
timestamp 1688980957
transform 1 0 39468 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_429
timestamp 1688980957
transform 1 0 40572 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_441
timestamp 1688980957
transform 1 0 41676 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_447
timestamp 1688980957
transform 1 0 42228 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_449
timestamp 1688980957
transform 1 0 42412 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_461
timestamp 1688980957
transform 1 0 43516 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_473
timestamp 1688980957
transform 1 0 44620 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_479
timestamp 1688980957
transform 1 0 45172 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 1688980957
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 1688980957
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1688980957
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 1688980957
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_41
timestamp 1688980957
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_53
timestamp 1688980957
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_65
timestamp 1688980957
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_77
timestamp 1688980957
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_83
timestamp 1688980957
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_85
timestamp 1688980957
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_97
timestamp 1688980957
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_109
timestamp 1688980957
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_121
timestamp 1688980957
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_133
timestamp 1688980957
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_139
timestamp 1688980957
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_141
timestamp 1688980957
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_153
timestamp 1688980957
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_165
timestamp 1688980957
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_177
timestamp 1688980957
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_189
timestamp 1688980957
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_195
timestamp 1688980957
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_197
timestamp 1688980957
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_209
timestamp 1688980957
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_221
timestamp 1688980957
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_233
timestamp 1688980957
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_245
timestamp 1688980957
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_251
timestamp 1688980957
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_253
timestamp 1688980957
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_265
timestamp 1688980957
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_277
timestamp 1688980957
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_289
timestamp 1688980957
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_301
timestamp 1688980957
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_307
timestamp 1688980957
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_309
timestamp 1688980957
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_321
timestamp 1688980957
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_333
timestamp 1688980957
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_345
timestamp 1688980957
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_357
timestamp 1688980957
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_363
timestamp 1688980957
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_365
timestamp 1688980957
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_377
timestamp 1688980957
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_389
timestamp 1688980957
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_401
timestamp 1688980957
transform 1 0 37996 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_413
timestamp 1688980957
transform 1 0 39100 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_419
timestamp 1688980957
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_421
timestamp 1688980957
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_433
timestamp 1688980957
transform 1 0 40940 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_445
timestamp 1688980957
transform 1 0 42044 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_457
timestamp 1688980957
transform 1 0 43148 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_469
timestamp 1688980957
transform 1 0 44252 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_475
timestamp 1688980957
transform 1 0 44804 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_477
timestamp 1688980957
transform 1 0 44988 0 1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 1688980957
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_15
timestamp 1688980957
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_27
timestamp 1688980957
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_39
timestamp 1688980957
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_51
timestamp 1688980957
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_55
timestamp 1688980957
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_57
timestamp 1688980957
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_69
timestamp 1688980957
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_81
timestamp 1688980957
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_93
timestamp 1688980957
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_105
timestamp 1688980957
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_111
timestamp 1688980957
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_113
timestamp 1688980957
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_125
timestamp 1688980957
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_137
timestamp 1688980957
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_149
timestamp 1688980957
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_161
timestamp 1688980957
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_167
timestamp 1688980957
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_169
timestamp 1688980957
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_181
timestamp 1688980957
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_193
timestamp 1688980957
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_205
timestamp 1688980957
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_217
timestamp 1688980957
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_223
timestamp 1688980957
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_225
timestamp 1688980957
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_237
timestamp 1688980957
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_249
timestamp 1688980957
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_261
timestamp 1688980957
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_273
timestamp 1688980957
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_279
timestamp 1688980957
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_281
timestamp 1688980957
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_293
timestamp 1688980957
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_305
timestamp 1688980957
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_317
timestamp 1688980957
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_329
timestamp 1688980957
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_335
timestamp 1688980957
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_337
timestamp 1688980957
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_349
timestamp 1688980957
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_361
timestamp 1688980957
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_373
timestamp 1688980957
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_385
timestamp 1688980957
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_391
timestamp 1688980957
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_393
timestamp 1688980957
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_405
timestamp 1688980957
transform 1 0 38364 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_417
timestamp 1688980957
transform 1 0 39468 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_429
timestamp 1688980957
transform 1 0 40572 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_441
timestamp 1688980957
transform 1 0 41676 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_447
timestamp 1688980957
transform 1 0 42228 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_449
timestamp 1688980957
transform 1 0 42412 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_461
timestamp 1688980957
transform 1 0 43516 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_473
timestamp 1688980957
transform 1 0 44620 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_9
timestamp 1688980957
transform 1 0 1932 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_21
timestamp 1688980957
transform 1 0 3036 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 1688980957
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_29
timestamp 1688980957
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_41
timestamp 1688980957
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_53
timestamp 1688980957
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_65
timestamp 1688980957
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_77
timestamp 1688980957
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_83
timestamp 1688980957
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_85
timestamp 1688980957
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_97
timestamp 1688980957
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_109
timestamp 1688980957
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_121
timestamp 1688980957
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_133
timestamp 1688980957
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_139
timestamp 1688980957
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_141
timestamp 1688980957
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_153
timestamp 1688980957
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_165
timestamp 1688980957
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_177
timestamp 1688980957
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_189
timestamp 1688980957
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_195
timestamp 1688980957
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_197
timestamp 1688980957
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_209
timestamp 1688980957
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_221
timestamp 1688980957
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_233
timestamp 1688980957
transform 1 0 22540 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_245
timestamp 1688980957
transform 1 0 23644 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_251
timestamp 1688980957
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_253
timestamp 1688980957
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_265
timestamp 1688980957
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_277
timestamp 1688980957
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_289
timestamp 1688980957
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_301
timestamp 1688980957
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_307
timestamp 1688980957
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_309
timestamp 1688980957
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_321
timestamp 1688980957
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_333
timestamp 1688980957
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_345
timestamp 1688980957
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_357
timestamp 1688980957
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_363
timestamp 1688980957
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_365
timestamp 1688980957
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_377
timestamp 1688980957
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_389
timestamp 1688980957
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_401
timestamp 1688980957
transform 1 0 37996 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_413
timestamp 1688980957
transform 1 0 39100 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_419
timestamp 1688980957
transform 1 0 39652 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_421
timestamp 1688980957
transform 1 0 39836 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_433
timestamp 1688980957
transform 1 0 40940 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_445
timestamp 1688980957
transform 1 0 42044 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_457
timestamp 1688980957
transform 1 0 43148 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_463
timestamp 1688980957
transform 1 0 43700 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_477
timestamp 1688980957
transform 1 0 44988 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_3
timestamp 1688980957
transform 1 0 1380 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_17
timestamp 1688980957
transform 1 0 2668 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_29
timestamp 1688980957
transform 1 0 3772 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_41
timestamp 1688980957
transform 1 0 4876 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_53
timestamp 1688980957
transform 1 0 5980 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_57
timestamp 1688980957
transform 1 0 6348 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_69
timestamp 1688980957
transform 1 0 7452 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_81
timestamp 1688980957
transform 1 0 8556 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_93
timestamp 1688980957
transform 1 0 9660 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_105
timestamp 1688980957
transform 1 0 10764 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_111
timestamp 1688980957
transform 1 0 11316 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_113
timestamp 1688980957
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_125
timestamp 1688980957
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_137
timestamp 1688980957
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_149
timestamp 1688980957
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_161
timestamp 1688980957
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_167
timestamp 1688980957
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_169
timestamp 1688980957
transform 1 0 16652 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_177
timestamp 1688980957
transform 1 0 17388 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_181
timestamp 1688980957
transform 1 0 17756 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_189
timestamp 1688980957
transform 1 0 18492 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_196
timestamp 1688980957
transform 1 0 19136 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_200
timestamp 1688980957
transform 1 0 19504 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_205
timestamp 1688980957
transform 1 0 19964 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_217
timestamp 1688980957
transform 1 0 21068 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_223
timestamp 1688980957
transform 1 0 21620 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_225
timestamp 1688980957
transform 1 0 21804 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_241
timestamp 1688980957
transform 1 0 23276 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_245
timestamp 1688980957
transform 1 0 23644 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_252
timestamp 1688980957
transform 1 0 24288 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_264
timestamp 1688980957
transform 1 0 25392 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_276
timestamp 1688980957
transform 1 0 26496 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_281
timestamp 1688980957
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_293
timestamp 1688980957
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_305
timestamp 1688980957
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_317
timestamp 1688980957
transform 1 0 30268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_329
timestamp 1688980957
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_335
timestamp 1688980957
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_337
timestamp 1688980957
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_349
timestamp 1688980957
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_361
timestamp 1688980957
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_373
timestamp 1688980957
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_385
timestamp 1688980957
transform 1 0 36524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_391
timestamp 1688980957
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_393
timestamp 1688980957
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_405
timestamp 1688980957
transform 1 0 38364 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_417
timestamp 1688980957
transform 1 0 39468 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_429
timestamp 1688980957
transform 1 0 40572 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_441
timestamp 1688980957
transform 1 0 41676 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_447
timestamp 1688980957
transform 1 0 42228 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_449
timestamp 1688980957
transform 1 0 42412 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_457
timestamp 1688980957
transform 1 0 43148 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_476
timestamp 1688980957
transform 1 0 44896 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_3
timestamp 1688980957
transform 1 0 1380 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_7
timestamp 1688980957
transform 1 0 1748 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_35
timestamp 1688980957
transform 1 0 4324 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_40
timestamp 1688980957
transform 1 0 4784 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_52
timestamp 1688980957
transform 1 0 5888 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_62
timestamp 1688980957
transform 1 0 6808 0 1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_72
timestamp 1688980957
transform 1 0 7728 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_91
timestamp 1688980957
transform 1 0 9476 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_95
timestamp 1688980957
transform 1 0 9844 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_100
timestamp 1688980957
transform 1 0 10304 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_122
timestamp 1688980957
transform 1 0 12328 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_132
timestamp 1688980957
transform 1 0 13248 0 1 7616
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_147
timestamp 1688980957
transform 1 0 14628 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_159
timestamp 1688980957
transform 1 0 15732 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_171
timestamp 1688980957
transform 1 0 16836 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_197
timestamp 1688980957
transform 1 0 19228 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_277
timestamp 1688980957
transform 1 0 26588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_281
timestamp 1688980957
transform 1 0 26956 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_285
timestamp 1688980957
transform 1 0 27324 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_301
timestamp 1688980957
transform 1 0 28796 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_307
timestamp 1688980957
transform 1 0 29348 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_309
timestamp 1688980957
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_321
timestamp 1688980957
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_333
timestamp 1688980957
transform 1 0 31740 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_345
timestamp 1688980957
transform 1 0 32844 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_357
timestamp 1688980957
transform 1 0 33948 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_363
timestamp 1688980957
transform 1 0 34500 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_365
timestamp 1688980957
transform 1 0 34684 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_377
timestamp 1688980957
transform 1 0 35788 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_389
timestamp 1688980957
transform 1 0 36892 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_401
timestamp 1688980957
transform 1 0 37996 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_413
timestamp 1688980957
transform 1 0 39100 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_419
timestamp 1688980957
transform 1 0 39652 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_421
timestamp 1688980957
transform 1 0 39836 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_437
timestamp 1688980957
transform 1 0 41308 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_449
timestamp 1688980957
transform 1 0 42412 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_474
timestamp 1688980957
transform 1 0 44712 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_477
timestamp 1688980957
transform 1 0 44988 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_3
timestamp 1688980957
transform 1 0 1380 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_8
timestamp 1688980957
transform 1 0 1840 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_14
timestamp 1688980957
transform 1 0 2392 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_29
timestamp 1688980957
transform 1 0 3772 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_34
timestamp 1688980957
transform 1 0 4232 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_61
timestamp 1688980957
transform 1 0 6716 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_68
timestamp 1688980957
transform 1 0 7360 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_85
timestamp 1688980957
transform 1 0 8924 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_96
timestamp 1688980957
transform 1 0 9936 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_113
timestamp 1688980957
transform 1 0 11500 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_128
timestamp 1688980957
transform 1 0 12880 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_141
timestamp 1688980957
transform 1 0 14076 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_175
timestamp 1688980957
transform 1 0 17204 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_194
timestamp 1688980957
transform 1 0 18952 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_197
timestamp 1688980957
transform 1 0 19228 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_208
timestamp 1688980957
transform 1 0 20240 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_240
timestamp 1688980957
transform 1 0 23184 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_245
timestamp 1688980957
transform 1 0 23644 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_253
timestamp 1688980957
transform 1 0 24380 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_269
timestamp 1688980957
transform 1 0 25852 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_273
timestamp 1688980957
transform 1 0 26220 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_277
timestamp 1688980957
transform 1 0 26588 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_293
timestamp 1688980957
transform 1 0 28060 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_297
timestamp 1688980957
transform 1 0 28428 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_301
timestamp 1688980957
transform 1 0 28796 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_305
timestamp 1688980957
transform 1 0 29164 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_321
timestamp 1688980957
transform 1 0 30636 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_325
timestamp 1688980957
transform 1 0 31004 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_329
timestamp 1688980957
transform 1 0 31372 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_333
timestamp 1688980957
transform 1 0 31740 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_349
timestamp 1688980957
transform 1 0 33212 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_353
timestamp 1688980957
transform 1 0 33580 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_357
timestamp 1688980957
transform 1 0 33948 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_361
timestamp 1688980957
transform 1 0 34316 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_377
timestamp 1688980957
transform 1 0 35788 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_381
timestamp 1688980957
transform 1 0 36156 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_385
timestamp 1688980957
transform 1 0 36524 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_389
timestamp 1688980957
transform 1 0 36892 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_405
timestamp 1688980957
transform 1 0 38364 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_409
timestamp 1688980957
transform 1 0 38732 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_443
timestamp 1688980957
transform 1 0 41860 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_447
timestamp 1688980957
transform 1 0 42228 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_473
timestamp 1688980957
transform 1 0 44620 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_477
timestamp 1688980957
transform 1 0 44988 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3772 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 25576 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1688980957
transform 1 0 27784 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1688980957
transform 1 0 29992 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1688980957
transform 1 0 32200 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1688980957
transform 1 0 34684 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1688980957
transform 1 0 36616 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1688980957
transform 1 0 38824 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1688980957
transform 1 0 41032 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1688980957
transform 1 0 43240 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1688980957
transform 1 0 44988 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input12
timestamp 1688980957
transform 1 0 5704 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input13
timestamp 1688980957
transform 1 0 7912 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input14
timestamp 1688980957
transform 1 0 10120 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input15
timestamp 1688980957
transform 1 0 12328 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1688980957
transform 1 0 14536 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1688980957
transform 1 0 16744 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1688980957
transform 1 0 19228 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1688980957
transform 1 0 21160 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1688980957
transform 1 0 23368 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1688980957
transform 1 0 19688 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1688980957
transform 1 0 19412 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1688980957
transform 1 0 20332 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 1688980957
transform 1 0 20608 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1688980957
transform 1 0 20884 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 1688980957
transform 1 0 21160 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1688980957
transform 1 0 21436 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1688980957
transform 1 0 21804 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1688980957
transform 1 0 22080 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1688980957
transform 1 0 22356 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1688980957
transform 1 0 23368 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 1688980957
transform 1 0 24012 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1688980957
transform 1 0 24748 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input34
timestamp 1688980957
transform 1 0 24472 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input35
timestamp 1688980957
transform 1 0 25024 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input36
timestamp 1688980957
transform 1 0 25300 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 1688980957
transform 1 0 25576 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input38
timestamp 1688980957
transform 1 0 25944 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input39
timestamp 1688980957
transform 1 0 26312 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input40
timestamp 1688980957
transform 1 0 26956 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input41
timestamp 1688980957
transform 1 0 27232 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input42
timestamp 1688980957
transform 1 0 30728 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input43
timestamp 1688980957
transform 1 0 31096 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input44
timestamp 1688980957
transform 1 0 31464 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input45
timestamp 1688980957
transform 1 0 32108 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input46
timestamp 1688980957
transform 1 0 32384 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input47
timestamp 1688980957
transform 1 0 32660 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input48
timestamp 1688980957
transform 1 0 27508 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input49
timestamp 1688980957
transform 1 0 27784 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input50
timestamp 1688980957
transform 1 0 28152 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input51
timestamp 1688980957
transform 1 0 28520 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input52
timestamp 1688980957
transform 1 0 28888 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input53
timestamp 1688980957
transform 1 0 29532 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input54
timestamp 1688980957
transform 1 0 29808 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input55
timestamp 1688980957
transform 1 0 30084 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input56
timestamp 1688980957
transform 1 0 30360 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input57
timestamp 1688980957
transform 1 0 32936 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input58
timestamp 1688980957
transform 1 0 36616 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input59
timestamp 1688980957
transform 1 0 37260 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input60
timestamp 1688980957
transform 1 0 37536 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input61
timestamp 1688980957
transform 1 0 37812 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input62
timestamp 1688980957
transform 1 0 38088 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input63
timestamp 1688980957
transform 1 0 38456 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input64
timestamp 1688980957
transform 1 0 33304 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input65
timestamp 1688980957
transform 1 0 33672 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input66
timestamp 1688980957
transform 1 0 34040 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input67
timestamp 1688980957
transform 1 0 34684 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input68
timestamp 1688980957
transform 1 0 34960 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input69
timestamp 1688980957
transform 1 0 35236 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input70
timestamp 1688980957
transform 1 0 35512 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input71
timestamp 1688980957
transform 1 0 35880 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input72
timestamp 1688980957
transform 1 0 36248 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input73
timestamp 1688980957
transform 1 0 1380 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  inst_clk_buf dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 19964 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_single2_switch_matrix__00_
timestamp 1688980957
transform 1 0 26036 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_single2_switch_matrix__01_
timestamp 1688980957
transform 1 0 25760 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_single2_switch_matrix__02_
timestamp 1688980957
transform 1 0 25484 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_single2_switch_matrix__03_
timestamp 1688980957
transform 1 0 25208 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_single2_switch_matrix__04_
timestamp 1688980957
transform 1 0 24932 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_single2_switch_matrix__05_
timestamp 1688980957
transform 1 0 24012 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_single2_switch_matrix__06_
timestamp 1688980957
transform 1 0 23736 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_single2_switch_matrix__07_
timestamp 1688980957
transform 1 0 22908 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_single2_switch_matrix__08_
timestamp 1688980957
transform 1 0 23000 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_single2_switch_matrix__09_
timestamp 1688980957
transform 1 0 22632 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_single2_switch_matrix__10_
timestamp 1688980957
transform 1 0 22172 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_single2_switch_matrix__11_
timestamp 1688980957
transform 1 0 21896 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_single2_switch_matrix__12_
timestamp 1688980957
transform 1 0 21252 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_single2_switch_matrix__13_
timestamp 1688980957
transform 1 0 20976 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_single2_switch_matrix__14_
timestamp 1688980957
transform 1 0 20700 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_single2_switch_matrix__15_
timestamp 1688980957
transform 1 0 20148 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_single2_switch_matrix__16_
timestamp 1688980957
transform 1 0 23368 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_single2_switch_matrix__17_
timestamp 1688980957
transform 1 0 23736 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_single2_switch_matrix__18_
timestamp 1688980957
transform 1 0 28244 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_single2_switch_matrix__19_
timestamp 1688980957
transform 1 0 27968 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_single2_switch_matrix__20_
timestamp 1688980957
transform 1 0 27416 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_single2_switch_matrix__21_
timestamp 1688980957
transform 1 0 27048 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_single2_switch_matrix__22_
timestamp 1688980957
transform 1 0 26680 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_single2_switch_matrix__23_
timestamp 1688980957
transform 1 0 26312 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_single2_switch_matrix__24_
timestamp 1688980957
transform 1 0 23184 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_single2_switch_matrix__25_
timestamp 1688980957
transform 1 0 23460 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_single2_switch_matrix__26_
timestamp 1688980957
transform 1 0 23736 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_single2_switch_matrix__27_
timestamp 1688980957
transform 1 0 24012 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_single2_switch_matrix__28_
timestamp 1688980957
transform 1 0 24380 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_single2_switch_matrix__29_
timestamp 1688980957
transform 1 0 24656 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_single2_switch_matrix__30_
timestamp 1688980957
transform 1 0 27692 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_single2_switch_matrix__31_
timestamp 1688980957
transform 1 0 28520 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_single2_switch_matrix__32_
timestamp 1688980957
transform 1 0 22908 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_single2_switch_matrix__33_
timestamp 1688980957
transform 1 0 22724 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_single2_switch_matrix__34_
timestamp 1688980957
transform 1 0 17480 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_single2_switch_matrix__35_
timestamp 1688980957
transform 1 0 17756 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_single2_switch_matrix__36_
timestamp 1688980957
transform 1 0 18032 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_single2_switch_matrix__37_
timestamp 1688980957
transform 1 0 18860 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_single2_switch_matrix__38_
timestamp 1688980957
transform 1 0 19228 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_single2_switch_matrix__39_
timestamp 1688980957
transform 1 0 18584 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_single2_switch_matrix__40_
timestamp 1688980957
transform 1 0 22632 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_single2_switch_matrix__41_
timestamp 1688980957
transform 1 0 22356 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_single2_switch_matrix__42_
timestamp 1688980957
transform 1 0 21804 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_single2_switch_matrix__43_
timestamp 1688980957
transform 1 0 22080 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_single2_switch_matrix__44_
timestamp 1688980957
transform 1 0 22448 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_single2_switch_matrix__45_
timestamp 1688980957
transform 1 0 21528 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_single2_switch_matrix__46_
timestamp 1688980957
transform 1 0 20424 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_single2_switch_matrix__47_
timestamp 1688980957
transform 1 0 17480 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_single2_switch_matrix__48_
timestamp 1688980957
transform 1 0 19872 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_single2_switch_matrix__49_
timestamp 1688980957
transform 1 0 18860 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_single2_switch_matrix__50_
timestamp 1688980957
transform 1 0 18308 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_single2_switch_matrix__51_
timestamp 1688980957
transform 1 0 18584 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output74 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 39376 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output75 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 43056 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output76
timestamp 1688980957
transform 1 0 43240 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output77
timestamp 1688980957
transform 1 0 43608 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output78
timestamp 1688980957
transform 1 0 44160 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output79
timestamp 1688980957
transform 1 0 42504 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output80
timestamp 1688980957
transform 1 0 44712 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output81
timestamp 1688980957
transform 1 0 44344 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output82
timestamp 1688980957
transform 1 0 44344 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output83
timestamp 1688980957
transform 1 0 43792 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output84
timestamp 1688980957
transform 1 0 43792 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output85
timestamp 1688980957
transform 1 0 39836 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output86
timestamp 1688980957
transform 1 0 40388 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output87
timestamp 1688980957
transform 1 0 40940 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output88
timestamp 1688980957
transform 1 0 40940 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output89
timestamp 1688980957
transform 1 0 41308 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output90
timestamp 1688980957
transform 1 0 42412 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output91
timestamp 1688980957
transform 1 0 42964 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output92
timestamp 1688980957
transform 1 0 43516 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output93
timestamp 1688980957
transform 1 0 44068 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output94
timestamp 1688980957
transform 1 0 2576 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output95
timestamp 1688980957
transform 1 0 1564 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output96
timestamp 1688980957
transform 1 0 1380 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output97
timestamp 1688980957
transform 1 0 2116 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output98
timestamp 1688980957
transform 1 0 1840 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output99
timestamp 1688980957
transform -1 0 2392 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output100
timestamp 1688980957
transform 1 0 2392 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output101
timestamp 1688980957
transform 1 0 2944 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output102
timestamp 1688980957
transform 1 0 3312 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output103
timestamp 1688980957
transform 1 0 3772 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output104
timestamp 1688980957
transform 1 0 3128 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output105
timestamp 1688980957
transform 1 0 4416 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output106
timestamp 1688980957
transform -1 0 4784 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output107
timestamp 1688980957
transform 1 0 4784 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output108
timestamp 1688980957
transform 1 0 5152 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output109
timestamp 1688980957
transform 1 0 6348 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output110
timestamp 1688980957
transform 1 0 6256 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output111
timestamp 1688980957
transform 1 0 5704 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output112
timestamp 1688980957
transform 1 0 6808 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output113
timestamp 1688980957
transform 1 0 7360 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output114
timestamp 1688980957
transform 1 0 7544 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output115
timestamp 1688980957
transform 1 0 11408 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output116
timestamp 1688980957
transform 1 0 11960 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output117
timestamp 1688980957
transform 1 0 11776 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output118
timestamp 1688980957
transform 1 0 12328 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output119
timestamp 1688980957
transform 1 0 12880 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output120
timestamp 1688980957
transform 1 0 13064 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output121
timestamp 1688980957
transform 1 0 7912 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output122
timestamp 1688980957
transform 1 0 8464 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output123
timestamp 1688980957
transform 1 0 8924 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output124
timestamp 1688980957
transform 1 0 9016 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output125
timestamp 1688980957
transform 1 0 9384 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output126
timestamp 1688980957
transform 1 0 9936 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output127
timestamp 1688980957
transform 1 0 10120 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output128
timestamp 1688980957
transform 1 0 10488 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output129
timestamp 1688980957
transform 1 0 10856 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output130
timestamp 1688980957
transform 1 0 13432 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output131
timestamp 1688980957
transform 1 0 17296 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output132
timestamp 1688980957
transform 1 0 17664 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output133
timestamp 1688980957
transform 1 0 18216 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output134
timestamp 1688980957
transform 1 0 18584 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output135
timestamp 1688980957
transform 1 0 19688 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output136
timestamp 1688980957
transform 1 0 19320 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output137
timestamp 1688980957
transform 1 0 14076 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output138
timestamp 1688980957
transform 1 0 14168 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output139
timestamp 1688980957
transform 1 0 14536 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output140
timestamp 1688980957
transform 1 0 14904 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output141
timestamp 1688980957
transform 1 0 15456 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output142
timestamp 1688980957
transform 1 0 15824 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output143
timestamp 1688980957
transform 1 0 16192 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output144
timestamp 1688980957
transform 1 0 16652 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output145
timestamp 1688980957
transform 1 0 17112 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output146
timestamp 1688980957
transform 1 0 38824 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1688980957
transform 1 0 1104 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1688980957
transform -1 0 45540 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1688980957
transform 1 0 1104 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1688980957
transform -1 0 45540 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1688980957
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1688980957
transform -1 0 45540 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1688980957
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1688980957
transform -1 0 45540 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1688980957
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1688980957
transform -1 0 45540 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1688980957
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1688980957
transform -1 0 45540 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1688980957
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1688980957
transform -1 0 45540 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1688980957
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1688980957
transform -1 0 45540 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1688980957
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1688980957
transform -1 0 45540 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1688980957
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1688980957
transform -1 0 45540 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1688980957
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1688980957
transform -1 0 45540 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1688980957
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1688980957
transform -1 0 45540 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1688980957
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1688980957
transform -1 0 45540 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1688980957
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1688980957
transform -1 0 45540 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_0__0_
timestamp 1688980957
transform 1 0 23368 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_1__0_
timestamp 1688980957
transform 1 0 21988 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_2__0_
timestamp 1688980957
transform 1 0 22540 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_3__0_
timestamp 1688980957
transform 1 0 23092 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_4__0_
timestamp 1688980957
transform 1 0 22264 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_5__0_
timestamp 1688980957
transform 1 0 22080 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_6__0_
timestamp 1688980957
transform 1 0 21160 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_7__0_
timestamp 1688980957
transform 1 0 19412 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_8__0_
timestamp 1688980957
transform 1 0 21436 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_9__0_
timestamp 1688980957
transform 1 0 23828 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_10__0_
timestamp 1688980957
transform 1 0 26036 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_11__0_
timestamp 1688980957
transform 1 0 28244 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_12__0_
timestamp 1688980957
transform 1 0 30452 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_13__0_
timestamp 1688980957
transform 1 0 32660 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_14__0_
timestamp 1688980957
transform 1 0 34868 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_15__0_
timestamp 1688980957
transform 1 0 37260 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_16__0_
timestamp 1688980957
transform 1 0 43424 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_17__0_
timestamp 1688980957
transform 1 0 41584 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_18__0_
timestamp 1688980957
transform 1 0 43884 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_19__0_
timestamp 1688980957
transform 1 0 44344 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  strobe_outbuf_0__0_
timestamp 1688980957
transform 1 0 23736 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  strobe_outbuf_1__0_
timestamp 1688980957
transform 1 0 22908 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  strobe_outbuf_2__0_
timestamp 1688980957
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  strobe_outbuf_3__0_
timestamp 1688980957
transform 1 0 23460 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  strobe_outbuf_4__0_
timestamp 1688980957
transform 1 0 23184 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  strobe_outbuf_5__0_
timestamp 1688980957
transform 1 0 22816 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  strobe_outbuf_6__0_
timestamp 1688980957
transform 1 0 22172 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  strobe_outbuf_7__0_
timestamp 1688980957
transform 1 0 20240 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  strobe_outbuf_8__0_
timestamp 1688980957
transform 1 0 22448 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  strobe_outbuf_9__0_
timestamp 1688980957
transform 1 0 24656 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  strobe_outbuf_10__0_
timestamp 1688980957
transform 1 0 26864 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  strobe_outbuf_11__0_
timestamp 1688980957
transform 1 0 29072 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  strobe_outbuf_12__0_
timestamp 1688980957
transform 1 0 31280 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  strobe_outbuf_13__0_
timestamp 1688980957
transform 1 0 33488 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  strobe_outbuf_14__0_
timestamp 1688980957
transform 1 0 35696 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  strobe_outbuf_15__0_
timestamp 1688980957
transform 1 0 37904 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_16__0_
timestamp 1688980957
transform 1 0 44160 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_17__0_
timestamp 1688980957
transform 1 0 44436 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_18__0_
timestamp 1688980957
transform 1 0 44988 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_19__0_
timestamp 1688980957
transform 1 0 43884 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_28 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3680 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_29
timestamp 1688980957
transform 1 0 6256 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_30
timestamp 1688980957
transform 1 0 8832 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_31
timestamp 1688980957
transform 1 0 11408 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_32
timestamp 1688980957
transform 1 0 13984 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_33
timestamp 1688980957
transform 1 0 16560 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_34
timestamp 1688980957
transform 1 0 19136 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_35
timestamp 1688980957
transform 1 0 21712 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_36
timestamp 1688980957
transform 1 0 24288 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_37
timestamp 1688980957
transform 1 0 26864 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_38
timestamp 1688980957
transform 1 0 29440 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_39
timestamp 1688980957
transform 1 0 32016 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_40
timestamp 1688980957
transform 1 0 34592 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_41
timestamp 1688980957
transform 1 0 37168 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_42
timestamp 1688980957
transform 1 0 39744 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_43
timestamp 1688980957
transform 1 0 42320 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_44
timestamp 1688980957
transform 1 0 44896 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_45
timestamp 1688980957
transform 1 0 6256 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_46
timestamp 1688980957
transform 1 0 11408 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_47
timestamp 1688980957
transform 1 0 16560 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_48
timestamp 1688980957
transform 1 0 21712 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_49
timestamp 1688980957
transform 1 0 26864 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_50
timestamp 1688980957
transform 1 0 32016 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_51
timestamp 1688980957
transform 1 0 37168 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_52
timestamp 1688980957
transform 1 0 42320 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_53
timestamp 1688980957
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_54
timestamp 1688980957
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_55
timestamp 1688980957
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56
timestamp 1688980957
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1688980957
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1688980957
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1688980957
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1688980957
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1688980957
transform 1 0 44896 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1688980957
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1688980957
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1688980957
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1688980957
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 1688980957
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 1688980957
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 1688980957
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1688980957
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1688980957
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1688980957
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1688980957
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1688980957
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1688980957
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1688980957
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1688980957
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1688980957
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1688980957
transform 1 0 44896 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1688980957
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1688980957
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1688980957
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1688980957
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1688980957
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1688980957
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1688980957
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1688980957
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1688980957
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1688980957
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1688980957
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1688980957
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1688980957
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1688980957
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1688980957
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1688980957
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1688980957
transform 1 0 44896 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1688980957
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1688980957
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1688980957
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1688980957
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1688980957
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1688980957
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1688980957
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1688980957
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1688980957
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1688980957
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1688980957
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1688980957
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1688980957
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1688980957
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1688980957
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1688980957
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1688980957
transform 1 0 44896 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1688980957
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1688980957
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1688980957
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1688980957
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1688980957
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1688980957
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1688980957
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1688980957
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1688980957
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1688980957
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1688980957
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1688980957
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1688980957
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1688980957
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1688980957
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1688980957
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1688980957
transform 1 0 44896 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1688980957
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1688980957
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1688980957
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1688980957
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1688980957
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1688980957
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1688980957
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1688980957
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1688980957
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1688980957
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1688980957
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1688980957
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1688980957
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1688980957
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1688980957
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1688980957
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1688980957
transform 1 0 44896 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1688980957
transform 1 0 3680 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1688980957
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1688980957
transform 1 0 8832 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1688980957
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1688980957
transform 1 0 13984 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1688980957
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1688980957
transform 1 0 19136 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1688980957
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1688980957
transform 1 0 24288 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156
timestamp 1688980957
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1688980957
transform 1 0 29440 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1688980957
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1688980957
transform 1 0 34592 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1688980957
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1688980957
transform 1 0 39744 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1688980957
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1688980957
transform 1 0 44896 0 -1 8704
box -38 -48 130 592
<< labels >>
flabel metal2 s 3422 -300 3478 160 0 FreeSans 224 90 0 0 FrameStrobe[0]
port 0 nsew signal input
flabel metal2 s 25502 -300 25558 160 0 FreeSans 224 90 0 0 FrameStrobe[10]
port 1 nsew signal input
flabel metal2 s 27710 -300 27766 160 0 FreeSans 224 90 0 0 FrameStrobe[11]
port 2 nsew signal input
flabel metal2 s 29918 -300 29974 160 0 FreeSans 224 90 0 0 FrameStrobe[12]
port 3 nsew signal input
flabel metal2 s 32126 -300 32182 160 0 FreeSans 224 90 0 0 FrameStrobe[13]
port 4 nsew signal input
flabel metal2 s 34334 -300 34390 160 0 FreeSans 224 90 0 0 FrameStrobe[14]
port 5 nsew signal input
flabel metal2 s 36542 -300 36598 160 0 FreeSans 224 90 0 0 FrameStrobe[15]
port 6 nsew signal input
flabel metal2 s 38750 -300 38806 160 0 FreeSans 224 90 0 0 FrameStrobe[16]
port 7 nsew signal input
flabel metal2 s 40958 -300 41014 160 0 FreeSans 224 90 0 0 FrameStrobe[17]
port 8 nsew signal input
flabel metal2 s 43166 -300 43222 160 0 FreeSans 224 90 0 0 FrameStrobe[18]
port 9 nsew signal input
flabel metal2 s 45374 -300 45430 160 0 FreeSans 224 90 0 0 FrameStrobe[19]
port 10 nsew signal input
flabel metal2 s 5630 -300 5686 160 0 FreeSans 224 90 0 0 FrameStrobe[1]
port 11 nsew signal input
flabel metal2 s 7838 -300 7894 160 0 FreeSans 224 90 0 0 FrameStrobe[2]
port 12 nsew signal input
flabel metal2 s 10046 -300 10102 160 0 FreeSans 224 90 0 0 FrameStrobe[3]
port 13 nsew signal input
flabel metal2 s 12254 -300 12310 160 0 FreeSans 224 90 0 0 FrameStrobe[4]
port 14 nsew signal input
flabel metal2 s 14462 -300 14518 160 0 FreeSans 224 90 0 0 FrameStrobe[5]
port 15 nsew signal input
flabel metal2 s 16670 -300 16726 160 0 FreeSans 224 90 0 0 FrameStrobe[6]
port 16 nsew signal input
flabel metal2 s 18878 -300 18934 160 0 FreeSans 224 90 0 0 FrameStrobe[7]
port 17 nsew signal input
flabel metal2 s 21086 -300 21142 160 0 FreeSans 224 90 0 0 FrameStrobe[8]
port 18 nsew signal input
flabel metal2 s 23294 -300 23350 160 0 FreeSans 224 90 0 0 FrameStrobe[9]
port 19 nsew signal input
flabel metal2 s 39118 9840 39174 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[0]
port 20 nsew signal tristate
flabel metal2 s 42798 9840 42854 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[10]
port 21 nsew signal tristate
flabel metal2 s 43166 9840 43222 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[11]
port 22 nsew signal tristate
flabel metal2 s 43534 9840 43590 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[12]
port 23 nsew signal tristate
flabel metal2 s 43902 9840 43958 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[13]
port 24 nsew signal tristate
flabel metal2 s 44270 9840 44326 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[14]
port 25 nsew signal tristate
flabel metal2 s 44638 9840 44694 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[15]
port 26 nsew signal tristate
flabel metal2 s 45006 9840 45062 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[16]
port 27 nsew signal tristate
flabel metal2 s 45374 9840 45430 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[17]
port 28 nsew signal tristate
flabel metal2 s 45742 9840 45798 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[18]
port 29 nsew signal tristate
flabel metal2 s 46110 9840 46166 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[19]
port 30 nsew signal tristate
flabel metal2 s 39486 9840 39542 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[1]
port 31 nsew signal tristate
flabel metal2 s 39854 9840 39910 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[2]
port 32 nsew signal tristate
flabel metal2 s 40222 9840 40278 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[3]
port 33 nsew signal tristate
flabel metal2 s 40590 9840 40646 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[4]
port 34 nsew signal tristate
flabel metal2 s 40958 9840 41014 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[5]
port 35 nsew signal tristate
flabel metal2 s 41326 9840 41382 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[6]
port 36 nsew signal tristate
flabel metal2 s 41694 9840 41750 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[7]
port 37 nsew signal tristate
flabel metal2 s 42062 9840 42118 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[8]
port 38 nsew signal tristate
flabel metal2 s 42430 9840 42486 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[9]
port 39 nsew signal tristate
flabel metal2 s 478 9840 534 10300 0 FreeSans 224 90 0 0 N1BEG[0]
port 40 nsew signal tristate
flabel metal2 s 846 9840 902 10300 0 FreeSans 224 90 0 0 N1BEG[1]
port 41 nsew signal tristate
flabel metal2 s 1214 9840 1270 10300 0 FreeSans 224 90 0 0 N1BEG[2]
port 42 nsew signal tristate
flabel metal2 s 1582 9840 1638 10300 0 FreeSans 224 90 0 0 N1BEG[3]
port 43 nsew signal tristate
flabel metal2 s 1950 9840 2006 10300 0 FreeSans 224 90 0 0 N2BEG[0]
port 44 nsew signal tristate
flabel metal2 s 2318 9840 2374 10300 0 FreeSans 224 90 0 0 N2BEG[1]
port 45 nsew signal tristate
flabel metal2 s 2686 9840 2742 10300 0 FreeSans 224 90 0 0 N2BEG[2]
port 46 nsew signal tristate
flabel metal2 s 3054 9840 3110 10300 0 FreeSans 224 90 0 0 N2BEG[3]
port 47 nsew signal tristate
flabel metal2 s 3422 9840 3478 10300 0 FreeSans 224 90 0 0 N2BEG[4]
port 48 nsew signal tristate
flabel metal2 s 3790 9840 3846 10300 0 FreeSans 224 90 0 0 N2BEG[5]
port 49 nsew signal tristate
flabel metal2 s 4158 9840 4214 10300 0 FreeSans 224 90 0 0 N2BEG[6]
port 50 nsew signal tristate
flabel metal2 s 4526 9840 4582 10300 0 FreeSans 224 90 0 0 N2BEG[7]
port 51 nsew signal tristate
flabel metal2 s 4894 9840 4950 10300 0 FreeSans 224 90 0 0 N2BEGb[0]
port 52 nsew signal tristate
flabel metal2 s 5262 9840 5318 10300 0 FreeSans 224 90 0 0 N2BEGb[1]
port 53 nsew signal tristate
flabel metal2 s 5630 9840 5686 10300 0 FreeSans 224 90 0 0 N2BEGb[2]
port 54 nsew signal tristate
flabel metal2 s 5998 9840 6054 10300 0 FreeSans 224 90 0 0 N2BEGb[3]
port 55 nsew signal tristate
flabel metal2 s 6366 9840 6422 10300 0 FreeSans 224 90 0 0 N2BEGb[4]
port 56 nsew signal tristate
flabel metal2 s 6734 9840 6790 10300 0 FreeSans 224 90 0 0 N2BEGb[5]
port 57 nsew signal tristate
flabel metal2 s 7102 9840 7158 10300 0 FreeSans 224 90 0 0 N2BEGb[6]
port 58 nsew signal tristate
flabel metal2 s 7470 9840 7526 10300 0 FreeSans 224 90 0 0 N2BEGb[7]
port 59 nsew signal tristate
flabel metal2 s 7838 9840 7894 10300 0 FreeSans 224 90 0 0 N4BEG[0]
port 60 nsew signal tristate
flabel metal2 s 11518 9840 11574 10300 0 FreeSans 224 90 0 0 N4BEG[10]
port 61 nsew signal tristate
flabel metal2 s 11886 9840 11942 10300 0 FreeSans 224 90 0 0 N4BEG[11]
port 62 nsew signal tristate
flabel metal2 s 12254 9840 12310 10300 0 FreeSans 224 90 0 0 N4BEG[12]
port 63 nsew signal tristate
flabel metal2 s 12622 9840 12678 10300 0 FreeSans 224 90 0 0 N4BEG[13]
port 64 nsew signal tristate
flabel metal2 s 12990 9840 13046 10300 0 FreeSans 224 90 0 0 N4BEG[14]
port 65 nsew signal tristate
flabel metal2 s 13358 9840 13414 10300 0 FreeSans 224 90 0 0 N4BEG[15]
port 66 nsew signal tristate
flabel metal2 s 8206 9840 8262 10300 0 FreeSans 224 90 0 0 N4BEG[1]
port 67 nsew signal tristate
flabel metal2 s 8574 9840 8630 10300 0 FreeSans 224 90 0 0 N4BEG[2]
port 68 nsew signal tristate
flabel metal2 s 8942 9840 8998 10300 0 FreeSans 224 90 0 0 N4BEG[3]
port 69 nsew signal tristate
flabel metal2 s 9310 9840 9366 10300 0 FreeSans 224 90 0 0 N4BEG[4]
port 70 nsew signal tristate
flabel metal2 s 9678 9840 9734 10300 0 FreeSans 224 90 0 0 N4BEG[5]
port 71 nsew signal tristate
flabel metal2 s 10046 9840 10102 10300 0 FreeSans 224 90 0 0 N4BEG[6]
port 72 nsew signal tristate
flabel metal2 s 10414 9840 10470 10300 0 FreeSans 224 90 0 0 N4BEG[7]
port 73 nsew signal tristate
flabel metal2 s 10782 9840 10838 10300 0 FreeSans 224 90 0 0 N4BEG[8]
port 74 nsew signal tristate
flabel metal2 s 11150 9840 11206 10300 0 FreeSans 224 90 0 0 N4BEG[9]
port 75 nsew signal tristate
flabel metal2 s 13726 9840 13782 10300 0 FreeSans 224 90 0 0 NN4BEG[0]
port 76 nsew signal tristate
flabel metal2 s 17406 9840 17462 10300 0 FreeSans 224 90 0 0 NN4BEG[10]
port 77 nsew signal tristate
flabel metal2 s 17774 9840 17830 10300 0 FreeSans 224 90 0 0 NN4BEG[11]
port 78 nsew signal tristate
flabel metal2 s 18142 9840 18198 10300 0 FreeSans 224 90 0 0 NN4BEG[12]
port 79 nsew signal tristate
flabel metal2 s 18510 9840 18566 10300 0 FreeSans 224 90 0 0 NN4BEG[13]
port 80 nsew signal tristate
flabel metal2 s 18878 9840 18934 10300 0 FreeSans 224 90 0 0 NN4BEG[14]
port 81 nsew signal tristate
flabel metal2 s 19246 9840 19302 10300 0 FreeSans 224 90 0 0 NN4BEG[15]
port 82 nsew signal tristate
flabel metal2 s 14094 9840 14150 10300 0 FreeSans 224 90 0 0 NN4BEG[1]
port 83 nsew signal tristate
flabel metal2 s 14462 9840 14518 10300 0 FreeSans 224 90 0 0 NN4BEG[2]
port 84 nsew signal tristate
flabel metal2 s 14830 9840 14886 10300 0 FreeSans 224 90 0 0 NN4BEG[3]
port 85 nsew signal tristate
flabel metal2 s 15198 9840 15254 10300 0 FreeSans 224 90 0 0 NN4BEG[4]
port 86 nsew signal tristate
flabel metal2 s 15566 9840 15622 10300 0 FreeSans 224 90 0 0 NN4BEG[5]
port 87 nsew signal tristate
flabel metal2 s 15934 9840 15990 10300 0 FreeSans 224 90 0 0 NN4BEG[6]
port 88 nsew signal tristate
flabel metal2 s 16302 9840 16358 10300 0 FreeSans 224 90 0 0 NN4BEG[7]
port 89 nsew signal tristate
flabel metal2 s 16670 9840 16726 10300 0 FreeSans 224 90 0 0 NN4BEG[8]
port 90 nsew signal tristate
flabel metal2 s 17038 9840 17094 10300 0 FreeSans 224 90 0 0 NN4BEG[9]
port 91 nsew signal tristate
flabel metal2 s 19614 9840 19670 10300 0 FreeSans 224 90 0 0 S1END[0]
port 92 nsew signal input
flabel metal2 s 19982 9840 20038 10300 0 FreeSans 224 90 0 0 S1END[1]
port 93 nsew signal input
flabel metal2 s 20350 9840 20406 10300 0 FreeSans 224 90 0 0 S1END[2]
port 94 nsew signal input
flabel metal2 s 20718 9840 20774 10300 0 FreeSans 224 90 0 0 S1END[3]
port 95 nsew signal input
flabel metal2 s 21086 9840 21142 10300 0 FreeSans 224 90 0 0 S2END[0]
port 96 nsew signal input
flabel metal2 s 21454 9840 21510 10300 0 FreeSans 224 90 0 0 S2END[1]
port 97 nsew signal input
flabel metal2 s 21822 9840 21878 10300 0 FreeSans 224 90 0 0 S2END[2]
port 98 nsew signal input
flabel metal2 s 22190 9840 22246 10300 0 FreeSans 224 90 0 0 S2END[3]
port 99 nsew signal input
flabel metal2 s 22558 9840 22614 10300 0 FreeSans 224 90 0 0 S2END[4]
port 100 nsew signal input
flabel metal2 s 22926 9840 22982 10300 0 FreeSans 224 90 0 0 S2END[5]
port 101 nsew signal input
flabel metal2 s 23294 9840 23350 10300 0 FreeSans 224 90 0 0 S2END[6]
port 102 nsew signal input
flabel metal2 s 23662 9840 23718 10300 0 FreeSans 224 90 0 0 S2END[7]
port 103 nsew signal input
flabel metal2 s 24030 9840 24086 10300 0 FreeSans 224 90 0 0 S2MID[0]
port 104 nsew signal input
flabel metal2 s 24398 9840 24454 10300 0 FreeSans 224 90 0 0 S2MID[1]
port 105 nsew signal input
flabel metal2 s 24766 9840 24822 10300 0 FreeSans 224 90 0 0 S2MID[2]
port 106 nsew signal input
flabel metal2 s 25134 9840 25190 10300 0 FreeSans 224 90 0 0 S2MID[3]
port 107 nsew signal input
flabel metal2 s 25502 9840 25558 10300 0 FreeSans 224 90 0 0 S2MID[4]
port 108 nsew signal input
flabel metal2 s 25870 9840 25926 10300 0 FreeSans 224 90 0 0 S2MID[5]
port 109 nsew signal input
flabel metal2 s 26238 9840 26294 10300 0 FreeSans 224 90 0 0 S2MID[6]
port 110 nsew signal input
flabel metal2 s 26606 9840 26662 10300 0 FreeSans 224 90 0 0 S2MID[7]
port 111 nsew signal input
flabel metal2 s 26974 9840 27030 10300 0 FreeSans 224 90 0 0 S4END[0]
port 112 nsew signal input
flabel metal2 s 30654 9840 30710 10300 0 FreeSans 224 90 0 0 S4END[10]
port 113 nsew signal input
flabel metal2 s 31022 9840 31078 10300 0 FreeSans 224 90 0 0 S4END[11]
port 114 nsew signal input
flabel metal2 s 31390 9840 31446 10300 0 FreeSans 224 90 0 0 S4END[12]
port 115 nsew signal input
flabel metal2 s 31758 9840 31814 10300 0 FreeSans 224 90 0 0 S4END[13]
port 116 nsew signal input
flabel metal2 s 32126 9840 32182 10300 0 FreeSans 224 90 0 0 S4END[14]
port 117 nsew signal input
flabel metal2 s 32494 9840 32550 10300 0 FreeSans 224 90 0 0 S4END[15]
port 118 nsew signal input
flabel metal2 s 27342 9840 27398 10300 0 FreeSans 224 90 0 0 S4END[1]
port 119 nsew signal input
flabel metal2 s 27710 9840 27766 10300 0 FreeSans 224 90 0 0 S4END[2]
port 120 nsew signal input
flabel metal2 s 28078 9840 28134 10300 0 FreeSans 224 90 0 0 S4END[3]
port 121 nsew signal input
flabel metal2 s 28446 9840 28502 10300 0 FreeSans 224 90 0 0 S4END[4]
port 122 nsew signal input
flabel metal2 s 28814 9840 28870 10300 0 FreeSans 224 90 0 0 S4END[5]
port 123 nsew signal input
flabel metal2 s 29182 9840 29238 10300 0 FreeSans 224 90 0 0 S4END[6]
port 124 nsew signal input
flabel metal2 s 29550 9840 29606 10300 0 FreeSans 224 90 0 0 S4END[7]
port 125 nsew signal input
flabel metal2 s 29918 9840 29974 10300 0 FreeSans 224 90 0 0 S4END[8]
port 126 nsew signal input
flabel metal2 s 30286 9840 30342 10300 0 FreeSans 224 90 0 0 S4END[9]
port 127 nsew signal input
flabel metal2 s 32862 9840 32918 10300 0 FreeSans 224 90 0 0 SS4END[0]
port 128 nsew signal input
flabel metal2 s 36542 9840 36598 10300 0 FreeSans 224 90 0 0 SS4END[10]
port 129 nsew signal input
flabel metal2 s 36910 9840 36966 10300 0 FreeSans 224 90 0 0 SS4END[11]
port 130 nsew signal input
flabel metal2 s 37278 9840 37334 10300 0 FreeSans 224 90 0 0 SS4END[12]
port 131 nsew signal input
flabel metal2 s 37646 9840 37702 10300 0 FreeSans 224 90 0 0 SS4END[13]
port 132 nsew signal input
flabel metal2 s 38014 9840 38070 10300 0 FreeSans 224 90 0 0 SS4END[14]
port 133 nsew signal input
flabel metal2 s 38382 9840 38438 10300 0 FreeSans 224 90 0 0 SS4END[15]
port 134 nsew signal input
flabel metal2 s 33230 9840 33286 10300 0 FreeSans 224 90 0 0 SS4END[1]
port 135 nsew signal input
flabel metal2 s 33598 9840 33654 10300 0 FreeSans 224 90 0 0 SS4END[2]
port 136 nsew signal input
flabel metal2 s 33966 9840 34022 10300 0 FreeSans 224 90 0 0 SS4END[3]
port 137 nsew signal input
flabel metal2 s 34334 9840 34390 10300 0 FreeSans 224 90 0 0 SS4END[4]
port 138 nsew signal input
flabel metal2 s 34702 9840 34758 10300 0 FreeSans 224 90 0 0 SS4END[5]
port 139 nsew signal input
flabel metal2 s 35070 9840 35126 10300 0 FreeSans 224 90 0 0 SS4END[6]
port 140 nsew signal input
flabel metal2 s 35438 9840 35494 10300 0 FreeSans 224 90 0 0 SS4END[7]
port 141 nsew signal input
flabel metal2 s 35806 9840 35862 10300 0 FreeSans 224 90 0 0 SS4END[8]
port 142 nsew signal input
flabel metal2 s 36174 9840 36230 10300 0 FreeSans 224 90 0 0 SS4END[9]
port 143 nsew signal input
flabel metal2 s 1214 -300 1270 160 0 FreeSans 224 90 0 0 UserCLK
port 144 nsew signal input
flabel metal2 s 38750 9840 38806 10300 0 FreeSans 224 90 0 0 UserCLKo
port 145 nsew signal tristate
flabel metal4 s 6498 1040 6818 8752 0 FreeSans 1920 90 0 0 vccd1
port 146 nsew power bidirectional
flabel metal4 s 17606 1040 17926 8752 0 FreeSans 1920 90 0 0 vccd1
port 146 nsew power bidirectional
flabel metal4 s 28714 1040 29034 8752 0 FreeSans 1920 90 0 0 vccd1
port 146 nsew power bidirectional
flabel metal4 s 39822 1040 40142 8752 0 FreeSans 1920 90 0 0 vccd1
port 146 nsew power bidirectional
flabel metal4 s 12052 1040 12372 8752 0 FreeSans 1920 90 0 0 vssd1
port 147 nsew ground bidirectional
flabel metal4 s 23160 1040 23480 8752 0 FreeSans 1920 90 0 0 vssd1
port 147 nsew ground bidirectional
flabel metal4 s 34268 1040 34588 8752 0 FreeSans 1920 90 0 0 vssd1
port 147 nsew ground bidirectional
flabel metal4 s 45376 1040 45696 8752 0 FreeSans 1920 90 0 0 vssd1
port 147 nsew ground bidirectional
rlabel metal1 23322 8160 23322 8160 0 vccd1
rlabel via1 23400 8704 23400 8704 0 vssd1
rlabel metal2 3641 68 3641 68 0 FrameStrobe[0]
rlabel metal2 25675 68 25675 68 0 FrameStrobe[10]
rlabel metal2 27883 68 27883 68 0 FrameStrobe[11]
rlabel metal2 30091 68 30091 68 0 FrameStrobe[12]
rlabel metal2 32299 68 32299 68 0 FrameStrobe[13]
rlabel metal2 34507 68 34507 68 0 FrameStrobe[14]
rlabel metal2 36715 68 36715 68 0 FrameStrobe[15]
rlabel metal2 38923 68 38923 68 0 FrameStrobe[16]
rlabel metal2 41131 68 41131 68 0 FrameStrobe[17]
rlabel metal2 43339 68 43339 68 0 FrameStrobe[18]
rlabel metal2 45303 68 45303 68 0 FrameStrobe[19]
rlabel metal2 5711 68 5711 68 0 FrameStrobe[1]
rlabel metal2 7919 68 7919 68 0 FrameStrobe[2]
rlabel metal2 10127 68 10127 68 0 FrameStrobe[3]
rlabel metal2 12137 68 12137 68 0 FrameStrobe[4]
rlabel metal2 14635 68 14635 68 0 FrameStrobe[5]
rlabel metal2 16843 68 16843 68 0 FrameStrobe[6]
rlabel metal2 19143 68 19143 68 0 FrameStrobe[7]
rlabel metal2 21259 68 21259 68 0 FrameStrobe[8]
rlabel metal2 23322 143 23322 143 0 FrameStrobe[9]
rlabel metal1 39376 8602 39376 8602 0 FrameStrobe_O[0]
rlabel metal2 42826 8952 42826 8952 0 FrameStrobe_O[10]
rlabel metal2 43194 8680 43194 8680 0 FrameStrobe_O[11]
rlabel metal2 43562 8952 43562 8952 0 FrameStrobe_O[12]
rlabel metal2 43930 8952 43930 8952 0 FrameStrobe_O[13]
rlabel metal1 43608 7990 43608 7990 0 FrameStrobe_O[14]
rlabel metal1 44804 6426 44804 6426 0 FrameStrobe_O[15]
rlabel metal1 44896 7514 44896 7514 0 FrameStrobe_O[16]
rlabel metal1 45034 6834 45034 6834 0 FrameStrobe_O[17]
rlabel metal1 45034 7446 45034 7446 0 FrameStrobe_O[18]
rlabel metal1 45218 6766 45218 6766 0 FrameStrobe_O[19]
rlabel metal2 39514 9836 39514 9836 0 FrameStrobe_O[1]
rlabel metal2 39882 9190 39882 9190 0 FrameStrobe_O[2]
rlabel metal1 40710 8330 40710 8330 0 FrameStrobe_O[3]
rlabel metal1 40894 8058 40894 8058 0 FrameStrobe_O[4]
rlabel metal2 40986 9224 40986 9224 0 FrameStrobe_O[5]
rlabel metal1 42642 8568 42642 8568 0 FrameStrobe_O[6]
rlabel metal2 41722 9088 41722 9088 0 FrameStrobe_O[7]
rlabel metal2 42090 9122 42090 9122 0 FrameStrobe_O[8]
rlabel metal2 42458 9785 42458 9785 0 FrameStrobe_O[9]
rlabel metal1 23598 2074 23598 2074 0 FrameStrobe_O_i\[0\]
rlabel metal2 26910 2244 26910 2244 0 FrameStrobe_O_i\[10\]
rlabel metal1 28704 2074 28704 2074 0 FrameStrobe_O_i\[11\]
rlabel metal1 30912 2074 30912 2074 0 FrameStrobe_O_i\[12\]
rlabel metal1 33120 2074 33120 2074 0 FrameStrobe_O_i\[13\]
rlabel metal1 35328 2074 35328 2074 0 FrameStrobe_O_i\[14\]
rlabel metal1 37628 2074 37628 2074 0 FrameStrobe_O_i\[15\]
rlabel metal2 43470 2210 43470 2210 0 FrameStrobe_O_i\[16\]
rlabel metal2 41630 2278 41630 2278 0 FrameStrobe_O_i\[17\]
rlabel metal1 43930 2040 43930 2040 0 FrameStrobe_O_i\[18\]
rlabel metal1 44252 2074 44252 2074 0 FrameStrobe_O_i\[19\]
rlabel metal1 22264 1802 22264 1802 0 FrameStrobe_O_i\[1\]
rlabel metal1 22586 2040 22586 2040 0 FrameStrobe_O_i\[2\]
rlabel metal1 23092 2074 23092 2074 0 FrameStrobe_O_i\[3\]
rlabel metal2 22310 2278 22310 2278 0 FrameStrobe_O_i\[4\]
rlabel metal1 22494 1530 22494 1530 0 FrameStrobe_O_i\[5\]
rlabel metal1 21712 2074 21712 2074 0 FrameStrobe_O_i\[6\]
rlabel metal1 19918 2074 19918 2074 0 FrameStrobe_O_i\[7\]
rlabel metal2 21482 2040 21482 2040 0 FrameStrobe_O_i\[8\]
rlabel metal1 24288 2074 24288 2074 0 FrameStrobe_O_i\[9\]
rlabel metal2 506 9785 506 9785 0 N1BEG[0]
rlabel metal2 874 8680 874 8680 0 N1BEG[1]
rlabel metal1 1518 6834 1518 6834 0 N1BEG[2]
rlabel metal2 1610 8646 1610 8646 0 N1BEG[3]
rlabel metal2 1978 9309 1978 9309 0 N2BEG[0]
rlabel metal1 2254 8602 2254 8602 0 N2BEG[1]
rlabel metal2 2714 9037 2714 9037 0 N2BEG[2]
rlabel metal1 3128 8058 3128 8058 0 N2BEG[3]
rlabel metal1 3496 8058 3496 8058 0 N2BEG[4]
rlabel metal2 3818 9785 3818 9785 0 N2BEG[5]
rlabel metal1 3864 8602 3864 8602 0 N2BEG[6]
rlabel metal1 4600 8058 4600 8058 0 N2BEG[7]
rlabel metal1 4738 8602 4738 8602 0 N2BEGb[0]
rlabel metal1 5152 8602 5152 8602 0 N2BEGb[1]
rlabel metal1 5612 8602 5612 8602 0 N2BEGb[2]
rlabel metal1 6302 8602 6302 8602 0 N2BEGb[3]
rlabel metal2 6394 8952 6394 8952 0 N2BEGb[4]
rlabel metal1 6486 8534 6486 8534 0 N2BEGb[5]
rlabel metal2 7130 9224 7130 9224 0 N2BEGb[6]
rlabel metal1 7544 8058 7544 8058 0 N2BEGb[7]
rlabel metal1 7820 8602 7820 8602 0 N4BEG[0]
rlabel metal2 11546 9309 11546 9309 0 N4BEG[10]
rlabel metal1 12052 8058 12052 8058 0 N4BEG[11]
rlabel metal2 12006 9231 12006 9231 0 N4BEG[12]
rlabel metal2 12650 9224 12650 9224 0 N4BEG[13]
rlabel metal1 13064 8058 13064 8058 0 N4BEG[14]
rlabel metal1 13340 8602 13340 8602 0 N4BEG[15]
rlabel metal2 8234 9224 8234 9224 0 N4BEG[1]
rlabel metal1 8648 8602 8648 8602 0 N4BEG[2]
rlabel metal2 8970 9836 8970 9836 0 N4BEG[3]
rlabel metal1 9292 8602 9292 8602 0 N4BEG[4]
rlabel metal2 9706 9224 9706 9224 0 N4BEG[5]
rlabel metal1 10120 8058 10120 8058 0 N4BEG[6]
rlabel metal1 10396 8602 10396 8602 0 N4BEG[7]
rlabel metal1 10764 8602 10764 8602 0 N4BEG[8]
rlabel metal2 11178 9224 11178 9224 0 N4BEG[9]
rlabel metal2 13754 9224 13754 9224 0 NN4BEG[0]
rlabel metal1 17480 8602 17480 8602 0 NN4BEG[10]
rlabel metal2 17802 9836 17802 9836 0 NN4BEG[11]
rlabel metal1 18308 8602 18308 8602 0 NN4BEG[12]
rlabel metal1 18676 8602 18676 8602 0 NN4BEG[13]
rlabel metal2 18906 9836 18906 9836 0 NN4BEG[14]
rlabel metal2 19274 8952 19274 8952 0 NN4BEG[15]
rlabel metal2 14122 9836 14122 9836 0 NN4BEG[1]
rlabel metal1 14444 8602 14444 8602 0 NN4BEG[2]
rlabel metal1 14812 8602 14812 8602 0 NN4BEG[3]
rlabel metal2 15226 9224 15226 9224 0 NN4BEG[4]
rlabel metal1 15640 8602 15640 8602 0 NN4BEG[5]
rlabel metal1 16008 8602 16008 8602 0 NN4BEG[6]
rlabel metal1 16376 8602 16376 8602 0 NN4BEG[7]
rlabel metal2 16698 9836 16698 9836 0 NN4BEG[8]
rlabel metal1 17204 8058 17204 8058 0 NN4BEG[9]
rlabel metal2 19642 9241 19642 9241 0 S1END[0]
rlabel metal2 20010 9785 20010 9785 0 S1END[1]
rlabel metal2 20378 9836 20378 9836 0 S1END[2]
rlabel metal2 20746 9156 20746 9156 0 S1END[3]
rlabel metal2 21114 9156 21114 9156 0 S2END[0]
rlabel metal2 21482 9156 21482 9156 0 S2END[1]
rlabel metal2 21850 9836 21850 9836 0 S2END[2]
rlabel metal2 21942 9163 21942 9163 0 S2END[3]
rlabel metal2 22586 9836 22586 9836 0 S2END[4]
rlabel metal2 22954 9836 22954 9836 0 S2END[5]
rlabel metal2 23322 9836 23322 9836 0 S2END[6]
rlabel metal2 23690 9581 23690 9581 0 S2END[7]
rlabel metal2 24058 9836 24058 9836 0 S2MID[0]
rlabel metal2 24426 9836 24426 9836 0 S2MID[1]
rlabel metal2 24794 9513 24794 9513 0 S2MID[2]
rlabel metal2 25162 9836 25162 9836 0 S2MID[3]
rlabel metal2 25530 9836 25530 9836 0 S2MID[4]
rlabel metal2 25898 9836 25898 9836 0 S2MID[5]
rlabel metal2 26266 9836 26266 9836 0 S2MID[6]
rlabel metal2 26634 9156 26634 9156 0 S2MID[7]
rlabel metal2 27002 9190 27002 9190 0 S4END[0]
rlabel metal2 30682 9836 30682 9836 0 S4END[10]
rlabel metal2 31050 9836 31050 9836 0 S4END[11]
rlabel metal2 31418 9836 31418 9836 0 S4END[12]
rlabel metal2 31786 9156 31786 9156 0 S4END[13]
rlabel metal2 32154 9156 32154 9156 0 S4END[14]
rlabel metal2 32522 9836 32522 9836 0 S4END[15]
rlabel metal2 27370 9836 27370 9836 0 S4END[1]
rlabel metal2 27738 9836 27738 9836 0 S4END[2]
rlabel metal2 28106 9836 28106 9836 0 S4END[3]
rlabel metal2 28474 9836 28474 9836 0 S4END[4]
rlabel metal2 28842 9156 28842 9156 0 S4END[5]
rlabel metal2 29210 9156 29210 9156 0 S4END[6]
rlabel metal2 29578 9190 29578 9190 0 S4END[7]
rlabel metal2 29946 9836 29946 9836 0 S4END[8]
rlabel metal2 30314 9224 30314 9224 0 S4END[9]
rlabel metal2 32890 9836 32890 9836 0 SS4END[0]
rlabel metal2 36570 9156 36570 9156 0 SS4END[10]
rlabel metal2 36938 9156 36938 9156 0 SS4END[11]
rlabel metal2 37306 9836 37306 9836 0 SS4END[12]
rlabel metal2 37674 9836 37674 9836 0 SS4END[13]
rlabel metal2 38042 9156 38042 9156 0 SS4END[14]
rlabel metal2 38410 9156 38410 9156 0 SS4END[15]
rlabel metal2 33258 9156 33258 9156 0 SS4END[1]
rlabel metal2 33626 9156 33626 9156 0 SS4END[2]
rlabel metal2 33994 9156 33994 9156 0 SS4END[3]
rlabel metal2 34362 9836 34362 9836 0 SS4END[4]
rlabel metal2 34730 9836 34730 9836 0 SS4END[5]
rlabel metal2 35098 9836 35098 9836 0 SS4END[6]
rlabel metal2 35466 9156 35466 9156 0 SS4END[7]
rlabel metal2 35834 9156 35834 9156 0 SS4END[8]
rlabel metal2 36202 9156 36202 9156 0 SS4END[9]
rlabel metal2 1242 704 1242 704 0 UserCLK
rlabel metal2 38778 9836 38778 9836 0 UserCLKo
rlabel metal2 4002 1088 4002 1088 0 net1
rlabel metal1 43700 1530 43700 1530 0 net10
rlabel metal2 2530 7072 2530 7072 0 net100
rlabel metal2 2990 7038 2990 7038 0 net101
rlabel metal2 3358 7242 3358 7242 0 net102
rlabel metal2 3910 7650 3910 7650 0 net103
rlabel metal1 3266 8908 3266 8908 0 net104
rlabel metal1 4462 7242 4462 7242 0 net105
rlabel metal1 4738 8500 4738 8500 0 net106
rlabel metal2 4830 8840 4830 8840 0 net107
rlabel metal1 5382 9826 5382 9826 0 net108
rlabel metal2 7406 8976 7406 8976 0 net109
rlabel metal1 44804 1530 44804 1530 0 net11
rlabel metal1 6394 7276 6394 7276 0 net110
rlabel metal2 5842 9078 5842 9078 0 net111
rlabel metal1 8878 9316 8878 9316 0 net112
rlabel metal2 19366 7854 19366 7854 0 net113
rlabel metal2 7590 9078 7590 9078 0 net114
rlabel metal2 28474 7361 28474 7361 0 net115
rlabel metal1 12006 7820 12006 7820 0 net116
rlabel metal1 11822 8840 11822 8840 0 net117
rlabel metal1 26266 8058 26266 8058 0 net118
rlabel metal1 21574 7276 21574 7276 0 net119
rlabel metal1 19550 1292 19550 1292 0 net12
rlabel metal1 13110 9316 13110 9316 0 net120
rlabel metal2 8050 9112 8050 9112 0 net121
rlabel metal1 8510 8874 8510 8874 0 net122
rlabel metal1 9062 7752 9062 7752 0 net123
rlabel metal2 9062 8840 9062 8840 0 net124
rlabel metal2 9522 9146 9522 9146 0 net125
rlabel metal2 9982 7412 9982 7412 0 net126
rlabel metal1 24656 7990 24656 7990 0 net127
rlabel metal2 10534 8772 10534 8772 0 net128
rlabel metal1 10994 8466 10994 8466 0 net129
rlabel metal2 21574 1190 21574 1190 0 net13
rlabel metal2 17802 8942 17802 8942 0 net130
rlabel metal1 17526 7752 17526 7752 0 net131
rlabel metal1 17664 8058 17664 8058 0 net132
rlabel metal1 18170 8058 18170 8058 0 net133
rlabel metal2 18906 7990 18906 7990 0 net134
rlabel metal1 19228 7514 19228 7514 0 net135
rlabel metal1 19044 7786 19044 7786 0 net136
rlabel metal2 14214 7378 14214 7378 0 net137
rlabel metal2 21666 7106 21666 7106 0 net138
rlabel metal1 19918 8466 19918 8466 0 net139
rlabel metal2 23046 1360 23046 1360 0 net14
rlabel metal2 21850 7616 21850 7616 0 net140
rlabel metal2 22034 7497 22034 7497 0 net141
rlabel metal2 20838 7905 20838 7905 0 net142
rlabel metal2 21574 8194 21574 8194 0 net143
rlabel metal2 20470 8466 20470 8466 0 net144
rlabel metal1 17342 7514 17342 7514 0 net145
rlabel metal1 20470 2006 20470 2006 0 net146
rlabel metal2 20838 1428 20838 1428 0 net15
rlabel metal1 22310 952 22310 952 0 net16
rlabel metal1 18768 1190 18768 1190 0 net17
rlabel metal1 19458 1530 19458 1530 0 net18
rlabel metal1 21436 1530 21436 1530 0 net19
rlabel metal2 26266 1564 26266 1564 0 net2
rlabel metal1 23736 1530 23736 1530 0 net20
rlabel metal1 18630 7412 18630 7412 0 net21
rlabel metal1 18354 7888 18354 7888 0 net22
rlabel metal1 19274 7854 19274 7854 0 net23
rlabel metal1 19918 7888 19918 7888 0 net24
rlabel metal1 20378 7854 20378 7854 0 net25
rlabel metal1 20746 7888 20746 7888 0 net26
rlabel metal1 21022 7820 21022 7820 0 net27
rlabel metal1 21298 7888 21298 7888 0 net28
rlabel metal2 21942 7854 21942 7854 0 net29
rlabel metal1 28152 1530 28152 1530 0 net3
rlabel metal1 22310 7378 22310 7378 0 net30
rlabel metal1 22678 8500 22678 8500 0 net31
rlabel metal2 23046 7888 23046 7888 0 net32
rlabel metal1 22954 7888 22954 7888 0 net33
rlabel metal1 23782 7412 23782 7412 0 net34
rlabel metal1 24196 7854 24196 7854 0 net35
rlabel metal1 25070 7854 25070 7854 0 net36
rlabel metal1 25346 7854 25346 7854 0 net37
rlabel metal1 25622 7854 25622 7854 0 net38
rlabel metal1 25852 7854 25852 7854 0 net39
rlabel metal1 30360 1190 30360 1190 0 net4
rlabel metal1 26128 7854 26128 7854 0 net40
rlabel metal1 26496 7854 26496 7854 0 net41
rlabel metal1 27416 7378 27416 7378 0 net42
rlabel metal1 23782 7820 23782 7820 0 net43
rlabel metal1 23598 7854 23598 7854 0 net44
rlabel metal2 32338 9146 32338 9146 0 net45
rlabel metal2 32430 8704 32430 8704 0 net46
rlabel metal2 23506 8483 23506 8483 0 net47
rlabel metal1 26726 7922 26726 7922 0 net48
rlabel metal1 27094 7888 27094 7888 0 net49
rlabel metal1 32568 1530 32568 1530 0 net5
rlabel metal1 27554 7854 27554 7854 0 net50
rlabel metal1 28014 7922 28014 7922 0 net51
rlabel metal1 28290 7888 28290 7888 0 net52
rlabel metal1 29072 7854 29072 7854 0 net53
rlabel metal1 27738 7820 27738 7820 0 net54
rlabel metal1 24702 7820 24702 7820 0 net55
rlabel metal1 24426 7786 24426 7786 0 net56
rlabel metal2 18814 8041 18814 8041 0 net57
rlabel metal1 36846 8398 36846 8398 0 net58
rlabel metal2 22034 7905 22034 7905 0 net59
rlabel metal1 34914 1530 34914 1530 0 net6
rlabel metal2 37766 7752 37766 7752 0 net60
rlabel metal2 27278 7922 27278 7922 0 net61
rlabel metal2 35926 8007 35926 8007 0 net62
rlabel metal2 38686 9044 38686 9044 0 net63
rlabel metal2 33534 8976 33534 8976 0 net64
rlabel metal2 19090 8092 19090 8092 0 net65
rlabel metal2 18354 8500 18354 8500 0 net66
rlabel metal2 18446 8874 18446 8874 0 net67
rlabel metal2 17710 9044 17710 9044 0 net68
rlabel metal1 35144 8602 35144 8602 0 net69
rlabel metal1 37076 1190 37076 1190 0 net7
rlabel metal2 20654 9163 20654 9163 0 net70
rlabel metal2 21758 7565 21758 7565 0 net71
rlabel metal1 36478 8432 36478 8432 0 net72
rlabel metal2 1610 1734 1610 1734 0 net73
rlabel metal2 37214 5882 37214 5882 0 net74
rlabel metal1 43010 7786 43010 7786 0 net75
rlabel metal2 43378 6086 43378 6086 0 net76
rlabel metal2 43378 7548 43378 7548 0 net77
rlabel metal1 44298 2584 44298 2584 0 net78
rlabel metal1 37812 2550 37812 2550 0 net79
rlabel metal2 43654 1598 43654 1598 0 net8
rlabel metal1 44850 2346 44850 2346 0 net80
rlabel metal1 44344 7378 44344 7378 0 net81
rlabel metal2 44482 4658 44482 4658 0 net82
rlabel metal1 44482 7310 44482 7310 0 net83
rlabel metal2 43930 4658 43930 4658 0 net84
rlabel metal1 23000 2278 23000 2278 0 net85
rlabel metal2 36018 7548 36018 7548 0 net86
rlabel metal2 33902 6290 33902 6290 0 net87
rlabel metal1 23230 2618 23230 2618 0 net88
rlabel metal1 22908 1734 22908 1734 0 net89
rlabel metal2 41814 1564 41814 1564 0 net9
rlabel metal1 22678 2618 22678 2618 0 net90
rlabel metal1 20516 2618 20516 2618 0 net91
rlabel metal2 43654 8840 43654 8840 0 net92
rlabel metal1 43746 8534 43746 8534 0 net93
rlabel metal1 2714 8432 2714 8432 0 net94
rlabel metal1 11730 7412 11730 7412 0 net95
rlabel metal1 1518 6358 1518 6358 0 net96
rlabel metal1 11638 7480 11638 7480 0 net97
rlabel metal1 3726 7718 3726 7718 0 net98
rlabel metal1 2346 8398 2346 8398 0 net99
<< properties >>
string FIXED_BBOX 0 0 46700 10000
<< end >>
