* NGSPICE file created from S_term_RAM_IO.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_ef_sc_hd__decap_12 abstract view
.subckt sky130_ef_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_1 abstract view
.subckt sky130_fd_sc_hd__buf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_4 abstract view
.subckt sky130_fd_sc_hd__clkbuf_4 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

.subckt S_term_RAM_IO FrameStrobe[0] FrameStrobe[10] FrameStrobe[11] FrameStrobe[12]
+ FrameStrobe[13] FrameStrobe[14] FrameStrobe[15] FrameStrobe[16] FrameStrobe[17]
+ FrameStrobe[18] FrameStrobe[19] FrameStrobe[1] FrameStrobe[2] FrameStrobe[3] FrameStrobe[4]
+ FrameStrobe[5] FrameStrobe[6] FrameStrobe[7] FrameStrobe[8] FrameStrobe[9] FrameStrobe_O[0]
+ FrameStrobe_O[10] FrameStrobe_O[11] FrameStrobe_O[12] FrameStrobe_O[13] FrameStrobe_O[14]
+ FrameStrobe_O[15] FrameStrobe_O[16] FrameStrobe_O[17] FrameStrobe_O[18] FrameStrobe_O[19]
+ FrameStrobe_O[1] FrameStrobe_O[2] FrameStrobe_O[3] FrameStrobe_O[4] FrameStrobe_O[5]
+ FrameStrobe_O[6] FrameStrobe_O[7] FrameStrobe_O[8] FrameStrobe_O[9] N1BEG[0] N1BEG[1]
+ N1BEG[2] N1BEG[3] N2BEG[0] N2BEG[1] N2BEG[2] N2BEG[3] N2BEG[4] N2BEG[5] N2BEG[6]
+ N2BEG[7] N2BEGb[0] N2BEGb[1] N2BEGb[2] N2BEGb[3] N2BEGb[4] N2BEGb[5] N2BEGb[6] N2BEGb[7]
+ N4BEG[0] N4BEG[10] N4BEG[11] N4BEG[12] N4BEG[13] N4BEG[14] N4BEG[15] N4BEG[1] N4BEG[2]
+ N4BEG[3] N4BEG[4] N4BEG[5] N4BEG[6] N4BEG[7] N4BEG[8] N4BEG[9] S1END[0] S1END[1]
+ S1END[2] S1END[3] S2END[0] S2END[1] S2END[2] S2END[3] S2END[4] S2END[5] S2END[6]
+ S2END[7] S2MID[0] S2MID[1] S2MID[2] S2MID[3] S2MID[4] S2MID[5] S2MID[6] S2MID[7]
+ S4END[0] S4END[10] S4END[11] S4END[12] S4END[13] S4END[14] S4END[15] S4END[1] S4END[2]
+ S4END[3] S4END[4] S4END[5] S4END[6] S4END[7] S4END[8] S4END[9] UserCLK UserCLKo
+ VGND VPWR
XFILLER_0_4_193 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_130 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_S_term_RAM_IO_switch_matrix__22_ net52 VGND VGND VPWR VPWR net99 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_6_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_S_term_RAM_IO_switch_matrix__05_ net39 VGND VGND VPWR VPWR net83 sky130_fd_sc_hd__buf_1
XFILLER_0_10_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_3_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_228 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput97 net97 VGND VGND VPWR VPWR N2BEGb[7] sky130_fd_sc_hd__clkbuf_4
Xoutput75 net75 VGND VGND VPWR VPWR FrameStrobe_O[7] sky130_fd_sc_hd__clkbuf_4
Xoutput86 net86 VGND VGND VPWR VPWR N2BEG[4] sky130_fd_sc_hd__clkbuf_4
Xoutput64 net64 VGND VGND VPWR VPWR FrameStrobe_O[15] sky130_fd_sc_hd__clkbuf_4
Xstrobe_outbuf_14__0_ FrameStrobe_O_i\[14\] VGND VGND VPWR VPWR net63 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_S_term_RAM_IO_switch_matrix__21_ net46 VGND VGND VPWR VPWR net105 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_6_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XInst_S_term_RAM_IO_switch_matrix__04_ net40 VGND VGND VPWR VPWR net82 sky130_fd_sc_hd__buf_1
Xstrobe_inbuf_11__0_ net3 VGND VGND VPWR VPWR FrameStrobe_O_i\[11\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xstrobe_outbuf_9__0_ FrameStrobe_O_i\[9\] VGND VGND VPWR VPWR net77 sky130_fd_sc_hd__buf_1
XFILLER_0_1_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_6_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput76 net76 VGND VGND VPWR VPWR FrameStrobe_O[8] sky130_fd_sc_hd__clkbuf_4
Xoutput98 net98 VGND VGND VPWR VPWR N4BEG[0] sky130_fd_sc_hd__clkbuf_4
Xoutput87 net87 VGND VGND VPWR VPWR N2BEG[5] sky130_fd_sc_hd__clkbuf_4
Xoutput65 net65 VGND VGND VPWR VPWR FrameStrobe_O[16] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_7_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_64 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_S_term_RAM_IO_switch_matrix__20_ net47 VGND VGND VPWR VPWR net98 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_S_term_RAM_IO_switch_matrix__03_ net21 VGND VGND VPWR VPWR net81 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_238 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xoutput99 net99 VGND VGND VPWR VPWR N4BEG[10] sky130_fd_sc_hd__clkbuf_4
Xoutput88 net88 VGND VGND VPWR VPWR N2BEG[6] sky130_fd_sc_hd__clkbuf_4
Xoutput77 net77 VGND VGND VPWR VPWR FrameStrobe_O[9] sky130_fd_sc_hd__clkbuf_4
Xoutput66 net66 VGND VGND VPWR VPWR FrameStrobe_O[17] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_7_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_185 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_7_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_1_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_144 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_S_term_RAM_IO_switch_matrix__02_ net22 VGND VGND VPWR VPWR net80 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xstrobe_inbuf_2__0_ net13 VGND VGND VPWR VPWR FrameStrobe_O_i\[2\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_209 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_12_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_12_145 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_134 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xstrobe_outbuf_17__0_ FrameStrobe_O_i\[17\] VGND VGND VPWR VPWR net66 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput78 net78 VGND VGND VPWR VPWR N1BEG[0] sky130_fd_sc_hd__clkbuf_4
Xoutput89 net89 VGND VGND VPWR VPWR N2BEG[7] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_7_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput67 net67 VGND VGND VPWR VPWR FrameStrobe_O[18] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_4_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_156 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xstrobe_inbuf_14__0_ net6 VGND VGND VPWR VPWR FrameStrobe_O_i\[14\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_S_term_RAM_IO_switch_matrix__01_ net23 VGND VGND VPWR VPWR net79 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_87 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_179 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput79 net79 VGND VGND VPWR VPWR N1BEG[1] sky130_fd_sc_hd__clkbuf_4
Xoutput68 net68 VGND VGND VPWR VPWR FrameStrobe_O[19] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_11_190 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_S_term_RAM_IO_switch_matrix__00_ net24 VGND VGND VPWR VPWR net78 sky130_fd_sc_hd__buf_1
XFILLER_0_10_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput69 net69 VGND VGND VPWR VPWR FrameStrobe_O[1] sky130_fd_sc_hd__clkbuf_4
Xoutput58 net58 VGND VGND VPWR VPWR FrameStrobe_O[0] sky130_fd_sc_hd__clkbuf_4
XPHY_0 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_4_177 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_4_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xstrobe_inbuf_5__0_ net16 VGND VGND VPWR VPWR FrameStrobe_O_i\[5\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput59 net59 VGND VGND VPWR VPWR FrameStrobe_O[10] sky130_fd_sc_hd__clkbuf_4
Xstrobe_outbuf_2__0_ FrameStrobe_O_i\[2\] VGND VGND VPWR VPWR net70 sky130_fd_sc_hd__buf_1
XPHY_1 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_126 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xstrobe_inbuf_17__0_ net9 VGND VGND VPWR VPWR FrameStrobe_O_i\[17\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_116 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_2 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_13_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_160 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_2_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_9 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xstrobe_outbuf_10__0_ FrameStrobe_O_i\[10\] VGND VGND VPWR VPWR net59 sky130_fd_sc_hd__buf_1
XFILLER_0_0_183 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_172 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_10_237 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xstrobe_inbuf_8__0_ net19 VGND VGND VPWR VPWR FrameStrobe_O_i\[8\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_5_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_1_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_60 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xstrobe_outbuf_5__0_ FrameStrobe_O_i\[5\] VGND VGND VPWR VPWR net73 sky130_fd_sc_hd__buf_1
XFILLER_0_7_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_4 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_50 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_5 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_119 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_4_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_84 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_1_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_6 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xstrobe_outbuf_13__0_ FrameStrobe_O_i\[13\] VGND VGND VPWR VPWR net62 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_153 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_197 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xstrobe_inbuf_10__0_ net2 VGND VGND VPWR VPWR FrameStrobe_O_i\[10\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_5_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_96 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_11_74 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XTAP_90 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xstrobe_outbuf_8__0_ FrameStrobe_O_i\[8\] VGND VGND VPWR VPWR net76 sky130_fd_sc_hd__buf_1
Xinput1 FrameStrobe[0] VGND VGND VPWR VPWR net1 sky130_fd_sc_hd__buf_1
XInst_S_term_RAM_IO_switch_matrix__19_ net25 VGND VGND VPWR VPWR net97 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_7_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_7_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_13_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_121 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_S_term_RAM_IO_switch_matrix__35_ net53 VGND VGND VPWR VPWR net113 sky130_fd_sc_hd__clkbuf_1
XTAP_91 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_80 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput2 FrameStrobe[10] VGND VGND VPWR VPWR net2 sky130_fd_sc_hd__clkbuf_1
XInst_S_term_RAM_IO_switch_matrix__18_ net26 VGND VGND VPWR VPWR net96 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_7_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_8 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_0_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_233 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xstrobe_inbuf_1__0_ net12 VGND VGND VPWR VPWR FrameStrobe_O_i\[1\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_5_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XInst_S_term_RAM_IO_switch_matrix__34_ net54 VGND VGND VPWR VPWR net112 sky130_fd_sc_hd__buf_1
XTAP_81 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_70 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput3 FrameStrobe[11] VGND VGND VPWR VPWR net3 sky130_fd_sc_hd__clkbuf_1
XInst_S_term_RAM_IO_switch_matrix__17_ net27 VGND VGND VPWR VPWR net95 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_178 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_101 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xstrobe_outbuf_16__0_ FrameStrobe_O_i\[16\] VGND VGND VPWR VPWR net65 sky130_fd_sc_hd__clkbuf_1
Xinst_clk_buf net57 VGND VGND VPWR VPWR net114 sky130_fd_sc_hd__buf_1
XFILLER_0_2_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_9 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xinput50 S4END[3] VGND VGND VPWR VPWR net50 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_245 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xstrobe_inbuf_13__0_ net5 VGND VGND VPWR VPWR FrameStrobe_O_i\[13\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_5_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_S_term_RAM_IO_switch_matrix__33_ net55 VGND VGND VPWR VPWR net111 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_82 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_11_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_71 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput4 FrameStrobe[12] VGND VGND VPWR VPWR net4 sky130_fd_sc_hd__clkbuf_1
XTAP_60 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_S_term_RAM_IO_switch_matrix__16_ net28 VGND VGND VPWR VPWR net94 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput51 S4END[4] VGND VGND VPWR VPWR net51 sky130_fd_sc_hd__clkbuf_1
Xinput40 S2MID[7] VGND VGND VPWR VPWR net40 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_113 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_1_230 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_S_term_RAM_IO_switch_matrix__32_ net56 VGND VGND VPWR VPWR net110 sky130_fd_sc_hd__buf_1
Xinput5 FrameStrobe[13] VGND VGND VPWR VPWR net5 sky130_fd_sc_hd__clkbuf_1
XTAP_83 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_72 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_50 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_61 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_S_term_RAM_IO_switch_matrix__15_ net29 VGND VGND VPWR VPWR net93 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_169 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_6_152 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput52 S4END[5] VGND VGND VPWR VPWR net52 sky130_fd_sc_hd__clkbuf_1
Xinput41 S4END[0] VGND VGND VPWR VPWR net41 sky130_fd_sc_hd__clkbuf_1
Xinput30 S2END[5] VGND VGND VPWR VPWR net30 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_147 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_0_125 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xstrobe_inbuf_4__0_ net15 VGND VGND VPWR VPWR FrameStrobe_O_i\[4\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_S_term_RAM_IO_switch_matrix__31_ net42 VGND VGND VPWR VPWR net109 sky130_fd_sc_hd__buf_1
XFILLER_0_11_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_84 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_73 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput6 FrameStrobe[14] VGND VGND VPWR VPWR net6 sky130_fd_sc_hd__clkbuf_1
XTAP_40 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xstrobe_outbuf_19__0_ FrameStrobe_O_i\[19\] VGND VGND VPWR VPWR net68 sky130_fd_sc_hd__clkbuf_1
XTAP_51 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_62 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_S_term_RAM_IO_switch_matrix__14_ net30 VGND VGND VPWR VPWR net92 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_9_161 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_164 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput31 S2END[6] VGND VGND VPWR VPWR net31 sky130_fd_sc_hd__clkbuf_1
Xstrobe_outbuf_1__0_ FrameStrobe_O_i\[1\] VGND VGND VPWR VPWR net69 sky130_fd_sc_hd__buf_1
Xinput20 FrameStrobe[9] VGND VGND VPWR VPWR net20 sky130_fd_sc_hd__clkbuf_1
Xinput42 S4END[10] VGND VGND VPWR VPWR net42 sky130_fd_sc_hd__clkbuf_1
Xinput53 S4END[6] VGND VGND VPWR VPWR net53 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xstrobe_inbuf_16__0_ net8 VGND VGND VPWR VPWR FrameStrobe_O_i\[16\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_8_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_S_term_RAM_IO_switch_matrix__30_ net43 VGND VGND VPWR VPWR net108 sky130_fd_sc_hd__buf_1
XFILLER_0_10_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_69 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_85 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_74 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_30 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput7 FrameStrobe[15] VGND VGND VPWR VPWR net7 sky130_fd_sc_hd__clkbuf_1
XTAP_41 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_52 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_63 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_S_term_RAM_IO_switch_matrix__13_ net31 VGND VGND VPWR VPWR net91 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_176 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput43 S4END[11] VGND VGND VPWR VPWR net43 sky130_fd_sc_hd__clkbuf_1
Xinput54 S4END[7] VGND VGND VPWR VPWR net54 sky130_fd_sc_hd__clkbuf_1
Xinput32 S2END[7] VGND VGND VPWR VPWR net32 sky130_fd_sc_hd__clkbuf_1
Xinput21 S1END[0] VGND VGND VPWR VPWR net21 sky130_fd_sc_hd__clkbuf_1
Xinput10 FrameStrobe[18] VGND VGND VPWR VPWR net10 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_138 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XTAP_86 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_75 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_31 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput8 FrameStrobe[16] VGND VGND VPWR VPWR net8 sky130_fd_sc_hd__clkbuf_1
XTAP_42 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_53 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_64 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_S_term_RAM_IO_switch_matrix__12_ net32 VGND VGND VPWR VPWR net90 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_10_172 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_6_188 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
Xinput44 S4END[12] VGND VGND VPWR VPWR net44 sky130_fd_sc_hd__buf_1
Xinput33 S2MID[0] VGND VGND VPWR VPWR net33 sky130_fd_sc_hd__clkbuf_1
Xinput55 S4END[8] VGND VGND VPWR VPWR net55 sky130_fd_sc_hd__clkbuf_1
Xinput22 S1END[1] VGND VGND VPWR VPWR net22 sky130_fd_sc_hd__clkbuf_1
Xinput11 FrameStrobe[19] VGND VGND VPWR VPWR net11 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xstrobe_inbuf_7__0_ net18 VGND VGND VPWR VPWR FrameStrobe_O_i\[7\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_87 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_76 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_32 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xinput9 FrameStrobe[17] VGND VGND VPWR VPWR net9 sky130_fd_sc_hd__clkbuf_1
XTAP_43 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_54 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_65 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_S_term_RAM_IO_switch_matrix__11_ net33 VGND VGND VPWR VPWR net89 sky130_fd_sc_hd__buf_1
Xoutput110 net110 VGND VGND VPWR VPWR N4BEG[6] sky130_fd_sc_hd__buf_2
XFILLER_0_12_70 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
Xstrobe_outbuf_4__0_ FrameStrobe_O_i\[4\] VGND VGND VPWR VPWR net72 sky130_fd_sc_hd__buf_1
XFILLER_0_10_184 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput34 S2MID[1] VGND VGND VPWR VPWR net34 sky130_fd_sc_hd__clkbuf_1
Xinput45 S4END[13] VGND VGND VPWR VPWR net45 sky130_fd_sc_hd__clkbuf_1
Xinput56 S4END[9] VGND VGND VPWR VPWR net56 sky130_fd_sc_hd__clkbuf_1
Xinput23 S1END[2] VGND VGND VPWR VPWR net23 sky130_fd_sc_hd__clkbuf_1
Xinput12 FrameStrobe[1] VGND VGND VPWR VPWR net12 sky130_fd_sc_hd__buf_1
Xstrobe_inbuf_19__0_ net11 VGND VGND VPWR VPWR FrameStrobe_O_i\[19\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_4_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_11_28 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_33 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_88 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_77 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_44 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_55 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_66 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XInst_S_term_RAM_IO_switch_matrix__10_ net34 VGND VGND VPWR VPWR net88 sky130_fd_sc_hd__buf_1
XFILLER_0_2_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput111 net111 VGND VGND VPWR VPWR N4BEG[7] sky130_fd_sc_hd__buf_2
Xoutput100 net100 VGND VGND VPWR VPWR N4BEG[11] sky130_fd_sc_hd__buf_2
XFILLER_0_10_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput35 S2MID[2] VGND VGND VPWR VPWR net35 sky130_fd_sc_hd__clkbuf_1
Xinput46 S4END[14] VGND VGND VPWR VPWR net46 sky130_fd_sc_hd__buf_1
Xinput24 S1END[3] VGND VGND VPWR VPWR net24 sky130_fd_sc_hd__clkbuf_1
Xinput13 FrameStrobe[2] VGND VGND VPWR VPWR net13 sky130_fd_sc_hd__clkbuf_1
Xinput57 UserCLK VGND VGND VPWR VPWR net57 sky130_fd_sc_hd__buf_1
XFILLER_0_3_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_3_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_92 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_4_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_8_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_7 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_5_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_89 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_78 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_34 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_45 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_56 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_67 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_11_109 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_2_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput101 net101 VGND VGND VPWR VPWR N4BEG[12] sky130_fd_sc_hd__buf_2
Xoutput112 net112 VGND VGND VPWR VPWR N4BEG[8] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_10_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput36 S2MID[3] VGND VGND VPWR VPWR net36 sky130_fd_sc_hd__clkbuf_1
Xinput25 S2END[0] VGND VGND VPWR VPWR net25 sky130_fd_sc_hd__clkbuf_1
Xstrobe_outbuf_12__0_ FrameStrobe_O_i\[12\] VGND VGND VPWR VPWR net61 sky130_fd_sc_hd__clkbuf_1
Xinput14 FrameStrobe[3] VGND VGND VPWR VPWR net14 sky130_fd_sc_hd__clkbuf_1
Xinput47 S4END[15] VGND VGND VPWR VPWR net47 sky130_fd_sc_hd__buf_1
XFILLER_0_3_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_71 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_5_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_79 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_35 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_46 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_57 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_68 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_167 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xstrobe_outbuf_7__0_ FrameStrobe_O_i\[7\] VGND VGND VPWR VPWR net75 sky130_fd_sc_hd__buf_1
Xoutput102 net102 VGND VGND VPWR VPWR N4BEG[13] sky130_fd_sc_hd__buf_2
Xoutput113 net113 VGND VGND VPWR VPWR N4BEG[9] sky130_fd_sc_hd__buf_2
XFILLER_0_10_165 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_10_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput48 S4END[1] VGND VGND VPWR VPWR net48 sky130_fd_sc_hd__clkbuf_1
Xinput37 S2MID[4] VGND VGND VPWR VPWR net37 sky130_fd_sc_hd__clkbuf_1
Xinput26 S2END[1] VGND VGND VPWR VPWR net26 sky130_fd_sc_hd__clkbuf_1
Xinput15 FrameStrobe[4] VGND VGND VPWR VPWR net15 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_81 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_39 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_69 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_36 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_47 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_58 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_20 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput114 net114 VGND VGND VPWR VPWR UserCLKo sky130_fd_sc_hd__buf_2
Xoutput103 net103 VGND VGND VPWR VPWR N4BEG[14] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_12_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_10_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xinput27 S2END[2] VGND VGND VPWR VPWR net27 sky130_fd_sc_hd__clkbuf_1
Xinput49 S4END[2] VGND VGND VPWR VPWR net49 sky130_fd_sc_hd__clkbuf_1
Xinput38 S2MID[5] VGND VGND VPWR VPWR net38 sky130_fd_sc_hd__clkbuf_1
Xinput16 FrameStrobe[5] VGND VGND VPWR VPWR net16 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_206 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_93 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_40 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_1_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xstrobe_inbuf_0__0_ net1 VGND VGND VPWR VPWR FrameStrobe_O_i\[0\] sky130_fd_sc_hd__clkbuf_1
XTAP_37 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_48 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_6_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XTAP_59 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_21 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput104 net104 VGND VGND VPWR VPWR N4BEG[15] sky130_fd_sc_hd__clkbuf_4
Xstrobe_outbuf_15__0_ FrameStrobe_O_i\[15\] VGND VGND VPWR VPWR net64 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_6_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xinput39 S2MID[6] VGND VGND VPWR VPWR net39 sky130_fd_sc_hd__clkbuf_1
Xinput28 S2END[3] VGND VGND VPWR VPWR net28 sky130_fd_sc_hd__clkbuf_1
Xinput17 FrameStrobe[6] VGND VGND VPWR VPWR net17 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_51 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_7_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_8_29 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xstrobe_inbuf_12__0_ net4 VGND VGND VPWR VPWR FrameStrobe_O_i\[12\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_0_85 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
XFILLER_0_0_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XTAP_38 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_49 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_137 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_11 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput105 net105 VGND VGND VPWR VPWR N4BEG[1] sky130_fd_sc_hd__clkbuf_4
Xinput29 S2END[4] VGND VGND VPWR VPWR net29 sky130_fd_sc_hd__clkbuf_1
Xinput18 FrameStrobe[7] VGND VGND VPWR VPWR net18 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_2_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XTAP_28 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XTAP_39 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_9_149 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_12 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_41 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_85 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_23 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput106 net106 VGND VGND VPWR VPWR N4BEG[2] sky130_fd_sc_hd__clkbuf_4
Xinput19 FrameStrobe[8] VGND VGND VPWR VPWR net19 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_2_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_2_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_225 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_10 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xstrobe_inbuf_3__0_ net14 VGND VGND VPWR VPWR FrameStrobe_O_i\[3\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_3_250 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XTAP_29 VGND VPWR sky130_fd_sc_hd__tapvpwrvgnd_1
Xstrobe_outbuf_18__0_ FrameStrobe_O_i\[18\] VGND VGND VPWR VPWR net67 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_6_53 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_97 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_24 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_4_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_13 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput107 net107 VGND VGND VPWR VPWR N4BEG[3] sky130_fd_sc_hd__buf_2
XFILLER_0_12_78 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xstrobe_outbuf_0__0_ FrameStrobe_O_i\[0\] VGND VGND VPWR VPWR net58 sky130_fd_sc_hd__buf_1
XFILLER_0_2_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xstrobe_inbuf_15__0_ net7 VGND VGND VPWR VPWR FrameStrobe_O_i\[15\] sky130_fd_sc_hd__clkbuf_1
XInst_S_term_RAM_IO_switch_matrix__29_ net44 VGND VGND VPWR VPWR net107 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_237 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_99 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_0_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_22 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_53 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_25 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_65 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_195 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput90 net90 VGND VGND VPWR VPWR N2BEGb[0] sky130_fd_sc_hd__buf_2
Xoutput108 net108 VGND VGND VPWR VPWR N4BEG[4] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_12_46 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_55 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_S_term_RAM_IO_switch_matrix__28_ net45 VGND VGND VPWR VPWR net106 sky130_fd_sc_hd__buf_1
XFILLER_0_7_205 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_7_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_11_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_9_21 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_222 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XPHY_26 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_77 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XPHY_15 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_141 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput109 net109 VGND VGND VPWR VPWR N4BEG[5] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_12_191 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_10_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput91 net91 VGND VGND VPWR VPWR N2BEGb[1] sky130_fd_sc_hd__buf_2
Xoutput80 net80 VGND VGND VPWR VPWR N1BEG[2] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_5_111 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_5_166 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XInst_S_term_RAM_IO_switch_matrix__27_ net41 VGND VGND VPWR VPWR net104 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_7_217 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xstrobe_inbuf_6__0_ net17 VGND VGND VPWR VPWR FrameStrobe_O_i\[6\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_4_209 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_0_57 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_33 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_13_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XPHY_16 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_153 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_197 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput70 net70 VGND VGND VPWR VPWR FrameStrobe_O[2] sky130_fd_sc_hd__buf_2
Xoutput92 net92 VGND VGND VPWR VPWR N2BEGb[2] sky130_fd_sc_hd__clkbuf_4
Xstrobe_outbuf_3__0_ FrameStrobe_O_i\[3\] VGND VGND VPWR VPWR net71 sky130_fd_sc_hd__buf_1
Xoutput81 net81 VGND VGND VPWR VPWR N1BEG[3] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_2_3 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xstrobe_inbuf_18__0_ net10 VGND VGND VPWR VPWR FrameStrobe_O_i\[18\] sky130_fd_sc_hd__clkbuf_1
XFILLER_0_1_181 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_S_term_RAM_IO_switch_matrix__26_ net48 VGND VGND VPWR VPWR net103 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_202 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_S_term_RAM_IO_switch_matrix__09_ net35 VGND VGND VPWR VPWR net87 sky130_fd_sc_hd__buf_1
XFILLER_0_0_14 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_9_45 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_0_235 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XANTENNA_1 net82 VGND VGND VPWR VPWR sky130_fd_sc_hd__diode_2
XPHY_17 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_8_121 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_165 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput71 net71 VGND VGND VPWR VPWR FrameStrobe_O[3] sky130_fd_sc_hd__clkbuf_4
Xoutput93 net93 VGND VGND VPWR VPWR N2BEGb[3] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_12_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput82 net82 VGND VGND VPWR VPWR N2BEG[0] sky130_fd_sc_hd__clkbuf_4
Xoutput60 net60 VGND VGND VPWR VPWR FrameStrobe_O[11] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_5_113 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_146 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_1_193 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_3_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_S_term_RAM_IO_switch_matrix__25_ net49 VGND VGND VPWR VPWR net102 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_225 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_214 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XInst_S_term_RAM_IO_switch_matrix__08_ net36 VGND VGND VPWR VPWR net86 sky130_fd_sc_hd__buf_1
XFILLER_0_0_48 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_233 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_3_244 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_9_57 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_8_133 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_8_177 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XPHY_18 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xoutput72 net72 VGND VGND VPWR VPWR FrameStrobe_O[4] sky130_fd_sc_hd__clkbuf_4
Xoutput94 net94 VGND VGND VPWR VPWR N2BEGb[4] sky130_fd_sc_hd__clkbuf_4
Xoutput83 net83 VGND VGND VPWR VPWR N2BEG[1] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_10_109 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xoutput61 net61 VGND VGND VPWR VPWR FrameStrobe_O[12] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_5_125 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_5_158 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_8
XFILLER_0_5_169 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
Xstrobe_outbuf_11__0_ FrameStrobe_O_i\[11\] VGND VGND VPWR VPWR net60 sky130_fd_sc_hd__buf_1
XFILLER_0_2_139 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_S_term_RAM_IO_switch_matrix__24_ net50 VGND VGND VPWR VPWR net101 sky130_fd_sc_hd__clkbuf_1
Xstrobe_inbuf_9__0_ net20 VGND VGND VPWR VPWR FrameStrobe_O_i\[9\] sky130_fd_sc_hd__clkbuf_1
XInst_S_term_RAM_IO_switch_matrix__07_ net37 VGND VGND VPWR VPWR net85 sky130_fd_sc_hd__buf_1
XFILLER_0_10_83 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_0_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_223 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_9_69 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_6_15 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_12_173 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XPHY_19 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
Xstrobe_outbuf_6__0_ FrameStrobe_O_i\[6\] VGND VGND VPWR VPWR net74 sky130_fd_sc_hd__buf_1
XFILLER_0_8_189 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
Xoutput73 net73 VGND VGND VPWR VPWR FrameStrobe_O[5] sky130_fd_sc_hd__clkbuf_4
Xoutput95 net95 VGND VGND VPWR VPWR N2BEGb[5] sky130_fd_sc_hd__buf_2
XFILLER_0_12_29 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
Xoutput84 net84 VGND VGND VPWR VPWR N2BEG[2] sky130_fd_sc_hd__clkbuf_4
Xoutput62 net62 VGND VGND VPWR VPWR FrameStrobe_O[13] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_5_137 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
XFILLER_0_11_3 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_4_181 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_3_27 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XFILLER_0_9_251 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_162 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XInst_S_term_RAM_IO_switch_matrix__23_ net51 VGND VGND VPWR VPWR net100 sky130_fd_sc_hd__clkbuf_1
XFILLER_0_11_249 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_3
XFILLER_0_6_221 VGND VGND VPWR VPWR sky130_ef_sc_hd__decap_12
XInst_S_term_RAM_IO_switch_matrix__06_ net38 VGND VGND VPWR VPWR net84 sky130_fd_sc_hd__buf_1
XFILLER_0_0_205 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_1_82 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_2
XFILLER_0_6_27 VGND VGND VPWR VPWR sky130_fd_sc_hd__fill_1
XFILLER_0_12_141 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_4
Xoutput96 net96 VGND VGND VPWR VPWR N2BEGb[6] sky130_fd_sc_hd__buf_2
Xoutput74 net74 VGND VGND VPWR VPWR FrameStrobe_O[6] sky130_fd_sc_hd__clkbuf_4
Xoutput85 net85 VGND VGND VPWR VPWR N2BEG[3] sky130_fd_sc_hd__clkbuf_4
Xoutput63 net63 VGND VGND VPWR VPWR FrameStrobe_O[14] sky130_fd_sc_hd__clkbuf_4
XFILLER_0_5_105 VGND VGND VPWR VPWR sky130_fd_sc_hd__decap_6
.ends

