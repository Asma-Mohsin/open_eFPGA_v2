// This is the unpowered netlist.
module BlockRAM_1KB (C0,
    C1,
    C2,
    C3,
    C4,
    C5,
    clk,
    rd_addr,
    rd_data,
    wr_addr,
    wr_data);
 input C0;
 input C1;
 input C2;
 input C3;
 input C4;
 input C5;
 input clk;
 input [7:0] rd_addr;
 output [31:0] rd_data;
 input [7:0] wr_addr;
 input [31:0] wr_data;

 wire _000_;
 wire _001_;
 wire _002_;
 wire _003_;
 wire _004_;
 wire _005_;
 wire _006_;
 wire _007_;
 wire _008_;
 wire _009_;
 wire _010_;
 wire _011_;
 wire _012_;
 wire _013_;
 wire _014_;
 wire _015_;
 wire _016_;
 wire _017_;
 wire _018_;
 wire _019_;
 wire _020_;
 wire _021_;
 wire _022_;
 wire _023_;
 wire _024_;
 wire _025_;
 wire _026_;
 wire _027_;
 wire _028_;
 wire _029_;
 wire _030_;
 wire _031_;
 wire _032_;
 wire _033_;
 wire _034_;
 wire _035_;
 wire _036_;
 wire _037_;
 wire _038_;
 wire _039_;
 wire _040_;
 wire _041_;
 wire _042_;
 wire _043_;
 wire _044_;
 wire _045_;
 wire _046_;
 wire _047_;
 wire _048_;
 wire _049_;
 wire _050_;
 wire _051_;
 wire _052_;
 wire _053_;
 wire _054_;
 wire _055_;
 wire _056_;
 wire _057_;
 wire _058_;
 wire _059_;
 wire _060_;
 wire _061_;
 wire _062_;
 wire _063_;
 wire _064_;
 wire _065_;
 wire _066_;
 wire _067_;
 wire _068_;
 wire _069_;
 wire _070_;
 wire _071_;
 wire _072_;
 wire _073_;
 wire _074_;
 wire _075_;
 wire _076_;
 wire _077_;
 wire _078_;
 wire _079_;
 wire _080_;
 wire _081_;
 wire _082_;
 wire _083_;
 wire _084_;
 wire _085_;
 wire _086_;
 wire _087_;
 wire _088_;
 wire _089_;
 wire _090_;
 wire _091_;
 wire _092_;
 wire _093_;
 wire _094_;
 wire _095_;
 wire _096_;
 wire _097_;
 wire _098_;
 wire _099_;
 wire _100_;
 wire _101_;
 wire _102_;
 wire _103_;
 wire _104_;
 wire _105_;
 wire _106_;
 wire _107_;
 wire _108_;
 wire _109_;
 wire _110_;
 wire _111_;
 wire _112_;
 wire _113_;
 wire _114_;
 wire _115_;
 wire _116_;
 wire _117_;
 wire _118_;
 wire _119_;
 wire _120_;
 wire _121_;
 wire _122_;
 wire _123_;
 wire _124_;
 wire _125_;
 wire _126_;
 wire _127_;
 wire _128_;
 wire _129_;
 wire _130_;
 wire _131_;
 wire _132_;
 wire _133_;
 wire _134_;
 wire _135_;
 wire _136_;
 wire _137_;
 wire _138_;
 wire _139_;
 wire _140_;
 wire _141_;
 wire _142_;
 wire _143_;
 wire _144_;
 wire _145_;
 wire _146_;
 wire _147_;
 wire _148_;
 wire _149_;
 wire _150_;
 wire _151_;
 wire _152_;
 wire _153_;
 wire _154_;
 wire _155_;
 wire _156_;
 wire _157_;
 wire _158_;
 wire _159_;
 wire _160_;
 wire _161_;
 wire _162_;
 wire _163_;
 wire _164_;
 wire _165_;
 wire _166_;
 wire _167_;
 wire _168_;
 wire _169_;
 wire _170_;
 wire _171_;
 wire clknet_0_clk;
 wire clknet_2_0__leaf_clk;
 wire clknet_2_1__leaf_clk;
 wire clknet_2_2__leaf_clk;
 wire clknet_2_3__leaf_clk;
 wire memWriteEnable;
 wire \mem_dout[0] ;
 wire \mem_dout[10] ;
 wire \mem_dout[11] ;
 wire \mem_dout[12] ;
 wire \mem_dout[13] ;
 wire \mem_dout[14] ;
 wire \mem_dout[15] ;
 wire \mem_dout[16] ;
 wire \mem_dout[17] ;
 wire \mem_dout[18] ;
 wire \mem_dout[19] ;
 wire \mem_dout[1] ;
 wire \mem_dout[20] ;
 wire \mem_dout[21] ;
 wire \mem_dout[22] ;
 wire \mem_dout[23] ;
 wire \mem_dout[24] ;
 wire \mem_dout[25] ;
 wire \mem_dout[26] ;
 wire \mem_dout[27] ;
 wire \mem_dout[28] ;
 wire \mem_dout[29] ;
 wire \mem_dout[2] ;
 wire \mem_dout[30] ;
 wire \mem_dout[31] ;
 wire \mem_dout[3] ;
 wire \mem_dout[4] ;
 wire \mem_dout[5] ;
 wire \mem_dout[6] ;
 wire \mem_dout[7] ;
 wire \mem_dout[8] ;
 wire \mem_dout[9] ;
 wire \mem_wr_mask[0] ;
 wire \mem_wr_mask[1] ;
 wire \mem_wr_mask[2] ;
 wire \mem_wr_mask[3] ;
 wire \muxedDataIn[10] ;
 wire \muxedDataIn[11] ;
 wire \muxedDataIn[12] ;
 wire \muxedDataIn[13] ;
 wire \muxedDataIn[14] ;
 wire \muxedDataIn[15] ;
 wire \muxedDataIn[16] ;
 wire \muxedDataIn[17] ;
 wire \muxedDataIn[18] ;
 wire \muxedDataIn[19] ;
 wire \muxedDataIn[20] ;
 wire \muxedDataIn[21] ;
 wire \muxedDataIn[22] ;
 wire \muxedDataIn[23] ;
 wire \muxedDataIn[24] ;
 wire \muxedDataIn[25] ;
 wire \muxedDataIn[26] ;
 wire \muxedDataIn[27] ;
 wire \muxedDataIn[28] ;
 wire \muxedDataIn[29] ;
 wire \muxedDataIn[30] ;
 wire \muxedDataIn[31] ;
 wire \muxedDataIn[8] ;
 wire \muxedDataIn[9] ;
 wire net1;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net18;
 wire net19;
 wire net2;
 wire net20;
 wire net21;
 wire net22;
 wire net23;
 wire net24;
 wire net25;
 wire net26;
 wire net27;
 wire net28;
 wire net29;
 wire net3;
 wire net30;
 wire net31;
 wire net32;
 wire net33;
 wire net34;
 wire net35;
 wire net36;
 wire net37;
 wire net38;
 wire net39;
 wire net4;
 wire net40;
 wire net41;
 wire net42;
 wire net43;
 wire net44;
 wire net45;
 wire net46;
 wire net47;
 wire net48;
 wire net49;
 wire net5;
 wire net50;
 wire net51;
 wire net52;
 wire net53;
 wire net54;
 wire net55;
 wire net56;
 wire net57;
 wire net58;
 wire net59;
 wire net6;
 wire net60;
 wire net61;
 wire net62;
 wire net63;
 wire net64;
 wire net65;
 wire net66;
 wire net67;
 wire net68;
 wire net69;
 wire net7;
 wire net70;
 wire net71;
 wire net72;
 wire net73;
 wire net74;
 wire net75;
 wire net76;
 wire net77;
 wire net78;
 wire net79;
 wire net8;
 wire net80;
 wire net81;
 wire net82;
 wire net83;
 wire net84;
 wire net85;
 wire net86;
 wire net87;
 wire net9;
 wire \rd_dout_additional_register[0] ;
 wire \rd_dout_additional_register[10] ;
 wire \rd_dout_additional_register[11] ;
 wire \rd_dout_additional_register[12] ;
 wire \rd_dout_additional_register[13] ;
 wire \rd_dout_additional_register[14] ;
 wire \rd_dout_additional_register[15] ;
 wire \rd_dout_additional_register[16] ;
 wire \rd_dout_additional_register[17] ;
 wire \rd_dout_additional_register[18] ;
 wire \rd_dout_additional_register[19] ;
 wire \rd_dout_additional_register[1] ;
 wire \rd_dout_additional_register[20] ;
 wire \rd_dout_additional_register[21] ;
 wire \rd_dout_additional_register[22] ;
 wire \rd_dout_additional_register[23] ;
 wire \rd_dout_additional_register[24] ;
 wire \rd_dout_additional_register[25] ;
 wire \rd_dout_additional_register[26] ;
 wire \rd_dout_additional_register[27] ;
 wire \rd_dout_additional_register[28] ;
 wire \rd_dout_additional_register[29] ;
 wire \rd_dout_additional_register[2] ;
 wire \rd_dout_additional_register[30] ;
 wire \rd_dout_additional_register[31] ;
 wire \rd_dout_additional_register[3] ;
 wire \rd_dout_additional_register[4] ;
 wire \rd_dout_additional_register[5] ;
 wire \rd_dout_additional_register[6] ;
 wire \rd_dout_additional_register[7] ;
 wire \rd_dout_additional_register[8] ;
 wire \rd_dout_additional_register[9] ;
 wire \rd_dout_muxed[0] ;
 wire \rd_dout_muxed[10] ;
 wire \rd_dout_muxed[11] ;
 wire \rd_dout_muxed[12] ;
 wire \rd_dout_muxed[13] ;
 wire \rd_dout_muxed[14] ;
 wire \rd_dout_muxed[15] ;
 wire \rd_dout_muxed[1] ;
 wire \rd_dout_muxed[2] ;
 wire \rd_dout_muxed[3] ;
 wire \rd_dout_muxed[4] ;
 wire \rd_dout_muxed[5] ;
 wire \rd_dout_muxed[6] ;
 wire \rd_dout_muxed[7] ;
 wire \rd_dout_muxed[8] ;
 wire \rd_dout_muxed[9] ;
 wire \rd_dout_sel[0] ;
 wire \rd_dout_sel[1] ;

 sky130_fd_sc_hd__diode_2 ANTENNA_1 (.DIODE(_164_));
 sky130_fd_sc_hd__diode_2 ANTENNA_10 (.DIODE(\mem_dout[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_11 (.DIODE(\mem_dout[5] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_12 (.DIODE(\mem_dout[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_13 (.DIODE(\mem_dout[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_14 (.DIODE(\mem_dout[8] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_15 (.DIODE(net32));
 sky130_fd_sc_hd__diode_2 ANTENNA_16 (.DIODE(net33));
 sky130_fd_sc_hd__diode_2 ANTENNA_17 (.DIODE(net48));
 sky130_fd_sc_hd__diode_2 ANTENNA_18 (.DIODE(_162_));
 sky130_fd_sc_hd__diode_2 ANTENNA_19 (.DIODE(\mem_dout[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_2 (.DIODE(_166_));
 sky130_fd_sc_hd__diode_2 ANTENNA_20 (.DIODE(\mem_dout[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_21 (.DIODE(\mem_dout[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_22 (.DIODE(\mem_dout[3] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_23 (.DIODE(\mem_dout[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_24 (.DIODE(\mem_dout[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_25 (.DIODE(\mem_dout[7] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_26 (.DIODE(\mem_dout[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_27 (.DIODE(net45));
 sky130_fd_sc_hd__diode_2 ANTENNA_28 (.DIODE(\mem_dout[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_29 (.DIODE(\mem_dout[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_3 (.DIODE(clk));
 sky130_fd_sc_hd__diode_2 ANTENNA_30 (.DIODE(\mem_dout[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_31 (.DIODE(\mem_dout[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_32 (.DIODE(\mem_dout[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_33 (.DIODE(\mem_dout[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_34 (.DIODE(\mem_dout[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_35 (.DIODE(\mem_dout[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_36 (.DIODE(\mem_dout[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_4 (.DIODE(\mem_dout[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_5 (.DIODE(\mem_dout[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_6 (.DIODE(\mem_dout[15] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_7 (.DIODE(\mem_dout[20] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_8 (.DIODE(\mem_dout[27] ));
 sky130_fd_sc_hd__diode_2 ANTENNA_9 (.DIODE(\mem_dout[5] ));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1089 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_1145 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_1149 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_1161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_193 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_209 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_221 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_225 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_233 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_243 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_251 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_257 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_269 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_0_275 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_279 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_285 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_300 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_313 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_317 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_323 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_335 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_0_347 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_363 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_375 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_379 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_391 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_393 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_405 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_409 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_417 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_421 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_433 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_445 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_449 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_461 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_473 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_477 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_489 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_501 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_505 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_517 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_529 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_533 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_545 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_557 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_561 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_573 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_585 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_589 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_601 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_641 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_657 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_669 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_100_47 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_100_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_100_63 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_100_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_100_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_101_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_101_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_72 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_101_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_101_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_101_92 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_102_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_102_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_102_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_48 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_60 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_102_68 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_102_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_102_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_102_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_103_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_103_78 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_103_90 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_104_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_104_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_104_61 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_104_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_104_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_104_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_105_39 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_105_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_105_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_105_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_105_92 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_106_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_106_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_106_63 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_106_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_106_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_106_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_32 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_36 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_107_40 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_107_46 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_107_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_107_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_107_69 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_108_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_108_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_108_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_108_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_108_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_109_30 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_109_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_109_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_109_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_109_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_110_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_110_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_110_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_111_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_111_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_111_7 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_111_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_112_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_112_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_112_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_112_59 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_112_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_112_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_21 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_33 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_113_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_44 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_113_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_113_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_113_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_114_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_114_57 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_114_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_114_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_114_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_115_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_115_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_115_78 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_115_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_49 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_116_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_116_74 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_116_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_117_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_117_40 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_44 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_117_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_117_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_78 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_117_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_118_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_118_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_68 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_118_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_118_80 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_118_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_119_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_119_39 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_119_43 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_119_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_119_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_119_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_11_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_120_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_29 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_120_43 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_120_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_120_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_120_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_121_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_121_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_121_33 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_121_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_67 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_71 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_121_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_43 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_122_63 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_122_7 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_122_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_122_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_122_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_123_31 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_39 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_123_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_57 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_123_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_123_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_124_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_124_3 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_51 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_55 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_124_75 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_124_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_124_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_125_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_125_66 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_125_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_125_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_125_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_126_3 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_126_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_126_81 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_126_85 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_126_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_127_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_127_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_127_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_127_79 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_128_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_128_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_128_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_69 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_128_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_129_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_129_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_129_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_12_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_29 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_56 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_130_7 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_130_74 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_130_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_130_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_130_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_131_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_131_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_55 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_131_73 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_131_91 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_132_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_41 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_47 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_132_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_132_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_71 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_132_81 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_132_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_133_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_55 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_133_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_133_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_133_78 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_133_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_134_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_134_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_134_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_134_77 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_135_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_135_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_135_69 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_135_75 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_136_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_136_7 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_136_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_136_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_137_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_137_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_138_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_138_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_138_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_138_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_139_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_139_7 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_139_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_13_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_13_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_140_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_140_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_140_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_140_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_141_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_141_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_142_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_142_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_142_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_142_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_143_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_143_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_144_7 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_144_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_144_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_144_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_145_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_145_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_145_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_146_7 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_146_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_146_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_146_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_147_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_147_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_147_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_148_7 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_148_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_148_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_148_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_149_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_149_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_149_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_14_85 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_150_7 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_150_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_150_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_150_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_151_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_151_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_152_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_152_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_152_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_152_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_153_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_153_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_154_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_154_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_154_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_154_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_155_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_155_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_155_81 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_1005 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1009 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1021 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_1033 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1037 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1049 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_1061 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1065 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1077 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_1089 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1093 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1105 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_1117 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1121 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_1133 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_1145 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_1149 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_1157 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_1163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_1167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_169 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_181 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_193 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_197 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_207 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_219 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_223 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_225 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_237 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_249 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_262 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_274 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_290 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_3 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_302 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_309 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_321 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_333 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_337 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_349 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_361 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_365 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_156_385 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_391 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_402 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_412 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_416 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_421 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_425 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_445 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_449 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_453 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_456 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_497 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_501 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_505 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_524 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_528 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_533 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_537 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_541 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_546 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_550 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_554 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_561 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_156_566 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_57 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_605 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_613 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_617 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_629 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_641 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_156_645 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_655 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_156_667 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_156_671 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_673 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_685 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_697 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_701 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_713 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_725 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_729 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_741 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_753 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_757 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_769 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_781 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_785 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_797 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_809 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_813 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_825 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_837 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_841 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_853 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_865 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_869 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_881 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_893 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_897 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_909 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_921 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_925 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_937 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_949 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_953 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_965 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_97 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_156_977 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_981 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_156_993 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_15_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_17_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_71 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_71 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_24_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_24_73 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_24_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_25_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_25_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_27_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_28_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_80 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_28_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_29_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_72 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_74 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_30_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_30_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_31_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_14 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_32_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_65 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_32_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_32_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_34_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_71 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_37_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_47 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_59 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_71 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_83 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_38_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_19 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_39_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_75 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_87 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_48 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_60 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_40_72 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_40_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_18 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_30 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_50 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_36 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_60 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_66 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_42_80 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_42_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_19 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_7 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_44_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_72 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_44_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_19 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_31 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_36 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_45_48 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_54 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_64 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_7 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_84 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_45_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_27 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_34 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_46 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_58 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_46_76 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_46_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_55 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_47_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_92 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_48_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_48_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_9 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_50_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_74 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_50_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_70 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_76 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_86 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_52_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_52_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_53_54 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_6 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_53_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_72 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_54_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_18 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_30 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_42 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_55_54 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_56_61 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_56_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_57_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_61 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_71 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_9 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_57_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_53 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_73 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_58_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_59_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_59_84 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_6 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_65 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_60_73 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_60_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_92 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_62_26 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_62_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_81 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_53 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_64_65 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_71 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_64_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_84 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_92 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_41 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_61 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_66_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_66_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_67_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_53 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_68_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_78 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_68_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_69_57 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_69_62 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_71_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_71_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_27 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_35 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_73 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_72_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_72_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_73_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_74_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_40 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_74_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_27 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_76_29 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_67 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_76_79 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_76_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_89 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_78_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_78_29 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_40 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_52 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_6 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_60 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_78_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_3 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_47 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_55 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_89 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_81 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_18 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_26 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_80_29 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_50 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_80_58 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_6 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_70 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_80_82 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_80_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_21 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_81_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_43 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_55 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_65 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_72 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_80 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_59 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_76 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_83 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_82_91 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_33 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_83_45 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_83_49 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_83_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_84_45 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_84_57 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_84_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_84_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_84_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_85_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_85_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_85_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_85_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_86_41 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_86_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_86_59 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_86_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_21 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_33 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_87_40 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_87_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_87_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_87_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_87_92 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_88_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_41 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_88_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_88_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_88_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_88_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_89_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_89_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_89_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_53 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_89_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_89_79 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_89_91 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_9 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_90_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_90_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_90_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_90_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_91_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_91_88 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_91_92 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_92_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_92_53 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_92_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_92_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_92_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_15 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_93_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_38 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_93_50 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_93_77 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_93_89 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_41 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_94_56 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_60 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_94_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_94_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_94_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_94_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_21 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_95_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_95_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_53 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_95_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_95_63 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_78 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_95_9 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_95_90 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_27 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_3 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_37 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_96_44 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_56 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_96_69 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_75 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_96_83 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_96_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_21 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_40 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_52 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_97_57 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_65 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_76 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_97_88 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_97_9 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_97_92 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_27 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_98_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_3 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_98_33 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_37 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_49 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_98_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_98_64 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_76 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_98_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_21 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_33 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_99_45 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_99_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_99_9 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_81 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_166 ();
 sky130_fd_sc_hd__decap_3 PHY_167 ();
 sky130_fd_sc_hd__decap_3 PHY_168 ();
 sky130_fd_sc_hd__decap_3 PHY_169 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_170 ();
 sky130_fd_sc_hd__decap_3 PHY_171 ();
 sky130_fd_sc_hd__decap_3 PHY_172 ();
 sky130_fd_sc_hd__decap_3 PHY_173 ();
 sky130_fd_sc_hd__decap_3 PHY_174 ();
 sky130_fd_sc_hd__decap_3 PHY_175 ();
 sky130_fd_sc_hd__decap_3 PHY_176 ();
 sky130_fd_sc_hd__decap_3 PHY_177 ();
 sky130_fd_sc_hd__decap_3 PHY_178 ();
 sky130_fd_sc_hd__decap_3 PHY_179 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_180 ();
 sky130_fd_sc_hd__decap_3 PHY_181 ();
 sky130_fd_sc_hd__decap_3 PHY_182 ();
 sky130_fd_sc_hd__decap_3 PHY_183 ();
 sky130_fd_sc_hd__decap_3 PHY_184 ();
 sky130_fd_sc_hd__decap_3 PHY_185 ();
 sky130_fd_sc_hd__decap_3 PHY_186 ();
 sky130_fd_sc_hd__decap_3 PHY_187 ();
 sky130_fd_sc_hd__decap_3 PHY_188 ();
 sky130_fd_sc_hd__decap_3 PHY_189 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_190 ();
 sky130_fd_sc_hd__decap_3 PHY_191 ();
 sky130_fd_sc_hd__decap_3 PHY_192 ();
 sky130_fd_sc_hd__decap_3 PHY_193 ();
 sky130_fd_sc_hd__decap_3 PHY_194 ();
 sky130_fd_sc_hd__decap_3 PHY_195 ();
 sky130_fd_sc_hd__decap_3 PHY_196 ();
 sky130_fd_sc_hd__decap_3 PHY_197 ();
 sky130_fd_sc_hd__decap_3 PHY_198 ();
 sky130_fd_sc_hd__decap_3 PHY_199 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_200 ();
 sky130_fd_sc_hd__decap_3 PHY_201 ();
 sky130_fd_sc_hd__decap_3 PHY_202 ();
 sky130_fd_sc_hd__decap_3 PHY_203 ();
 sky130_fd_sc_hd__decap_3 PHY_204 ();
 sky130_fd_sc_hd__decap_3 PHY_205 ();
 sky130_fd_sc_hd__decap_3 PHY_206 ();
 sky130_fd_sc_hd__decap_3 PHY_207 ();
 sky130_fd_sc_hd__decap_3 PHY_208 ();
 sky130_fd_sc_hd__decap_3 PHY_209 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_210 ();
 sky130_fd_sc_hd__decap_3 PHY_211 ();
 sky130_fd_sc_hd__decap_3 PHY_212 ();
 sky130_fd_sc_hd__decap_3 PHY_213 ();
 sky130_fd_sc_hd__decap_3 PHY_214 ();
 sky130_fd_sc_hd__decap_3 PHY_215 ();
 sky130_fd_sc_hd__decap_3 PHY_216 ();
 sky130_fd_sc_hd__decap_3 PHY_217 ();
 sky130_fd_sc_hd__decap_3 PHY_218 ();
 sky130_fd_sc_hd__decap_3 PHY_219 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_220 ();
 sky130_fd_sc_hd__decap_3 PHY_221 ();
 sky130_fd_sc_hd__decap_3 PHY_222 ();
 sky130_fd_sc_hd__decap_3 PHY_223 ();
 sky130_fd_sc_hd__decap_3 PHY_224 ();
 sky130_fd_sc_hd__decap_3 PHY_225 ();
 sky130_fd_sc_hd__decap_3 PHY_226 ();
 sky130_fd_sc_hd__decap_3 PHY_227 ();
 sky130_fd_sc_hd__decap_3 PHY_228 ();
 sky130_fd_sc_hd__decap_3 PHY_229 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_230 ();
 sky130_fd_sc_hd__decap_3 PHY_231 ();
 sky130_fd_sc_hd__decap_3 PHY_232 ();
 sky130_fd_sc_hd__decap_3 PHY_233 ();
 sky130_fd_sc_hd__decap_3 PHY_234 ();
 sky130_fd_sc_hd__decap_3 PHY_235 ();
 sky130_fd_sc_hd__decap_3 PHY_236 ();
 sky130_fd_sc_hd__decap_3 PHY_237 ();
 sky130_fd_sc_hd__decap_3 PHY_238 ();
 sky130_fd_sc_hd__decap_3 PHY_239 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_240 ();
 sky130_fd_sc_hd__decap_3 PHY_241 ();
 sky130_fd_sc_hd__decap_3 PHY_242 ();
 sky130_fd_sc_hd__decap_3 PHY_243 ();
 sky130_fd_sc_hd__decap_3 PHY_244 ();
 sky130_fd_sc_hd__decap_3 PHY_245 ();
 sky130_fd_sc_hd__decap_3 PHY_246 ();
 sky130_fd_sc_hd__decap_3 PHY_247 ();
 sky130_fd_sc_hd__decap_3 PHY_248 ();
 sky130_fd_sc_hd__decap_3 PHY_249 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_250 ();
 sky130_fd_sc_hd__decap_3 PHY_251 ();
 sky130_fd_sc_hd__decap_3 PHY_252 ();
 sky130_fd_sc_hd__decap_3 PHY_253 ();
 sky130_fd_sc_hd__decap_3 PHY_254 ();
 sky130_fd_sc_hd__decap_3 PHY_255 ();
 sky130_fd_sc_hd__decap_3 PHY_256 ();
 sky130_fd_sc_hd__decap_3 PHY_257 ();
 sky130_fd_sc_hd__decap_3 PHY_258 ();
 sky130_fd_sc_hd__decap_3 PHY_259 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_260 ();
 sky130_fd_sc_hd__decap_3 PHY_261 ();
 sky130_fd_sc_hd__decap_3 PHY_262 ();
 sky130_fd_sc_hd__decap_3 PHY_263 ();
 sky130_fd_sc_hd__decap_3 PHY_264 ();
 sky130_fd_sc_hd__decap_3 PHY_265 ();
 sky130_fd_sc_hd__decap_3 PHY_266 ();
 sky130_fd_sc_hd__decap_3 PHY_267 ();
 sky130_fd_sc_hd__decap_3 PHY_268 ();
 sky130_fd_sc_hd__decap_3 PHY_269 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_270 ();
 sky130_fd_sc_hd__decap_3 PHY_271 ();
 sky130_fd_sc_hd__decap_3 PHY_272 ();
 sky130_fd_sc_hd__decap_3 PHY_273 ();
 sky130_fd_sc_hd__decap_3 PHY_274 ();
 sky130_fd_sc_hd__decap_3 PHY_275 ();
 sky130_fd_sc_hd__decap_3 PHY_276 ();
 sky130_fd_sc_hd__decap_3 PHY_277 ();
 sky130_fd_sc_hd__decap_3 PHY_278 ();
 sky130_fd_sc_hd__decap_3 PHY_279 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_280 ();
 sky130_fd_sc_hd__decap_3 PHY_281 ();
 sky130_fd_sc_hd__decap_3 PHY_282 ();
 sky130_fd_sc_hd__decap_3 PHY_283 ();
 sky130_fd_sc_hd__decap_3 PHY_284 ();
 sky130_fd_sc_hd__decap_3 PHY_285 ();
 sky130_fd_sc_hd__decap_3 PHY_286 ();
 sky130_fd_sc_hd__decap_3 PHY_287 ();
 sky130_fd_sc_hd__decap_3 PHY_288 ();
 sky130_fd_sc_hd__decap_3 PHY_289 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_290 ();
 sky130_fd_sc_hd__decap_3 PHY_291 ();
 sky130_fd_sc_hd__decap_3 PHY_292 ();
 sky130_fd_sc_hd__decap_3 PHY_293 ();
 sky130_fd_sc_hd__decap_3 PHY_294 ();
 sky130_fd_sc_hd__decap_3 PHY_295 ();
 sky130_fd_sc_hd__decap_3 PHY_296 ();
 sky130_fd_sc_hd__decap_3 PHY_297 ();
 sky130_fd_sc_hd__decap_3 PHY_298 ();
 sky130_fd_sc_hd__decap_3 PHY_299 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_300 ();
 sky130_fd_sc_hd__decap_3 PHY_301 ();
 sky130_fd_sc_hd__decap_3 PHY_302 ();
 sky130_fd_sc_hd__decap_3 PHY_303 ();
 sky130_fd_sc_hd__decap_3 PHY_304 ();
 sky130_fd_sc_hd__decap_3 PHY_305 ();
 sky130_fd_sc_hd__decap_3 PHY_306 ();
 sky130_fd_sc_hd__decap_3 PHY_307 ();
 sky130_fd_sc_hd__decap_3 PHY_308 ();
 sky130_fd_sc_hd__decap_3 PHY_309 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_310 ();
 sky130_fd_sc_hd__decap_3 PHY_311 ();
 sky130_fd_sc_hd__decap_3 PHY_312 ();
 sky130_fd_sc_hd__decap_3 PHY_313 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_421 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_422 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_423 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_424 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_425 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_426 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_427 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_428 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_429 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_430 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_431 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_432 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_433 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_434 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_435 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_436 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_437 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_438 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_439 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_440 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_441 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_442 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_443 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_444 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_445 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_446 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_447 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_448 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_449 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_450 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_451 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_452 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_453 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_454 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_455 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_456 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_457 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_458 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_459 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_460 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_461 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_462 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_463 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_464 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_465 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_466 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_467 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_468 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_469 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_470 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_471 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_472 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_473 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_474 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_475 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_476 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_477 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_478 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_479 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_480 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_481 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_482 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_483 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_484 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_485 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_486 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_487 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_488 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_489 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_490 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_491 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_492 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_493 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_494 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_495 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_496 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_497 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_498 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_499 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_500 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_501 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_502 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_503 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_504 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_505 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_506 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_507 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_508 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_509 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_510 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_511 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_512 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_513 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_514 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_515 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_516 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_517 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_518 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_519 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_520 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_521 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_522 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_523 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_524 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_525 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_526 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_527 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_528 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_529 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_530 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_531 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_532 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_533 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_534 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_535 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_536 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_537 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_538 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_539 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_540 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_541 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_542 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_543 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_544 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_545 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_546 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_547 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_548 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_549 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_550 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_551 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_552 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_553 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_554 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_555 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_556 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_557 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_558 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_559 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_560 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_561 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_562 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_563 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_564 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_565 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_566 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_567 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_568 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_569 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_570 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_571 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_572 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_573 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_574 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_575 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_576 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_577 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_578 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_579 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_580 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_581 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_582 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_583 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_584 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_585 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_586 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_587 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_588 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_589 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_590 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_591 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_592 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_593 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_594 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_595 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_596 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_597 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_598 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_599 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_600 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_601 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_602 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_603 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_604 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_605 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_606 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_607 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_608 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_609 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_610 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_611 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_612 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_613 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_614 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_615 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_616 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_617 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_618 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_619 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_620 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_621 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_622 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_623 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_624 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_625 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_626 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_627 ();
 sky130_fd_sc_hd__or2_1 _173_ (.A(_065_),
    .B(_069_),
    .X(_070_));
 sky130_fd_sc_hd__clkbuf_1 _174_ (.A(_070_),
    .X(\rd_dout_muxed[4] ));
 sky130_fd_sc_hd__or2b_1 _175_ (.A(\rd_dout_additional_register[4] ),
    .B_N(_054_),
    .X(_071_));
 sky130_fd_sc_hd__o31a_1 _176_ (.A1(_031_),
    .A2(_065_),
    .A3(_069_),
    .B1(_071_),
    .X(net81));
 sky130_fd_sc_hd__mux2_1 _177_ (.A0(\mem_dout[5] ),
    .A1(\mem_dout[21] ),
    .S(_007_),
    .X(_072_));
 sky130_fd_sc_hd__and2_1 _178_ (.A(_005_),
    .B(_072_),
    .X(_073_));
 sky130_fd_sc_hd__or3b_1 _179_ (.A(_037_),
    .B(\mem_dout[21] ),
    .C_N(_013_),
    .X(_074_));
 sky130_fd_sc_hd__o211a_1 _180_ (.A1(\mem_dout[29] ),
    .A2(_019_),
    .B1(_074_),
    .C1(_023_),
    .X(_075_));
 sky130_fd_sc_hd__a211o_1 _181_ (.A1(\mem_dout[13] ),
    .A2(_040_),
    .B1(_041_),
    .C1(_042_),
    .X(_076_));
 sky130_fd_sc_hd__o221a_2 _182_ (.A1(\mem_dout[5] ),
    .A2(_015_),
    .B1(_075_),
    .B2(_076_),
    .C1(_026_),
    .X(_077_));
 sky130_fd_sc_hd__or2_1 _183_ (.A(_073_),
    .B(_077_),
    .X(_078_));
 sky130_fd_sc_hd__clkbuf_1 _184_ (.A(_078_),
    .X(\rd_dout_muxed[5] ));
 sky130_fd_sc_hd__or2b_1 _185_ (.A(\rd_dout_additional_register[5] ),
    .B_N(_054_),
    .X(_079_));
 sky130_fd_sc_hd__o31a_1 _186_ (.A1(_033_),
    .A2(_073_),
    .A3(_077_),
    .B1(_079_),
    .X(net82));
 sky130_fd_sc_hd__mux2_1 _187_ (.A0(\mem_dout[6] ),
    .A1(\mem_dout[22] ),
    .S(_007_),
    .X(_080_));
 sky130_fd_sc_hd__and2_1 _188_ (.A(_005_),
    .B(_080_),
    .X(_081_));
 sky130_fd_sc_hd__or3b_1 _189_ (.A(_012_),
    .B(\mem_dout[22] ),
    .C_N(_013_),
    .X(_082_));
 sky130_fd_sc_hd__o211a_1 _190_ (.A1(\mem_dout[30] ),
    .A2(_019_),
    .B1(_082_),
    .C1(_023_),
    .X(_083_));
 sky130_fd_sc_hd__a211o_1 _191_ (.A1(\mem_dout[14] ),
    .A2(_017_),
    .B1(_014_),
    .C1(_011_),
    .X(_084_));
 sky130_fd_sc_hd__o221a_1 _192_ (.A1(\mem_dout[6] ),
    .A2(_015_),
    .B1(_083_),
    .B2(_084_),
    .C1(_026_),
    .X(_085_));
 sky130_fd_sc_hd__or2_1 _193_ (.A(_081_),
    .B(_085_),
    .X(_086_));
 sky130_fd_sc_hd__clkbuf_1 _194_ (.A(_086_),
    .X(\rd_dout_muxed[6] ));
 sky130_fd_sc_hd__or2b_1 _195_ (.A(\rd_dout_additional_register[6] ),
    .B_N(_054_),
    .X(_087_));
 sky130_fd_sc_hd__o31a_1 _196_ (.A1(_033_),
    .A2(_081_),
    .A3(_085_),
    .B1(_087_),
    .X(net83));
 sky130_fd_sc_hd__mux2_1 _197_ (.A0(\mem_dout[7] ),
    .A1(\mem_dout[23] ),
    .S(_007_),
    .X(_088_));
 sky130_fd_sc_hd__and2_1 _198_ (.A(_005_),
    .B(_088_),
    .X(_089_));
 sky130_fd_sc_hd__or3b_1 _199_ (.A(_012_),
    .B(\mem_dout[23] ),
    .C_N(_013_),
    .X(_090_));
 sky130_fd_sc_hd__o211a_1 _200_ (.A1(\mem_dout[31] ),
    .A2(_019_),
    .B1(_090_),
    .C1(_023_),
    .X(_091_));
 sky130_fd_sc_hd__a211o_1 _201_ (.A1(\mem_dout[15] ),
    .A2(_017_),
    .B1(_014_),
    .C1(_011_),
    .X(_092_));
 sky130_fd_sc_hd__o221a_1 _202_ (.A1(\mem_dout[7] ),
    .A2(_015_),
    .B1(_091_),
    .B2(_092_),
    .C1(_026_),
    .X(_093_));
 sky130_fd_sc_hd__or2_1 _203_ (.A(_089_),
    .B(_093_),
    .X(_094_));
 sky130_fd_sc_hd__clkbuf_1 _204_ (.A(_094_),
    .X(\rd_dout_muxed[7] ));
 sky130_fd_sc_hd__or2b_1 _205_ (.A(\rd_dout_additional_register[7] ),
    .B_N(_030_),
    .X(_095_));
 sky130_fd_sc_hd__o31a_1 _206_ (.A1(_033_),
    .A2(_089_),
    .A3(_093_),
    .B1(_095_),
    .X(net84));
 sky130_fd_sc_hd__and2_2 _207_ (.A(_012_),
    .B(_005_),
    .X(_096_));
 sky130_fd_sc_hd__buf_2 _208_ (.A(_096_),
    .X(_097_));
 sky130_fd_sc_hd__mux2_1 _209_ (.A0(\mem_dout[8] ),
    .A1(\mem_dout[24] ),
    .S(_097_),
    .X(_098_));
 sky130_fd_sc_hd__buf_1 _210_ (.A(_098_),
    .X(\rd_dout_muxed[8] ));
 sky130_fd_sc_hd__mux2_1 _211_ (.A0(\rd_dout_muxed[8] ),
    .A1(\rd_dout_additional_register[8] ),
    .S(_030_),
    .X(_099_));
 sky130_fd_sc_hd__buf_1 _212_ (.A(_099_),
    .X(net85));
 sky130_fd_sc_hd__mux2_1 _213_ (.A0(\mem_dout[9] ),
    .A1(\mem_dout[25] ),
    .S(_097_),
    .X(_100_));
 sky130_fd_sc_hd__buf_1 _214_ (.A(_100_),
    .X(\rd_dout_muxed[9] ));
 sky130_fd_sc_hd__mux2_1 _215_ (.A0(\rd_dout_muxed[9] ),
    .A1(\rd_dout_additional_register[9] ),
    .S(_030_),
    .X(_101_));
 sky130_fd_sc_hd__buf_1 _216_ (.A(_101_),
    .X(net86));
 sky130_fd_sc_hd__mux2_1 _217_ (.A0(\mem_dout[10] ),
    .A1(\mem_dout[26] ),
    .S(_097_),
    .X(_102_));
 sky130_fd_sc_hd__buf_1 _218_ (.A(_102_),
    .X(\rd_dout_muxed[10] ));
 sky130_fd_sc_hd__mux2_1 _219_ (.A0(\rd_dout_muxed[10] ),
    .A1(\rd_dout_additional_register[10] ),
    .S(_030_),
    .X(_103_));
 sky130_fd_sc_hd__buf_1 _220_ (.A(_103_),
    .X(net56));
 sky130_fd_sc_hd__mux2_1 _221_ (.A0(\mem_dout[11] ),
    .A1(\mem_dout[27] ),
    .S(_097_),
    .X(_104_));
 sky130_fd_sc_hd__buf_1 _222_ (.A(_104_),
    .X(\rd_dout_muxed[11] ));
 sky130_fd_sc_hd__clkbuf_2 _223_ (.A(_032_),
    .X(_105_));
 sky130_fd_sc_hd__mux2_1 _224_ (.A0(\rd_dout_muxed[11] ),
    .A1(\rd_dout_additional_register[11] ),
    .S(_105_),
    .X(_106_));
 sky130_fd_sc_hd__buf_1 _225_ (.A(_106_),
    .X(net57));
 sky130_fd_sc_hd__mux2_2 _226_ (.A0(\mem_dout[12] ),
    .A1(\mem_dout[28] ),
    .S(_097_),
    .X(_107_));
 sky130_fd_sc_hd__buf_1 _227_ (.A(_107_),
    .X(\rd_dout_muxed[12] ));
 sky130_fd_sc_hd__mux2_1 _228_ (.A0(\rd_dout_muxed[12] ),
    .A1(\rd_dout_additional_register[12] ),
    .S(_105_),
    .X(_108_));
 sky130_fd_sc_hd__buf_1 _229_ (.A(_108_),
    .X(net58));
 sky130_fd_sc_hd__mux2_1 _230_ (.A0(\mem_dout[13] ),
    .A1(\mem_dout[29] ),
    .S(_096_),
    .X(_109_));
 sky130_fd_sc_hd__buf_1 _231_ (.A(_109_),
    .X(\rd_dout_muxed[13] ));
 sky130_fd_sc_hd__mux2_1 _232_ (.A0(\rd_dout_muxed[13] ),
    .A1(\rd_dout_additional_register[13] ),
    .S(_105_),
    .X(_110_));
 sky130_fd_sc_hd__buf_1 _233_ (.A(_110_),
    .X(net59));
 sky130_fd_sc_hd__mux2_1 _234_ (.A0(\mem_dout[14] ),
    .A1(\mem_dout[30] ),
    .S(_096_),
    .X(_111_));
 sky130_fd_sc_hd__buf_1 _235_ (.A(_111_),
    .X(\rd_dout_muxed[14] ));
 sky130_fd_sc_hd__mux2_1 _236_ (.A0(\rd_dout_muxed[14] ),
    .A1(\rd_dout_additional_register[14] ),
    .S(_105_),
    .X(_112_));
 sky130_fd_sc_hd__buf_1 _237_ (.A(_112_),
    .X(net60));
 sky130_fd_sc_hd__mux2_1 _238_ (.A0(\mem_dout[15] ),
    .A1(\mem_dout[31] ),
    .S(_096_),
    .X(_113_));
 sky130_fd_sc_hd__buf_1 _239_ (.A(_113_),
    .X(\rd_dout_muxed[15] ));
 sky130_fd_sc_hd__mux2_1 _240_ (.A0(\rd_dout_muxed[15] ),
    .A1(\rd_dout_additional_register[15] ),
    .S(_105_),
    .X(_114_));
 sky130_fd_sc_hd__buf_1 _241_ (.A(_114_),
    .X(net61));
 sky130_fd_sc_hd__clkbuf_2 _242_ (.A(_032_),
    .X(_115_));
 sky130_fd_sc_hd__mux2_1 _243_ (.A0(\mem_dout[16] ),
    .A1(\rd_dout_additional_register[16] ),
    .S(_115_),
    .X(_116_));
 sky130_fd_sc_hd__buf_1 _244_ (.A(_116_),
    .X(net62));
 sky130_fd_sc_hd__mux2_1 _245_ (.A0(\mem_dout[17] ),
    .A1(\rd_dout_additional_register[17] ),
    .S(_115_),
    .X(_117_));
 sky130_fd_sc_hd__buf_1 _246_ (.A(_117_),
    .X(net63));
 sky130_fd_sc_hd__mux2_1 _247_ (.A0(\mem_dout[18] ),
    .A1(\rd_dout_additional_register[18] ),
    .S(_115_),
    .X(_118_));
 sky130_fd_sc_hd__clkbuf_1 _248_ (.A(_118_),
    .X(net64));
 sky130_fd_sc_hd__mux2_1 _249_ (.A0(\mem_dout[19] ),
    .A1(\rd_dout_additional_register[19] ),
    .S(_115_),
    .X(_119_));
 sky130_fd_sc_hd__clkbuf_1 _250_ (.A(_119_),
    .X(net65));
 sky130_fd_sc_hd__mux2_1 _251_ (.A0(\mem_dout[20] ),
    .A1(\rd_dout_additional_register[20] ),
    .S(_115_),
    .X(_120_));
 sky130_fd_sc_hd__buf_1 _252_ (.A(_120_),
    .X(net67));
 sky130_fd_sc_hd__clkbuf_2 _253_ (.A(net6),
    .X(_121_));
 sky130_fd_sc_hd__mux2_1 _254_ (.A0(\mem_dout[21] ),
    .A1(\rd_dout_additional_register[21] ),
    .S(_121_),
    .X(_122_));
 sky130_fd_sc_hd__buf_1 _255_ (.A(_122_),
    .X(net68));
 sky130_fd_sc_hd__mux2_1 _256_ (.A0(\mem_dout[22] ),
    .A1(\rd_dout_additional_register[22] ),
    .S(_121_),
    .X(_123_));
 sky130_fd_sc_hd__clkbuf_1 _257_ (.A(_123_),
    .X(net69));
 sky130_fd_sc_hd__mux2_1 _258_ (.A0(\mem_dout[23] ),
    .A1(\rd_dout_additional_register[23] ),
    .S(_121_),
    .X(_124_));
 sky130_fd_sc_hd__clkbuf_1 _259_ (.A(_124_),
    .X(net70));
 sky130_fd_sc_hd__mux2_1 _260_ (.A0(\mem_dout[24] ),
    .A1(\rd_dout_additional_register[24] ),
    .S(_121_),
    .X(_125_));
 sky130_fd_sc_hd__clkbuf_1 _261_ (.A(_125_),
    .X(net71));
 sky130_fd_sc_hd__mux2_1 _262_ (.A0(\mem_dout[25] ),
    .A1(\rd_dout_additional_register[25] ),
    .S(_121_),
    .X(_126_));
 sky130_fd_sc_hd__clkbuf_1 _263_ (.A(_126_),
    .X(net72));
 sky130_fd_sc_hd__clkbuf_4 _264_ (.A(net6),
    .X(_127_));
 sky130_fd_sc_hd__mux2_2 _265_ (.A0(\mem_dout[26] ),
    .A1(\rd_dout_additional_register[26] ),
    .S(_127_),
    .X(_128_));
 sky130_fd_sc_hd__buf_1 _266_ (.A(_128_),
    .X(net73));
 sky130_fd_sc_hd__mux2_2 _267_ (.A0(\mem_dout[27] ),
    .A1(\rd_dout_additional_register[27] ),
    .S(_127_),
    .X(_129_));
 sky130_fd_sc_hd__buf_1 _268_ (.A(_129_),
    .X(net74));
 sky130_fd_sc_hd__mux2_2 _269_ (.A0(\mem_dout[28] ),
    .A1(\rd_dout_additional_register[28] ),
    .S(_127_),
    .X(_130_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _270_ (.A(_130_),
    .X(net75));
 sky130_fd_sc_hd__mux2_2 _271_ (.A0(\mem_dout[29] ),
    .A1(\rd_dout_additional_register[29] ),
    .S(_127_),
    .X(_131_));
 sky130_fd_sc_hd__buf_1 _272_ (.A(_131_),
    .X(net76));
 sky130_fd_sc_hd__mux2_2 _273_ (.A0(\mem_dout[30] ),
    .A1(\rd_dout_additional_register[30] ),
    .S(_127_),
    .X(_132_));
 sky130_fd_sc_hd__buf_1 _274_ (.A(_132_),
    .X(net78));
 sky130_fd_sc_hd__mux2_1 _275_ (.A0(\mem_dout[31] ),
    .A1(\rd_dout_additional_register[31] ),
    .S(_032_),
    .X(_133_));
 sky130_fd_sc_hd__clkbuf_1 _276_ (.A(_133_),
    .X(net79));
 sky130_fd_sc_hd__clkbuf_2 _277_ (.A(net1),
    .X(_134_));
 sky130_fd_sc_hd__mux2_1 _278_ (.A0(net53),
    .A1(net23),
    .S(_134_),
    .X(_135_));
 sky130_fd_sc_hd__buf_2 _279_ (.A(_135_),
    .X(\muxedDataIn[8] ));
 sky130_fd_sc_hd__clkbuf_2 _280_ (.A(net1),
    .X(_136_));
 sky130_fd_sc_hd__mux2_1 _281_ (.A0(net54),
    .A1(net34),
    .S(_136_),
    .X(_137_));
 sky130_fd_sc_hd__buf_2 _282_ (.A(_137_),
    .X(\muxedDataIn[9] ));
 sky130_fd_sc_hd__mux2_1 _283_ (.A0(net24),
    .A1(net45),
    .S(_136_),
    .X(_138_));
 sky130_fd_sc_hd__buf_2 _284_ (.A(_138_),
    .X(\muxedDataIn[10] ));
 sky130_fd_sc_hd__mux2_1 _285_ (.A0(net25),
    .A1(net48),
    .S(_136_),
    .X(_139_));
 sky130_fd_sc_hd__buf_2 _286_ (.A(_139_),
    .X(\muxedDataIn[11] ));
 sky130_fd_sc_hd__mux2_1 _287_ (.A0(net26),
    .A1(net49),
    .S(_136_),
    .X(_140_));
 sky130_fd_sc_hd__clkbuf_4 _288_ (.A(_140_),
    .X(\muxedDataIn[12] ));
 sky130_fd_sc_hd__mux2_1 _289_ (.A0(net27),
    .A1(net50),
    .S(_136_),
    .X(_141_));
 sky130_fd_sc_hd__clkbuf_4 _290_ (.A(_141_),
    .X(\muxedDataIn[13] ));
 sky130_fd_sc_hd__mux2_1 _291_ (.A0(net28),
    .A1(net51),
    .S(net1),
    .X(_142_));
 sky130_fd_sc_hd__clkbuf_4 _292_ (.A(_142_),
    .X(\muxedDataIn[14] ));
 sky130_fd_sc_hd__mux2_1 _293_ (.A0(net29),
    .A1(net52),
    .S(net1),
    .X(_143_));
 sky130_fd_sc_hd__clkbuf_4 _294_ (.A(_143_),
    .X(\muxedDataIn[15] ));
 sky130_fd_sc_hd__clkbuf_2 _295_ (.A(net30),
    .X(_144_));
 sky130_fd_sc_hd__nor2_1 _296_ (.A(net2),
    .B(net1),
    .Y(_145_));
 sky130_fd_sc_hd__clkbuf_2 _297_ (.A(_145_),
    .X(_146_));
 sky130_fd_sc_hd__mux2_2 _298_ (.A0(net23),
    .A1(_144_),
    .S(_146_),
    .X(_147_));
 sky130_fd_sc_hd__buf_1 _299_ (.A(_147_),
    .X(\muxedDataIn[16] ));
 sky130_fd_sc_hd__clkbuf_2 _300_ (.A(net31),
    .X(_148_));
 sky130_fd_sc_hd__mux2_2 _301_ (.A0(net34),
    .A1(_148_),
    .S(_146_),
    .X(_149_));
 sky130_fd_sc_hd__buf_1 _302_ (.A(_149_),
    .X(\muxedDataIn[17] ));
 sky130_fd_sc_hd__clkbuf_2 _303_ (.A(_145_),
    .X(_150_));
 sky130_fd_sc_hd__clkbuf_2 _304_ (.A(_150_),
    .X(_151_));
 sky130_fd_sc_hd__mux2_1 _305_ (.A0(net45),
    .A1(net32),
    .S(_151_),
    .X(_152_));
 sky130_fd_sc_hd__buf_2 _306_ (.A(_152_),
    .X(\muxedDataIn[18] ));
 sky130_fd_sc_hd__mux2_1 _307_ (.A0(net48),
    .A1(net33),
    .S(_151_),
    .X(_153_));
 sky130_fd_sc_hd__buf_2 _308_ (.A(_153_),
    .X(\muxedDataIn[19] ));
 sky130_fd_sc_hd__mux2_2 _309_ (.A0(net49),
    .A1(net35),
    .S(_151_),
    .X(_154_));
 sky130_fd_sc_hd__clkbuf_2 _310_ (.A(_154_),
    .X(\muxedDataIn[20] ));
 sky130_fd_sc_hd__mux2_1 _311_ (.A0(net50),
    .A1(net36),
    .S(_151_),
    .X(_155_));
 sky130_fd_sc_hd__buf_2 _312_ (.A(_155_),
    .X(\muxedDataIn[21] ));
 sky130_fd_sc_hd__mux2_2 _313_ (.A0(net51),
    .A1(net37),
    .S(_151_),
    .X(_156_));
 sky130_fd_sc_hd__clkbuf_2 _314_ (.A(_156_),
    .X(\muxedDataIn[22] ));
 sky130_fd_sc_hd__clkbuf_2 _315_ (.A(_145_),
    .X(_157_));
 sky130_fd_sc_hd__mux2_2 _316_ (.A0(net52),
    .A1(net38),
    .S(_157_),
    .X(_158_));
 sky130_fd_sc_hd__clkbuf_2 _317_ (.A(_158_),
    .X(\muxedDataIn[23] ));
 sky130_fd_sc_hd__mux2_2 _318_ (.A0(\muxedDataIn[8] ),
    .A1(net39),
    .S(_157_),
    .X(_159_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _319_ (.A(_159_),
    .X(\muxedDataIn[24] ));
 sky130_fd_sc_hd__mux2_2 _320_ (.A0(\muxedDataIn[9] ),
    .A1(net40),
    .S(_157_),
    .X(_160_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _321_ (.A(_160_),
    .X(\muxedDataIn[25] ));
 sky130_fd_sc_hd__mux2_2 _322_ (.A0(\muxedDataIn[10] ),
    .A1(net41),
    .S(_157_),
    .X(_161_));
 sky130_fd_sc_hd__clkbuf_2 _323_ (.A(_161_),
    .X(\muxedDataIn[26] ));
 sky130_fd_sc_hd__mux2_2 _324_ (.A0(\muxedDataIn[11] ),
    .A1(net42),
    .S(_157_),
    .X(_162_));
 sky130_fd_sc_hd__clkbuf_2 _325_ (.A(_162_),
    .X(\muxedDataIn[27] ));
 sky130_fd_sc_hd__mux2_2 _326_ (.A0(\muxedDataIn[12] ),
    .A1(net43),
    .S(_150_),
    .X(_163_));
 sky130_fd_sc_hd__clkbuf_2 _327_ (.A(_163_),
    .X(\muxedDataIn[28] ));
 sky130_fd_sc_hd__mux2_2 _328_ (.A0(\muxedDataIn[13] ),
    .A1(net44),
    .S(_150_),
    .X(_164_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _329_ (.A(_164_),
    .X(\muxedDataIn[29] ));
 sky130_fd_sc_hd__mux2_2 _330_ (.A0(\muxedDataIn[14] ),
    .A1(net46),
    .S(_150_),
    .X(_165_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _331_ (.A(_165_),
    .X(\muxedDataIn[30] ));
 sky130_fd_sc_hd__mux2_4 _332_ (.A0(\muxedDataIn[15] ),
    .A1(net47),
    .S(_150_),
    .X(_166_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _333_ (.A(_166_),
    .X(\muxedDataIn[31] ));
 sky130_fd_sc_hd__o21bai_1 _334_ (.A1(_144_),
    .A2(_148_),
    .B1_N(_146_),
    .Y(_000_));
 sky130_fd_sc_hd__or2b_1 _335_ (.A(net31),
    .B_N(net30),
    .X(_167_));
 sky130_fd_sc_hd__inv_2 _336_ (.A(_134_),
    .Y(_168_));
 sky130_fd_sc_hd__o211a_1 _337_ (.A1(net30),
    .A2(_148_),
    .B1(net2),
    .C1(_168_),
    .X(_169_));
 sky130_fd_sc_hd__a21oi_1 _338_ (.A1(_134_),
    .A2(_167_),
    .B1(_169_),
    .Y(_001_));
 sky130_fd_sc_hd__nand2_1 _339_ (.A(_134_),
    .B(_144_),
    .Y(_170_));
 sky130_fd_sc_hd__o31a_1 _340_ (.A1(_144_),
    .A2(_148_),
    .A3(_146_),
    .B1(_170_),
    .X(_002_));
 sky130_fd_sc_hd__a211o_1 _341_ (.A1(_144_),
    .A2(_148_),
    .B1(_146_),
    .C1(_169_),
    .X(_003_));
 sky130_fd_sc_hd__nor2_2 _342_ (.A(net35),
    .B(net5),
    .Y(memWriteEnable));
 sky130_fd_sc_hd__and2_1 _343_ (.A(net2),
    .B(_134_),
    .X(_171_));
 sky130_fd_sc_hd__buf_1 _344_ (.A(_171_),
    .X(_004_));
 sky130_fd_sc_hd__and2b_1 _345_ (.A_N(net3),
    .B(net4),
    .X(_005_));
 sky130_fd_sc_hd__buf_1 _346_ (.A(_005_),
    .X(_006_));
 sky130_fd_sc_hd__clkbuf_2 _347_ (.A(\rd_dout_sel[0] ),
    .X(_007_));
 sky130_fd_sc_hd__clkbuf_2 _348_ (.A(_007_),
    .X(_008_));
 sky130_fd_sc_hd__mux2_1 _349_ (.A0(\mem_dout[0] ),
    .A1(\mem_dout[16] ),
    .S(_008_),
    .X(_009_));
 sky130_fd_sc_hd__and2_1 _350_ (.A(_006_),
    .B(_009_),
    .X(_010_));
 sky130_fd_sc_hd__clkbuf_2 _351_ (.A(net4),
    .X(_011_));
 sky130_fd_sc_hd__clkbuf_2 _352_ (.A(\rd_dout_sel[0] ),
    .X(_012_));
 sky130_fd_sc_hd__clkbuf_2 _353_ (.A(\rd_dout_sel[1] ),
    .X(_013_));
 sky130_fd_sc_hd__o21ai_4 _354_ (.A1(_012_),
    .A2(_013_),
    .B1(net3),
    .Y(_014_));
 sky130_fd_sc_hd__nor2_1 _355_ (.A(_011_),
    .B(_014_),
    .Y(_015_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _356_ (.A(_015_),
    .X(_016_));
 sky130_fd_sc_hd__and2b_1 _357_ (.A_N(\rd_dout_sel[1] ),
    .B(\rd_dout_sel[0] ),
    .X(_017_));
 sky130_fd_sc_hd__a211o_1 _358_ (.A1(\mem_dout[8] ),
    .A2(_017_),
    .B1(_014_),
    .C1(_011_),
    .X(_018_));
 sky130_fd_sc_hd__and2b_1 _359_ (.A_N(\rd_dout_sel[0] ),
    .B(\rd_dout_sel[1] ),
    .X(_019_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _360_ (.A(_019_),
    .X(_020_));
 sky130_fd_sc_hd__buf_1 _361_ (.A(\rd_dout_sel[1] ),
    .X(_021_));
 sky130_fd_sc_hd__or3b_1 _362_ (.A(\mem_dout[16] ),
    .B(_007_),
    .C_N(_021_),
    .X(_022_));
 sky130_fd_sc_hd__or2b_1 _363_ (.A(_013_),
    .B_N(_012_),
    .X(_023_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _364_ (.A(_023_),
    .X(_024_));
 sky130_fd_sc_hd__o211a_1 _365_ (.A1(\mem_dout[24] ),
    .A2(_020_),
    .B1(_022_),
    .C1(_024_),
    .X(_025_));
 sky130_fd_sc_hd__or2b_2 _366_ (.A(net3),
    .B_N(_011_),
    .X(_026_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _367_ (.A(_026_),
    .X(_027_));
 sky130_fd_sc_hd__o221a_2 _368_ (.A1(\mem_dout[0] ),
    .A2(_016_),
    .B1(_018_),
    .B2(_025_),
    .C1(_027_),
    .X(_028_));
 sky130_fd_sc_hd__or2_1 _369_ (.A(_010_),
    .B(_028_),
    .X(_029_));
 sky130_fd_sc_hd__clkbuf_1 _370_ (.A(_029_),
    .X(\rd_dout_muxed[0] ));
 sky130_fd_sc_hd__clkbuf_2 _371_ (.A(net6),
    .X(_030_));
 sky130_fd_sc_hd__buf_1 _372_ (.A(_030_),
    .X(_031_));
 sky130_fd_sc_hd__clkbuf_2 _373_ (.A(net6),
    .X(_032_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _374_ (.A(_032_),
    .X(_033_));
 sky130_fd_sc_hd__or2b_1 _375_ (.A(\rd_dout_additional_register[0] ),
    .B_N(_033_),
    .X(_034_));
 sky130_fd_sc_hd__o31a_1 _376_ (.A1(_031_),
    .A2(_010_),
    .A3(_028_),
    .B1(_034_),
    .X(net55));
 sky130_fd_sc_hd__mux2_1 _377_ (.A0(\mem_dout[1] ),
    .A1(\mem_dout[17] ),
    .S(_008_),
    .X(_035_));
 sky130_fd_sc_hd__and2_1 _378_ (.A(_006_),
    .B(_035_),
    .X(_036_));
 sky130_fd_sc_hd__buf_1 _379_ (.A(\rd_dout_sel[0] ),
    .X(_037_));
 sky130_fd_sc_hd__or3b_1 _380_ (.A(_037_),
    .B(\mem_dout[17] ),
    .C_N(_021_),
    .X(_038_));
 sky130_fd_sc_hd__o211a_1 _381_ (.A1(\mem_dout[25] ),
    .A2(_020_),
    .B1(_038_),
    .C1(_024_),
    .X(_039_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _382_ (.A(_017_),
    .X(_040_));
 sky130_fd_sc_hd__dlymetal6s2s_1 _383_ (.A(_014_),
    .X(_041_));
 sky130_fd_sc_hd__clkbuf_2 _384_ (.A(net4),
    .X(_042_));
 sky130_fd_sc_hd__a211o_1 _385_ (.A1(\mem_dout[9] ),
    .A2(_040_),
    .B1(_041_),
    .C1(_042_),
    .X(_043_));
 sky130_fd_sc_hd__o221a_2 _386_ (.A1(\mem_dout[1] ),
    .A2(_016_),
    .B1(_039_),
    .B2(_043_),
    .C1(_027_),
    .X(_044_));
 sky130_fd_sc_hd__or2_1 _387_ (.A(_036_),
    .B(_044_),
    .X(_045_));
 sky130_fd_sc_hd__clkbuf_1 _388_ (.A(_045_),
    .X(\rd_dout_muxed[1] ));
 sky130_fd_sc_hd__or2b_1 _389_ (.A(\rd_dout_additional_register[1] ),
    .B_N(_033_),
    .X(_046_));
 sky130_fd_sc_hd__o31a_1 _390_ (.A1(_031_),
    .A2(_036_),
    .A3(_044_),
    .B1(_046_),
    .X(net66));
 sky130_fd_sc_hd__mux2_1 _391_ (.A0(\mem_dout[2] ),
    .A1(\mem_dout[18] ),
    .S(_008_),
    .X(_047_));
 sky130_fd_sc_hd__and2_1 _392_ (.A(_006_),
    .B(_047_),
    .X(_048_));
 sky130_fd_sc_hd__or3b_1 _393_ (.A(_037_),
    .B(\mem_dout[18] ),
    .C_N(_021_),
    .X(_049_));
 sky130_fd_sc_hd__o211a_1 _394_ (.A1(\mem_dout[26] ),
    .A2(_020_),
    .B1(_049_),
    .C1(_024_),
    .X(_050_));
 sky130_fd_sc_hd__a211o_1 _395_ (.A1(\mem_dout[10] ),
    .A2(_040_),
    .B1(_041_),
    .C1(_042_),
    .X(_051_));
 sky130_fd_sc_hd__o221a_2 _396_ (.A1(\mem_dout[2] ),
    .A2(_016_),
    .B1(_050_),
    .B2(_051_),
    .C1(_027_),
    .X(_052_));
 sky130_fd_sc_hd__or2_1 _397_ (.A(_048_),
    .B(_052_),
    .X(_053_));
 sky130_fd_sc_hd__clkbuf_1 _398_ (.A(_053_),
    .X(\rd_dout_muxed[2] ));
 sky130_fd_sc_hd__buf_1 _399_ (.A(_032_),
    .X(_054_));
 sky130_fd_sc_hd__or2b_1 _400_ (.A(\rd_dout_additional_register[2] ),
    .B_N(_054_),
    .X(_055_));
 sky130_fd_sc_hd__o31a_1 _401_ (.A1(_031_),
    .A2(_048_),
    .A3(_052_),
    .B1(_055_),
    .X(net77));
 sky130_fd_sc_hd__mux2_1 _402_ (.A0(\mem_dout[3] ),
    .A1(\mem_dout[19] ),
    .S(_008_),
    .X(_056_));
 sky130_fd_sc_hd__and2_1 _403_ (.A(_006_),
    .B(_056_),
    .X(_057_));
 sky130_fd_sc_hd__or3b_1 _404_ (.A(_037_),
    .B(\mem_dout[19] ),
    .C_N(_021_),
    .X(_058_));
 sky130_fd_sc_hd__o211a_1 _405_ (.A1(\mem_dout[27] ),
    .A2(_020_),
    .B1(_058_),
    .C1(_024_),
    .X(_059_));
 sky130_fd_sc_hd__a211o_1 _406_ (.A1(\mem_dout[11] ),
    .A2(_040_),
    .B1(_041_),
    .C1(_042_),
    .X(_060_));
 sky130_fd_sc_hd__o221a_2 _407_ (.A1(\mem_dout[3] ),
    .A2(_016_),
    .B1(_059_),
    .B2(_060_),
    .C1(_027_),
    .X(_061_));
 sky130_fd_sc_hd__or2_1 _408_ (.A(_057_),
    .B(_061_),
    .X(_062_));
 sky130_fd_sc_hd__clkbuf_1 _409_ (.A(_062_),
    .X(\rd_dout_muxed[3] ));
 sky130_fd_sc_hd__or2b_1 _410_ (.A(\rd_dout_additional_register[3] ),
    .B_N(_054_),
    .X(_063_));
 sky130_fd_sc_hd__o31a_1 _411_ (.A1(_031_),
    .A2(_057_),
    .A3(_061_),
    .B1(_063_),
    .X(net80));
 sky130_fd_sc_hd__mux2_1 _412_ (.A0(\mem_dout[4] ),
    .A1(\mem_dout[20] ),
    .S(_008_),
    .X(_064_));
 sky130_fd_sc_hd__and2_1 _413_ (.A(_006_),
    .B(_064_),
    .X(_065_));
 sky130_fd_sc_hd__or3b_1 _414_ (.A(_037_),
    .B(\mem_dout[20] ),
    .C_N(_021_),
    .X(_066_));
 sky130_fd_sc_hd__o211a_1 _415_ (.A1(\mem_dout[28] ),
    .A2(_020_),
    .B1(_066_),
    .C1(_024_),
    .X(_067_));
 sky130_fd_sc_hd__a211o_1 _416_ (.A1(\mem_dout[12] ),
    .A2(_040_),
    .B1(_041_),
    .C1(_042_),
    .X(_068_));
 sky130_fd_sc_hd__o221a_2 _417_ (.A1(\mem_dout[4] ),
    .A2(_016_),
    .B1(_067_),
    .B2(_068_),
    .C1(_027_),
    .X(_069_));
 sky130_fd_sc_hd__dlxtn_1 _418_ (.D(_000_),
    .GATE_N(_004_),
    .Q(\mem_wr_mask[0] ));
 sky130_fd_sc_hd__dlxtn_1 _419_ (.D(_001_),
    .GATE_N(_004_),
    .Q(\mem_wr_mask[1] ));
 sky130_fd_sc_hd__dlxtn_1 _420_ (.D(_002_),
    .GATE_N(_004_),
    .Q(\mem_wr_mask[2] ));
 sky130_fd_sc_hd__dlxtn_1 _421_ (.D(_003_),
    .GATE_N(_004_),
    .Q(\mem_wr_mask[3] ));
 sky130_fd_sc_hd__dfxtp_1 _422_ (.CLK(clknet_2_1__leaf_clk),
    .D(\rd_dout_muxed[0] ),
    .Q(\rd_dout_additional_register[0] ));
 sky130_fd_sc_hd__dfxtp_1 _423_ (.CLK(clknet_2_1__leaf_clk),
    .D(\rd_dout_muxed[1] ),
    .Q(\rd_dout_additional_register[1] ));
 sky130_fd_sc_hd__dfxtp_1 _424_ (.CLK(clknet_2_1__leaf_clk),
    .D(\rd_dout_muxed[2] ),
    .Q(\rd_dout_additional_register[2] ));
 sky130_fd_sc_hd__dfxtp_1 _425_ (.CLK(clknet_2_1__leaf_clk),
    .D(\rd_dout_muxed[3] ),
    .Q(\rd_dout_additional_register[3] ));
 sky130_fd_sc_hd__dfxtp_1 _426_ (.CLK(clknet_2_1__leaf_clk),
    .D(\rd_dout_muxed[4] ),
    .Q(\rd_dout_additional_register[4] ));
 sky130_fd_sc_hd__dfxtp_1 _427_ (.CLK(clknet_2_1__leaf_clk),
    .D(\rd_dout_muxed[5] ),
    .Q(\rd_dout_additional_register[5] ));
 sky130_fd_sc_hd__dfxtp_1 _428_ (.CLK(clknet_2_1__leaf_clk),
    .D(\rd_dout_muxed[6] ),
    .Q(\rd_dout_additional_register[6] ));
 sky130_fd_sc_hd__dfxtp_1 _429_ (.CLK(clknet_2_1__leaf_clk),
    .D(\rd_dout_muxed[7] ),
    .Q(\rd_dout_additional_register[7] ));
 sky130_fd_sc_hd__dfxtp_1 _430_ (.CLK(clknet_2_0__leaf_clk),
    .D(\rd_dout_muxed[8] ),
    .Q(\rd_dout_additional_register[8] ));
 sky130_fd_sc_hd__dfxtp_1 _431_ (.CLK(clknet_2_0__leaf_clk),
    .D(\rd_dout_muxed[9] ),
    .Q(\rd_dout_additional_register[9] ));
 sky130_fd_sc_hd__dfxtp_1 _432_ (.CLK(clknet_2_1__leaf_clk),
    .D(\rd_dout_muxed[10] ),
    .Q(\rd_dout_additional_register[10] ));
 sky130_fd_sc_hd__dfxtp_1 _433_ (.CLK(clknet_2_1__leaf_clk),
    .D(\rd_dout_muxed[11] ),
    .Q(\rd_dout_additional_register[11] ));
 sky130_fd_sc_hd__dfxtp_1 _434_ (.CLK(clknet_2_0__leaf_clk),
    .D(\rd_dout_muxed[12] ),
    .Q(\rd_dout_additional_register[12] ));
 sky130_fd_sc_hd__dfxtp_1 _435_ (.CLK(clknet_2_0__leaf_clk),
    .D(\rd_dout_muxed[13] ),
    .Q(\rd_dout_additional_register[13] ));
 sky130_fd_sc_hd__dfxtp_1 _436_ (.CLK(clknet_2_0__leaf_clk),
    .D(\rd_dout_muxed[14] ),
    .Q(\rd_dout_additional_register[14] ));
 sky130_fd_sc_hd__dfxtp_1 _437_ (.CLK(clknet_2_0__leaf_clk),
    .D(\rd_dout_muxed[15] ),
    .Q(\rd_dout_additional_register[15] ));
 sky130_fd_sc_hd__dfxtp_1 _438_ (.CLK(clknet_2_2__leaf_clk),
    .D(\mem_dout[16] ),
    .Q(\rd_dout_additional_register[16] ));
 sky130_fd_sc_hd__dfxtp_1 _439_ (.CLK(clknet_2_2__leaf_clk),
    .D(\mem_dout[17] ),
    .Q(\rd_dout_additional_register[17] ));
 sky130_fd_sc_hd__dfxtp_1 _440_ (.CLK(clknet_2_2__leaf_clk),
    .D(\mem_dout[18] ),
    .Q(\rd_dout_additional_register[18] ));
 sky130_fd_sc_hd__dfxtp_1 _441_ (.CLK(clknet_2_2__leaf_clk),
    .D(\mem_dout[19] ),
    .Q(\rd_dout_additional_register[19] ));
 sky130_fd_sc_hd__dfxtp_1 _442_ (.CLK(clknet_2_2__leaf_clk),
    .D(\mem_dout[20] ),
    .Q(\rd_dout_additional_register[20] ));
 sky130_fd_sc_hd__dfxtp_1 _443_ (.CLK(clknet_2_2__leaf_clk),
    .D(\mem_dout[21] ),
    .Q(\rd_dout_additional_register[21] ));
 sky130_fd_sc_hd__dfxtp_1 _444_ (.CLK(clknet_2_2__leaf_clk),
    .D(\mem_dout[22] ),
    .Q(\rd_dout_additional_register[22] ));
 sky130_fd_sc_hd__dfxtp_1 _445_ (.CLK(clknet_2_2__leaf_clk),
    .D(\mem_dout[23] ),
    .Q(\rd_dout_additional_register[23] ));
 sky130_fd_sc_hd__dfxtp_1 _446_ (.CLK(clknet_2_2__leaf_clk),
    .D(\mem_dout[24] ),
    .Q(\rd_dout_additional_register[24] ));
 sky130_fd_sc_hd__dfxtp_1 _447_ (.CLK(clknet_2_3__leaf_clk),
    .D(\mem_dout[25] ),
    .Q(\rd_dout_additional_register[25] ));
 sky130_fd_sc_hd__dfxtp_1 _448_ (.CLK(clknet_2_3__leaf_clk),
    .D(\mem_dout[26] ),
    .Q(\rd_dout_additional_register[26] ));
 sky130_fd_sc_hd__dfxtp_1 _449_ (.CLK(clknet_2_3__leaf_clk),
    .D(\mem_dout[27] ),
    .Q(\rd_dout_additional_register[27] ));
 sky130_fd_sc_hd__dfxtp_1 _450_ (.CLK(clknet_2_3__leaf_clk),
    .D(\mem_dout[28] ),
    .Q(\rd_dout_additional_register[28] ));
 sky130_fd_sc_hd__dfxtp_1 _451_ (.CLK(clknet_2_3__leaf_clk),
    .D(\mem_dout[29] ),
    .Q(\rd_dout_additional_register[29] ));
 sky130_fd_sc_hd__dfxtp_1 _452_ (.CLK(clknet_2_3__leaf_clk),
    .D(\mem_dout[30] ),
    .Q(\rd_dout_additional_register[30] ));
 sky130_fd_sc_hd__dfxtp_1 _453_ (.CLK(clknet_2_2__leaf_clk),
    .D(\mem_dout[31] ),
    .Q(\rd_dout_additional_register[31] ));
 sky130_fd_sc_hd__dfxtp_1 _454_ (.CLK(clknet_2_2__leaf_clk),
    .D(net39),
    .Q(\rd_dout_sel[0] ));
 sky130_fd_sc_hd__dfxtp_1 _455_ (.CLK(clknet_2_2__leaf_clk),
    .D(net40),
    .Q(\rd_dout_sel[1] ));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_clk (.A(clk),
    .X(clknet_0_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_0__f_clk (.A(clknet_0_clk),
    .X(clknet_2_0__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_1__f_clk (.A(clknet_0_clk),
    .X(clknet_2_1__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_2__f_clk (.A(clknet_0_clk),
    .X(clknet_2_2__leaf_clk));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_2_3__f_clk (.A(clknet_0_clk),
    .X(clknet_2_3__leaf_clk));
 sky130_fd_sc_hd__clkbuf_2 input1 (.A(C0),
    .X(net1));
 sky130_fd_sc_hd__buf_4 input10 (.A(rd_addr[3]),
    .X(net10));
 sky130_fd_sc_hd__buf_4 input11 (.A(rd_addr[4]),
    .X(net11));
 sky130_fd_sc_hd__buf_4 input12 (.A(rd_addr[5]),
    .X(net12));
 sky130_fd_sc_hd__buf_4 input13 (.A(rd_addr[6]),
    .X(net13));
 sky130_fd_sc_hd__buf_4 input14 (.A(rd_addr[7]),
    .X(net14));
 sky130_fd_sc_hd__clkbuf_4 input15 (.A(wr_addr[0]),
    .X(net15));
 sky130_fd_sc_hd__clkbuf_2 input16 (.A(wr_addr[1]),
    .X(net16));
 sky130_fd_sc_hd__clkbuf_2 input17 (.A(wr_addr[2]),
    .X(net17));
 sky130_fd_sc_hd__clkbuf_2 input18 (.A(wr_addr[3]),
    .X(net18));
 sky130_fd_sc_hd__clkbuf_2 input19 (.A(wr_addr[4]),
    .X(net19));
 sky130_fd_sc_hd__buf_1 input2 (.A(C1),
    .X(net2));
 sky130_fd_sc_hd__clkbuf_2 input20 (.A(wr_addr[5]),
    .X(net20));
 sky130_fd_sc_hd__clkbuf_2 input21 (.A(wr_addr[6]),
    .X(net21));
 sky130_fd_sc_hd__clkbuf_2 input22 (.A(wr_addr[7]),
    .X(net22));
 sky130_fd_sc_hd__clkbuf_4 input23 (.A(wr_data[0]),
    .X(net23));
 sky130_fd_sc_hd__clkbuf_1 input24 (.A(wr_data[10]),
    .X(net24));
 sky130_fd_sc_hd__clkbuf_1 input25 (.A(wr_data[11]),
    .X(net25));
 sky130_fd_sc_hd__clkbuf_1 input26 (.A(wr_data[12]),
    .X(net26));
 sky130_fd_sc_hd__clkbuf_1 input27 (.A(wr_data[13]),
    .X(net27));
 sky130_fd_sc_hd__buf_1 input28 (.A(wr_data[14]),
    .X(net28));
 sky130_fd_sc_hd__buf_1 input29 (.A(wr_data[15]),
    .X(net29));
 sky130_fd_sc_hd__buf_2 input3 (.A(C2),
    .X(net3));
 sky130_fd_sc_hd__buf_2 input30 (.A(wr_data[16]),
    .X(net30));
 sky130_fd_sc_hd__clkbuf_2 input31 (.A(wr_data[17]),
    .X(net31));
 sky130_fd_sc_hd__clkbuf_2 input32 (.A(wr_data[18]),
    .X(net32));
 sky130_fd_sc_hd__clkbuf_2 input33 (.A(wr_data[19]),
    .X(net33));
 sky130_fd_sc_hd__clkbuf_4 input34 (.A(wr_data[1]),
    .X(net34));
 sky130_fd_sc_hd__buf_2 input35 (.A(wr_data[20]),
    .X(net35));
 sky130_fd_sc_hd__clkbuf_2 input36 (.A(wr_data[21]),
    .X(net36));
 sky130_fd_sc_hd__clkbuf_2 input37 (.A(wr_data[22]),
    .X(net37));
 sky130_fd_sc_hd__clkbuf_2 input38 (.A(wr_data[23]),
    .X(net38));
 sky130_fd_sc_hd__buf_2 input39 (.A(wr_data[24]),
    .X(net39));
 sky130_fd_sc_hd__clkbuf_2 input4 (.A(C3),
    .X(net4));
 sky130_fd_sc_hd__buf_2 input40 (.A(wr_data[25]),
    .X(net40));
 sky130_fd_sc_hd__clkbuf_2 input41 (.A(wr_data[26]),
    .X(net41));
 sky130_fd_sc_hd__clkbuf_2 input42 (.A(wr_data[27]),
    .X(net42));
 sky130_fd_sc_hd__clkbuf_2 input43 (.A(wr_data[28]),
    .X(net43));
 sky130_fd_sc_hd__clkbuf_2 input44 (.A(wr_data[29]),
    .X(net44));
 sky130_fd_sc_hd__clkbuf_4 input45 (.A(wr_data[2]),
    .X(net45));
 sky130_fd_sc_hd__clkbuf_2 input46 (.A(wr_data[30]),
    .X(net46));
 sky130_fd_sc_hd__clkbuf_2 input47 (.A(wr_data[31]),
    .X(net47));
 sky130_fd_sc_hd__clkbuf_4 input48 (.A(wr_data[3]),
    .X(net48));
 sky130_fd_sc_hd__clkbuf_4 input49 (.A(wr_data[4]),
    .X(net49));
 sky130_fd_sc_hd__buf_1 input5 (.A(C4),
    .X(net5));
 sky130_fd_sc_hd__clkbuf_4 input50 (.A(wr_data[5]),
    .X(net50));
 sky130_fd_sc_hd__clkbuf_4 input51 (.A(wr_data[6]),
    .X(net51));
 sky130_fd_sc_hd__clkbuf_4 input52 (.A(wr_data[7]),
    .X(net52));
 sky130_fd_sc_hd__buf_1 input53 (.A(wr_data[8]),
    .X(net53));
 sky130_fd_sc_hd__buf_1 input54 (.A(wr_data[9]),
    .X(net54));
 sky130_fd_sc_hd__clkbuf_2 input6 (.A(C5),
    .X(net6));
 sky130_fd_sc_hd__clkbuf_8 input7 (.A(rd_addr[0]),
    .X(net7));
 sky130_fd_sc_hd__buf_4 input8 (.A(rd_addr[1]),
    .X(net8));
 sky130_fd_sc_hd__buf_4 input9 (.A(rd_addr[2]),
    .X(net9));
 sky130_sram_1kbyte_1rw1r_32x256_8 memory_cell (.csb0(memWriteEnable),
    .csb1(net87),
    .web0(memWriteEnable),
    .clk0(clknet_2_0__leaf_clk),
    .clk1(clknet_2_3__leaf_clk),
    .addr0({net22,
    net21,
    net20,
    net19,
    net18,
    net17,
    net16,
    net15}),
    .addr1({net14,
    net13,
    net12,
    net11,
    net10,
    net9,
    net8,
    net7}),
    .din0({\muxedDataIn[31] ,
    \muxedDataIn[30] ,
    \muxedDataIn[29] ,
    \muxedDataIn[28] ,
    \muxedDataIn[27] ,
    \muxedDataIn[26] ,
    \muxedDataIn[25] ,
    \muxedDataIn[24] ,
    \muxedDataIn[23] ,
    \muxedDataIn[22] ,
    \muxedDataIn[21] ,
    \muxedDataIn[20] ,
    \muxedDataIn[19] ,
    \muxedDataIn[18] ,
    \muxedDataIn[17] ,
    \muxedDataIn[16] ,
    \muxedDataIn[15] ,
    \muxedDataIn[14] ,
    \muxedDataIn[13] ,
    \muxedDataIn[12] ,
    \muxedDataIn[11] ,
    \muxedDataIn[10] ,
    \muxedDataIn[9] ,
    \muxedDataIn[8] ,
    net52,
    net51,
    net50,
    net49,
    net48,
    net45,
    net34,
    net23}),
    .dout0({_NC1,
    _NC2,
    _NC3,
    _NC4,
    _NC5,
    _NC6,
    _NC7,
    _NC8,
    _NC9,
    _NC10,
    _NC11,
    _NC12,
    _NC13,
    _NC14,
    _NC15,
    _NC16,
    _NC17,
    _NC18,
    _NC19,
    _NC20,
    _NC21,
    _NC22,
    _NC23,
    _NC24,
    _NC25,
    _NC26,
    _NC27,
    _NC28,
    _NC29,
    _NC30,
    _NC31,
    _NC32}),
    .dout1({\mem_dout[31] ,
    \mem_dout[30] ,
    \mem_dout[29] ,
    \mem_dout[28] ,
    \mem_dout[27] ,
    \mem_dout[26] ,
    \mem_dout[25] ,
    \mem_dout[24] ,
    \mem_dout[23] ,
    \mem_dout[22] ,
    \mem_dout[21] ,
    \mem_dout[20] ,
    \mem_dout[19] ,
    \mem_dout[18] ,
    \mem_dout[17] ,
    \mem_dout[16] ,
    \mem_dout[15] ,
    \mem_dout[14] ,
    \mem_dout[13] ,
    \mem_dout[12] ,
    \mem_dout[11] ,
    \mem_dout[10] ,
    \mem_dout[9] ,
    \mem_dout[8] ,
    \mem_dout[7] ,
    \mem_dout[6] ,
    \mem_dout[5] ,
    \mem_dout[4] ,
    \mem_dout[3] ,
    \mem_dout[2] ,
    \mem_dout[1] ,
    \mem_dout[0] }),
    .wmask0({\mem_wr_mask[3] ,
    \mem_wr_mask[2] ,
    \mem_wr_mask[1] ,
    \mem_wr_mask[0] }));
 sky130_fd_sc_hd__conb_1 memory_cell_87 (.LO(net87));
 sky130_fd_sc_hd__clkbuf_4 output55 (.A(net55),
    .X(rd_data[0]));
 sky130_fd_sc_hd__clkbuf_4 output56 (.A(net56),
    .X(rd_data[10]));
 sky130_fd_sc_hd__clkbuf_4 output57 (.A(net57),
    .X(rd_data[11]));
 sky130_fd_sc_hd__clkbuf_4 output58 (.A(net58),
    .X(rd_data[12]));
 sky130_fd_sc_hd__clkbuf_4 output59 (.A(net59),
    .X(rd_data[13]));
 sky130_fd_sc_hd__clkbuf_4 output60 (.A(net60),
    .X(rd_data[14]));
 sky130_fd_sc_hd__clkbuf_4 output61 (.A(net61),
    .X(rd_data[15]));
 sky130_fd_sc_hd__clkbuf_4 output62 (.A(net62),
    .X(rd_data[16]));
 sky130_fd_sc_hd__clkbuf_4 output63 (.A(net63),
    .X(rd_data[17]));
 sky130_fd_sc_hd__clkbuf_4 output64 (.A(net64),
    .X(rd_data[18]));
 sky130_fd_sc_hd__clkbuf_4 output65 (.A(net65),
    .X(rd_data[19]));
 sky130_fd_sc_hd__clkbuf_4 output66 (.A(net66),
    .X(rd_data[1]));
 sky130_fd_sc_hd__clkbuf_4 output67 (.A(net67),
    .X(rd_data[20]));
 sky130_fd_sc_hd__clkbuf_4 output68 (.A(net68),
    .X(rd_data[21]));
 sky130_fd_sc_hd__clkbuf_4 output69 (.A(net69),
    .X(rd_data[22]));
 sky130_fd_sc_hd__clkbuf_4 output70 (.A(net70),
    .X(rd_data[23]));
 sky130_fd_sc_hd__clkbuf_4 output71 (.A(net71),
    .X(rd_data[24]));
 sky130_fd_sc_hd__clkbuf_4 output72 (.A(net72),
    .X(rd_data[25]));
 sky130_fd_sc_hd__clkbuf_4 output73 (.A(net73),
    .X(rd_data[26]));
 sky130_fd_sc_hd__clkbuf_4 output74 (.A(net74),
    .X(rd_data[27]));
 sky130_fd_sc_hd__clkbuf_4 output75 (.A(net75),
    .X(rd_data[28]));
 sky130_fd_sc_hd__clkbuf_4 output76 (.A(net76),
    .X(rd_data[29]));
 sky130_fd_sc_hd__clkbuf_4 output77 (.A(net77),
    .X(rd_data[2]));
 sky130_fd_sc_hd__clkbuf_4 output78 (.A(net78),
    .X(rd_data[30]));
 sky130_fd_sc_hd__clkbuf_4 output79 (.A(net79),
    .X(rd_data[31]));
 sky130_fd_sc_hd__clkbuf_4 output80 (.A(net80),
    .X(rd_data[3]));
 sky130_fd_sc_hd__clkbuf_4 output81 (.A(net81),
    .X(rd_data[4]));
 sky130_fd_sc_hd__clkbuf_4 output82 (.A(net82),
    .X(rd_data[5]));
 sky130_fd_sc_hd__clkbuf_4 output83 (.A(net83),
    .X(rd_data[6]));
 sky130_fd_sc_hd__clkbuf_4 output84 (.A(net84),
    .X(rd_data[7]));
 sky130_fd_sc_hd__clkbuf_4 output85 (.A(net85),
    .X(rd_data[8]));
 sky130_fd_sc_hd__clkbuf_4 output86 (.A(net86),
    .X(rd_data[9]));
endmodule

