magic
tech sky130A
magscale 1 2
timestamp 1733619021
<< viali >>
rect 2053 8585 2087 8619
rect 2789 8585 2823 8619
rect 3157 8585 3191 8619
rect 4261 8585 4295 8619
rect 4629 8585 4663 8619
rect 5181 8585 5215 8619
rect 5733 8585 5767 8619
rect 6101 8585 6135 8619
rect 6837 8585 6871 8619
rect 7389 8585 7423 8619
rect 7757 8585 7791 8619
rect 8309 8585 8343 8619
rect 8677 8585 8711 8619
rect 9321 8585 9355 8619
rect 9689 8585 9723 8619
rect 10241 8585 10275 8619
rect 13185 8585 13219 8619
rect 13737 8585 13771 8619
rect 14565 8585 14599 8619
rect 14841 8585 14875 8619
rect 16681 8585 16715 8619
rect 16957 8585 16991 8619
rect 17233 8585 17267 8619
rect 17509 8585 17543 8619
rect 17785 8585 17819 8619
rect 18245 8585 18279 8619
rect 18337 8585 18371 8619
rect 20269 8585 20303 8619
rect 20637 8585 20671 8619
rect 22017 8585 22051 8619
rect 22569 8585 22603 8619
rect 23673 8585 23707 8619
rect 3985 8517 4019 8551
rect 6561 8517 6595 8551
rect 8033 8517 8067 8551
rect 9597 8517 9631 8551
rect 10149 8517 10183 8551
rect 20545 8517 20579 8551
rect 1501 8449 1535 8483
rect 1961 8449 1995 8483
rect 2513 8449 2547 8483
rect 3065 8449 3099 8483
rect 4445 8449 4479 8483
rect 4905 8449 4939 8483
rect 5457 8449 5491 8483
rect 5917 8449 5951 8483
rect 7205 8449 7239 8483
rect 7573 8449 7607 8483
rect 8493 8449 8527 8483
rect 9137 8449 9171 8483
rect 10793 8449 10827 8483
rect 11069 8449 11103 8483
rect 11345 8449 11379 8483
rect 11713 8449 11747 8483
rect 11989 8449 12023 8483
rect 12265 8449 12299 8483
rect 12541 8449 12575 8483
rect 12633 8449 12667 8483
rect 12909 8449 12943 8483
rect 13369 8449 13403 8483
rect 13461 8449 13495 8483
rect 13921 8449 13955 8483
rect 14289 8449 14323 8483
rect 14381 8449 14415 8483
rect 14657 8449 14691 8483
rect 15117 8449 15151 8483
rect 15209 8449 15243 8483
rect 15485 8449 15519 8483
rect 15761 8449 15795 8483
rect 16221 8449 16255 8483
rect 16497 8449 16531 8483
rect 16865 8449 16899 8483
rect 17141 8449 17175 8483
rect 17417 8449 17451 8483
rect 17693 8449 17727 8483
rect 17969 8449 18003 8483
rect 18061 8449 18095 8483
rect 18521 8449 18555 8483
rect 18613 8449 18647 8483
rect 18889 8449 18923 8483
rect 19441 8449 19475 8483
rect 19717 8449 19751 8483
rect 19809 8449 19843 8483
rect 20085 8449 20119 8483
rect 21097 8449 21131 8483
rect 21925 8449 21959 8483
rect 22477 8449 22511 8483
rect 23029 8449 23063 8483
rect 23581 8449 23615 8483
rect 1685 8313 1719 8347
rect 10609 8313 10643 8347
rect 10885 8313 10919 8347
rect 11161 8313 11195 8347
rect 11529 8313 11563 8347
rect 12357 8313 12391 8347
rect 12817 8313 12851 8347
rect 13093 8313 13127 8347
rect 13645 8313 13679 8347
rect 14105 8313 14139 8347
rect 14933 8313 14967 8347
rect 16313 8313 16347 8347
rect 18797 8313 18831 8347
rect 19073 8313 19107 8347
rect 19257 8313 19291 8347
rect 19993 8313 20027 8347
rect 21281 8313 21315 8347
rect 23213 8313 23247 8347
rect 11805 8245 11839 8279
rect 12081 8245 12115 8279
rect 15393 8245 15427 8279
rect 15669 8245 15703 8279
rect 15945 8245 15979 8279
rect 16037 8245 16071 8279
rect 19533 8245 19567 8279
rect 1777 8041 1811 8075
rect 2329 8041 2363 8075
rect 3249 8041 3283 8075
rect 4629 8041 4663 8075
rect 5181 8041 5215 8075
rect 5733 8041 5767 8075
rect 6285 8041 6319 8075
rect 7389 8041 7423 8075
rect 7941 8041 7975 8075
rect 8677 8041 8711 8075
rect 9321 8041 9355 8075
rect 9597 8041 9631 8075
rect 11253 8041 11287 8075
rect 12357 8041 12391 8075
rect 12633 8041 12667 8075
rect 12909 8041 12943 8075
rect 13185 8041 13219 8075
rect 14565 8041 14599 8075
rect 14841 8041 14875 8075
rect 15393 8041 15427 8075
rect 15669 8041 15703 8075
rect 16221 8041 16255 8075
rect 18153 8041 18187 8075
rect 21281 8041 21315 8075
rect 22201 8041 22235 8075
rect 22753 8041 22787 8075
rect 23489 8041 23523 8075
rect 23857 8041 23891 8075
rect 2789 7973 2823 8007
rect 4169 7973 4203 8007
rect 6929 7973 6963 8007
rect 9045 7973 9079 8007
rect 10701 7973 10735 8007
rect 10977 7973 11011 8007
rect 12081 7973 12115 8007
rect 15117 7973 15151 8007
rect 15945 7973 15979 8007
rect 19257 7973 19291 8007
rect 1501 7837 1535 7871
rect 2605 7837 2639 7871
rect 3157 7837 3191 7871
rect 4997 7837 5031 7871
rect 7205 7837 7239 7871
rect 8493 7837 8527 7871
rect 9229 7837 9263 7871
rect 9505 7837 9539 7871
rect 9781 7837 9815 7871
rect 9873 7837 9907 7871
rect 10333 7837 10367 7871
rect 10609 7837 10643 7871
rect 10885 7837 10919 7871
rect 11161 7837 11195 7871
rect 11437 7837 11471 7871
rect 11713 7837 11747 7871
rect 12265 7837 12299 7871
rect 12541 7837 12575 7871
rect 12817 7837 12851 7871
rect 13093 7837 13127 7871
rect 13369 7837 13403 7871
rect 14749 7837 14783 7871
rect 15025 7837 15059 7871
rect 15301 7837 15335 7871
rect 15577 7837 15611 7871
rect 15853 7837 15887 7871
rect 16129 7837 16163 7871
rect 16405 7837 16439 7871
rect 16957 7837 16991 7871
rect 17509 7837 17543 7871
rect 18061 7837 18095 7871
rect 18337 7837 18371 7871
rect 18429 7837 18463 7871
rect 18889 7837 18923 7871
rect 19441 7837 19475 7871
rect 19533 7837 19567 7871
rect 19809 7837 19843 7871
rect 21097 7837 21131 7871
rect 21925 7837 21959 7871
rect 2053 7769 2087 7803
rect 3985 7769 4019 7803
rect 4537 7769 4571 7803
rect 5641 7769 5675 7803
rect 6193 7769 6227 7803
rect 6745 7769 6779 7803
rect 7849 7769 7883 7803
rect 21557 7769 21591 7803
rect 22109 7769 22143 7803
rect 22661 7769 22695 7803
rect 23213 7769 23247 7803
rect 23765 7769 23799 7803
rect 10057 7701 10091 7735
rect 10149 7701 10183 7735
rect 10425 7701 10459 7735
rect 11529 7701 11563 7735
rect 16773 7701 16807 7735
rect 17325 7701 17359 7735
rect 17877 7701 17911 7735
rect 18613 7701 18647 7735
rect 19073 7701 19107 7735
rect 19717 7701 19751 7735
rect 19993 7701 20027 7735
rect 1685 7497 1719 7531
rect 2237 7497 2271 7531
rect 3525 7497 3559 7531
rect 5457 7497 5491 7531
rect 6377 7497 6411 7531
rect 7665 7497 7699 7531
rect 8309 7497 8343 7531
rect 8585 7497 8619 7531
rect 23857 7497 23891 7531
rect 23397 7429 23431 7463
rect 1593 7361 1627 7395
rect 2145 7361 2179 7395
rect 2697 7361 2731 7395
rect 3341 7361 3375 7395
rect 5641 7361 5675 7395
rect 6193 7361 6227 7395
rect 6561 7361 6595 7395
rect 7389 7361 7423 7395
rect 7849 7361 7883 7395
rect 8493 7365 8527 7399
rect 8769 7361 8803 7395
rect 10333 7361 10367 7395
rect 17417 7361 17451 7395
rect 22477 7361 22511 7395
rect 23029 7361 23063 7395
rect 23581 7361 23615 7395
rect 22753 7293 22787 7327
rect 7205 7225 7239 7259
rect 2789 7157 2823 7191
rect 6009 7157 6043 7191
rect 10149 7157 10183 7191
rect 17233 7157 17267 7191
rect 16681 6953 16715 6987
rect 23949 6817 23983 6851
rect 1961 6749 1995 6783
rect 16865 6749 16899 6783
rect 23489 6749 23523 6783
rect 1685 6681 1719 6715
rect 2329 6681 2363 6715
rect 23121 6681 23155 6715
rect 23673 6681 23707 6715
rect 1593 6409 1627 6443
rect 23305 6409 23339 6443
rect 23857 6409 23891 6443
rect 1501 6341 1535 6375
rect 23765 6341 23799 6375
rect 23213 6273 23247 6307
rect 24133 5865 24167 5899
rect 23857 5593 23891 5627
rect 14841 4573 14875 4607
rect 15025 4437 15059 4471
rect 14289 4233 14323 4267
rect 14473 4097 14507 4131
rect 23305 3689 23339 3723
rect 18061 3485 18095 3519
rect 23489 3485 23523 3519
rect 17877 3349 17911 3383
rect 23305 3145 23339 3179
rect 23857 3145 23891 3179
rect 22937 3009 22971 3043
rect 23489 3009 23523 3043
rect 24041 3009 24075 3043
rect 22753 2873 22787 2907
rect 23857 2601 23891 2635
rect 24041 2397 24075 2431
rect 9045 2057 9079 2091
rect 10425 2057 10459 2091
rect 10701 2057 10735 2091
rect 11713 2057 11747 2091
rect 12633 2057 12667 2091
rect 13001 2057 13035 2091
rect 13829 2057 13863 2091
rect 14289 2057 14323 2091
rect 22017 2057 22051 2091
rect 23397 2057 23431 2091
rect 23673 2057 23707 2091
rect 23949 2057 23983 2091
rect 7665 1921 7699 1955
rect 8861 1921 8895 1955
rect 10241 1921 10275 1955
rect 10517 1921 10551 1955
rect 11529 1921 11563 1955
rect 11805 1921 11839 1955
rect 12449 1921 12483 1955
rect 12817 1921 12851 1955
rect 13645 1921 13679 1955
rect 14105 1921 14139 1955
rect 16129 1921 16163 1955
rect 22201 1921 22235 1955
rect 23581 1921 23615 1955
rect 23857 1921 23891 1955
rect 24133 1921 24167 1955
rect 7849 1785 7883 1819
rect 11989 1785 12023 1819
rect 16313 1717 16347 1751
rect 7113 1513 7147 1547
rect 8309 1513 8343 1547
rect 9689 1513 9723 1547
rect 11069 1513 11103 1547
rect 12357 1513 12391 1547
rect 13093 1513 13127 1547
rect 15577 1513 15611 1547
rect 21833 1513 21867 1547
rect 22845 1513 22879 1547
rect 23121 1513 23155 1547
rect 23397 1513 23431 1547
rect 23673 1513 23707 1547
rect 9965 1445 9999 1479
rect 21281 1445 21315 1479
rect 1409 1309 1443 1343
rect 2145 1309 2179 1343
rect 3341 1309 3375 1343
rect 4721 1309 4755 1343
rect 5917 1309 5951 1343
rect 7297 1309 7331 1343
rect 7573 1309 7607 1343
rect 8493 1309 8527 1343
rect 8769 1309 8803 1343
rect 9505 1309 9539 1343
rect 9873 1309 9907 1343
rect 10149 1309 10183 1343
rect 10701 1309 10735 1343
rect 10977 1309 11011 1343
rect 11253 1309 11287 1343
rect 11897 1309 11931 1343
rect 12173 1309 12207 1343
rect 12541 1309 12575 1343
rect 13001 1309 13035 1343
rect 13277 1309 13311 1343
rect 13737 1309 13771 1343
rect 14289 1309 14323 1343
rect 14381 1309 14415 1343
rect 15485 1309 15519 1343
rect 15761 1309 15795 1343
rect 16865 1309 16899 1343
rect 17877 1309 17911 1343
rect 19073 1309 19107 1343
rect 20269 1309 20303 1343
rect 21465 1309 21499 1343
rect 22017 1309 22051 1343
rect 22661 1309 22695 1343
rect 23029 1309 23063 1343
rect 23305 1309 23339 1343
rect 23581 1309 23615 1343
rect 23857 1309 23891 1343
rect 24133 1309 24167 1343
rect 1593 1173 1627 1207
rect 2329 1173 2363 1207
rect 3525 1173 3559 1207
rect 4537 1173 4571 1207
rect 5733 1173 5767 1207
rect 7389 1173 7423 1207
rect 8585 1173 8619 1207
rect 9321 1173 9355 1207
rect 10517 1173 10551 1207
rect 10793 1173 10827 1207
rect 11713 1173 11747 1207
rect 11989 1173 12023 1207
rect 12817 1173 12851 1207
rect 13553 1173 13587 1207
rect 14105 1173 14139 1207
rect 14565 1173 14599 1207
rect 15301 1173 15335 1207
rect 16681 1173 16715 1207
rect 17693 1173 17727 1207
rect 18889 1173 18923 1207
rect 20085 1173 20119 1207
rect 22477 1173 22511 1207
rect 23949 1173 23983 1207
<< metal1 >>
rect 2222 9936 2228 9988
rect 2280 9976 2286 9988
rect 11790 9976 11796 9988
rect 2280 9948 11796 9976
rect 2280 9936 2286 9948
rect 11790 9936 11796 9948
rect 11848 9936 11854 9988
rect 11882 9936 11888 9988
rect 11940 9976 11946 9988
rect 17862 9976 17868 9988
rect 11940 9948 17868 9976
rect 11940 9936 11946 9948
rect 17862 9936 17868 9948
rect 17920 9936 17926 9988
rect 14274 9908 14280 9920
rect 2746 9880 14280 9908
rect 1578 9800 1584 9852
rect 1636 9840 1642 9852
rect 2746 9840 2774 9880
rect 14274 9868 14280 9880
rect 14332 9868 14338 9920
rect 1636 9812 2774 9840
rect 1636 9800 1642 9812
rect 5994 9800 6000 9852
rect 6052 9840 6058 9852
rect 14642 9840 14648 9852
rect 6052 9812 14648 9840
rect 6052 9800 6058 9812
rect 14642 9800 14648 9812
rect 14700 9800 14706 9852
rect 2424 9744 6684 9772
rect 2424 9716 2452 9744
rect 2406 9664 2412 9716
rect 2464 9664 2470 9716
rect 6656 9704 6684 9744
rect 7650 9732 7656 9784
rect 7708 9772 7714 9784
rect 7708 9744 18184 9772
rect 7708 9732 7714 9744
rect 18156 9716 18184 9744
rect 14826 9704 14832 9716
rect 6656 9676 14832 9704
rect 14826 9664 14832 9676
rect 14884 9664 14890 9716
rect 18138 9664 18144 9716
rect 18196 9664 18202 9716
rect 9490 9596 9496 9648
rect 9548 9636 9554 9648
rect 10134 9636 10140 9648
rect 9548 9608 10140 9636
rect 9548 9596 9554 9608
rect 10134 9596 10140 9608
rect 10192 9596 10198 9648
rect 11514 9596 11520 9648
rect 11572 9636 11578 9648
rect 19610 9636 19616 9648
rect 11572 9608 19616 9636
rect 11572 9596 11578 9608
rect 19610 9596 19616 9608
rect 19668 9596 19674 9648
rect 18966 9568 18972 9580
rect 6564 9540 18972 9568
rect 6564 9512 6592 9540
rect 18966 9528 18972 9540
rect 19024 9528 19030 9580
rect 6546 9460 6552 9512
rect 6604 9460 6610 9512
rect 7926 9460 7932 9512
rect 7984 9500 7990 9512
rect 11882 9500 11888 9512
rect 7984 9472 11888 9500
rect 7984 9460 7990 9472
rect 11882 9460 11888 9472
rect 11940 9460 11946 9512
rect 11238 9432 11244 9444
rect 6380 9404 11244 9432
rect 6380 9376 6408 9404
rect 11238 9392 11244 9404
rect 11296 9392 11302 9444
rect 6362 9324 6368 9376
rect 6420 9324 6426 9376
rect 8202 9324 8208 9376
rect 8260 9364 8266 9376
rect 12066 9364 12072 9376
rect 8260 9336 12072 9364
rect 8260 9324 8266 9336
rect 12066 9324 12072 9336
rect 12124 9324 12130 9376
rect 9030 9296 9036 9308
rect 1964 9268 9036 9296
rect 1964 9240 1992 9268
rect 9030 9256 9036 9268
rect 9088 9256 9094 9308
rect 9582 9256 9588 9308
rect 9640 9296 9646 9308
rect 15378 9296 15384 9308
rect 9640 9268 15384 9296
rect 9640 9256 9646 9268
rect 15378 9256 15384 9268
rect 15436 9256 15442 9308
rect 1946 9188 1952 9240
rect 2004 9188 2010 9240
rect 2498 9188 2504 9240
rect 2556 9228 2562 9240
rect 13446 9228 13452 9240
rect 2556 9200 13452 9228
rect 2556 9188 2562 9200
rect 13446 9188 13452 9200
rect 13504 9188 13510 9240
rect 7742 9120 7748 9172
rect 7800 9160 7806 9172
rect 11146 9160 11152 9172
rect 7800 9132 11152 9160
rect 7800 9120 7806 9132
rect 11146 9120 11152 9132
rect 11204 9120 11210 9172
rect 11238 9120 11244 9172
rect 11296 9120 11302 9172
rect 11790 9120 11796 9172
rect 11848 9160 11854 9172
rect 14550 9160 14556 9172
rect 11848 9132 14556 9160
rect 11848 9120 11854 9132
rect 14550 9120 14556 9132
rect 14608 9120 14614 9172
rect 4154 9052 4160 9104
rect 4212 9092 4218 9104
rect 11256 9092 11284 9120
rect 19334 9092 19340 9104
rect 4212 9064 11008 9092
rect 11256 9064 19340 9092
rect 4212 9052 4218 9064
rect 5534 8984 5540 9036
rect 5592 9024 5598 9036
rect 10870 9024 10876 9036
rect 5592 8996 10876 9024
rect 5592 8984 5598 8996
rect 10870 8984 10876 8996
rect 10928 8984 10934 9036
rect 10980 9024 11008 9064
rect 19334 9052 19340 9064
rect 19392 9052 19398 9104
rect 12342 9024 12348 9036
rect 10980 8996 12348 9024
rect 12342 8984 12348 8996
rect 12400 8984 12406 9036
rect 10042 8956 10048 8968
rect 4448 8928 10048 8956
rect 4448 8832 4476 8928
rect 10042 8916 10048 8928
rect 10100 8916 10106 8968
rect 16206 8956 16212 8968
rect 10336 8928 16212 8956
rect 9398 8888 9404 8900
rect 4908 8860 9404 8888
rect 4908 8832 4936 8860
rect 9398 8848 9404 8860
rect 9456 8848 9462 8900
rect 9950 8848 9956 8900
rect 10008 8888 10014 8900
rect 10336 8888 10364 8928
rect 16206 8916 16212 8928
rect 16264 8916 16270 8968
rect 10008 8860 10364 8888
rect 10008 8848 10014 8860
rect 10410 8848 10416 8900
rect 10468 8888 10474 8900
rect 16942 8888 16948 8900
rect 10468 8860 16948 8888
rect 10468 8848 10474 8860
rect 16942 8848 16948 8860
rect 17000 8848 17006 8900
rect 18874 8848 18880 8900
rect 18932 8888 18938 8900
rect 19794 8888 19800 8900
rect 18932 8860 19800 8888
rect 18932 8848 18938 8860
rect 19794 8848 19800 8860
rect 19852 8848 19858 8900
rect 106 8780 112 8832
rect 164 8820 170 8832
rect 2958 8820 2964 8832
rect 164 8792 2964 8820
rect 164 8780 170 8792
rect 2958 8780 2964 8792
rect 3016 8780 3022 8832
rect 4430 8780 4436 8832
rect 4488 8780 4494 8832
rect 4890 8780 4896 8832
rect 4948 8780 4954 8832
rect 8018 8780 8024 8832
rect 8076 8820 8082 8832
rect 17310 8820 17316 8832
rect 8076 8792 17316 8820
rect 8076 8780 8082 8792
rect 17310 8780 17316 8792
rect 17368 8780 17374 8832
rect 18598 8780 18604 8832
rect 18656 8820 18662 8832
rect 19518 8820 19524 8832
rect 18656 8792 19524 8820
rect 18656 8780 18662 8792
rect 19518 8780 19524 8792
rect 19576 8780 19582 8832
rect 1104 8730 24723 8752
rect 1104 8678 6814 8730
rect 6866 8678 6878 8730
rect 6930 8678 6942 8730
rect 6994 8678 7006 8730
rect 7058 8678 7070 8730
rect 7122 8678 12679 8730
rect 12731 8678 12743 8730
rect 12795 8678 12807 8730
rect 12859 8678 12871 8730
rect 12923 8678 12935 8730
rect 12987 8678 18544 8730
rect 18596 8678 18608 8730
rect 18660 8678 18672 8730
rect 18724 8678 18736 8730
rect 18788 8678 18800 8730
rect 18852 8678 24409 8730
rect 24461 8678 24473 8730
rect 24525 8678 24537 8730
rect 24589 8678 24601 8730
rect 24653 8678 24665 8730
rect 24717 8678 24723 8730
rect 1104 8656 24723 8678
rect 566 8576 572 8628
rect 624 8616 630 8628
rect 2041 8619 2099 8625
rect 2041 8616 2053 8619
rect 624 8588 2053 8616
rect 624 8576 630 8588
rect 2041 8585 2053 8588
rect 2087 8585 2099 8619
rect 2041 8579 2099 8585
rect 2777 8619 2835 8625
rect 2777 8585 2789 8619
rect 2823 8616 2835 8619
rect 2866 8616 2872 8628
rect 2823 8588 2872 8616
rect 2823 8585 2835 8588
rect 2777 8579 2835 8585
rect 2866 8576 2872 8588
rect 2924 8576 2930 8628
rect 2958 8576 2964 8628
rect 3016 8616 3022 8628
rect 3145 8619 3203 8625
rect 3145 8616 3157 8619
rect 3016 8588 3157 8616
rect 3016 8576 3022 8588
rect 3145 8585 3157 8588
rect 3191 8585 3203 8619
rect 4154 8616 4160 8628
rect 3145 8579 3203 8585
rect 3896 8588 4160 8616
rect 3896 8548 3924 8588
rect 4154 8576 4160 8588
rect 4212 8576 4218 8628
rect 4246 8576 4252 8628
rect 4304 8576 4310 8628
rect 4617 8619 4675 8625
rect 4617 8585 4629 8619
rect 4663 8616 4675 8619
rect 5074 8616 5080 8628
rect 4663 8588 5080 8616
rect 4663 8585 4675 8588
rect 4617 8579 4675 8585
rect 5074 8576 5080 8588
rect 5132 8576 5138 8628
rect 5169 8619 5227 8625
rect 5169 8585 5181 8619
rect 5215 8616 5227 8619
rect 5350 8616 5356 8628
rect 5215 8588 5356 8616
rect 5215 8585 5227 8588
rect 5169 8579 5227 8585
rect 5350 8576 5356 8588
rect 5408 8576 5414 8628
rect 5721 8619 5779 8625
rect 5721 8585 5733 8619
rect 5767 8616 5779 8619
rect 5902 8616 5908 8628
rect 5767 8588 5908 8616
rect 5767 8585 5779 8588
rect 5721 8579 5779 8585
rect 5902 8576 5908 8588
rect 5960 8576 5966 8628
rect 6089 8619 6147 8625
rect 6089 8585 6101 8619
rect 6135 8616 6147 8619
rect 6454 8616 6460 8628
rect 6135 8588 6460 8616
rect 6135 8585 6147 8588
rect 6089 8579 6147 8585
rect 6454 8576 6460 8588
rect 6512 8576 6518 8628
rect 6825 8619 6883 8625
rect 6825 8585 6837 8619
rect 6871 8616 6883 8619
rect 7190 8616 7196 8628
rect 6871 8588 7196 8616
rect 6871 8585 6883 8588
rect 6825 8579 6883 8585
rect 7190 8576 7196 8588
rect 7248 8576 7254 8628
rect 7377 8619 7435 8625
rect 7377 8585 7389 8619
rect 7423 8616 7435 8619
rect 7558 8616 7564 8628
rect 7423 8588 7564 8616
rect 7423 8585 7435 8588
rect 7377 8579 7435 8585
rect 7558 8576 7564 8588
rect 7616 8576 7622 8628
rect 7745 8619 7803 8625
rect 7745 8585 7757 8619
rect 7791 8616 7803 8619
rect 8110 8616 8116 8628
rect 7791 8588 8116 8616
rect 7791 8585 7803 8588
rect 7745 8579 7803 8585
rect 8110 8576 8116 8588
rect 8168 8576 8174 8628
rect 8297 8619 8355 8625
rect 8297 8585 8309 8619
rect 8343 8616 8355 8619
rect 8386 8616 8392 8628
rect 8343 8588 8392 8616
rect 8343 8585 8355 8588
rect 8297 8579 8355 8585
rect 8386 8576 8392 8588
rect 8444 8576 8450 8628
rect 8665 8619 8723 8625
rect 8665 8585 8677 8619
rect 8711 8616 8723 8619
rect 8938 8616 8944 8628
rect 8711 8588 8944 8616
rect 8711 8585 8723 8588
rect 8665 8579 8723 8585
rect 8938 8576 8944 8588
rect 8996 8576 9002 8628
rect 9214 8576 9220 8628
rect 9272 8616 9278 8628
rect 9309 8619 9367 8625
rect 9309 8616 9321 8619
rect 9272 8588 9321 8616
rect 9272 8576 9278 8588
rect 9309 8585 9321 8588
rect 9355 8585 9367 8619
rect 9309 8579 9367 8585
rect 9674 8576 9680 8628
rect 9732 8576 9738 8628
rect 9950 8576 9956 8628
rect 10008 8616 10014 8628
rect 10008 8588 10180 8616
rect 10008 8576 10014 8588
rect 1504 8520 3924 8548
rect 3973 8551 4031 8557
rect 1504 8489 1532 8520
rect 3973 8517 3985 8551
rect 4019 8548 4031 8551
rect 4019 8520 6500 8548
rect 4019 8517 4031 8520
rect 3973 8511 4031 8517
rect 1489 8483 1547 8489
rect 1489 8449 1501 8483
rect 1535 8449 1547 8483
rect 1489 8443 1547 8449
rect 1946 8440 1952 8492
rect 2004 8440 2010 8492
rect 2498 8440 2504 8492
rect 2556 8440 2562 8492
rect 3053 8483 3111 8489
rect 3053 8449 3065 8483
rect 3099 8449 3111 8483
rect 3053 8443 3111 8449
rect 3068 8412 3096 8443
rect 4430 8440 4436 8492
rect 4488 8440 4494 8492
rect 4890 8440 4896 8492
rect 4948 8440 4954 8492
rect 5445 8483 5503 8489
rect 5445 8449 5457 8483
rect 5491 8480 5503 8483
rect 5810 8480 5816 8492
rect 5491 8452 5816 8480
rect 5491 8449 5503 8452
rect 5445 8443 5503 8449
rect 5810 8440 5816 8452
rect 5868 8440 5874 8492
rect 5902 8440 5908 8492
rect 5960 8440 5966 8492
rect 6472 8480 6500 8520
rect 6546 8508 6552 8560
rect 6604 8508 6610 8560
rect 7116 8520 7696 8548
rect 7116 8480 7144 8520
rect 6472 8452 7144 8480
rect 7190 8440 7196 8492
rect 7248 8440 7254 8492
rect 7561 8483 7619 8489
rect 7561 8449 7573 8483
rect 7607 8449 7619 8483
rect 7668 8480 7696 8520
rect 8018 8508 8024 8560
rect 8076 8508 8082 8560
rect 8128 8520 9260 8548
rect 8128 8480 8156 8520
rect 7668 8452 8156 8480
rect 8481 8483 8539 8489
rect 7561 8443 7619 8449
rect 8481 8449 8493 8483
rect 8527 8449 8539 8483
rect 8481 8443 8539 8449
rect 9125 8483 9183 8489
rect 9125 8449 9137 8483
rect 9171 8449 9183 8483
rect 9232 8480 9260 8520
rect 9582 8508 9588 8560
rect 9640 8508 9646 8560
rect 10152 8557 10180 8588
rect 10226 8576 10232 8628
rect 10284 8576 10290 8628
rect 12894 8616 12900 8628
rect 12544 8588 12900 8616
rect 10137 8551 10195 8557
rect 10137 8517 10149 8551
rect 10183 8517 10195 8551
rect 10137 8511 10195 8517
rect 10428 8520 10732 8548
rect 10428 8480 10456 8520
rect 9232 8452 10456 8480
rect 9125 8443 9183 8449
rect 7374 8412 7380 8424
rect 3068 8384 7380 8412
rect 7374 8372 7380 8384
rect 7432 8372 7438 8424
rect 7576 8412 7604 8443
rect 8294 8412 8300 8424
rect 7576 8384 8300 8412
rect 8294 8372 8300 8384
rect 8352 8372 8358 8424
rect 1673 8347 1731 8353
rect 1673 8313 1685 8347
rect 1719 8344 1731 8347
rect 3418 8344 3424 8356
rect 1719 8316 3424 8344
rect 1719 8313 1731 8316
rect 1673 8307 1731 8313
rect 3418 8304 3424 8316
rect 3476 8304 3482 8356
rect 6638 8304 6644 8356
rect 6696 8344 6702 8356
rect 8496 8344 8524 8443
rect 9140 8412 9168 8443
rect 10226 8412 10232 8424
rect 9140 8384 10232 8412
rect 10226 8372 10232 8384
rect 10284 8372 10290 8424
rect 10410 8344 10416 8356
rect 6696 8316 8432 8344
rect 8496 8316 10416 8344
rect 6696 8304 6702 8316
rect 8404 8276 8432 8316
rect 10410 8304 10416 8316
rect 10468 8304 10474 8356
rect 10597 8347 10655 8353
rect 10597 8344 10609 8347
rect 10520 8316 10609 8344
rect 10520 8276 10548 8316
rect 10597 8313 10609 8316
rect 10643 8313 10655 8347
rect 10597 8307 10655 8313
rect 8404 8248 10548 8276
rect 10704 8276 10732 8520
rect 11146 8508 11152 8560
rect 11204 8548 11210 8560
rect 12544 8548 12572 8588
rect 12894 8576 12900 8588
rect 12952 8576 12958 8628
rect 13173 8619 13231 8625
rect 13173 8585 13185 8619
rect 13219 8585 13231 8619
rect 13725 8619 13783 8625
rect 13725 8616 13737 8619
rect 13173 8579 13231 8585
rect 13280 8588 13737 8616
rect 13188 8548 13216 8579
rect 11204 8520 11928 8548
rect 11204 8508 11210 8520
rect 10781 8483 10839 8489
rect 10781 8449 10793 8483
rect 10827 8449 10839 8483
rect 10781 8443 10839 8449
rect 10796 8412 10824 8443
rect 11054 8440 11060 8492
rect 11112 8440 11118 8492
rect 11333 8483 11391 8489
rect 11333 8449 11345 8483
rect 11379 8480 11391 8483
rect 11514 8480 11520 8492
rect 11379 8452 11520 8480
rect 11379 8449 11391 8452
rect 11333 8443 11391 8449
rect 11514 8440 11520 8452
rect 11572 8440 11578 8492
rect 11698 8440 11704 8492
rect 11756 8440 11762 8492
rect 10796 8384 11560 8412
rect 10870 8304 10876 8356
rect 10928 8304 10934 8356
rect 11532 8353 11560 8384
rect 11149 8347 11207 8353
rect 11149 8313 11161 8347
rect 11195 8313 11207 8347
rect 11149 8307 11207 8313
rect 11517 8347 11575 8353
rect 11517 8313 11529 8347
rect 11563 8313 11575 8347
rect 11900 8344 11928 8520
rect 12406 8520 12572 8548
rect 12636 8520 13216 8548
rect 11977 8483 12035 8489
rect 11977 8449 11989 8483
rect 12023 8449 12035 8483
rect 11977 8443 12035 8449
rect 12253 8483 12311 8489
rect 12253 8449 12265 8483
rect 12299 8480 12311 8483
rect 12406 8480 12434 8520
rect 12636 8489 12664 8520
rect 12299 8452 12434 8480
rect 12529 8483 12587 8489
rect 12299 8449 12311 8452
rect 12253 8443 12311 8449
rect 12529 8449 12541 8483
rect 12575 8449 12587 8483
rect 12529 8443 12587 8449
rect 12621 8483 12679 8489
rect 12621 8449 12633 8483
rect 12667 8449 12679 8483
rect 12621 8443 12679 8449
rect 12897 8483 12955 8489
rect 12897 8449 12909 8483
rect 12943 8480 12955 8483
rect 13280 8480 13308 8588
rect 13725 8585 13737 8588
rect 13771 8585 13783 8619
rect 13725 8579 13783 8585
rect 14550 8576 14556 8628
rect 14608 8576 14614 8628
rect 14826 8576 14832 8628
rect 14884 8576 14890 8628
rect 15010 8576 15016 8628
rect 15068 8616 15074 8628
rect 16669 8619 16727 8625
rect 16669 8616 16681 8619
rect 15068 8588 16681 8616
rect 15068 8576 15074 8588
rect 16669 8585 16681 8588
rect 16715 8585 16727 8619
rect 16669 8579 16727 8585
rect 16942 8576 16948 8628
rect 17000 8576 17006 8628
rect 17221 8619 17279 8625
rect 17221 8585 17233 8619
rect 17267 8585 17279 8619
rect 17221 8579 17279 8585
rect 14182 8508 14188 8560
rect 14240 8548 14246 8560
rect 14240 8520 15148 8548
rect 14240 8508 14246 8520
rect 12943 8452 13308 8480
rect 12943 8449 12955 8452
rect 12897 8443 12955 8449
rect 11992 8412 12020 8443
rect 12434 8412 12440 8424
rect 11992 8384 12440 8412
rect 12434 8372 12440 8384
rect 12492 8372 12498 8424
rect 12544 8412 12572 8443
rect 13354 8440 13360 8492
rect 13412 8440 13418 8492
rect 13449 8483 13507 8489
rect 13449 8449 13461 8483
rect 13495 8449 13507 8483
rect 13449 8443 13507 8449
rect 13170 8412 13176 8424
rect 12544 8384 13176 8412
rect 13170 8372 13176 8384
rect 13228 8372 13234 8424
rect 13464 8412 13492 8443
rect 13630 8440 13636 8492
rect 13688 8480 13694 8492
rect 13909 8483 13967 8489
rect 13909 8480 13921 8483
rect 13688 8452 13921 8480
rect 13688 8440 13694 8452
rect 13909 8449 13921 8452
rect 13955 8449 13967 8483
rect 13909 8443 13967 8449
rect 13998 8440 14004 8492
rect 14056 8480 14062 8492
rect 14277 8483 14335 8489
rect 14277 8480 14289 8483
rect 14056 8452 14289 8480
rect 14056 8440 14062 8452
rect 14277 8449 14289 8452
rect 14323 8449 14335 8483
rect 14277 8443 14335 8449
rect 14369 8483 14427 8489
rect 14369 8449 14381 8483
rect 14415 8449 14427 8483
rect 14369 8443 14427 8449
rect 14384 8412 14412 8443
rect 14642 8440 14648 8492
rect 14700 8440 14706 8492
rect 14734 8440 14740 8492
rect 14792 8480 14798 8492
rect 15120 8489 15148 8520
rect 15378 8508 15384 8560
rect 15436 8548 15442 8560
rect 15436 8520 15884 8548
rect 15436 8508 15442 8520
rect 15105 8483 15163 8489
rect 14792 8452 15056 8480
rect 14792 8440 14798 8452
rect 13464 8384 14136 8412
rect 14384 8384 14964 8412
rect 11900 8316 12296 8344
rect 11517 8307 11575 8313
rect 11164 8276 11192 8307
rect 10704 8248 11192 8276
rect 11790 8236 11796 8288
rect 11848 8236 11854 8288
rect 12066 8236 12072 8288
rect 12124 8236 12130 8288
rect 12268 8276 12296 8316
rect 12342 8304 12348 8356
rect 12400 8304 12406 8356
rect 12805 8347 12863 8353
rect 12805 8344 12817 8347
rect 12452 8316 12817 8344
rect 12452 8276 12480 8316
rect 12805 8313 12817 8316
rect 12851 8313 12863 8347
rect 12805 8307 12863 8313
rect 13081 8347 13139 8353
rect 13081 8313 13093 8347
rect 13127 8344 13139 8347
rect 13446 8344 13452 8356
rect 13127 8316 13452 8344
rect 13127 8313 13139 8316
rect 13081 8307 13139 8313
rect 13446 8304 13452 8316
rect 13504 8304 13510 8356
rect 13630 8304 13636 8356
rect 13688 8304 13694 8356
rect 14108 8353 14136 8384
rect 14093 8347 14151 8353
rect 14093 8313 14105 8347
rect 14139 8313 14151 8347
rect 14093 8307 14151 8313
rect 14274 8304 14280 8356
rect 14332 8344 14338 8356
rect 14936 8353 14964 8384
rect 14921 8347 14979 8353
rect 14332 8316 14872 8344
rect 14332 8304 14338 8316
rect 12268 8248 12480 8276
rect 14844 8276 14872 8316
rect 14921 8313 14933 8347
rect 14967 8313 14979 8347
rect 15028 8344 15056 8452
rect 15105 8449 15117 8483
rect 15151 8449 15163 8483
rect 15105 8443 15163 8449
rect 15194 8440 15200 8492
rect 15252 8440 15258 8492
rect 15286 8440 15292 8492
rect 15344 8480 15350 8492
rect 15473 8483 15531 8489
rect 15473 8480 15485 8483
rect 15344 8452 15485 8480
rect 15344 8440 15350 8452
rect 15473 8449 15485 8452
rect 15519 8449 15531 8483
rect 15473 8443 15531 8449
rect 15749 8483 15807 8489
rect 15749 8449 15761 8483
rect 15795 8449 15807 8483
rect 15749 8443 15807 8449
rect 15378 8372 15384 8424
rect 15436 8412 15442 8424
rect 15764 8412 15792 8443
rect 15436 8384 15792 8412
rect 15856 8412 15884 8520
rect 16114 8440 16120 8492
rect 16172 8480 16178 8492
rect 16209 8483 16267 8489
rect 16209 8480 16221 8483
rect 16172 8452 16221 8480
rect 16172 8440 16178 8452
rect 16209 8449 16221 8452
rect 16255 8449 16267 8483
rect 16209 8443 16267 8449
rect 16482 8440 16488 8492
rect 16540 8440 16546 8492
rect 16850 8440 16856 8492
rect 16908 8440 16914 8492
rect 17129 8483 17187 8489
rect 17129 8449 17141 8483
rect 17175 8480 17187 8483
rect 17236 8480 17264 8579
rect 17310 8576 17316 8628
rect 17368 8616 17374 8628
rect 17497 8619 17555 8625
rect 17497 8616 17509 8619
rect 17368 8588 17509 8616
rect 17368 8576 17374 8588
rect 17497 8585 17509 8588
rect 17543 8585 17555 8619
rect 17497 8579 17555 8585
rect 17773 8619 17831 8625
rect 17773 8585 17785 8619
rect 17819 8585 17831 8619
rect 17773 8579 17831 8585
rect 17175 8452 17264 8480
rect 17405 8483 17463 8489
rect 17175 8449 17187 8452
rect 17129 8443 17187 8449
rect 17405 8449 17417 8483
rect 17451 8449 17463 8483
rect 17405 8443 17463 8449
rect 17681 8483 17739 8489
rect 17681 8449 17693 8483
rect 17727 8480 17739 8483
rect 17788 8480 17816 8579
rect 17862 8576 17868 8628
rect 17920 8616 17926 8628
rect 18233 8619 18291 8625
rect 18233 8616 18245 8619
rect 17920 8588 18245 8616
rect 17920 8576 17926 8588
rect 18233 8585 18245 8588
rect 18279 8585 18291 8619
rect 18233 8579 18291 8585
rect 18325 8619 18383 8625
rect 18325 8585 18337 8619
rect 18371 8585 18383 8619
rect 18325 8579 18383 8585
rect 17727 8452 17816 8480
rect 17727 8449 17739 8452
rect 17681 8443 17739 8449
rect 15856 8384 16160 8412
rect 15436 8372 15442 8384
rect 15028 8316 15700 8344
rect 14921 8307 14979 8313
rect 15672 8285 15700 8316
rect 15381 8279 15439 8285
rect 15381 8276 15393 8279
rect 14844 8248 15393 8276
rect 15381 8245 15393 8248
rect 15427 8245 15439 8279
rect 15381 8239 15439 8245
rect 15657 8279 15715 8285
rect 15657 8245 15669 8279
rect 15703 8245 15715 8279
rect 15657 8239 15715 8245
rect 15838 8236 15844 8288
rect 15896 8276 15902 8288
rect 15933 8279 15991 8285
rect 15933 8276 15945 8279
rect 15896 8248 15945 8276
rect 15896 8236 15902 8248
rect 15933 8245 15945 8248
rect 15979 8245 15991 8279
rect 15933 8239 15991 8245
rect 16025 8279 16083 8285
rect 16025 8245 16037 8279
rect 16071 8276 16083 8279
rect 16132 8276 16160 8384
rect 16574 8372 16580 8424
rect 16632 8412 16638 8424
rect 17420 8412 17448 8443
rect 17862 8440 17868 8492
rect 17920 8480 17926 8492
rect 17957 8483 18015 8489
rect 17957 8480 17969 8483
rect 17920 8452 17969 8480
rect 17920 8440 17926 8452
rect 17957 8449 17969 8452
rect 18003 8449 18015 8483
rect 17957 8443 18015 8449
rect 18049 8483 18107 8489
rect 18049 8449 18061 8483
rect 18095 8480 18107 8483
rect 18340 8480 18368 8579
rect 18414 8576 18420 8628
rect 18472 8616 18478 8628
rect 18472 8588 19472 8616
rect 18472 8576 18478 8588
rect 18095 8452 18368 8480
rect 18509 8483 18567 8489
rect 18095 8449 18107 8452
rect 18049 8443 18107 8449
rect 18509 8449 18521 8483
rect 18555 8449 18567 8483
rect 18509 8443 18567 8449
rect 16632 8384 17448 8412
rect 16632 8372 16638 8384
rect 17494 8372 17500 8424
rect 17552 8412 17558 8424
rect 18524 8412 18552 8443
rect 18598 8440 18604 8492
rect 18656 8440 18662 8492
rect 18877 8483 18935 8489
rect 18877 8449 18889 8483
rect 18923 8480 18935 8483
rect 18923 8452 19288 8480
rect 18923 8449 18935 8452
rect 18877 8443 18935 8449
rect 17552 8384 18552 8412
rect 17552 8372 17558 8384
rect 18966 8372 18972 8424
rect 19024 8372 19030 8424
rect 16206 8304 16212 8356
rect 16264 8344 16270 8356
rect 16301 8347 16359 8353
rect 16301 8344 16313 8347
rect 16264 8316 16313 8344
rect 16264 8304 16270 8316
rect 16301 8313 16313 8316
rect 16347 8313 16359 8347
rect 16301 8307 16359 8313
rect 17126 8304 17132 8356
rect 17184 8344 17190 8356
rect 17862 8344 17868 8356
rect 17184 8316 17868 8344
rect 17184 8304 17190 8316
rect 17862 8304 17868 8316
rect 17920 8304 17926 8356
rect 18138 8304 18144 8356
rect 18196 8344 18202 8356
rect 18785 8347 18843 8353
rect 18785 8344 18797 8347
rect 18196 8316 18797 8344
rect 18196 8304 18202 8316
rect 18785 8313 18797 8316
rect 18831 8313 18843 8347
rect 18984 8344 19012 8372
rect 19260 8353 19288 8452
rect 19334 8440 19340 8492
rect 19392 8440 19398 8492
rect 19444 8489 19472 8588
rect 19610 8576 19616 8628
rect 19668 8616 19674 8628
rect 19668 8588 19932 8616
rect 19668 8576 19674 8588
rect 19904 8548 19932 8588
rect 19978 8576 19984 8628
rect 20036 8616 20042 8628
rect 20257 8619 20315 8625
rect 20257 8616 20269 8619
rect 20036 8588 20269 8616
rect 20036 8576 20042 8588
rect 20257 8585 20269 8588
rect 20303 8585 20315 8619
rect 20257 8579 20315 8585
rect 20346 8576 20352 8628
rect 20404 8616 20410 8628
rect 20625 8619 20683 8625
rect 20625 8616 20637 8619
rect 20404 8588 20637 8616
rect 20404 8576 20410 8588
rect 20625 8585 20637 8588
rect 20671 8585 20683 8619
rect 20625 8579 20683 8585
rect 21082 8576 21088 8628
rect 21140 8616 21146 8628
rect 22005 8619 22063 8625
rect 22005 8616 22017 8619
rect 21140 8588 22017 8616
rect 21140 8576 21146 8588
rect 22005 8585 22017 8588
rect 22051 8585 22063 8619
rect 22005 8579 22063 8585
rect 22557 8619 22615 8625
rect 22557 8585 22569 8619
rect 22603 8585 22615 8619
rect 22557 8579 22615 8585
rect 20533 8551 20591 8557
rect 20533 8548 20545 8551
rect 19904 8520 20545 8548
rect 20533 8517 20545 8520
rect 20579 8517 20591 8551
rect 20533 8511 20591 8517
rect 21358 8508 21364 8560
rect 21416 8548 21422 8560
rect 22572 8548 22600 8579
rect 23198 8576 23204 8628
rect 23256 8616 23262 8628
rect 23661 8619 23719 8625
rect 23661 8616 23673 8619
rect 23256 8588 23673 8616
rect 23256 8576 23262 8588
rect 23661 8585 23673 8588
rect 23707 8585 23719 8619
rect 23661 8579 23719 8585
rect 21416 8520 22600 8548
rect 21416 8508 21422 8520
rect 19429 8483 19487 8489
rect 19429 8449 19441 8483
rect 19475 8449 19487 8483
rect 19429 8443 19487 8449
rect 19518 8440 19524 8492
rect 19576 8480 19582 8492
rect 19705 8483 19763 8489
rect 19705 8480 19717 8483
rect 19576 8452 19717 8480
rect 19576 8440 19582 8452
rect 19705 8449 19717 8452
rect 19751 8449 19763 8483
rect 19705 8443 19763 8449
rect 19794 8440 19800 8492
rect 19852 8440 19858 8492
rect 20070 8440 20076 8492
rect 20128 8440 20134 8492
rect 20714 8440 20720 8492
rect 20772 8480 20778 8492
rect 21085 8483 21143 8489
rect 21085 8480 21097 8483
rect 20772 8452 21097 8480
rect 20772 8440 20778 8452
rect 21085 8449 21097 8452
rect 21131 8449 21143 8483
rect 21085 8443 21143 8449
rect 21174 8440 21180 8492
rect 21232 8480 21238 8492
rect 21913 8483 21971 8489
rect 21913 8480 21925 8483
rect 21232 8452 21925 8480
rect 21232 8440 21238 8452
rect 21913 8449 21925 8452
rect 21959 8449 21971 8483
rect 21913 8443 21971 8449
rect 22462 8440 22468 8492
rect 22520 8440 22526 8492
rect 23014 8440 23020 8492
rect 23072 8440 23078 8492
rect 23566 8440 23572 8492
rect 23624 8440 23630 8492
rect 19061 8347 19119 8353
rect 19061 8344 19073 8347
rect 18984 8316 19073 8344
rect 18785 8307 18843 8313
rect 19061 8313 19073 8316
rect 19107 8313 19119 8347
rect 19061 8307 19119 8313
rect 19245 8347 19303 8353
rect 19245 8313 19257 8347
rect 19291 8313 19303 8347
rect 19352 8344 19380 8440
rect 19981 8347 20039 8353
rect 19981 8344 19993 8347
rect 19352 8316 19993 8344
rect 19245 8307 19303 8313
rect 19981 8313 19993 8316
rect 20027 8313 20039 8347
rect 19981 8307 20039 8313
rect 20530 8304 20536 8356
rect 20588 8344 20594 8356
rect 21269 8347 21327 8353
rect 21269 8344 21281 8347
rect 20588 8316 21281 8344
rect 20588 8304 20594 8316
rect 21269 8313 21281 8316
rect 21315 8313 21327 8347
rect 21269 8307 21327 8313
rect 21634 8304 21640 8356
rect 21692 8344 21698 8356
rect 23201 8347 23259 8353
rect 23201 8344 23213 8347
rect 21692 8316 23213 8344
rect 21692 8304 21698 8316
rect 23201 8313 23213 8316
rect 23247 8313 23259 8347
rect 23201 8307 23259 8313
rect 16071 8248 16160 8276
rect 16071 8245 16083 8248
rect 16025 8239 16083 8245
rect 19518 8236 19524 8288
rect 19576 8236 19582 8288
rect 1104 8186 24564 8208
rect 1104 8134 3882 8186
rect 3934 8134 3946 8186
rect 3998 8134 4010 8186
rect 4062 8134 4074 8186
rect 4126 8134 4138 8186
rect 4190 8134 9747 8186
rect 9799 8134 9811 8186
rect 9863 8134 9875 8186
rect 9927 8134 9939 8186
rect 9991 8134 10003 8186
rect 10055 8134 15612 8186
rect 15664 8134 15676 8186
rect 15728 8134 15740 8186
rect 15792 8134 15804 8186
rect 15856 8134 15868 8186
rect 15920 8134 21477 8186
rect 21529 8134 21541 8186
rect 21593 8134 21605 8186
rect 21657 8134 21669 8186
rect 21721 8134 21733 8186
rect 21785 8134 24564 8186
rect 1104 8112 24564 8134
rect 1765 8075 1823 8081
rect 1765 8041 1777 8075
rect 1811 8072 1823 8075
rect 2038 8072 2044 8084
rect 1811 8044 2044 8072
rect 1811 8041 1823 8044
rect 1765 8035 1823 8041
rect 2038 8032 2044 8044
rect 2096 8032 2102 8084
rect 2314 8032 2320 8084
rect 2372 8032 2378 8084
rect 3234 8032 3240 8084
rect 3292 8032 3298 8084
rect 4614 8032 4620 8084
rect 4672 8032 4678 8084
rect 4798 8032 4804 8084
rect 4856 8072 4862 8084
rect 5169 8075 5227 8081
rect 5169 8072 5181 8075
rect 4856 8044 5181 8072
rect 4856 8032 4862 8044
rect 5169 8041 5181 8044
rect 5215 8041 5227 8075
rect 5169 8035 5227 8041
rect 5718 8032 5724 8084
rect 5776 8032 5782 8084
rect 6270 8032 6276 8084
rect 6328 8032 6334 8084
rect 6840 8044 7236 8072
rect 2774 7964 2780 8016
rect 2832 7964 2838 8016
rect 4154 7964 4160 8016
rect 4212 7964 4218 8016
rect 6840 8004 6868 8044
rect 5368 7976 6868 8004
rect 5368 7936 5396 7976
rect 6914 7964 6920 8016
rect 6972 7964 6978 8016
rect 7208 8004 7236 8044
rect 7282 8032 7288 8084
rect 7340 8072 7346 8084
rect 7377 8075 7435 8081
rect 7377 8072 7389 8075
rect 7340 8044 7389 8072
rect 7340 8032 7346 8044
rect 7377 8041 7389 8044
rect 7423 8041 7435 8075
rect 7377 8035 7435 8041
rect 7926 8032 7932 8084
rect 7984 8032 7990 8084
rect 8662 8032 8668 8084
rect 8720 8032 8726 8084
rect 9309 8075 9367 8081
rect 9309 8072 9321 8075
rect 8772 8044 9321 8072
rect 7742 8004 7748 8016
rect 7208 7976 7748 8004
rect 7742 7964 7748 7976
rect 7800 7964 7806 8016
rect 3160 7908 5396 7936
rect 1489 7871 1547 7877
rect 1489 7837 1501 7871
rect 1535 7868 1547 7871
rect 2406 7868 2412 7880
rect 1535 7840 2412 7868
rect 1535 7837 1547 7840
rect 1489 7831 1547 7837
rect 2406 7828 2412 7840
rect 2464 7828 2470 7880
rect 2590 7828 2596 7880
rect 2648 7828 2654 7880
rect 3160 7877 3188 7908
rect 5442 7896 5448 7948
rect 5500 7936 5506 7948
rect 8772 7936 8800 8044
rect 9309 8041 9321 8044
rect 9355 8041 9367 8075
rect 9309 8035 9367 8041
rect 9398 8032 9404 8084
rect 9456 8072 9462 8084
rect 9585 8075 9643 8081
rect 9585 8072 9597 8075
rect 9456 8044 9597 8072
rect 9456 8032 9462 8044
rect 9585 8041 9597 8044
rect 9631 8041 9643 8075
rect 9585 8035 9643 8041
rect 9766 8032 9772 8084
rect 9824 8072 9830 8084
rect 11241 8075 11299 8081
rect 11241 8072 11253 8075
rect 9824 8044 11253 8072
rect 9824 8032 9830 8044
rect 11241 8041 11253 8044
rect 11287 8041 11299 8075
rect 11241 8035 11299 8041
rect 11514 8032 11520 8084
rect 11572 8072 11578 8084
rect 12345 8075 12403 8081
rect 12345 8072 12357 8075
rect 11572 8044 12357 8072
rect 11572 8032 11578 8044
rect 12345 8041 12357 8044
rect 12391 8041 12403 8075
rect 12345 8035 12403 8041
rect 12434 8032 12440 8084
rect 12492 8072 12498 8084
rect 12621 8075 12679 8081
rect 12621 8072 12633 8075
rect 12492 8044 12633 8072
rect 12492 8032 12498 8044
rect 12621 8041 12633 8044
rect 12667 8041 12679 8075
rect 12621 8035 12679 8041
rect 12894 8032 12900 8084
rect 12952 8032 12958 8084
rect 13170 8032 13176 8084
rect 13228 8032 13234 8084
rect 14553 8075 14611 8081
rect 14553 8041 14565 8075
rect 14599 8072 14611 8075
rect 14642 8072 14648 8084
rect 14599 8044 14648 8072
rect 14599 8041 14611 8044
rect 14553 8035 14611 8041
rect 14642 8032 14648 8044
rect 14700 8032 14706 8084
rect 14829 8075 14887 8081
rect 14829 8041 14841 8075
rect 14875 8072 14887 8075
rect 15194 8072 15200 8084
rect 14875 8044 15200 8072
rect 14875 8041 14887 8044
rect 14829 8035 14887 8041
rect 15194 8032 15200 8044
rect 15252 8032 15258 8084
rect 15286 8032 15292 8084
rect 15344 8032 15350 8084
rect 15378 8032 15384 8084
rect 15436 8032 15442 8084
rect 15657 8075 15715 8081
rect 15657 8041 15669 8075
rect 15703 8072 15715 8075
rect 16114 8072 16120 8084
rect 15703 8044 16120 8072
rect 15703 8041 15715 8044
rect 15657 8035 15715 8041
rect 16114 8032 16120 8044
rect 16172 8032 16178 8084
rect 16209 8075 16267 8081
rect 16209 8041 16221 8075
rect 16255 8072 16267 8075
rect 16850 8072 16856 8084
rect 16255 8044 16856 8072
rect 16255 8041 16267 8044
rect 16209 8035 16267 8041
rect 16850 8032 16856 8044
rect 16908 8032 16914 8084
rect 18141 8075 18199 8081
rect 18141 8041 18153 8075
rect 18187 8072 18199 8075
rect 18598 8072 18604 8084
rect 18187 8044 18604 8072
rect 18187 8041 18199 8044
rect 18141 8035 18199 8041
rect 18598 8032 18604 8044
rect 18656 8032 18662 8084
rect 19518 8072 19524 8084
rect 18800 8044 19524 8072
rect 9030 7964 9036 8016
rect 9088 7964 9094 8016
rect 10689 8007 10747 8013
rect 10689 8004 10701 8007
rect 9784 7976 10701 8004
rect 9784 7936 9812 7976
rect 10689 7973 10701 7976
rect 10735 7973 10747 8007
rect 10689 7967 10747 7973
rect 10965 8007 11023 8013
rect 10965 7973 10977 8007
rect 11011 7973 11023 8007
rect 10965 7967 11023 7973
rect 10980 7936 11008 7967
rect 11054 7964 11060 8016
rect 11112 8004 11118 8016
rect 12069 8007 12127 8013
rect 12069 8004 12081 8007
rect 11112 7976 12081 8004
rect 11112 7964 11118 7976
rect 12069 7973 12081 7976
rect 12115 7973 12127 8007
rect 12069 7967 12127 7973
rect 15105 8007 15163 8013
rect 15105 7973 15117 8007
rect 15151 8004 15163 8007
rect 15304 8004 15332 8032
rect 15151 7976 15332 8004
rect 15933 8007 15991 8013
rect 15151 7973 15163 7976
rect 15105 7967 15163 7973
rect 15933 7973 15945 8007
rect 15979 8004 15991 8007
rect 16482 8004 16488 8016
rect 15979 7976 16488 8004
rect 15979 7973 15991 7976
rect 15933 7967 15991 7973
rect 16482 7964 16488 7976
rect 16540 7964 16546 8016
rect 5500 7908 8800 7936
rect 9232 7908 9812 7936
rect 9876 7908 11008 7936
rect 5500 7896 5506 7908
rect 3145 7871 3203 7877
rect 3145 7837 3157 7871
rect 3191 7837 3203 7871
rect 3145 7831 3203 7837
rect 4985 7871 5043 7877
rect 4985 7837 4997 7871
rect 5031 7868 5043 7871
rect 6638 7868 6644 7880
rect 5031 7840 6644 7868
rect 5031 7837 5043 7840
rect 4985 7831 5043 7837
rect 6638 7828 6644 7840
rect 6696 7828 6702 7880
rect 7193 7871 7251 7877
rect 7193 7837 7205 7871
rect 7239 7837 7251 7871
rect 7193 7831 7251 7837
rect 2041 7803 2099 7809
rect 2041 7769 2053 7803
rect 2087 7800 2099 7803
rect 2222 7800 2228 7812
rect 2087 7772 2228 7800
rect 2087 7769 2099 7772
rect 2041 7763 2099 7769
rect 2222 7760 2228 7772
rect 2280 7760 2286 7812
rect 3973 7803 4031 7809
rect 3973 7769 3985 7803
rect 4019 7769 4031 7803
rect 3973 7763 4031 7769
rect 4525 7803 4583 7809
rect 4525 7769 4537 7803
rect 4571 7800 4583 7803
rect 5534 7800 5540 7812
rect 4571 7772 5540 7800
rect 4571 7769 4583 7772
rect 4525 7763 4583 7769
rect 3988 7732 4016 7763
rect 5534 7760 5540 7772
rect 5592 7760 5598 7812
rect 5626 7760 5632 7812
rect 5684 7760 5690 7812
rect 6181 7803 6239 7809
rect 6181 7769 6193 7803
rect 6227 7800 6239 7803
rect 6546 7800 6552 7812
rect 6227 7772 6552 7800
rect 6227 7769 6239 7772
rect 6181 7763 6239 7769
rect 6546 7760 6552 7772
rect 6604 7760 6610 7812
rect 6730 7760 6736 7812
rect 6788 7760 6794 7812
rect 7208 7800 7236 7831
rect 7374 7828 7380 7880
rect 7432 7868 7438 7880
rect 7432 7840 7972 7868
rect 7432 7828 7438 7840
rect 7650 7800 7656 7812
rect 7208 7772 7656 7800
rect 7650 7760 7656 7772
rect 7708 7760 7714 7812
rect 7834 7760 7840 7812
rect 7892 7760 7898 7812
rect 7944 7800 7972 7840
rect 8478 7828 8484 7880
rect 8536 7828 8542 7880
rect 9232 7877 9260 7908
rect 9217 7871 9275 7877
rect 8588 7840 8984 7868
rect 8588 7800 8616 7840
rect 7944 7772 8616 7800
rect 8846 7732 8852 7744
rect 3988 7704 8852 7732
rect 8846 7692 8852 7704
rect 8904 7692 8910 7744
rect 8956 7732 8984 7840
rect 9217 7837 9229 7871
rect 9263 7837 9275 7871
rect 9217 7831 9275 7837
rect 9493 7871 9551 7877
rect 9493 7837 9505 7871
rect 9539 7868 9551 7871
rect 9582 7868 9588 7880
rect 9539 7840 9588 7868
rect 9539 7837 9551 7840
rect 9493 7831 9551 7837
rect 9582 7828 9588 7840
rect 9640 7828 9646 7880
rect 9766 7828 9772 7880
rect 9824 7828 9830 7880
rect 9876 7877 9904 7908
rect 16206 7896 16212 7948
rect 16264 7936 16270 7948
rect 16264 7908 18184 7936
rect 16264 7896 16270 7908
rect 9861 7871 9919 7877
rect 9861 7837 9873 7871
rect 9907 7837 9919 7871
rect 9861 7831 9919 7837
rect 10321 7871 10379 7877
rect 10321 7837 10333 7871
rect 10367 7837 10379 7871
rect 10321 7831 10379 7837
rect 9030 7760 9036 7812
rect 9088 7800 9094 7812
rect 10336 7800 10364 7831
rect 10594 7828 10600 7880
rect 10652 7828 10658 7880
rect 10870 7828 10876 7880
rect 10928 7828 10934 7880
rect 11146 7828 11152 7880
rect 11204 7828 11210 7880
rect 11422 7828 11428 7880
rect 11480 7828 11486 7880
rect 11698 7828 11704 7880
rect 11756 7828 11762 7880
rect 11974 7828 11980 7880
rect 12032 7868 12038 7880
rect 12253 7871 12311 7877
rect 12253 7868 12265 7871
rect 12032 7840 12265 7868
rect 12032 7828 12038 7840
rect 12253 7837 12265 7840
rect 12299 7837 12311 7871
rect 12253 7831 12311 7837
rect 12526 7828 12532 7880
rect 12584 7828 12590 7880
rect 12802 7828 12808 7880
rect 12860 7828 12866 7880
rect 13078 7828 13084 7880
rect 13136 7828 13142 7880
rect 13354 7828 13360 7880
rect 13412 7828 13418 7880
rect 14458 7828 14464 7880
rect 14516 7868 14522 7880
rect 14737 7871 14795 7877
rect 14737 7868 14749 7871
rect 14516 7840 14749 7868
rect 14516 7828 14522 7840
rect 14737 7837 14749 7840
rect 14783 7837 14795 7871
rect 14737 7831 14795 7837
rect 15010 7828 15016 7880
rect 15068 7828 15074 7880
rect 15286 7828 15292 7880
rect 15344 7828 15350 7880
rect 15562 7828 15568 7880
rect 15620 7828 15626 7880
rect 15838 7828 15844 7880
rect 15896 7828 15902 7880
rect 16114 7828 16120 7880
rect 16172 7828 16178 7880
rect 16390 7828 16396 7880
rect 16448 7828 16454 7880
rect 16666 7828 16672 7880
rect 16724 7868 16730 7880
rect 16945 7871 17003 7877
rect 16945 7868 16957 7871
rect 16724 7840 16957 7868
rect 16724 7828 16730 7840
rect 16945 7837 16957 7840
rect 16991 7837 17003 7871
rect 16945 7831 17003 7837
rect 17218 7828 17224 7880
rect 17276 7868 17282 7880
rect 17497 7871 17555 7877
rect 17497 7868 17509 7871
rect 17276 7840 17509 7868
rect 17276 7828 17282 7840
rect 17497 7837 17509 7840
rect 17543 7837 17555 7871
rect 17497 7831 17555 7837
rect 17770 7828 17776 7880
rect 17828 7868 17834 7880
rect 18049 7871 18107 7877
rect 18049 7868 18061 7871
rect 17828 7840 18061 7868
rect 17828 7828 17834 7840
rect 18049 7837 18061 7840
rect 18095 7837 18107 7871
rect 18049 7831 18107 7837
rect 18156 7800 18184 7908
rect 18322 7828 18328 7880
rect 18380 7828 18386 7880
rect 18417 7871 18475 7877
rect 18417 7837 18429 7871
rect 18463 7868 18475 7871
rect 18800 7868 18828 8044
rect 19518 8032 19524 8044
rect 19576 8032 19582 8084
rect 20806 8032 20812 8084
rect 20864 8072 20870 8084
rect 21269 8075 21327 8081
rect 21269 8072 21281 8075
rect 20864 8044 21281 8072
rect 20864 8032 20870 8044
rect 21269 8041 21281 8044
rect 21315 8041 21327 8075
rect 21269 8035 21327 8041
rect 21910 8032 21916 8084
rect 21968 8072 21974 8084
rect 22189 8075 22247 8081
rect 22189 8072 22201 8075
rect 21968 8044 22201 8072
rect 21968 8032 21974 8044
rect 22189 8041 22201 8044
rect 22235 8041 22247 8075
rect 22189 8035 22247 8041
rect 22278 8032 22284 8084
rect 22336 8072 22342 8084
rect 22741 8075 22799 8081
rect 22741 8072 22753 8075
rect 22336 8044 22753 8072
rect 22336 8032 22342 8044
rect 22741 8041 22753 8044
rect 22787 8041 22799 8075
rect 22741 8035 22799 8041
rect 22830 8032 22836 8084
rect 22888 8072 22894 8084
rect 23477 8075 23535 8081
rect 23477 8072 23489 8075
rect 22888 8044 23489 8072
rect 22888 8032 22894 8044
rect 23477 8041 23489 8044
rect 23523 8041 23535 8075
rect 23477 8035 23535 8041
rect 23845 8075 23903 8081
rect 23845 8041 23857 8075
rect 23891 8041 23903 8075
rect 23845 8035 23903 8041
rect 19245 8007 19303 8013
rect 19245 7973 19257 8007
rect 19291 7973 19303 8007
rect 19245 7967 19303 7973
rect 18463 7840 18828 7868
rect 18877 7871 18935 7877
rect 18463 7837 18475 7840
rect 18417 7831 18475 7837
rect 18877 7837 18889 7871
rect 18923 7868 18935 7871
rect 19260 7868 19288 7967
rect 23198 7964 23204 8016
rect 23256 8004 23262 8016
rect 23860 8004 23888 8035
rect 23256 7976 23888 8004
rect 23256 7964 23262 7976
rect 18923 7840 19288 7868
rect 18923 7837 18935 7840
rect 18877 7831 18935 7837
rect 19334 7828 19340 7880
rect 19392 7868 19398 7880
rect 19429 7871 19487 7877
rect 19429 7868 19441 7871
rect 19392 7840 19441 7868
rect 19392 7828 19398 7840
rect 19429 7837 19441 7840
rect 19475 7837 19487 7871
rect 19429 7831 19487 7837
rect 19518 7828 19524 7880
rect 19576 7828 19582 7880
rect 19794 7828 19800 7880
rect 19852 7828 19858 7880
rect 21085 7871 21143 7877
rect 21085 7837 21097 7871
rect 21131 7837 21143 7871
rect 21085 7831 21143 7837
rect 21913 7871 21971 7877
rect 21913 7837 21925 7871
rect 21959 7868 21971 7871
rect 25498 7868 25504 7880
rect 21959 7840 25504 7868
rect 21959 7837 21971 7840
rect 21913 7831 21971 7837
rect 21100 7800 21128 7831
rect 25498 7828 25504 7840
rect 25556 7828 25562 7880
rect 9088 7772 10272 7800
rect 10336 7772 11560 7800
rect 9088 7760 9094 7772
rect 10045 7735 10103 7741
rect 10045 7732 10057 7735
rect 8956 7704 10057 7732
rect 10045 7701 10057 7704
rect 10091 7701 10103 7735
rect 10045 7695 10103 7701
rect 10134 7692 10140 7744
rect 10192 7692 10198 7744
rect 10244 7732 10272 7772
rect 11532 7741 11560 7772
rect 12406 7772 17908 7800
rect 18156 7772 21128 7800
rect 21545 7803 21603 7809
rect 10413 7735 10471 7741
rect 10413 7732 10425 7735
rect 10244 7704 10425 7732
rect 10413 7701 10425 7704
rect 10459 7701 10471 7735
rect 10413 7695 10471 7701
rect 11517 7735 11575 7741
rect 11517 7701 11529 7735
rect 11563 7701 11575 7735
rect 11517 7695 11575 7701
rect 11606 7692 11612 7744
rect 11664 7732 11670 7744
rect 12406 7732 12434 7772
rect 11664 7704 12434 7732
rect 11664 7692 11670 7704
rect 16758 7692 16764 7744
rect 16816 7692 16822 7744
rect 17310 7692 17316 7744
rect 17368 7692 17374 7744
rect 17880 7741 17908 7772
rect 21545 7769 21557 7803
rect 21591 7800 21603 7803
rect 21591 7772 21956 7800
rect 21591 7769 21603 7772
rect 21545 7763 21603 7769
rect 17865 7735 17923 7741
rect 17865 7701 17877 7735
rect 17911 7701 17923 7735
rect 17865 7695 17923 7701
rect 18598 7692 18604 7744
rect 18656 7692 18662 7744
rect 19058 7692 19064 7744
rect 19116 7692 19122 7744
rect 19702 7692 19708 7744
rect 19760 7692 19766 7744
rect 19978 7692 19984 7744
rect 20036 7692 20042 7744
rect 21928 7732 21956 7772
rect 22094 7760 22100 7812
rect 22152 7760 22158 7812
rect 22646 7760 22652 7812
rect 22704 7760 22710 7812
rect 22738 7760 22744 7812
rect 22796 7800 22802 7812
rect 23201 7803 23259 7809
rect 23201 7800 23213 7803
rect 22796 7772 23213 7800
rect 22796 7760 22802 7772
rect 23201 7769 23213 7772
rect 23247 7769 23259 7803
rect 23201 7763 23259 7769
rect 23750 7760 23756 7812
rect 23808 7760 23814 7812
rect 22830 7732 22836 7744
rect 21928 7704 22836 7732
rect 22830 7692 22836 7704
rect 22888 7692 22894 7744
rect 1104 7642 24723 7664
rect 1104 7590 6814 7642
rect 6866 7590 6878 7642
rect 6930 7590 6942 7642
rect 6994 7590 7006 7642
rect 7058 7590 7070 7642
rect 7122 7590 12679 7642
rect 12731 7590 12743 7642
rect 12795 7590 12807 7642
rect 12859 7590 12871 7642
rect 12923 7590 12935 7642
rect 12987 7590 18544 7642
rect 18596 7590 18608 7642
rect 18660 7590 18672 7642
rect 18724 7590 18736 7642
rect 18788 7590 18800 7642
rect 18852 7590 24409 7642
rect 24461 7590 24473 7642
rect 24525 7590 24537 7642
rect 24589 7590 24601 7642
rect 24653 7590 24665 7642
rect 24717 7590 24723 7642
rect 1104 7568 24723 7590
rect 1670 7488 1676 7540
rect 1728 7488 1734 7540
rect 2225 7531 2283 7537
rect 2225 7497 2237 7531
rect 2271 7497 2283 7531
rect 2225 7491 2283 7497
rect 3513 7531 3571 7537
rect 3513 7497 3525 7531
rect 3559 7528 3571 7531
rect 3694 7528 3700 7540
rect 3559 7500 3700 7528
rect 3559 7497 3571 7500
rect 3513 7491 3571 7497
rect 1486 7420 1492 7472
rect 1544 7460 1550 7472
rect 2240 7460 2268 7491
rect 3694 7488 3700 7500
rect 3752 7488 3758 7540
rect 5445 7531 5503 7537
rect 5445 7497 5457 7531
rect 5491 7528 5503 7531
rect 5626 7528 5632 7540
rect 5491 7500 5632 7528
rect 5491 7497 5503 7500
rect 5445 7491 5503 7497
rect 5626 7488 5632 7500
rect 5684 7488 5690 7540
rect 5902 7488 5908 7540
rect 5960 7528 5966 7540
rect 6365 7531 6423 7537
rect 6365 7528 6377 7531
rect 5960 7500 6377 7528
rect 5960 7488 5966 7500
rect 6365 7497 6377 7500
rect 6411 7497 6423 7531
rect 6365 7491 6423 7497
rect 7190 7488 7196 7540
rect 7248 7528 7254 7540
rect 7653 7531 7711 7537
rect 7653 7528 7665 7531
rect 7248 7500 7665 7528
rect 7248 7488 7254 7500
rect 7653 7497 7665 7500
rect 7699 7497 7711 7531
rect 7653 7491 7711 7497
rect 8294 7488 8300 7540
rect 8352 7488 8358 7540
rect 8478 7488 8484 7540
rect 8536 7528 8542 7540
rect 8573 7531 8631 7537
rect 8573 7528 8585 7531
rect 8536 7500 8585 7528
rect 8536 7488 8542 7500
rect 8573 7497 8585 7500
rect 8619 7497 8631 7531
rect 16758 7528 16764 7540
rect 8573 7491 8631 7497
rect 8772 7500 16764 7528
rect 5994 7460 6000 7472
rect 1544 7432 2268 7460
rect 2608 7432 6000 7460
rect 1544 7420 1550 7432
rect 1578 7352 1584 7404
rect 1636 7352 1642 7404
rect 2133 7395 2191 7401
rect 2133 7361 2145 7395
rect 2179 7392 2191 7395
rect 2608 7392 2636 7432
rect 5994 7420 6000 7432
rect 6052 7420 6058 7472
rect 8496 7405 8616 7416
rect 2179 7364 2636 7392
rect 2685 7395 2743 7401
rect 2179 7361 2191 7364
rect 2133 7355 2191 7361
rect 2685 7361 2697 7395
rect 2731 7361 2743 7395
rect 2685 7355 2743 7361
rect 3329 7395 3387 7401
rect 3329 7361 3341 7395
rect 3375 7361 3387 7395
rect 3329 7355 3387 7361
rect 2700 7324 2728 7355
rect 3344 7324 3372 7355
rect 5626 7352 5632 7404
rect 5684 7352 5690 7404
rect 6178 7352 6184 7404
rect 6236 7352 6242 7404
rect 6362 7352 6368 7404
rect 6420 7392 6426 7404
rect 6549 7395 6607 7401
rect 6549 7392 6561 7395
rect 6420 7364 6561 7392
rect 6420 7352 6426 7364
rect 6549 7361 6561 7364
rect 6595 7361 6607 7395
rect 6549 7355 6607 7361
rect 7374 7352 7380 7404
rect 7432 7352 7438 7404
rect 7837 7395 7895 7401
rect 7837 7361 7849 7395
rect 7883 7392 7895 7395
rect 8386 7392 8392 7404
rect 7883 7364 8392 7392
rect 7883 7361 7895 7364
rect 7837 7355 7895 7361
rect 8386 7352 8392 7364
rect 8444 7352 8450 7404
rect 8481 7399 8616 7405
rect 8481 7365 8493 7399
rect 8527 7388 8616 7399
rect 8527 7365 8539 7388
rect 8481 7359 8539 7365
rect 8202 7324 8208 7336
rect 2700 7296 2774 7324
rect 3344 7296 8208 7324
rect 2746 7256 2774 7296
rect 8202 7284 8208 7296
rect 8260 7284 8266 7336
rect 7193 7259 7251 7265
rect 7193 7256 7205 7259
rect 2746 7228 7205 7256
rect 7193 7225 7205 7228
rect 7239 7225 7251 7259
rect 8588 7256 8616 7388
rect 8662 7352 8668 7404
rect 8720 7352 8726 7404
rect 8772 7401 8800 7500
rect 16758 7488 16764 7500
rect 16816 7488 16822 7540
rect 17310 7488 17316 7540
rect 17368 7488 17374 7540
rect 23845 7531 23903 7537
rect 23845 7497 23857 7531
rect 23891 7528 23903 7531
rect 24118 7528 24124 7540
rect 23891 7500 24124 7528
rect 23891 7497 23903 7500
rect 23845 7491 23903 7497
rect 24118 7488 24124 7500
rect 24176 7488 24182 7540
rect 24762 7488 24768 7540
rect 24820 7488 24826 7540
rect 8846 7420 8852 7472
rect 8904 7460 8910 7472
rect 11790 7460 11796 7472
rect 8904 7432 11796 7460
rect 8904 7420 8910 7432
rect 11790 7420 11796 7432
rect 11848 7420 11854 7472
rect 8757 7395 8815 7401
rect 8757 7361 8769 7395
rect 8803 7361 8815 7395
rect 8757 7355 8815 7361
rect 9232 7392 9352 7396
rect 9508 7392 9674 7396
rect 9232 7368 9674 7392
rect 8680 7324 8708 7352
rect 9232 7324 9260 7368
rect 9324 7364 9536 7368
rect 8680 7296 9260 7324
rect 9646 7324 9674 7368
rect 10318 7352 10324 7404
rect 10376 7352 10382 7404
rect 11606 7324 11612 7336
rect 9646 7296 11612 7324
rect 11606 7284 11612 7296
rect 11664 7284 11670 7336
rect 9306 7256 9312 7268
rect 8588 7228 9312 7256
rect 7193 7219 7251 7225
rect 9306 7216 9312 7228
rect 9364 7216 9370 7268
rect 9490 7216 9496 7268
rect 9548 7256 9554 7268
rect 17328 7256 17356 7488
rect 23385 7463 23443 7469
rect 23385 7429 23397 7463
rect 23431 7460 23443 7463
rect 24780 7460 24808 7488
rect 23431 7432 24808 7460
rect 23431 7429 23443 7432
rect 23385 7423 23443 7429
rect 17402 7352 17408 7404
rect 17460 7352 17466 7404
rect 22462 7352 22468 7404
rect 22520 7352 22526 7404
rect 23014 7352 23020 7404
rect 23072 7352 23078 7404
rect 23566 7352 23572 7404
rect 23624 7352 23630 7404
rect 22741 7327 22799 7333
rect 22741 7293 22753 7327
rect 22787 7324 22799 7327
rect 24946 7324 24952 7336
rect 22787 7296 24952 7324
rect 22787 7293 22799 7296
rect 22741 7287 22799 7293
rect 24946 7284 24952 7296
rect 25004 7284 25010 7336
rect 9548 7228 17356 7256
rect 9548 7216 9554 7228
rect 2774 7148 2780 7200
rect 2832 7148 2838 7200
rect 5810 7148 5816 7200
rect 5868 7188 5874 7200
rect 5997 7191 6055 7197
rect 5997 7188 6009 7191
rect 5868 7160 6009 7188
rect 5868 7148 5874 7160
rect 5997 7157 6009 7160
rect 6043 7157 6055 7191
rect 5997 7151 6055 7157
rect 7374 7148 7380 7200
rect 7432 7188 7438 7200
rect 9030 7188 9036 7200
rect 7432 7160 9036 7188
rect 7432 7148 7438 7160
rect 9030 7148 9036 7160
rect 9088 7148 9094 7200
rect 9628 7148 9634 7200
rect 9686 7188 9692 7200
rect 10137 7191 10195 7197
rect 10137 7188 10149 7191
rect 9686 7160 10149 7188
rect 9686 7148 9692 7160
rect 10137 7157 10149 7160
rect 10183 7157 10195 7191
rect 10137 7151 10195 7157
rect 17221 7191 17279 7197
rect 17221 7157 17233 7191
rect 17267 7188 17279 7191
rect 22094 7188 22100 7200
rect 17267 7160 22100 7188
rect 17267 7157 17279 7160
rect 17221 7151 17279 7157
rect 22094 7148 22100 7160
rect 22152 7148 22158 7200
rect 1104 7098 24564 7120
rect 1104 7046 3882 7098
rect 3934 7046 3946 7098
rect 3998 7046 4010 7098
rect 4062 7046 4074 7098
rect 4126 7046 4138 7098
rect 4190 7046 9747 7098
rect 9799 7046 9811 7098
rect 9863 7046 9875 7098
rect 9927 7046 9939 7098
rect 9991 7046 10003 7098
rect 10055 7046 15612 7098
rect 15664 7046 15676 7098
rect 15728 7046 15740 7098
rect 15792 7046 15804 7098
rect 15856 7046 15868 7098
rect 15920 7046 21477 7098
rect 21529 7046 21541 7098
rect 21593 7046 21605 7098
rect 21657 7046 21669 7098
rect 21721 7046 21733 7098
rect 21785 7046 24564 7098
rect 1104 7024 24564 7046
rect 6546 6944 6552 6996
rect 6604 6984 6610 6996
rect 16669 6987 16727 6993
rect 6604 6956 12434 6984
rect 6604 6944 6610 6956
rect 12406 6916 12434 6956
rect 16669 6953 16681 6987
rect 16715 6984 16727 6987
rect 17402 6984 17408 6996
rect 16715 6956 17408 6984
rect 16715 6953 16727 6956
rect 16669 6947 16727 6953
rect 17402 6944 17408 6956
rect 17460 6944 17466 6996
rect 19058 6944 19064 6996
rect 19116 6944 19122 6996
rect 19076 6916 19104 6944
rect 12406 6888 19104 6916
rect 658 6808 664 6860
rect 716 6848 722 6860
rect 2774 6848 2780 6860
rect 716 6820 2780 6848
rect 716 6808 722 6820
rect 2774 6808 2780 6820
rect 2832 6808 2838 6860
rect 23937 6851 23995 6857
rect 23937 6817 23949 6851
rect 23983 6848 23995 6851
rect 24302 6848 24308 6860
rect 23983 6820 24308 6848
rect 23983 6817 23995 6820
rect 23937 6811 23995 6817
rect 24302 6808 24308 6820
rect 24360 6808 24366 6860
rect 1210 6740 1216 6792
rect 1268 6780 1274 6792
rect 1949 6783 2007 6789
rect 1949 6780 1961 6783
rect 1268 6752 1961 6780
rect 1268 6740 1274 6752
rect 1949 6749 1961 6752
rect 1995 6749 2007 6783
rect 1949 6743 2007 6749
rect 16850 6740 16856 6792
rect 16908 6740 16914 6792
rect 23477 6783 23535 6789
rect 23477 6749 23489 6783
rect 23523 6780 23535 6783
rect 23523 6752 23980 6780
rect 23523 6749 23535 6752
rect 23477 6743 23535 6749
rect 23952 6724 23980 6752
rect 1673 6715 1731 6721
rect 1673 6681 1685 6715
rect 1719 6712 1731 6715
rect 2317 6715 2375 6721
rect 2317 6712 2329 6715
rect 1719 6684 2329 6712
rect 1719 6681 1731 6684
rect 1673 6675 1731 6681
rect 2317 6681 2329 6684
rect 2363 6712 2375 6715
rect 2682 6712 2688 6724
rect 2363 6684 2688 6712
rect 2363 6681 2375 6684
rect 2317 6675 2375 6681
rect 2682 6672 2688 6684
rect 2740 6672 2746 6724
rect 23106 6672 23112 6724
rect 23164 6672 23170 6724
rect 23382 6672 23388 6724
rect 23440 6712 23446 6724
rect 23661 6715 23719 6721
rect 23661 6712 23673 6715
rect 23440 6684 23673 6712
rect 23440 6672 23446 6684
rect 23661 6681 23673 6684
rect 23707 6681 23719 6715
rect 23661 6675 23719 6681
rect 23934 6672 23940 6724
rect 23992 6672 23998 6724
rect 1104 6554 24723 6576
rect 1104 6502 6814 6554
rect 6866 6502 6878 6554
rect 6930 6502 6942 6554
rect 6994 6502 7006 6554
rect 7058 6502 7070 6554
rect 7122 6502 12679 6554
rect 12731 6502 12743 6554
rect 12795 6502 12807 6554
rect 12859 6502 12871 6554
rect 12923 6502 12935 6554
rect 12987 6502 18544 6554
rect 18596 6502 18608 6554
rect 18660 6502 18672 6554
rect 18724 6502 18736 6554
rect 18788 6502 18800 6554
rect 18852 6502 24409 6554
rect 24461 6502 24473 6554
rect 24525 6502 24537 6554
rect 24589 6502 24601 6554
rect 24653 6502 24665 6554
rect 24717 6502 24723 6554
rect 1104 6480 24723 6502
rect 934 6400 940 6452
rect 992 6440 998 6452
rect 1581 6443 1639 6449
rect 1581 6440 1593 6443
rect 992 6412 1593 6440
rect 992 6400 998 6412
rect 1581 6409 1593 6412
rect 1627 6409 1639 6443
rect 1581 6403 1639 6409
rect 23290 6400 23296 6452
rect 23348 6400 23354 6452
rect 23842 6400 23848 6452
rect 23900 6400 23906 6452
rect 1489 6375 1547 6381
rect 1489 6341 1501 6375
rect 1535 6372 1547 6375
rect 5442 6372 5448 6384
rect 1535 6344 5448 6372
rect 1535 6341 1547 6344
rect 1489 6335 1547 6341
rect 5442 6332 5448 6344
rect 5500 6332 5506 6384
rect 22094 6332 22100 6384
rect 22152 6372 22158 6384
rect 23753 6375 23811 6381
rect 23753 6372 23765 6375
rect 22152 6344 23765 6372
rect 22152 6332 22158 6344
rect 23753 6341 23765 6344
rect 23799 6341 23811 6375
rect 23753 6335 23811 6341
rect 23198 6264 23204 6316
rect 23256 6264 23262 6316
rect 1104 6010 24564 6032
rect 1104 5958 3882 6010
rect 3934 5958 3946 6010
rect 3998 5958 4010 6010
rect 4062 5958 4074 6010
rect 4126 5958 4138 6010
rect 4190 5958 9747 6010
rect 9799 5958 9811 6010
rect 9863 5958 9875 6010
rect 9927 5958 9939 6010
rect 9991 5958 10003 6010
rect 10055 5958 15612 6010
rect 15664 5958 15676 6010
rect 15728 5958 15740 6010
rect 15792 5958 15804 6010
rect 15856 5958 15868 6010
rect 15920 5958 21477 6010
rect 21529 5958 21541 6010
rect 21593 5958 21605 6010
rect 21657 5958 21669 6010
rect 21721 5958 21733 6010
rect 21785 5958 24564 6010
rect 1104 5936 24564 5958
rect 24121 5899 24179 5905
rect 24121 5865 24133 5899
rect 24167 5896 24179 5899
rect 25222 5896 25228 5908
rect 24167 5868 25228 5896
rect 24167 5865 24179 5868
rect 24121 5859 24179 5865
rect 25222 5856 25228 5868
rect 25280 5856 25286 5908
rect 23842 5584 23848 5636
rect 23900 5584 23906 5636
rect 1104 5466 24723 5488
rect 1104 5414 6814 5466
rect 6866 5414 6878 5466
rect 6930 5414 6942 5466
rect 6994 5414 7006 5466
rect 7058 5414 7070 5466
rect 7122 5414 12679 5466
rect 12731 5414 12743 5466
rect 12795 5414 12807 5466
rect 12859 5414 12871 5466
rect 12923 5414 12935 5466
rect 12987 5414 18544 5466
rect 18596 5414 18608 5466
rect 18660 5414 18672 5466
rect 18724 5414 18736 5466
rect 18788 5414 18800 5466
rect 18852 5414 24409 5466
rect 24461 5414 24473 5466
rect 24525 5414 24537 5466
rect 24589 5414 24601 5466
rect 24653 5414 24665 5466
rect 24717 5414 24723 5466
rect 1104 5392 24723 5414
rect 1104 4922 24564 4944
rect 1104 4870 3882 4922
rect 3934 4870 3946 4922
rect 3998 4870 4010 4922
rect 4062 4870 4074 4922
rect 4126 4870 4138 4922
rect 4190 4870 9747 4922
rect 9799 4870 9811 4922
rect 9863 4870 9875 4922
rect 9927 4870 9939 4922
rect 9991 4870 10003 4922
rect 10055 4870 15612 4922
rect 15664 4870 15676 4922
rect 15728 4870 15740 4922
rect 15792 4870 15804 4922
rect 15856 4870 15868 4922
rect 15920 4870 21477 4922
rect 21529 4870 21541 4922
rect 21593 4870 21605 4922
rect 21657 4870 21669 4922
rect 21721 4870 21733 4922
rect 21785 4870 24564 4922
rect 1104 4848 24564 4870
rect 14826 4564 14832 4616
rect 14884 4564 14890 4616
rect 15013 4471 15071 4477
rect 15013 4437 15025 4471
rect 15059 4468 15071 4471
rect 23474 4468 23480 4480
rect 15059 4440 23480 4468
rect 15059 4437 15071 4440
rect 15013 4431 15071 4437
rect 23474 4428 23480 4440
rect 23532 4428 23538 4480
rect 1104 4378 24723 4400
rect 1104 4326 6814 4378
rect 6866 4326 6878 4378
rect 6930 4326 6942 4378
rect 6994 4326 7006 4378
rect 7058 4326 7070 4378
rect 7122 4326 12679 4378
rect 12731 4326 12743 4378
rect 12795 4326 12807 4378
rect 12859 4326 12871 4378
rect 12923 4326 12935 4378
rect 12987 4326 18544 4378
rect 18596 4326 18608 4378
rect 18660 4326 18672 4378
rect 18724 4326 18736 4378
rect 18788 4326 18800 4378
rect 18852 4326 24409 4378
rect 24461 4326 24473 4378
rect 24525 4326 24537 4378
rect 24589 4326 24601 4378
rect 24653 4326 24665 4378
rect 24717 4326 24723 4378
rect 1104 4304 24723 4326
rect 14277 4267 14335 4273
rect 14277 4233 14289 4267
rect 14323 4264 14335 4267
rect 14826 4264 14832 4276
rect 14323 4236 14832 4264
rect 14323 4233 14335 4236
rect 14277 4227 14335 4233
rect 14826 4224 14832 4236
rect 14884 4224 14890 4276
rect 14458 4088 14464 4140
rect 14516 4088 14522 4140
rect 1104 3834 24564 3856
rect 1104 3782 3882 3834
rect 3934 3782 3946 3834
rect 3998 3782 4010 3834
rect 4062 3782 4074 3834
rect 4126 3782 4138 3834
rect 4190 3782 9747 3834
rect 9799 3782 9811 3834
rect 9863 3782 9875 3834
rect 9927 3782 9939 3834
rect 9991 3782 10003 3834
rect 10055 3782 15612 3834
rect 15664 3782 15676 3834
rect 15728 3782 15740 3834
rect 15792 3782 15804 3834
rect 15856 3782 15868 3834
rect 15920 3782 21477 3834
rect 21529 3782 21541 3834
rect 21593 3782 21605 3834
rect 21657 3782 21669 3834
rect 21721 3782 21733 3834
rect 21785 3782 24564 3834
rect 1104 3760 24564 3782
rect 23106 3680 23112 3732
rect 23164 3720 23170 3732
rect 23293 3723 23351 3729
rect 23293 3720 23305 3723
rect 23164 3692 23305 3720
rect 23164 3680 23170 3692
rect 23293 3689 23305 3692
rect 23339 3689 23351 3723
rect 23293 3683 23351 3689
rect 17770 3476 17776 3528
rect 17828 3516 17834 3528
rect 18049 3519 18107 3525
rect 18049 3516 18061 3519
rect 17828 3488 18061 3516
rect 17828 3476 17834 3488
rect 18049 3485 18061 3488
rect 18095 3485 18107 3519
rect 18049 3479 18107 3485
rect 23477 3519 23535 3525
rect 23477 3485 23489 3519
rect 23523 3485 23535 3519
rect 23477 3479 23535 3485
rect 23492 3448 23520 3479
rect 22066 3420 23520 3448
rect 17865 3383 17923 3389
rect 17865 3349 17877 3383
rect 17911 3380 17923 3383
rect 22066 3380 22094 3420
rect 17911 3352 22094 3380
rect 17911 3349 17923 3352
rect 17865 3343 17923 3349
rect 1104 3290 24723 3312
rect 1104 3238 6814 3290
rect 6866 3238 6878 3290
rect 6930 3238 6942 3290
rect 6994 3238 7006 3290
rect 7058 3238 7070 3290
rect 7122 3238 12679 3290
rect 12731 3238 12743 3290
rect 12795 3238 12807 3290
rect 12859 3238 12871 3290
rect 12923 3238 12935 3290
rect 12987 3238 18544 3290
rect 18596 3238 18608 3290
rect 18660 3238 18672 3290
rect 18724 3238 18736 3290
rect 18788 3238 18800 3290
rect 18852 3238 24409 3290
rect 24461 3238 24473 3290
rect 24525 3238 24537 3290
rect 24589 3238 24601 3290
rect 24653 3238 24665 3290
rect 24717 3238 24723 3290
rect 1104 3216 24723 3238
rect 22462 3136 22468 3188
rect 22520 3176 22526 3188
rect 23293 3179 23351 3185
rect 23293 3176 23305 3179
rect 22520 3148 23305 3176
rect 22520 3136 22526 3148
rect 23293 3145 23305 3148
rect 23339 3145 23351 3179
rect 23293 3139 23351 3145
rect 23845 3179 23903 3185
rect 23845 3145 23857 3179
rect 23891 3145 23903 3179
rect 23845 3139 23903 3145
rect 22830 3068 22836 3120
rect 22888 3108 22894 3120
rect 23860 3108 23888 3139
rect 22888 3080 23888 3108
rect 22888 3068 22894 3080
rect 22462 3000 22468 3052
rect 22520 3040 22526 3052
rect 22925 3043 22983 3049
rect 22925 3040 22937 3043
rect 22520 3012 22937 3040
rect 22520 3000 22526 3012
rect 22925 3009 22937 3012
rect 22971 3009 22983 3043
rect 22925 3003 22983 3009
rect 23477 3043 23535 3049
rect 23477 3009 23489 3043
rect 23523 3009 23535 3043
rect 23477 3003 23535 3009
rect 23492 2972 23520 3003
rect 24026 3000 24032 3052
rect 24084 3000 24090 3052
rect 22756 2944 23520 2972
rect 22756 2913 22784 2944
rect 22741 2907 22799 2913
rect 22741 2873 22753 2907
rect 22787 2873 22799 2907
rect 22741 2867 22799 2873
rect 1104 2746 24564 2768
rect 1104 2694 3882 2746
rect 3934 2694 3946 2746
rect 3998 2694 4010 2746
rect 4062 2694 4074 2746
rect 4126 2694 4138 2746
rect 4190 2694 9747 2746
rect 9799 2694 9811 2746
rect 9863 2694 9875 2746
rect 9927 2694 9939 2746
rect 9991 2694 10003 2746
rect 10055 2694 15612 2746
rect 15664 2694 15676 2746
rect 15728 2694 15740 2746
rect 15792 2694 15804 2746
rect 15856 2694 15868 2746
rect 15920 2694 21477 2746
rect 21529 2694 21541 2746
rect 21593 2694 21605 2746
rect 21657 2694 21669 2746
rect 21721 2694 21733 2746
rect 21785 2694 24564 2746
rect 1104 2672 24564 2694
rect 23845 2635 23903 2641
rect 23845 2601 23857 2635
rect 23891 2632 23903 2635
rect 24026 2632 24032 2644
rect 23891 2604 24032 2632
rect 23891 2601 23903 2604
rect 23845 2595 23903 2601
rect 24026 2592 24032 2604
rect 24084 2592 24090 2644
rect 23290 2388 23296 2440
rect 23348 2428 23354 2440
rect 24029 2431 24087 2437
rect 24029 2428 24041 2431
rect 23348 2400 24041 2428
rect 23348 2388 23354 2400
rect 24029 2397 24041 2400
rect 24075 2397 24087 2431
rect 24029 2391 24087 2397
rect 13814 2320 13820 2372
rect 13872 2360 13878 2372
rect 23750 2360 23756 2372
rect 13872 2332 23756 2360
rect 13872 2320 13878 2332
rect 23750 2320 23756 2332
rect 23808 2320 23814 2372
rect 10410 2252 10416 2304
rect 10468 2292 10474 2304
rect 21174 2292 21180 2304
rect 10468 2264 21180 2292
rect 10468 2252 10474 2264
rect 21174 2252 21180 2264
rect 21232 2252 21238 2304
rect 1104 2202 24723 2224
rect 1104 2150 6814 2202
rect 6866 2150 6878 2202
rect 6930 2150 6942 2202
rect 6994 2150 7006 2202
rect 7058 2150 7070 2202
rect 7122 2150 12679 2202
rect 12731 2150 12743 2202
rect 12795 2150 12807 2202
rect 12859 2150 12871 2202
rect 12923 2150 12935 2202
rect 12987 2150 18544 2202
rect 18596 2150 18608 2202
rect 18660 2150 18672 2202
rect 18724 2150 18736 2202
rect 18788 2150 18800 2202
rect 18852 2150 24409 2202
rect 24461 2150 24473 2202
rect 24525 2150 24537 2202
rect 24589 2150 24601 2202
rect 24653 2150 24665 2202
rect 24717 2150 24723 2202
rect 1104 2128 24723 2150
rect 9030 2048 9036 2100
rect 9088 2048 9094 2100
rect 10410 2048 10416 2100
rect 10468 2048 10474 2100
rect 10686 2048 10692 2100
rect 10744 2048 10750 2100
rect 11514 2048 11520 2100
rect 11572 2088 11578 2100
rect 11701 2091 11759 2097
rect 11701 2088 11713 2091
rect 11572 2060 11713 2088
rect 11572 2048 11578 2060
rect 11701 2057 11713 2060
rect 11747 2057 11759 2091
rect 11701 2051 11759 2057
rect 12621 2091 12679 2097
rect 12621 2057 12633 2091
rect 12667 2057 12679 2091
rect 12621 2051 12679 2057
rect 12989 2091 13047 2097
rect 12989 2057 13001 2091
rect 13035 2057 13047 2091
rect 12989 2051 13047 2057
rect 7650 1912 7656 1964
rect 7708 1912 7714 1964
rect 8846 1912 8852 1964
rect 8904 1912 8910 1964
rect 10226 1912 10232 1964
rect 10284 1912 10290 1964
rect 10502 1912 10508 1964
rect 10560 1912 10566 1964
rect 11514 1912 11520 1964
rect 11572 1912 11578 1964
rect 11790 1912 11796 1964
rect 11848 1912 11854 1964
rect 12434 1912 12440 1964
rect 12492 1912 12498 1964
rect 12636 1884 12664 2051
rect 13004 2020 13032 2051
rect 13814 2048 13820 2100
rect 13872 2048 13878 2100
rect 14277 2091 14335 2097
rect 14277 2057 14289 2091
rect 14323 2088 14335 2091
rect 20714 2088 20720 2100
rect 14323 2060 20720 2088
rect 14323 2057 14335 2060
rect 14277 2051 14335 2057
rect 20714 2048 20720 2060
rect 20772 2048 20778 2100
rect 22005 2091 22063 2097
rect 22005 2057 22017 2091
rect 22051 2088 22063 2091
rect 23014 2088 23020 2100
rect 22051 2060 23020 2088
rect 22051 2057 22063 2060
rect 22005 2051 22063 2057
rect 23014 2048 23020 2060
rect 23072 2048 23078 2100
rect 23198 2048 23204 2100
rect 23256 2048 23262 2100
rect 23382 2048 23388 2100
rect 23440 2048 23446 2100
rect 23566 2048 23572 2100
rect 23624 2088 23630 2100
rect 23661 2091 23719 2097
rect 23661 2088 23673 2091
rect 23624 2060 23673 2088
rect 23624 2048 23630 2060
rect 23661 2057 23673 2060
rect 23707 2057 23719 2091
rect 23661 2051 23719 2057
rect 23842 2048 23848 2100
rect 23900 2088 23906 2100
rect 23937 2091 23995 2097
rect 23937 2088 23949 2091
rect 23900 2060 23949 2088
rect 23900 2048 23906 2060
rect 23937 2057 23949 2060
rect 23983 2057 23995 2091
rect 23937 2051 23995 2057
rect 16206 2020 16212 2032
rect 13004 1992 16212 2020
rect 16206 1980 16212 1992
rect 16264 1980 16270 2032
rect 23216 2020 23244 2048
rect 16546 1992 23244 2020
rect 12802 1912 12808 1964
rect 12860 1912 12866 1964
rect 13630 1912 13636 1964
rect 13688 1912 13694 1964
rect 14090 1912 14096 1964
rect 14148 1912 14154 1964
rect 16114 1912 16120 1964
rect 16172 1912 16178 1964
rect 16298 1912 16304 1964
rect 16356 1952 16362 1964
rect 16546 1952 16574 1992
rect 16356 1924 16574 1952
rect 16356 1912 16362 1924
rect 22186 1912 22192 1964
rect 22244 1912 22250 1964
rect 22830 1912 22836 1964
rect 22888 1952 22894 1964
rect 23569 1955 23627 1961
rect 23569 1952 23581 1955
rect 22888 1924 23581 1952
rect 22888 1912 22894 1924
rect 23569 1921 23581 1924
rect 23615 1921 23627 1955
rect 23569 1915 23627 1921
rect 23845 1955 23903 1961
rect 23845 1921 23857 1955
rect 23891 1921 23903 1955
rect 23845 1915 23903 1921
rect 22738 1884 22744 1896
rect 12636 1856 22744 1884
rect 22738 1844 22744 1856
rect 22796 1844 22802 1896
rect 23106 1844 23112 1896
rect 23164 1884 23170 1896
rect 23860 1884 23888 1915
rect 24118 1912 24124 1964
rect 24176 1912 24182 1964
rect 23164 1856 23888 1884
rect 23164 1844 23170 1856
rect 7834 1776 7840 1828
rect 7892 1776 7898 1828
rect 11977 1819 12035 1825
rect 11977 1785 11989 1819
rect 12023 1816 12035 1819
rect 22646 1816 22652 1828
rect 12023 1788 22652 1816
rect 12023 1785 12035 1788
rect 11977 1779 12035 1785
rect 22646 1776 22652 1788
rect 22704 1776 22710 1828
rect 16298 1708 16304 1760
rect 16356 1708 16362 1760
rect 1104 1658 24564 1680
rect 1104 1606 3882 1658
rect 3934 1606 3946 1658
rect 3998 1606 4010 1658
rect 4062 1606 4074 1658
rect 4126 1606 4138 1658
rect 4190 1606 9747 1658
rect 9799 1606 9811 1658
rect 9863 1606 9875 1658
rect 9927 1606 9939 1658
rect 9991 1606 10003 1658
rect 10055 1606 15612 1658
rect 15664 1606 15676 1658
rect 15728 1606 15740 1658
rect 15792 1606 15804 1658
rect 15856 1606 15868 1658
rect 15920 1606 21477 1658
rect 21529 1606 21541 1658
rect 21593 1606 21605 1658
rect 21657 1606 21669 1658
rect 21721 1606 21733 1658
rect 21785 1606 24564 1658
rect 1104 1584 24564 1606
rect 7101 1547 7159 1553
rect 7101 1513 7113 1547
rect 7147 1544 7159 1547
rect 7650 1544 7656 1556
rect 7147 1516 7656 1544
rect 7147 1513 7159 1516
rect 7101 1507 7159 1513
rect 7650 1504 7656 1516
rect 7708 1504 7714 1556
rect 8297 1547 8355 1553
rect 8297 1513 8309 1547
rect 8343 1544 8355 1547
rect 8846 1544 8852 1556
rect 8343 1516 8852 1544
rect 8343 1513 8355 1516
rect 8297 1507 8355 1513
rect 8846 1504 8852 1516
rect 8904 1504 8910 1556
rect 9677 1547 9735 1553
rect 9677 1513 9689 1547
rect 9723 1544 9735 1547
rect 10226 1544 10232 1556
rect 9723 1516 10232 1544
rect 9723 1513 9735 1516
rect 9677 1507 9735 1513
rect 10226 1504 10232 1516
rect 10284 1504 10290 1556
rect 10502 1504 10508 1556
rect 10560 1504 10566 1556
rect 11057 1547 11115 1553
rect 11057 1513 11069 1547
rect 11103 1544 11115 1547
rect 11514 1544 11520 1556
rect 11103 1516 11520 1544
rect 11103 1513 11115 1516
rect 11057 1507 11115 1513
rect 11514 1504 11520 1516
rect 11572 1504 11578 1556
rect 12345 1547 12403 1553
rect 12345 1513 12357 1547
rect 12391 1544 12403 1547
rect 12802 1544 12808 1556
rect 12391 1516 12808 1544
rect 12391 1513 12403 1516
rect 12345 1507 12403 1513
rect 12802 1504 12808 1516
rect 12860 1504 12866 1556
rect 13081 1547 13139 1553
rect 13081 1513 13093 1547
rect 13127 1544 13139 1547
rect 13630 1544 13636 1556
rect 13127 1516 13636 1544
rect 13127 1513 13139 1516
rect 13081 1507 13139 1513
rect 13630 1504 13636 1516
rect 13688 1504 13694 1556
rect 15565 1547 15623 1553
rect 15565 1513 15577 1547
rect 15611 1544 15623 1547
rect 16114 1544 16120 1556
rect 15611 1516 16120 1544
rect 15611 1513 15623 1516
rect 15565 1507 15623 1513
rect 16114 1504 16120 1516
rect 16172 1504 16178 1556
rect 21821 1547 21879 1553
rect 21821 1513 21833 1547
rect 21867 1544 21879 1547
rect 22186 1544 22192 1556
rect 21867 1516 22192 1544
rect 21867 1513 21879 1516
rect 21821 1507 21879 1513
rect 22186 1504 22192 1516
rect 22244 1504 22250 1556
rect 22830 1504 22836 1556
rect 22888 1504 22894 1556
rect 23106 1504 23112 1556
rect 23164 1504 23170 1556
rect 23290 1504 23296 1556
rect 23348 1544 23354 1556
rect 23385 1547 23443 1553
rect 23385 1544 23397 1547
rect 23348 1516 23397 1544
rect 23348 1504 23354 1516
rect 23385 1513 23397 1516
rect 23431 1513 23443 1547
rect 23385 1507 23443 1513
rect 23661 1547 23719 1553
rect 23661 1513 23673 1547
rect 23707 1544 23719 1547
rect 24118 1544 24124 1556
rect 23707 1516 24124 1544
rect 23707 1513 23719 1516
rect 23661 1507 23719 1513
rect 24118 1504 24124 1516
rect 24176 1504 24182 1556
rect 9953 1479 10011 1485
rect 9953 1445 9965 1479
rect 9999 1476 10011 1479
rect 10520 1476 10548 1504
rect 9999 1448 10548 1476
rect 21269 1479 21327 1485
rect 9999 1445 10011 1448
rect 9953 1439 10011 1445
rect 21269 1445 21281 1479
rect 21315 1445 21327 1479
rect 21269 1439 21327 1445
rect 842 1300 848 1352
rect 900 1340 906 1352
rect 1397 1343 1455 1349
rect 1397 1340 1409 1343
rect 900 1312 1409 1340
rect 900 1300 906 1312
rect 1397 1309 1409 1312
rect 1443 1309 1455 1343
rect 1397 1303 1455 1309
rect 2130 1300 2136 1352
rect 2188 1300 2194 1352
rect 3326 1300 3332 1352
rect 3384 1300 3390 1352
rect 4706 1300 4712 1352
rect 4764 1300 4770 1352
rect 5902 1300 5908 1352
rect 5960 1300 5966 1352
rect 7285 1343 7343 1349
rect 7285 1309 7297 1343
rect 7331 1340 7343 1343
rect 7331 1312 7420 1340
rect 7331 1309 7343 1312
rect 7285 1303 7343 1309
rect 3528 1244 6914 1272
rect 1578 1164 1584 1216
rect 1636 1164 1642 1216
rect 2314 1164 2320 1216
rect 2372 1164 2378 1216
rect 3528 1213 3556 1244
rect 3513 1207 3571 1213
rect 3513 1173 3525 1207
rect 3559 1173 3571 1207
rect 3513 1167 3571 1173
rect 4522 1164 4528 1216
rect 4580 1164 4586 1216
rect 5718 1164 5724 1216
rect 5776 1164 5782 1216
rect 6886 1204 6914 1244
rect 7282 1204 7288 1216
rect 6886 1176 7288 1204
rect 7282 1164 7288 1176
rect 7340 1164 7346 1216
rect 7392 1213 7420 1312
rect 7558 1300 7564 1352
rect 7616 1300 7622 1352
rect 8481 1343 8539 1349
rect 8481 1309 8493 1343
rect 8527 1340 8539 1343
rect 8527 1312 8616 1340
rect 8527 1309 8539 1312
rect 8481 1303 8539 1309
rect 8588 1213 8616 1312
rect 8754 1300 8760 1352
rect 8812 1300 8818 1352
rect 9490 1300 9496 1352
rect 9548 1300 9554 1352
rect 9858 1300 9864 1352
rect 9916 1300 9922 1352
rect 10137 1343 10195 1349
rect 10137 1309 10149 1343
rect 10183 1309 10195 1343
rect 10137 1303 10195 1309
rect 10152 1272 10180 1303
rect 10686 1300 10692 1352
rect 10744 1300 10750 1352
rect 10965 1343 11023 1349
rect 10965 1309 10977 1343
rect 11011 1309 11023 1343
rect 10965 1303 11023 1309
rect 10980 1272 11008 1303
rect 11238 1300 11244 1352
rect 11296 1300 11302 1352
rect 11790 1340 11796 1352
rect 11348 1312 11796 1340
rect 9324 1244 10180 1272
rect 10520 1244 11008 1272
rect 9324 1213 9352 1244
rect 10520 1213 10548 1244
rect 7377 1207 7435 1213
rect 7377 1173 7389 1207
rect 7423 1173 7435 1207
rect 7377 1167 7435 1173
rect 8573 1207 8631 1213
rect 8573 1173 8585 1207
rect 8619 1173 8631 1207
rect 8573 1167 8631 1173
rect 9309 1207 9367 1213
rect 9309 1173 9321 1207
rect 9355 1173 9367 1207
rect 9309 1167 9367 1173
rect 10505 1207 10563 1213
rect 10505 1173 10517 1207
rect 10551 1173 10563 1207
rect 10505 1167 10563 1173
rect 10781 1207 10839 1213
rect 10781 1173 10793 1207
rect 10827 1204 10839 1207
rect 11348 1204 11376 1312
rect 11790 1300 11796 1312
rect 11848 1300 11854 1352
rect 11882 1300 11888 1352
rect 11940 1300 11946 1352
rect 12161 1343 12219 1349
rect 12161 1309 12173 1343
rect 12207 1309 12219 1343
rect 12434 1340 12440 1352
rect 12161 1303 12219 1309
rect 12268 1312 12440 1340
rect 12176 1272 12204 1303
rect 11716 1244 12204 1272
rect 11716 1213 11744 1244
rect 10827 1176 11376 1204
rect 11701 1207 11759 1213
rect 10827 1173 10839 1176
rect 10781 1167 10839 1173
rect 11701 1173 11713 1207
rect 11747 1173 11759 1207
rect 11701 1167 11759 1173
rect 11977 1207 12035 1213
rect 11977 1173 11989 1207
rect 12023 1204 12035 1207
rect 12268 1204 12296 1312
rect 12434 1300 12440 1312
rect 12492 1300 12498 1352
rect 12526 1300 12532 1352
rect 12584 1300 12590 1352
rect 12986 1300 12992 1352
rect 13044 1300 13050 1352
rect 13265 1343 13323 1349
rect 13265 1309 13277 1343
rect 13311 1309 13323 1343
rect 13265 1303 13323 1309
rect 13280 1272 13308 1303
rect 13722 1300 13728 1352
rect 13780 1300 13786 1352
rect 14090 1300 14096 1352
rect 14148 1300 14154 1352
rect 14274 1300 14280 1352
rect 14332 1300 14338 1352
rect 14366 1300 14372 1352
rect 14424 1300 14430 1352
rect 14458 1300 14464 1352
rect 14516 1300 14522 1352
rect 15470 1300 15476 1352
rect 15528 1300 15534 1352
rect 15749 1343 15807 1349
rect 15749 1309 15761 1343
rect 15795 1309 15807 1343
rect 15749 1303 15807 1309
rect 14108 1272 14136 1300
rect 12820 1244 13308 1272
rect 13556 1244 14136 1272
rect 12820 1213 12848 1244
rect 13556 1213 13584 1244
rect 12023 1176 12296 1204
rect 12805 1207 12863 1213
rect 12023 1173 12035 1176
rect 11977 1167 12035 1173
rect 12805 1173 12817 1207
rect 12851 1173 12863 1207
rect 12805 1167 12863 1173
rect 13541 1207 13599 1213
rect 13541 1173 13553 1207
rect 13587 1173 13599 1207
rect 13541 1167 13599 1173
rect 14093 1207 14151 1213
rect 14093 1173 14105 1207
rect 14139 1204 14151 1207
rect 14476 1204 14504 1300
rect 15764 1272 15792 1303
rect 16666 1300 16672 1352
rect 16724 1340 16730 1352
rect 16853 1343 16911 1349
rect 16853 1340 16865 1343
rect 16724 1312 16865 1340
rect 16724 1300 16730 1312
rect 16853 1309 16865 1312
rect 16899 1309 16911 1343
rect 16853 1303 16911 1309
rect 17862 1300 17868 1352
rect 17920 1300 17926 1352
rect 19058 1300 19064 1352
rect 19116 1300 19122 1352
rect 20254 1300 20260 1352
rect 20312 1300 20318 1352
rect 15304 1244 15792 1272
rect 14139 1176 14504 1204
rect 14139 1173 14151 1176
rect 14093 1167 14151 1173
rect 14550 1164 14556 1216
rect 14608 1164 14614 1216
rect 15304 1213 15332 1244
rect 16758 1232 16764 1284
rect 16816 1232 16822 1284
rect 17770 1232 17776 1284
rect 17828 1232 17834 1284
rect 21284 1272 21312 1439
rect 21450 1300 21456 1352
rect 21508 1300 21514 1352
rect 22005 1343 22063 1349
rect 22005 1309 22017 1343
rect 22051 1309 22063 1343
rect 22005 1303 22063 1309
rect 22020 1272 22048 1303
rect 22646 1300 22652 1352
rect 22704 1300 22710 1352
rect 23017 1343 23075 1349
rect 23017 1309 23029 1343
rect 23063 1309 23075 1343
rect 23017 1303 23075 1309
rect 23293 1343 23351 1349
rect 23293 1309 23305 1343
rect 23339 1309 23351 1343
rect 23293 1303 23351 1309
rect 23032 1272 23060 1303
rect 21284 1244 22048 1272
rect 22388 1244 23060 1272
rect 15289 1207 15347 1213
rect 15289 1173 15301 1207
rect 15335 1173 15347 1207
rect 15289 1167 15347 1173
rect 16669 1207 16727 1213
rect 16669 1173 16681 1207
rect 16715 1204 16727 1207
rect 16776 1204 16804 1232
rect 16715 1176 16804 1204
rect 17681 1207 17739 1213
rect 16715 1173 16727 1176
rect 16669 1167 16727 1173
rect 17681 1173 17693 1207
rect 17727 1204 17739 1207
rect 17788 1204 17816 1232
rect 17727 1176 17816 1204
rect 18877 1207 18935 1213
rect 17727 1173 17739 1176
rect 17681 1167 17739 1173
rect 18877 1173 18889 1207
rect 18923 1204 18935 1207
rect 19978 1204 19984 1216
rect 18923 1176 19984 1204
rect 18923 1173 18935 1176
rect 18877 1167 18935 1173
rect 19978 1164 19984 1176
rect 20036 1164 20042 1216
rect 20073 1207 20131 1213
rect 20073 1173 20085 1207
rect 20119 1204 20131 1207
rect 22388 1204 22416 1244
rect 20119 1176 22416 1204
rect 20119 1173 20131 1176
rect 20073 1167 20131 1173
rect 22462 1164 22468 1216
rect 22520 1164 22526 1216
rect 22554 1164 22560 1216
rect 22612 1204 22618 1216
rect 23308 1204 23336 1303
rect 23566 1300 23572 1352
rect 23624 1300 23630 1352
rect 23845 1343 23903 1349
rect 23845 1309 23857 1343
rect 23891 1340 23903 1343
rect 23891 1312 23980 1340
rect 23891 1309 23903 1312
rect 23845 1303 23903 1309
rect 23952 1213 23980 1312
rect 24118 1300 24124 1352
rect 24176 1300 24182 1352
rect 22612 1176 23336 1204
rect 23937 1207 23995 1213
rect 22612 1164 22618 1176
rect 23937 1173 23949 1207
rect 23983 1173 23995 1207
rect 23937 1167 23995 1173
rect 1104 1114 24723 1136
rect 1104 1062 6814 1114
rect 6866 1062 6878 1114
rect 6930 1062 6942 1114
rect 6994 1062 7006 1114
rect 7058 1062 7070 1114
rect 7122 1062 12679 1114
rect 12731 1062 12743 1114
rect 12795 1062 12807 1114
rect 12859 1062 12871 1114
rect 12923 1062 12935 1114
rect 12987 1062 18544 1114
rect 18596 1062 18608 1114
rect 18660 1062 18672 1114
rect 18724 1062 18736 1114
rect 18788 1062 18800 1114
rect 18852 1062 24409 1114
rect 24461 1062 24473 1114
rect 24525 1062 24537 1114
rect 24589 1062 24601 1114
rect 24653 1062 24665 1114
rect 24717 1062 24723 1114
rect 1104 1040 24723 1062
rect 1578 960 1584 1012
rect 1636 960 1642 1012
rect 4522 960 4528 1012
rect 4580 960 4586 1012
rect 5718 960 5724 1012
rect 5776 1000 5782 1012
rect 9858 1000 9864 1012
rect 5776 972 9864 1000
rect 5776 960 5782 972
rect 9858 960 9864 972
rect 9916 960 9922 1012
rect 13722 960 13728 1012
rect 13780 960 13786 1012
rect 14366 960 14372 1012
rect 14424 960 14430 1012
rect 14550 960 14556 1012
rect 14608 1000 14614 1012
rect 19886 1000 19892 1012
rect 14608 972 19892 1000
rect 14608 960 14614 972
rect 19886 960 19892 972
rect 19944 960 19950 1012
rect 19978 960 19984 1012
rect 20036 1000 20042 1012
rect 22554 1000 22560 1012
rect 20036 972 22560 1000
rect 20036 960 20042 972
rect 22554 960 22560 972
rect 22612 960 22618 1012
rect 1596 864 1624 960
rect 4540 932 4568 960
rect 4540 904 7236 932
rect 7208 864 7236 904
rect 7282 892 7288 944
rect 7340 932 7346 944
rect 13740 932 13768 960
rect 7340 904 13768 932
rect 7340 892 7346 904
rect 12526 864 12532 876
rect 1596 836 7052 864
rect 7208 836 12532 864
rect 2314 756 2320 808
rect 2372 796 2378 808
rect 2372 768 6960 796
rect 2372 756 2378 768
rect 6932 660 6960 768
rect 7024 728 7052 836
rect 12526 824 12532 836
rect 12584 824 12590 876
rect 14384 728 14412 960
rect 7024 700 14412 728
rect 23566 688 23572 740
rect 23624 728 23630 740
rect 24762 728 24768 740
rect 23624 700 24768 728
rect 23624 688 23630 700
rect 24762 688 24768 700
rect 24820 688 24826 740
rect 11238 660 11244 672
rect 6932 632 11244 660
rect 11238 620 11244 632
rect 11296 620 11302 672
rect 6914 552 6920 604
rect 6972 592 6978 604
rect 7558 592 7564 604
rect 6972 564 7564 592
rect 6972 552 6978 564
rect 7558 552 7564 564
rect 7616 552 7622 604
<< via1 >>
rect 2228 9936 2280 9988
rect 11796 9936 11848 9988
rect 11888 9936 11940 9988
rect 17868 9936 17920 9988
rect 1584 9800 1636 9852
rect 14280 9868 14332 9920
rect 6000 9800 6052 9852
rect 14648 9800 14700 9852
rect 2412 9664 2464 9716
rect 7656 9732 7708 9784
rect 14832 9664 14884 9716
rect 18144 9664 18196 9716
rect 9496 9596 9548 9648
rect 10140 9596 10192 9648
rect 11520 9596 11572 9648
rect 19616 9596 19668 9648
rect 18972 9528 19024 9580
rect 6552 9460 6604 9512
rect 7932 9460 7984 9512
rect 11888 9460 11940 9512
rect 11244 9392 11296 9444
rect 6368 9324 6420 9376
rect 8208 9324 8260 9376
rect 12072 9324 12124 9376
rect 9036 9256 9088 9308
rect 9588 9256 9640 9308
rect 15384 9256 15436 9308
rect 1952 9188 2004 9240
rect 2504 9188 2556 9240
rect 13452 9188 13504 9240
rect 7748 9120 7800 9172
rect 11152 9120 11204 9172
rect 11244 9120 11296 9172
rect 11796 9120 11848 9172
rect 14556 9120 14608 9172
rect 4160 9052 4212 9104
rect 5540 8984 5592 9036
rect 10876 8984 10928 9036
rect 19340 9052 19392 9104
rect 12348 8984 12400 9036
rect 10048 8916 10100 8968
rect 9404 8848 9456 8900
rect 9956 8848 10008 8900
rect 16212 8916 16264 8968
rect 10416 8848 10468 8900
rect 16948 8848 17000 8900
rect 18880 8848 18932 8900
rect 19800 8848 19852 8900
rect 112 8780 164 8832
rect 2964 8780 3016 8832
rect 4436 8780 4488 8832
rect 4896 8780 4948 8832
rect 8024 8780 8076 8832
rect 17316 8780 17368 8832
rect 18604 8780 18656 8832
rect 19524 8780 19576 8832
rect 6814 8678 6866 8730
rect 6878 8678 6930 8730
rect 6942 8678 6994 8730
rect 7006 8678 7058 8730
rect 7070 8678 7122 8730
rect 12679 8678 12731 8730
rect 12743 8678 12795 8730
rect 12807 8678 12859 8730
rect 12871 8678 12923 8730
rect 12935 8678 12987 8730
rect 18544 8678 18596 8730
rect 18608 8678 18660 8730
rect 18672 8678 18724 8730
rect 18736 8678 18788 8730
rect 18800 8678 18852 8730
rect 24409 8678 24461 8730
rect 24473 8678 24525 8730
rect 24537 8678 24589 8730
rect 24601 8678 24653 8730
rect 24665 8678 24717 8730
rect 572 8576 624 8628
rect 2872 8576 2924 8628
rect 2964 8576 3016 8628
rect 4160 8576 4212 8628
rect 4252 8619 4304 8628
rect 4252 8585 4261 8619
rect 4261 8585 4295 8619
rect 4295 8585 4304 8619
rect 4252 8576 4304 8585
rect 5080 8576 5132 8628
rect 5356 8576 5408 8628
rect 5908 8576 5960 8628
rect 6460 8576 6512 8628
rect 7196 8576 7248 8628
rect 7564 8576 7616 8628
rect 8116 8576 8168 8628
rect 8392 8576 8444 8628
rect 8944 8576 8996 8628
rect 9220 8576 9272 8628
rect 9680 8619 9732 8628
rect 9680 8585 9689 8619
rect 9689 8585 9723 8619
rect 9723 8585 9732 8619
rect 9680 8576 9732 8585
rect 9956 8576 10008 8628
rect 1952 8483 2004 8492
rect 1952 8449 1961 8483
rect 1961 8449 1995 8483
rect 1995 8449 2004 8483
rect 1952 8440 2004 8449
rect 2504 8483 2556 8492
rect 2504 8449 2513 8483
rect 2513 8449 2547 8483
rect 2547 8449 2556 8483
rect 2504 8440 2556 8449
rect 4436 8483 4488 8492
rect 4436 8449 4445 8483
rect 4445 8449 4479 8483
rect 4479 8449 4488 8483
rect 4436 8440 4488 8449
rect 4896 8483 4948 8492
rect 4896 8449 4905 8483
rect 4905 8449 4939 8483
rect 4939 8449 4948 8483
rect 4896 8440 4948 8449
rect 5816 8440 5868 8492
rect 5908 8483 5960 8492
rect 5908 8449 5917 8483
rect 5917 8449 5951 8483
rect 5951 8449 5960 8483
rect 5908 8440 5960 8449
rect 6552 8551 6604 8560
rect 6552 8517 6561 8551
rect 6561 8517 6595 8551
rect 6595 8517 6604 8551
rect 6552 8508 6604 8517
rect 7196 8483 7248 8492
rect 7196 8449 7205 8483
rect 7205 8449 7239 8483
rect 7239 8449 7248 8483
rect 7196 8440 7248 8449
rect 8024 8551 8076 8560
rect 8024 8517 8033 8551
rect 8033 8517 8067 8551
rect 8067 8517 8076 8551
rect 8024 8508 8076 8517
rect 9588 8551 9640 8560
rect 9588 8517 9597 8551
rect 9597 8517 9631 8551
rect 9631 8517 9640 8551
rect 9588 8508 9640 8517
rect 10232 8619 10284 8628
rect 10232 8585 10241 8619
rect 10241 8585 10275 8619
rect 10275 8585 10284 8619
rect 10232 8576 10284 8585
rect 7380 8372 7432 8424
rect 8300 8372 8352 8424
rect 3424 8304 3476 8356
rect 6644 8304 6696 8356
rect 10232 8372 10284 8424
rect 10416 8304 10468 8356
rect 11152 8508 11204 8560
rect 12900 8576 12952 8628
rect 11060 8483 11112 8492
rect 11060 8449 11069 8483
rect 11069 8449 11103 8483
rect 11103 8449 11112 8483
rect 11060 8440 11112 8449
rect 11520 8440 11572 8492
rect 11704 8483 11756 8492
rect 11704 8449 11713 8483
rect 11713 8449 11747 8483
rect 11747 8449 11756 8483
rect 11704 8440 11756 8449
rect 10876 8347 10928 8356
rect 10876 8313 10885 8347
rect 10885 8313 10919 8347
rect 10919 8313 10928 8347
rect 10876 8304 10928 8313
rect 14556 8619 14608 8628
rect 14556 8585 14565 8619
rect 14565 8585 14599 8619
rect 14599 8585 14608 8619
rect 14556 8576 14608 8585
rect 14832 8619 14884 8628
rect 14832 8585 14841 8619
rect 14841 8585 14875 8619
rect 14875 8585 14884 8619
rect 14832 8576 14884 8585
rect 15016 8576 15068 8628
rect 16948 8619 17000 8628
rect 16948 8585 16957 8619
rect 16957 8585 16991 8619
rect 16991 8585 17000 8619
rect 16948 8576 17000 8585
rect 14188 8508 14240 8560
rect 12440 8372 12492 8424
rect 13360 8483 13412 8492
rect 13360 8449 13369 8483
rect 13369 8449 13403 8483
rect 13403 8449 13412 8483
rect 13360 8440 13412 8449
rect 13176 8372 13228 8424
rect 13636 8440 13688 8492
rect 14004 8440 14056 8492
rect 14648 8483 14700 8492
rect 14648 8449 14657 8483
rect 14657 8449 14691 8483
rect 14691 8449 14700 8483
rect 14648 8440 14700 8449
rect 14740 8440 14792 8492
rect 15384 8508 15436 8560
rect 11796 8279 11848 8288
rect 11796 8245 11805 8279
rect 11805 8245 11839 8279
rect 11839 8245 11848 8279
rect 11796 8236 11848 8245
rect 12072 8279 12124 8288
rect 12072 8245 12081 8279
rect 12081 8245 12115 8279
rect 12115 8245 12124 8279
rect 12072 8236 12124 8245
rect 12348 8347 12400 8356
rect 12348 8313 12357 8347
rect 12357 8313 12391 8347
rect 12391 8313 12400 8347
rect 12348 8304 12400 8313
rect 13452 8304 13504 8356
rect 13636 8347 13688 8356
rect 13636 8313 13645 8347
rect 13645 8313 13679 8347
rect 13679 8313 13688 8347
rect 13636 8304 13688 8313
rect 14280 8304 14332 8356
rect 15200 8483 15252 8492
rect 15200 8449 15209 8483
rect 15209 8449 15243 8483
rect 15243 8449 15252 8483
rect 15200 8440 15252 8449
rect 15292 8440 15344 8492
rect 15384 8372 15436 8424
rect 16120 8440 16172 8492
rect 16488 8483 16540 8492
rect 16488 8449 16497 8483
rect 16497 8449 16531 8483
rect 16531 8449 16540 8483
rect 16488 8440 16540 8449
rect 16856 8483 16908 8492
rect 16856 8449 16865 8483
rect 16865 8449 16899 8483
rect 16899 8449 16908 8483
rect 16856 8440 16908 8449
rect 17316 8576 17368 8628
rect 17868 8576 17920 8628
rect 15844 8236 15896 8288
rect 16580 8372 16632 8424
rect 17868 8440 17920 8492
rect 18420 8576 18472 8628
rect 17500 8372 17552 8424
rect 18604 8483 18656 8492
rect 18604 8449 18613 8483
rect 18613 8449 18647 8483
rect 18647 8449 18656 8483
rect 18604 8440 18656 8449
rect 18972 8372 19024 8424
rect 16212 8304 16264 8356
rect 17132 8304 17184 8356
rect 17868 8304 17920 8356
rect 18144 8304 18196 8356
rect 19340 8440 19392 8492
rect 19616 8576 19668 8628
rect 19984 8576 20036 8628
rect 20352 8576 20404 8628
rect 21088 8576 21140 8628
rect 21364 8508 21416 8560
rect 23204 8576 23256 8628
rect 19524 8440 19576 8492
rect 19800 8483 19852 8492
rect 19800 8449 19809 8483
rect 19809 8449 19843 8483
rect 19843 8449 19852 8483
rect 19800 8440 19852 8449
rect 20076 8483 20128 8492
rect 20076 8449 20085 8483
rect 20085 8449 20119 8483
rect 20119 8449 20128 8483
rect 20076 8440 20128 8449
rect 20720 8440 20772 8492
rect 21180 8440 21232 8492
rect 22468 8483 22520 8492
rect 22468 8449 22477 8483
rect 22477 8449 22511 8483
rect 22511 8449 22520 8483
rect 22468 8440 22520 8449
rect 23020 8483 23072 8492
rect 23020 8449 23029 8483
rect 23029 8449 23063 8483
rect 23063 8449 23072 8483
rect 23020 8440 23072 8449
rect 23572 8483 23624 8492
rect 23572 8449 23581 8483
rect 23581 8449 23615 8483
rect 23615 8449 23624 8483
rect 23572 8440 23624 8449
rect 20536 8304 20588 8356
rect 21640 8304 21692 8356
rect 19524 8279 19576 8288
rect 19524 8245 19533 8279
rect 19533 8245 19567 8279
rect 19567 8245 19576 8279
rect 19524 8236 19576 8245
rect 3882 8134 3934 8186
rect 3946 8134 3998 8186
rect 4010 8134 4062 8186
rect 4074 8134 4126 8186
rect 4138 8134 4190 8186
rect 9747 8134 9799 8186
rect 9811 8134 9863 8186
rect 9875 8134 9927 8186
rect 9939 8134 9991 8186
rect 10003 8134 10055 8186
rect 15612 8134 15664 8186
rect 15676 8134 15728 8186
rect 15740 8134 15792 8186
rect 15804 8134 15856 8186
rect 15868 8134 15920 8186
rect 21477 8134 21529 8186
rect 21541 8134 21593 8186
rect 21605 8134 21657 8186
rect 21669 8134 21721 8186
rect 21733 8134 21785 8186
rect 2044 8032 2096 8084
rect 2320 8075 2372 8084
rect 2320 8041 2329 8075
rect 2329 8041 2363 8075
rect 2363 8041 2372 8075
rect 2320 8032 2372 8041
rect 3240 8075 3292 8084
rect 3240 8041 3249 8075
rect 3249 8041 3283 8075
rect 3283 8041 3292 8075
rect 3240 8032 3292 8041
rect 4620 8075 4672 8084
rect 4620 8041 4629 8075
rect 4629 8041 4663 8075
rect 4663 8041 4672 8075
rect 4620 8032 4672 8041
rect 4804 8032 4856 8084
rect 5724 8075 5776 8084
rect 5724 8041 5733 8075
rect 5733 8041 5767 8075
rect 5767 8041 5776 8075
rect 5724 8032 5776 8041
rect 6276 8075 6328 8084
rect 6276 8041 6285 8075
rect 6285 8041 6319 8075
rect 6319 8041 6328 8075
rect 6276 8032 6328 8041
rect 2780 8007 2832 8016
rect 2780 7973 2789 8007
rect 2789 7973 2823 8007
rect 2823 7973 2832 8007
rect 2780 7964 2832 7973
rect 4160 8007 4212 8016
rect 4160 7973 4169 8007
rect 4169 7973 4203 8007
rect 4203 7973 4212 8007
rect 4160 7964 4212 7973
rect 6920 8007 6972 8016
rect 6920 7973 6929 8007
rect 6929 7973 6963 8007
rect 6963 7973 6972 8007
rect 6920 7964 6972 7973
rect 7288 8032 7340 8084
rect 7932 8075 7984 8084
rect 7932 8041 7941 8075
rect 7941 8041 7975 8075
rect 7975 8041 7984 8075
rect 7932 8032 7984 8041
rect 8668 8075 8720 8084
rect 8668 8041 8677 8075
rect 8677 8041 8711 8075
rect 8711 8041 8720 8075
rect 8668 8032 8720 8041
rect 7748 7964 7800 8016
rect 2412 7828 2464 7880
rect 2596 7871 2648 7880
rect 2596 7837 2605 7871
rect 2605 7837 2639 7871
rect 2639 7837 2648 7871
rect 2596 7828 2648 7837
rect 5448 7896 5500 7948
rect 9404 8032 9456 8084
rect 9772 8032 9824 8084
rect 11520 8032 11572 8084
rect 12440 8032 12492 8084
rect 12900 8075 12952 8084
rect 12900 8041 12909 8075
rect 12909 8041 12943 8075
rect 12943 8041 12952 8075
rect 12900 8032 12952 8041
rect 13176 8075 13228 8084
rect 13176 8041 13185 8075
rect 13185 8041 13219 8075
rect 13219 8041 13228 8075
rect 13176 8032 13228 8041
rect 14648 8032 14700 8084
rect 15200 8032 15252 8084
rect 15292 8032 15344 8084
rect 15384 8075 15436 8084
rect 15384 8041 15393 8075
rect 15393 8041 15427 8075
rect 15427 8041 15436 8075
rect 15384 8032 15436 8041
rect 16120 8032 16172 8084
rect 16856 8032 16908 8084
rect 18604 8032 18656 8084
rect 9036 8007 9088 8016
rect 9036 7973 9045 8007
rect 9045 7973 9079 8007
rect 9079 7973 9088 8007
rect 9036 7964 9088 7973
rect 11060 7964 11112 8016
rect 16488 7964 16540 8016
rect 6644 7828 6696 7880
rect 2228 7760 2280 7812
rect 5540 7760 5592 7812
rect 5632 7803 5684 7812
rect 5632 7769 5641 7803
rect 5641 7769 5675 7803
rect 5675 7769 5684 7803
rect 5632 7760 5684 7769
rect 6552 7760 6604 7812
rect 6736 7803 6788 7812
rect 6736 7769 6745 7803
rect 6745 7769 6779 7803
rect 6779 7769 6788 7803
rect 6736 7760 6788 7769
rect 7380 7828 7432 7880
rect 7656 7760 7708 7812
rect 7840 7803 7892 7812
rect 7840 7769 7849 7803
rect 7849 7769 7883 7803
rect 7883 7769 7892 7803
rect 7840 7760 7892 7769
rect 8484 7871 8536 7880
rect 8484 7837 8493 7871
rect 8493 7837 8527 7871
rect 8527 7837 8536 7871
rect 8484 7828 8536 7837
rect 8852 7692 8904 7744
rect 9588 7828 9640 7880
rect 9772 7871 9824 7880
rect 9772 7837 9781 7871
rect 9781 7837 9815 7871
rect 9815 7837 9824 7871
rect 9772 7828 9824 7837
rect 16212 7896 16264 7948
rect 9036 7760 9088 7812
rect 10600 7871 10652 7880
rect 10600 7837 10609 7871
rect 10609 7837 10643 7871
rect 10643 7837 10652 7871
rect 10600 7828 10652 7837
rect 10876 7871 10928 7880
rect 10876 7837 10885 7871
rect 10885 7837 10919 7871
rect 10919 7837 10928 7871
rect 10876 7828 10928 7837
rect 11152 7871 11204 7880
rect 11152 7837 11161 7871
rect 11161 7837 11195 7871
rect 11195 7837 11204 7871
rect 11152 7828 11204 7837
rect 11428 7871 11480 7880
rect 11428 7837 11437 7871
rect 11437 7837 11471 7871
rect 11471 7837 11480 7871
rect 11428 7828 11480 7837
rect 11704 7871 11756 7880
rect 11704 7837 11713 7871
rect 11713 7837 11747 7871
rect 11747 7837 11756 7871
rect 11704 7828 11756 7837
rect 11980 7828 12032 7880
rect 12532 7871 12584 7880
rect 12532 7837 12541 7871
rect 12541 7837 12575 7871
rect 12575 7837 12584 7871
rect 12532 7828 12584 7837
rect 12808 7871 12860 7880
rect 12808 7837 12817 7871
rect 12817 7837 12851 7871
rect 12851 7837 12860 7871
rect 12808 7828 12860 7837
rect 13084 7871 13136 7880
rect 13084 7837 13093 7871
rect 13093 7837 13127 7871
rect 13127 7837 13136 7871
rect 13084 7828 13136 7837
rect 13360 7871 13412 7880
rect 13360 7837 13369 7871
rect 13369 7837 13403 7871
rect 13403 7837 13412 7871
rect 13360 7828 13412 7837
rect 14464 7828 14516 7880
rect 15016 7871 15068 7880
rect 15016 7837 15025 7871
rect 15025 7837 15059 7871
rect 15059 7837 15068 7871
rect 15016 7828 15068 7837
rect 15292 7871 15344 7880
rect 15292 7837 15301 7871
rect 15301 7837 15335 7871
rect 15335 7837 15344 7871
rect 15292 7828 15344 7837
rect 15568 7871 15620 7880
rect 15568 7837 15577 7871
rect 15577 7837 15611 7871
rect 15611 7837 15620 7871
rect 15568 7828 15620 7837
rect 15844 7871 15896 7880
rect 15844 7837 15853 7871
rect 15853 7837 15887 7871
rect 15887 7837 15896 7871
rect 15844 7828 15896 7837
rect 16120 7871 16172 7880
rect 16120 7837 16129 7871
rect 16129 7837 16163 7871
rect 16163 7837 16172 7871
rect 16120 7828 16172 7837
rect 16396 7871 16448 7880
rect 16396 7837 16405 7871
rect 16405 7837 16439 7871
rect 16439 7837 16448 7871
rect 16396 7828 16448 7837
rect 16672 7828 16724 7880
rect 17224 7828 17276 7880
rect 17776 7828 17828 7880
rect 18328 7871 18380 7880
rect 18328 7837 18337 7871
rect 18337 7837 18371 7871
rect 18371 7837 18380 7871
rect 18328 7828 18380 7837
rect 19524 8032 19576 8084
rect 20812 8032 20864 8084
rect 21916 8032 21968 8084
rect 22284 8032 22336 8084
rect 22836 8032 22888 8084
rect 23204 7964 23256 8016
rect 19340 7828 19392 7880
rect 19524 7871 19576 7880
rect 19524 7837 19533 7871
rect 19533 7837 19567 7871
rect 19567 7837 19576 7871
rect 19524 7828 19576 7837
rect 19800 7871 19852 7880
rect 19800 7837 19809 7871
rect 19809 7837 19843 7871
rect 19843 7837 19852 7871
rect 19800 7828 19852 7837
rect 25504 7828 25556 7880
rect 10140 7735 10192 7744
rect 10140 7701 10149 7735
rect 10149 7701 10183 7735
rect 10183 7701 10192 7735
rect 10140 7692 10192 7701
rect 11612 7692 11664 7744
rect 16764 7735 16816 7744
rect 16764 7701 16773 7735
rect 16773 7701 16807 7735
rect 16807 7701 16816 7735
rect 16764 7692 16816 7701
rect 17316 7735 17368 7744
rect 17316 7701 17325 7735
rect 17325 7701 17359 7735
rect 17359 7701 17368 7735
rect 17316 7692 17368 7701
rect 18604 7735 18656 7744
rect 18604 7701 18613 7735
rect 18613 7701 18647 7735
rect 18647 7701 18656 7735
rect 18604 7692 18656 7701
rect 19064 7735 19116 7744
rect 19064 7701 19073 7735
rect 19073 7701 19107 7735
rect 19107 7701 19116 7735
rect 19064 7692 19116 7701
rect 19708 7735 19760 7744
rect 19708 7701 19717 7735
rect 19717 7701 19751 7735
rect 19751 7701 19760 7735
rect 19708 7692 19760 7701
rect 19984 7735 20036 7744
rect 19984 7701 19993 7735
rect 19993 7701 20027 7735
rect 20027 7701 20036 7735
rect 19984 7692 20036 7701
rect 22100 7803 22152 7812
rect 22100 7769 22109 7803
rect 22109 7769 22143 7803
rect 22143 7769 22152 7803
rect 22100 7760 22152 7769
rect 22652 7803 22704 7812
rect 22652 7769 22661 7803
rect 22661 7769 22695 7803
rect 22695 7769 22704 7803
rect 22652 7760 22704 7769
rect 22744 7760 22796 7812
rect 23756 7803 23808 7812
rect 23756 7769 23765 7803
rect 23765 7769 23799 7803
rect 23799 7769 23808 7803
rect 23756 7760 23808 7769
rect 22836 7692 22888 7744
rect 6814 7590 6866 7642
rect 6878 7590 6930 7642
rect 6942 7590 6994 7642
rect 7006 7590 7058 7642
rect 7070 7590 7122 7642
rect 12679 7590 12731 7642
rect 12743 7590 12795 7642
rect 12807 7590 12859 7642
rect 12871 7590 12923 7642
rect 12935 7590 12987 7642
rect 18544 7590 18596 7642
rect 18608 7590 18660 7642
rect 18672 7590 18724 7642
rect 18736 7590 18788 7642
rect 18800 7590 18852 7642
rect 24409 7590 24461 7642
rect 24473 7590 24525 7642
rect 24537 7590 24589 7642
rect 24601 7590 24653 7642
rect 24665 7590 24717 7642
rect 1676 7531 1728 7540
rect 1676 7497 1685 7531
rect 1685 7497 1719 7531
rect 1719 7497 1728 7531
rect 1676 7488 1728 7497
rect 1492 7420 1544 7472
rect 3700 7488 3752 7540
rect 5632 7488 5684 7540
rect 5908 7488 5960 7540
rect 7196 7488 7248 7540
rect 8300 7531 8352 7540
rect 8300 7497 8309 7531
rect 8309 7497 8343 7531
rect 8343 7497 8352 7531
rect 8300 7488 8352 7497
rect 8484 7488 8536 7540
rect 1584 7395 1636 7404
rect 1584 7361 1593 7395
rect 1593 7361 1627 7395
rect 1627 7361 1636 7395
rect 1584 7352 1636 7361
rect 6000 7420 6052 7472
rect 5632 7395 5684 7404
rect 5632 7361 5641 7395
rect 5641 7361 5675 7395
rect 5675 7361 5684 7395
rect 5632 7352 5684 7361
rect 6184 7395 6236 7404
rect 6184 7361 6193 7395
rect 6193 7361 6227 7395
rect 6227 7361 6236 7395
rect 6184 7352 6236 7361
rect 6368 7352 6420 7404
rect 7380 7395 7432 7404
rect 7380 7361 7389 7395
rect 7389 7361 7423 7395
rect 7423 7361 7432 7395
rect 7380 7352 7432 7361
rect 8392 7352 8444 7404
rect 8208 7284 8260 7336
rect 8668 7352 8720 7404
rect 16764 7488 16816 7540
rect 17316 7488 17368 7540
rect 24124 7488 24176 7540
rect 24768 7488 24820 7540
rect 8852 7420 8904 7472
rect 11796 7420 11848 7472
rect 10324 7395 10376 7404
rect 10324 7361 10333 7395
rect 10333 7361 10367 7395
rect 10367 7361 10376 7395
rect 10324 7352 10376 7361
rect 11612 7284 11664 7336
rect 9312 7216 9364 7268
rect 9496 7216 9548 7268
rect 17408 7395 17460 7404
rect 17408 7361 17417 7395
rect 17417 7361 17451 7395
rect 17451 7361 17460 7395
rect 17408 7352 17460 7361
rect 22468 7395 22520 7404
rect 22468 7361 22477 7395
rect 22477 7361 22511 7395
rect 22511 7361 22520 7395
rect 22468 7352 22520 7361
rect 23020 7395 23072 7404
rect 23020 7361 23029 7395
rect 23029 7361 23063 7395
rect 23063 7361 23072 7395
rect 23020 7352 23072 7361
rect 23572 7395 23624 7404
rect 23572 7361 23581 7395
rect 23581 7361 23615 7395
rect 23615 7361 23624 7395
rect 23572 7352 23624 7361
rect 24952 7284 25004 7336
rect 2780 7191 2832 7200
rect 2780 7157 2789 7191
rect 2789 7157 2823 7191
rect 2823 7157 2832 7191
rect 2780 7148 2832 7157
rect 5816 7148 5868 7200
rect 7380 7148 7432 7200
rect 9036 7148 9088 7200
rect 9634 7148 9686 7200
rect 22100 7148 22152 7200
rect 3882 7046 3934 7098
rect 3946 7046 3998 7098
rect 4010 7046 4062 7098
rect 4074 7046 4126 7098
rect 4138 7046 4190 7098
rect 9747 7046 9799 7098
rect 9811 7046 9863 7098
rect 9875 7046 9927 7098
rect 9939 7046 9991 7098
rect 10003 7046 10055 7098
rect 15612 7046 15664 7098
rect 15676 7046 15728 7098
rect 15740 7046 15792 7098
rect 15804 7046 15856 7098
rect 15868 7046 15920 7098
rect 21477 7046 21529 7098
rect 21541 7046 21593 7098
rect 21605 7046 21657 7098
rect 21669 7046 21721 7098
rect 21733 7046 21785 7098
rect 6552 6944 6604 6996
rect 17408 6944 17460 6996
rect 19064 6944 19116 6996
rect 664 6808 716 6860
rect 2780 6808 2832 6860
rect 24308 6808 24360 6860
rect 1216 6740 1268 6792
rect 16856 6783 16908 6792
rect 16856 6749 16865 6783
rect 16865 6749 16899 6783
rect 16899 6749 16908 6783
rect 16856 6740 16908 6749
rect 2688 6672 2740 6724
rect 23112 6715 23164 6724
rect 23112 6681 23121 6715
rect 23121 6681 23155 6715
rect 23155 6681 23164 6715
rect 23112 6672 23164 6681
rect 23388 6672 23440 6724
rect 23940 6672 23992 6724
rect 6814 6502 6866 6554
rect 6878 6502 6930 6554
rect 6942 6502 6994 6554
rect 7006 6502 7058 6554
rect 7070 6502 7122 6554
rect 12679 6502 12731 6554
rect 12743 6502 12795 6554
rect 12807 6502 12859 6554
rect 12871 6502 12923 6554
rect 12935 6502 12987 6554
rect 18544 6502 18596 6554
rect 18608 6502 18660 6554
rect 18672 6502 18724 6554
rect 18736 6502 18788 6554
rect 18800 6502 18852 6554
rect 24409 6502 24461 6554
rect 24473 6502 24525 6554
rect 24537 6502 24589 6554
rect 24601 6502 24653 6554
rect 24665 6502 24717 6554
rect 940 6400 992 6452
rect 23296 6443 23348 6452
rect 23296 6409 23305 6443
rect 23305 6409 23339 6443
rect 23339 6409 23348 6443
rect 23296 6400 23348 6409
rect 23848 6443 23900 6452
rect 23848 6409 23857 6443
rect 23857 6409 23891 6443
rect 23891 6409 23900 6443
rect 23848 6400 23900 6409
rect 5448 6332 5500 6384
rect 22100 6332 22152 6384
rect 23204 6307 23256 6316
rect 23204 6273 23213 6307
rect 23213 6273 23247 6307
rect 23247 6273 23256 6307
rect 23204 6264 23256 6273
rect 3882 5958 3934 6010
rect 3946 5958 3998 6010
rect 4010 5958 4062 6010
rect 4074 5958 4126 6010
rect 4138 5958 4190 6010
rect 9747 5958 9799 6010
rect 9811 5958 9863 6010
rect 9875 5958 9927 6010
rect 9939 5958 9991 6010
rect 10003 5958 10055 6010
rect 15612 5958 15664 6010
rect 15676 5958 15728 6010
rect 15740 5958 15792 6010
rect 15804 5958 15856 6010
rect 15868 5958 15920 6010
rect 21477 5958 21529 6010
rect 21541 5958 21593 6010
rect 21605 5958 21657 6010
rect 21669 5958 21721 6010
rect 21733 5958 21785 6010
rect 25228 5856 25280 5908
rect 23848 5627 23900 5636
rect 23848 5593 23857 5627
rect 23857 5593 23891 5627
rect 23891 5593 23900 5627
rect 23848 5584 23900 5593
rect 6814 5414 6866 5466
rect 6878 5414 6930 5466
rect 6942 5414 6994 5466
rect 7006 5414 7058 5466
rect 7070 5414 7122 5466
rect 12679 5414 12731 5466
rect 12743 5414 12795 5466
rect 12807 5414 12859 5466
rect 12871 5414 12923 5466
rect 12935 5414 12987 5466
rect 18544 5414 18596 5466
rect 18608 5414 18660 5466
rect 18672 5414 18724 5466
rect 18736 5414 18788 5466
rect 18800 5414 18852 5466
rect 24409 5414 24461 5466
rect 24473 5414 24525 5466
rect 24537 5414 24589 5466
rect 24601 5414 24653 5466
rect 24665 5414 24717 5466
rect 3882 4870 3934 4922
rect 3946 4870 3998 4922
rect 4010 4870 4062 4922
rect 4074 4870 4126 4922
rect 4138 4870 4190 4922
rect 9747 4870 9799 4922
rect 9811 4870 9863 4922
rect 9875 4870 9927 4922
rect 9939 4870 9991 4922
rect 10003 4870 10055 4922
rect 15612 4870 15664 4922
rect 15676 4870 15728 4922
rect 15740 4870 15792 4922
rect 15804 4870 15856 4922
rect 15868 4870 15920 4922
rect 21477 4870 21529 4922
rect 21541 4870 21593 4922
rect 21605 4870 21657 4922
rect 21669 4870 21721 4922
rect 21733 4870 21785 4922
rect 14832 4607 14884 4616
rect 14832 4573 14841 4607
rect 14841 4573 14875 4607
rect 14875 4573 14884 4607
rect 14832 4564 14884 4573
rect 23480 4428 23532 4480
rect 6814 4326 6866 4378
rect 6878 4326 6930 4378
rect 6942 4326 6994 4378
rect 7006 4326 7058 4378
rect 7070 4326 7122 4378
rect 12679 4326 12731 4378
rect 12743 4326 12795 4378
rect 12807 4326 12859 4378
rect 12871 4326 12923 4378
rect 12935 4326 12987 4378
rect 18544 4326 18596 4378
rect 18608 4326 18660 4378
rect 18672 4326 18724 4378
rect 18736 4326 18788 4378
rect 18800 4326 18852 4378
rect 24409 4326 24461 4378
rect 24473 4326 24525 4378
rect 24537 4326 24589 4378
rect 24601 4326 24653 4378
rect 24665 4326 24717 4378
rect 14832 4224 14884 4276
rect 14464 4131 14516 4140
rect 14464 4097 14473 4131
rect 14473 4097 14507 4131
rect 14507 4097 14516 4131
rect 14464 4088 14516 4097
rect 3882 3782 3934 3834
rect 3946 3782 3998 3834
rect 4010 3782 4062 3834
rect 4074 3782 4126 3834
rect 4138 3782 4190 3834
rect 9747 3782 9799 3834
rect 9811 3782 9863 3834
rect 9875 3782 9927 3834
rect 9939 3782 9991 3834
rect 10003 3782 10055 3834
rect 15612 3782 15664 3834
rect 15676 3782 15728 3834
rect 15740 3782 15792 3834
rect 15804 3782 15856 3834
rect 15868 3782 15920 3834
rect 21477 3782 21529 3834
rect 21541 3782 21593 3834
rect 21605 3782 21657 3834
rect 21669 3782 21721 3834
rect 21733 3782 21785 3834
rect 23112 3680 23164 3732
rect 17776 3476 17828 3528
rect 6814 3238 6866 3290
rect 6878 3238 6930 3290
rect 6942 3238 6994 3290
rect 7006 3238 7058 3290
rect 7070 3238 7122 3290
rect 12679 3238 12731 3290
rect 12743 3238 12795 3290
rect 12807 3238 12859 3290
rect 12871 3238 12923 3290
rect 12935 3238 12987 3290
rect 18544 3238 18596 3290
rect 18608 3238 18660 3290
rect 18672 3238 18724 3290
rect 18736 3238 18788 3290
rect 18800 3238 18852 3290
rect 24409 3238 24461 3290
rect 24473 3238 24525 3290
rect 24537 3238 24589 3290
rect 24601 3238 24653 3290
rect 24665 3238 24717 3290
rect 22468 3136 22520 3188
rect 22836 3068 22888 3120
rect 22468 3000 22520 3052
rect 24032 3043 24084 3052
rect 24032 3009 24041 3043
rect 24041 3009 24075 3043
rect 24075 3009 24084 3043
rect 24032 3000 24084 3009
rect 3882 2694 3934 2746
rect 3946 2694 3998 2746
rect 4010 2694 4062 2746
rect 4074 2694 4126 2746
rect 4138 2694 4190 2746
rect 9747 2694 9799 2746
rect 9811 2694 9863 2746
rect 9875 2694 9927 2746
rect 9939 2694 9991 2746
rect 10003 2694 10055 2746
rect 15612 2694 15664 2746
rect 15676 2694 15728 2746
rect 15740 2694 15792 2746
rect 15804 2694 15856 2746
rect 15868 2694 15920 2746
rect 21477 2694 21529 2746
rect 21541 2694 21593 2746
rect 21605 2694 21657 2746
rect 21669 2694 21721 2746
rect 21733 2694 21785 2746
rect 24032 2592 24084 2644
rect 23296 2388 23348 2440
rect 13820 2320 13872 2372
rect 23756 2320 23808 2372
rect 10416 2252 10468 2304
rect 21180 2252 21232 2304
rect 6814 2150 6866 2202
rect 6878 2150 6930 2202
rect 6942 2150 6994 2202
rect 7006 2150 7058 2202
rect 7070 2150 7122 2202
rect 12679 2150 12731 2202
rect 12743 2150 12795 2202
rect 12807 2150 12859 2202
rect 12871 2150 12923 2202
rect 12935 2150 12987 2202
rect 18544 2150 18596 2202
rect 18608 2150 18660 2202
rect 18672 2150 18724 2202
rect 18736 2150 18788 2202
rect 18800 2150 18852 2202
rect 24409 2150 24461 2202
rect 24473 2150 24525 2202
rect 24537 2150 24589 2202
rect 24601 2150 24653 2202
rect 24665 2150 24717 2202
rect 9036 2091 9088 2100
rect 9036 2057 9045 2091
rect 9045 2057 9079 2091
rect 9079 2057 9088 2091
rect 9036 2048 9088 2057
rect 10416 2091 10468 2100
rect 10416 2057 10425 2091
rect 10425 2057 10459 2091
rect 10459 2057 10468 2091
rect 10416 2048 10468 2057
rect 10692 2091 10744 2100
rect 10692 2057 10701 2091
rect 10701 2057 10735 2091
rect 10735 2057 10744 2091
rect 10692 2048 10744 2057
rect 11520 2048 11572 2100
rect 7656 1955 7708 1964
rect 7656 1921 7665 1955
rect 7665 1921 7699 1955
rect 7699 1921 7708 1955
rect 7656 1912 7708 1921
rect 8852 1955 8904 1964
rect 8852 1921 8861 1955
rect 8861 1921 8895 1955
rect 8895 1921 8904 1955
rect 8852 1912 8904 1921
rect 10232 1955 10284 1964
rect 10232 1921 10241 1955
rect 10241 1921 10275 1955
rect 10275 1921 10284 1955
rect 10232 1912 10284 1921
rect 10508 1955 10560 1964
rect 10508 1921 10517 1955
rect 10517 1921 10551 1955
rect 10551 1921 10560 1955
rect 10508 1912 10560 1921
rect 11520 1955 11572 1964
rect 11520 1921 11529 1955
rect 11529 1921 11563 1955
rect 11563 1921 11572 1955
rect 11520 1912 11572 1921
rect 11796 1955 11848 1964
rect 11796 1921 11805 1955
rect 11805 1921 11839 1955
rect 11839 1921 11848 1955
rect 11796 1912 11848 1921
rect 12440 1955 12492 1964
rect 12440 1921 12449 1955
rect 12449 1921 12483 1955
rect 12483 1921 12492 1955
rect 12440 1912 12492 1921
rect 13820 2091 13872 2100
rect 13820 2057 13829 2091
rect 13829 2057 13863 2091
rect 13863 2057 13872 2091
rect 13820 2048 13872 2057
rect 20720 2048 20772 2100
rect 23020 2048 23072 2100
rect 23204 2048 23256 2100
rect 23388 2091 23440 2100
rect 23388 2057 23397 2091
rect 23397 2057 23431 2091
rect 23431 2057 23440 2091
rect 23388 2048 23440 2057
rect 23572 2048 23624 2100
rect 23848 2048 23900 2100
rect 16212 1980 16264 2032
rect 12808 1955 12860 1964
rect 12808 1921 12817 1955
rect 12817 1921 12851 1955
rect 12851 1921 12860 1955
rect 12808 1912 12860 1921
rect 13636 1955 13688 1964
rect 13636 1921 13645 1955
rect 13645 1921 13679 1955
rect 13679 1921 13688 1955
rect 13636 1912 13688 1921
rect 14096 1955 14148 1964
rect 14096 1921 14105 1955
rect 14105 1921 14139 1955
rect 14139 1921 14148 1955
rect 14096 1912 14148 1921
rect 16120 1955 16172 1964
rect 16120 1921 16129 1955
rect 16129 1921 16163 1955
rect 16163 1921 16172 1955
rect 16120 1912 16172 1921
rect 16304 1912 16356 1964
rect 22192 1955 22244 1964
rect 22192 1921 22201 1955
rect 22201 1921 22235 1955
rect 22235 1921 22244 1955
rect 22192 1912 22244 1921
rect 22836 1912 22888 1964
rect 22744 1844 22796 1896
rect 23112 1844 23164 1896
rect 24124 1955 24176 1964
rect 24124 1921 24133 1955
rect 24133 1921 24167 1955
rect 24167 1921 24176 1955
rect 24124 1912 24176 1921
rect 7840 1819 7892 1828
rect 7840 1785 7849 1819
rect 7849 1785 7883 1819
rect 7883 1785 7892 1819
rect 7840 1776 7892 1785
rect 22652 1776 22704 1828
rect 16304 1751 16356 1760
rect 16304 1717 16313 1751
rect 16313 1717 16347 1751
rect 16347 1717 16356 1751
rect 16304 1708 16356 1717
rect 3882 1606 3934 1658
rect 3946 1606 3998 1658
rect 4010 1606 4062 1658
rect 4074 1606 4126 1658
rect 4138 1606 4190 1658
rect 9747 1606 9799 1658
rect 9811 1606 9863 1658
rect 9875 1606 9927 1658
rect 9939 1606 9991 1658
rect 10003 1606 10055 1658
rect 15612 1606 15664 1658
rect 15676 1606 15728 1658
rect 15740 1606 15792 1658
rect 15804 1606 15856 1658
rect 15868 1606 15920 1658
rect 21477 1606 21529 1658
rect 21541 1606 21593 1658
rect 21605 1606 21657 1658
rect 21669 1606 21721 1658
rect 21733 1606 21785 1658
rect 7656 1504 7708 1556
rect 8852 1504 8904 1556
rect 10232 1504 10284 1556
rect 10508 1504 10560 1556
rect 11520 1504 11572 1556
rect 12808 1504 12860 1556
rect 13636 1504 13688 1556
rect 16120 1504 16172 1556
rect 22192 1504 22244 1556
rect 22836 1547 22888 1556
rect 22836 1513 22845 1547
rect 22845 1513 22879 1547
rect 22879 1513 22888 1547
rect 22836 1504 22888 1513
rect 23112 1547 23164 1556
rect 23112 1513 23121 1547
rect 23121 1513 23155 1547
rect 23155 1513 23164 1547
rect 23112 1504 23164 1513
rect 23296 1504 23348 1556
rect 24124 1504 24176 1556
rect 848 1300 900 1352
rect 2136 1343 2188 1352
rect 2136 1309 2145 1343
rect 2145 1309 2179 1343
rect 2179 1309 2188 1343
rect 2136 1300 2188 1309
rect 3332 1343 3384 1352
rect 3332 1309 3341 1343
rect 3341 1309 3375 1343
rect 3375 1309 3384 1343
rect 3332 1300 3384 1309
rect 4712 1343 4764 1352
rect 4712 1309 4721 1343
rect 4721 1309 4755 1343
rect 4755 1309 4764 1343
rect 4712 1300 4764 1309
rect 5908 1343 5960 1352
rect 5908 1309 5917 1343
rect 5917 1309 5951 1343
rect 5951 1309 5960 1343
rect 5908 1300 5960 1309
rect 1584 1207 1636 1216
rect 1584 1173 1593 1207
rect 1593 1173 1627 1207
rect 1627 1173 1636 1207
rect 1584 1164 1636 1173
rect 2320 1207 2372 1216
rect 2320 1173 2329 1207
rect 2329 1173 2363 1207
rect 2363 1173 2372 1207
rect 2320 1164 2372 1173
rect 4528 1207 4580 1216
rect 4528 1173 4537 1207
rect 4537 1173 4571 1207
rect 4571 1173 4580 1207
rect 4528 1164 4580 1173
rect 5724 1207 5776 1216
rect 5724 1173 5733 1207
rect 5733 1173 5767 1207
rect 5767 1173 5776 1207
rect 5724 1164 5776 1173
rect 7288 1164 7340 1216
rect 7564 1343 7616 1352
rect 7564 1309 7573 1343
rect 7573 1309 7607 1343
rect 7607 1309 7616 1343
rect 7564 1300 7616 1309
rect 8760 1343 8812 1352
rect 8760 1309 8769 1343
rect 8769 1309 8803 1343
rect 8803 1309 8812 1343
rect 8760 1300 8812 1309
rect 9496 1343 9548 1352
rect 9496 1309 9505 1343
rect 9505 1309 9539 1343
rect 9539 1309 9548 1343
rect 9496 1300 9548 1309
rect 9864 1343 9916 1352
rect 9864 1309 9873 1343
rect 9873 1309 9907 1343
rect 9907 1309 9916 1343
rect 9864 1300 9916 1309
rect 10692 1343 10744 1352
rect 10692 1309 10701 1343
rect 10701 1309 10735 1343
rect 10735 1309 10744 1343
rect 10692 1300 10744 1309
rect 11244 1343 11296 1352
rect 11244 1309 11253 1343
rect 11253 1309 11287 1343
rect 11287 1309 11296 1343
rect 11244 1300 11296 1309
rect 11796 1300 11848 1352
rect 11888 1343 11940 1352
rect 11888 1309 11897 1343
rect 11897 1309 11931 1343
rect 11931 1309 11940 1343
rect 11888 1300 11940 1309
rect 12440 1300 12492 1352
rect 12532 1343 12584 1352
rect 12532 1309 12541 1343
rect 12541 1309 12575 1343
rect 12575 1309 12584 1343
rect 12532 1300 12584 1309
rect 12992 1343 13044 1352
rect 12992 1309 13001 1343
rect 13001 1309 13035 1343
rect 13035 1309 13044 1343
rect 12992 1300 13044 1309
rect 13728 1343 13780 1352
rect 13728 1309 13737 1343
rect 13737 1309 13771 1343
rect 13771 1309 13780 1343
rect 13728 1300 13780 1309
rect 14096 1300 14148 1352
rect 14280 1343 14332 1352
rect 14280 1309 14289 1343
rect 14289 1309 14323 1343
rect 14323 1309 14332 1343
rect 14280 1300 14332 1309
rect 14372 1343 14424 1352
rect 14372 1309 14381 1343
rect 14381 1309 14415 1343
rect 14415 1309 14424 1343
rect 14372 1300 14424 1309
rect 14464 1300 14516 1352
rect 15476 1343 15528 1352
rect 15476 1309 15485 1343
rect 15485 1309 15519 1343
rect 15519 1309 15528 1343
rect 15476 1300 15528 1309
rect 16672 1300 16724 1352
rect 17868 1343 17920 1352
rect 17868 1309 17877 1343
rect 17877 1309 17911 1343
rect 17911 1309 17920 1343
rect 17868 1300 17920 1309
rect 19064 1343 19116 1352
rect 19064 1309 19073 1343
rect 19073 1309 19107 1343
rect 19107 1309 19116 1343
rect 19064 1300 19116 1309
rect 20260 1343 20312 1352
rect 20260 1309 20269 1343
rect 20269 1309 20303 1343
rect 20303 1309 20312 1343
rect 20260 1300 20312 1309
rect 14556 1207 14608 1216
rect 14556 1173 14565 1207
rect 14565 1173 14599 1207
rect 14599 1173 14608 1207
rect 14556 1164 14608 1173
rect 16764 1232 16816 1284
rect 17776 1232 17828 1284
rect 21456 1343 21508 1352
rect 21456 1309 21465 1343
rect 21465 1309 21499 1343
rect 21499 1309 21508 1343
rect 21456 1300 21508 1309
rect 22652 1343 22704 1352
rect 22652 1309 22661 1343
rect 22661 1309 22695 1343
rect 22695 1309 22704 1343
rect 22652 1300 22704 1309
rect 19984 1164 20036 1216
rect 22468 1207 22520 1216
rect 22468 1173 22477 1207
rect 22477 1173 22511 1207
rect 22511 1173 22520 1207
rect 22468 1164 22520 1173
rect 22560 1164 22612 1216
rect 23572 1343 23624 1352
rect 23572 1309 23581 1343
rect 23581 1309 23615 1343
rect 23615 1309 23624 1343
rect 23572 1300 23624 1309
rect 24124 1343 24176 1352
rect 24124 1309 24133 1343
rect 24133 1309 24167 1343
rect 24167 1309 24176 1343
rect 24124 1300 24176 1309
rect 6814 1062 6866 1114
rect 6878 1062 6930 1114
rect 6942 1062 6994 1114
rect 7006 1062 7058 1114
rect 7070 1062 7122 1114
rect 12679 1062 12731 1114
rect 12743 1062 12795 1114
rect 12807 1062 12859 1114
rect 12871 1062 12923 1114
rect 12935 1062 12987 1114
rect 18544 1062 18596 1114
rect 18608 1062 18660 1114
rect 18672 1062 18724 1114
rect 18736 1062 18788 1114
rect 18800 1062 18852 1114
rect 24409 1062 24461 1114
rect 24473 1062 24525 1114
rect 24537 1062 24589 1114
rect 24601 1062 24653 1114
rect 24665 1062 24717 1114
rect 1584 960 1636 1012
rect 4528 960 4580 1012
rect 5724 960 5776 1012
rect 9864 960 9916 1012
rect 13728 960 13780 1012
rect 14372 960 14424 1012
rect 14556 960 14608 1012
rect 19892 960 19944 1012
rect 19984 960 20036 1012
rect 22560 960 22612 1012
rect 7288 892 7340 944
rect 2320 756 2372 808
rect 12532 824 12584 876
rect 23572 688 23624 740
rect 24768 688 24820 740
rect 11244 620 11296 672
rect 6920 552 6972 604
rect 7564 552 7616 604
<< metal2 >>
rect 110 9840 166 10300
rect 386 9840 442 10300
rect 662 9840 718 10300
rect 938 9840 994 10300
rect 1214 9840 1270 10300
rect 1490 9840 1546 10300
rect 1584 9852 1636 9858
rect 124 8838 152 9840
rect 112 8832 164 8838
rect 112 8774 164 8780
rect 400 8616 428 9840
rect 572 8628 624 8634
rect 400 8588 572 8616
rect 572 8570 624 8576
rect 676 6866 704 9840
rect 664 6860 716 6866
rect 664 6802 716 6808
rect 952 6458 980 9840
rect 1228 6798 1256 9840
rect 1504 7478 1532 9840
rect 1766 9840 1822 10300
rect 2042 9840 2098 10300
rect 2228 9988 2280 9994
rect 2228 9930 2280 9936
rect 1584 9794 1636 9800
rect 1492 7472 1544 7478
rect 1492 7414 1544 7420
rect 1596 7410 1624 9794
rect 1676 7540 1728 7546
rect 1780 7528 1808 9840
rect 1952 9240 2004 9246
rect 1952 9182 2004 9188
rect 1964 8498 1992 9182
rect 1952 8492 2004 8498
rect 1952 8434 2004 8440
rect 2056 8090 2084 9840
rect 2044 8084 2096 8090
rect 2044 8026 2096 8032
rect 2240 7818 2268 9930
rect 2318 9840 2374 10300
rect 2594 9840 2650 10300
rect 2870 9840 2926 10300
rect 3146 9840 3202 10300
rect 3422 9840 3478 10300
rect 3698 9840 3754 10300
rect 3974 9840 4030 10300
rect 4250 9840 4306 10300
rect 4526 9840 4582 10300
rect 4802 9840 4858 10300
rect 5078 9840 5134 10300
rect 5354 9840 5410 10300
rect 5630 9840 5686 10300
rect 5906 9840 5962 10300
rect 6000 9852 6052 9858
rect 2332 8090 2360 9840
rect 2412 9716 2464 9722
rect 2412 9658 2464 9664
rect 2320 8084 2372 8090
rect 2320 8026 2372 8032
rect 2424 7886 2452 9658
rect 2504 9240 2556 9246
rect 2504 9182 2556 9188
rect 2516 8498 2544 9182
rect 2504 8492 2556 8498
rect 2504 8434 2556 8440
rect 2608 8004 2636 9840
rect 2884 8634 2912 9840
rect 2964 8832 3016 8838
rect 2964 8774 3016 8780
rect 2976 8634 3004 8774
rect 2872 8628 2924 8634
rect 2872 8570 2924 8576
rect 2964 8628 3016 8634
rect 2964 8570 3016 8576
rect 3160 8072 3188 9840
rect 3436 8362 3464 9840
rect 3424 8356 3476 8362
rect 3424 8298 3476 8304
rect 3240 8084 3292 8090
rect 3160 8044 3240 8072
rect 3240 8026 3292 8032
rect 2780 8016 2832 8022
rect 2608 7976 2780 8004
rect 2780 7958 2832 7964
rect 2412 7880 2464 7886
rect 2596 7880 2648 7886
rect 2412 7822 2464 7828
rect 2594 7848 2596 7857
rect 2648 7848 2650 7857
rect 2228 7812 2280 7818
rect 2594 7783 2650 7792
rect 2228 7754 2280 7760
rect 3712 7546 3740 9840
rect 3988 8378 4016 9840
rect 4160 9104 4212 9110
rect 4160 9046 4212 9052
rect 4172 8634 4200 9046
rect 4264 8634 4292 9840
rect 4436 8832 4488 8838
rect 4436 8774 4488 8780
rect 4160 8628 4212 8634
rect 4160 8570 4212 8576
rect 4252 8628 4304 8634
rect 4252 8570 4304 8576
rect 4448 8498 4476 8774
rect 4436 8492 4488 8498
rect 4436 8434 4488 8440
rect 3988 8350 4292 8378
rect 3882 8188 4190 8197
rect 3882 8186 3888 8188
rect 3944 8186 3968 8188
rect 4024 8186 4048 8188
rect 4104 8186 4128 8188
rect 4184 8186 4190 8188
rect 3944 8134 3946 8186
rect 4126 8134 4128 8186
rect 3882 8132 3888 8134
rect 3944 8132 3968 8134
rect 4024 8132 4048 8134
rect 4104 8132 4128 8134
rect 4184 8132 4190 8134
rect 3882 8123 4190 8132
rect 4160 8016 4212 8022
rect 4264 8004 4292 8350
rect 4540 8072 4568 9840
rect 4816 8090 4844 9840
rect 4896 8832 4948 8838
rect 4896 8774 4948 8780
rect 4908 8498 4936 8774
rect 5092 8634 5120 9840
rect 5368 8634 5396 9840
rect 5540 9036 5592 9042
rect 5540 8978 5592 8984
rect 5080 8628 5132 8634
rect 5080 8570 5132 8576
rect 5356 8628 5408 8634
rect 5356 8570 5408 8576
rect 4896 8492 4948 8498
rect 4896 8434 4948 8440
rect 4620 8084 4672 8090
rect 4540 8044 4620 8072
rect 4620 8026 4672 8032
rect 4804 8084 4856 8090
rect 4804 8026 4856 8032
rect 4212 7976 4292 8004
rect 4160 7958 4212 7964
rect 5448 7948 5500 7954
rect 5448 7890 5500 7896
rect 1728 7500 1808 7528
rect 3700 7540 3752 7546
rect 1676 7482 1728 7488
rect 3700 7482 3752 7488
rect 1584 7404 1636 7410
rect 1584 7346 1636 7352
rect 2780 7200 2832 7206
rect 2780 7142 2832 7148
rect 2792 6866 2820 7142
rect 3882 7100 4190 7109
rect 3882 7098 3888 7100
rect 3944 7098 3968 7100
rect 4024 7098 4048 7100
rect 4104 7098 4128 7100
rect 4184 7098 4190 7100
rect 3944 7046 3946 7098
rect 4126 7046 4128 7098
rect 3882 7044 3888 7046
rect 3944 7044 3968 7046
rect 4024 7044 4048 7046
rect 4104 7044 4128 7046
rect 4184 7044 4190 7046
rect 3882 7035 4190 7044
rect 2780 6860 2832 6866
rect 2780 6802 2832 6808
rect 1216 6792 1268 6798
rect 1216 6734 1268 6740
rect 2686 6760 2742 6769
rect 2686 6695 2688 6704
rect 2740 6695 2742 6704
rect 2688 6666 2740 6672
rect 940 6452 992 6458
rect 940 6394 992 6400
rect 5460 6390 5488 7890
rect 5552 7818 5580 8978
rect 5644 8072 5672 9840
rect 5920 8634 5948 9840
rect 6182 9840 6238 10300
rect 6458 9840 6514 10300
rect 6734 9840 6790 10300
rect 7010 9840 7066 10300
rect 7116 9846 7236 9874
rect 7116 9840 7144 9846
rect 6000 9794 6052 9800
rect 5908 8628 5960 8634
rect 5908 8570 5960 8576
rect 5816 8492 5868 8498
rect 5816 8434 5868 8440
rect 5908 8492 5960 8498
rect 5908 8434 5960 8440
rect 5724 8084 5776 8090
rect 5644 8044 5724 8072
rect 5724 8026 5776 8032
rect 5540 7812 5592 7818
rect 5540 7754 5592 7760
rect 5632 7812 5684 7818
rect 5632 7754 5684 7760
rect 5644 7546 5672 7754
rect 5632 7540 5684 7546
rect 5632 7482 5684 7488
rect 5630 7440 5686 7449
rect 5630 7375 5632 7384
rect 5684 7375 5686 7384
rect 5632 7346 5684 7352
rect 5828 7206 5856 8434
rect 5920 7546 5948 8434
rect 5908 7540 5960 7546
rect 5908 7482 5960 7488
rect 6012 7478 6040 9794
rect 6196 8072 6224 9840
rect 6368 9376 6420 9382
rect 6368 9318 6420 9324
rect 6276 8084 6328 8090
rect 6196 8044 6276 8072
rect 6276 8026 6328 8032
rect 6000 7472 6052 7478
rect 6000 7414 6052 7420
rect 6380 7410 6408 9318
rect 6472 8634 6500 9840
rect 6552 9512 6604 9518
rect 6552 9454 6604 9460
rect 6460 8628 6512 8634
rect 6460 8570 6512 8576
rect 6564 8566 6592 9454
rect 6552 8560 6604 8566
rect 6552 8502 6604 8508
rect 6644 8356 6696 8362
rect 6644 8298 6696 8304
rect 6656 7886 6684 8298
rect 6748 8004 6776 9840
rect 7024 9812 7144 9840
rect 6814 8732 7122 8741
rect 6814 8730 6820 8732
rect 6876 8730 6900 8732
rect 6956 8730 6980 8732
rect 7036 8730 7060 8732
rect 7116 8730 7122 8732
rect 6876 8678 6878 8730
rect 7058 8678 7060 8730
rect 6814 8676 6820 8678
rect 6876 8676 6900 8678
rect 6956 8676 6980 8678
rect 7036 8676 7060 8678
rect 7116 8676 7122 8678
rect 6814 8667 7122 8676
rect 7208 8634 7236 9846
rect 7286 9840 7342 10300
rect 7562 9840 7618 10300
rect 7838 9840 7894 10300
rect 8114 9840 8170 10300
rect 8390 9840 8446 10300
rect 8666 9840 8722 10300
rect 8942 9840 8998 10300
rect 9218 9840 9274 10300
rect 9494 9840 9550 10300
rect 9770 9840 9826 10300
rect 10046 9840 10102 10300
rect 10152 9846 10272 9874
rect 10152 9840 10180 9846
rect 7196 8628 7248 8634
rect 7196 8570 7248 8576
rect 7196 8492 7248 8498
rect 7196 8434 7248 8440
rect 6920 8016 6972 8022
rect 6748 7976 6920 8004
rect 6920 7958 6972 7964
rect 6644 7880 6696 7886
rect 6644 7822 6696 7828
rect 6734 7848 6790 7857
rect 6552 7812 6604 7818
rect 6734 7783 6736 7792
rect 6552 7754 6604 7760
rect 6788 7783 6790 7792
rect 6736 7754 6788 7760
rect 6184 7404 6236 7410
rect 6184 7346 6236 7352
rect 6368 7404 6420 7410
rect 6368 7346 6420 7352
rect 6196 7313 6224 7346
rect 6182 7304 6238 7313
rect 6182 7239 6238 7248
rect 5816 7200 5868 7206
rect 5816 7142 5868 7148
rect 6564 7002 6592 7754
rect 6814 7644 7122 7653
rect 6814 7642 6820 7644
rect 6876 7642 6900 7644
rect 6956 7642 6980 7644
rect 7036 7642 7060 7644
rect 7116 7642 7122 7644
rect 6876 7590 6878 7642
rect 7058 7590 7060 7642
rect 6814 7588 6820 7590
rect 6876 7588 6900 7590
rect 6956 7588 6980 7590
rect 7036 7588 7060 7590
rect 7116 7588 7122 7590
rect 6814 7579 7122 7588
rect 7208 7546 7236 8434
rect 7300 8090 7328 9840
rect 7576 8634 7604 9840
rect 7656 9784 7708 9790
rect 7656 9726 7708 9732
rect 7564 8628 7616 8634
rect 7564 8570 7616 8576
rect 7380 8424 7432 8430
rect 7380 8366 7432 8372
rect 7288 8084 7340 8090
rect 7288 8026 7340 8032
rect 7392 7886 7420 8366
rect 7380 7880 7432 7886
rect 7380 7822 7432 7828
rect 7668 7818 7696 9726
rect 7748 9172 7800 9178
rect 7748 9114 7800 9120
rect 7760 8022 7788 9114
rect 7852 8072 7880 9840
rect 7932 9512 7984 9518
rect 7932 9454 7984 9460
rect 7944 8412 7972 9454
rect 8024 8832 8076 8838
rect 8024 8774 8076 8780
rect 8036 8566 8064 8774
rect 8128 8634 8156 9840
rect 8208 9376 8260 9382
rect 8208 9318 8260 9324
rect 8116 8628 8168 8634
rect 8116 8570 8168 8576
rect 8024 8560 8076 8566
rect 8024 8502 8076 8508
rect 7944 8384 8064 8412
rect 7932 8084 7984 8090
rect 7852 8044 7932 8072
rect 7932 8026 7984 8032
rect 7748 8016 7800 8022
rect 8036 7970 8064 8384
rect 7748 7958 7800 7964
rect 7852 7942 8064 7970
rect 7852 7818 7880 7942
rect 7656 7812 7708 7818
rect 7656 7754 7708 7760
rect 7840 7812 7892 7818
rect 7840 7754 7892 7760
rect 7196 7540 7248 7546
rect 7196 7482 7248 7488
rect 7380 7404 7432 7410
rect 7380 7346 7432 7352
rect 7392 7206 7420 7346
rect 8220 7342 8248 9318
rect 8404 8634 8432 9840
rect 8392 8628 8444 8634
rect 8392 8570 8444 8576
rect 8300 8424 8352 8430
rect 8300 8366 8352 8372
rect 8312 7546 8340 8366
rect 8680 8090 8708 9840
rect 8956 8634 8984 9840
rect 9036 9308 9088 9314
rect 9036 9250 9088 9256
rect 8944 8628 8996 8634
rect 8944 8570 8996 8576
rect 8668 8084 8720 8090
rect 8668 8026 8720 8032
rect 9048 8022 9076 9250
rect 9232 8634 9260 9840
rect 9508 9654 9536 9840
rect 9496 9648 9548 9654
rect 9496 9590 9548 9596
rect 9588 9308 9640 9314
rect 9588 9250 9640 9256
rect 9404 8900 9456 8906
rect 9404 8842 9456 8848
rect 9220 8628 9272 8634
rect 9220 8570 9272 8576
rect 9416 8090 9444 8842
rect 9600 8566 9628 9250
rect 9680 8628 9732 8634
rect 9784 8616 9812 9840
rect 10060 9812 10180 9840
rect 10140 9648 10192 9654
rect 10140 9590 10192 9596
rect 10152 9330 10180 9590
rect 10244 9466 10272 9846
rect 10322 9840 10378 10300
rect 10428 9846 10548 9874
rect 10428 9840 10456 9846
rect 10336 9812 10456 9840
rect 10244 9438 10364 9466
rect 10152 9302 10272 9330
rect 10048 8968 10100 8974
rect 10048 8910 10100 8916
rect 9956 8900 10008 8906
rect 9956 8842 10008 8848
rect 9968 8634 9996 8842
rect 9732 8588 9812 8616
rect 9956 8628 10008 8634
rect 9680 8570 9732 8576
rect 9956 8570 10008 8576
rect 9588 8560 9640 8566
rect 9588 8502 9640 8508
rect 10060 8378 10088 8910
rect 10244 8634 10272 9302
rect 10232 8628 10284 8634
rect 10232 8570 10284 8576
rect 10230 8528 10286 8537
rect 10230 8463 10286 8472
rect 10244 8430 10272 8463
rect 10232 8424 10284 8430
rect 10060 8350 10180 8378
rect 10232 8366 10284 8372
rect 9747 8188 10055 8197
rect 9747 8186 9753 8188
rect 9809 8186 9833 8188
rect 9889 8186 9913 8188
rect 9969 8186 9993 8188
rect 10049 8186 10055 8188
rect 9809 8134 9811 8186
rect 9991 8134 9993 8186
rect 9747 8132 9753 8134
rect 9809 8132 9833 8134
rect 9889 8132 9913 8134
rect 9969 8132 9993 8134
rect 10049 8132 10055 8134
rect 9747 8123 10055 8132
rect 9404 8084 9456 8090
rect 9404 8026 9456 8032
rect 9772 8084 9824 8090
rect 9772 8026 9824 8032
rect 9036 8016 9088 8022
rect 9036 7958 9088 7964
rect 9784 7886 9812 8026
rect 8484 7880 8536 7886
rect 8484 7822 8536 7828
rect 9588 7880 9640 7886
rect 9588 7822 9640 7828
rect 9772 7880 9824 7886
rect 9772 7822 9824 7828
rect 8496 7546 8524 7822
rect 9036 7812 9088 7818
rect 9036 7754 9088 7760
rect 8852 7744 8904 7750
rect 8852 7686 8904 7692
rect 8300 7540 8352 7546
rect 8300 7482 8352 7488
rect 8484 7540 8536 7546
rect 8484 7482 8536 7488
rect 8864 7478 8892 7686
rect 8852 7472 8904 7478
rect 8852 7414 8904 7420
rect 8392 7404 8444 7410
rect 8668 7404 8720 7410
rect 8444 7364 8668 7392
rect 8392 7346 8444 7352
rect 8668 7346 8720 7352
rect 8208 7336 8260 7342
rect 8208 7278 8260 7284
rect 9048 7206 9076 7754
rect 9600 7392 9628 7822
rect 10152 7750 10180 8350
rect 10140 7744 10192 7750
rect 10140 7686 10192 7692
rect 10336 7410 10364 9438
rect 10416 8900 10468 8906
rect 10416 8842 10468 8848
rect 10428 8362 10456 8842
rect 10416 8356 10468 8362
rect 10416 8298 10468 8304
rect 10520 7868 10548 9846
rect 10598 9840 10654 10300
rect 10704 9846 10824 9874
rect 10704 9840 10732 9846
rect 10612 9812 10732 9840
rect 10600 7880 10652 7886
rect 10520 7840 10600 7868
rect 10796 7868 10824 9846
rect 10874 9840 10930 10300
rect 11150 9840 11206 10300
rect 11256 9846 11376 9874
rect 11256 9840 11284 9846
rect 10888 9330 10916 9840
rect 11164 9812 11284 9840
rect 11244 9444 11296 9450
rect 11244 9386 11296 9392
rect 10888 9302 11008 9330
rect 10876 9036 10928 9042
rect 10876 8978 10928 8984
rect 10888 8362 10916 8978
rect 10876 8356 10928 8362
rect 10876 8298 10928 8304
rect 10876 7880 10928 7886
rect 10796 7840 10876 7868
rect 10600 7822 10652 7828
rect 10980 7868 11008 9302
rect 11256 9178 11284 9386
rect 11152 9172 11204 9178
rect 11152 9114 11204 9120
rect 11244 9172 11296 9178
rect 11244 9114 11296 9120
rect 11164 8566 11192 9114
rect 11152 8560 11204 8566
rect 11152 8502 11204 8508
rect 11060 8492 11112 8498
rect 11060 8434 11112 8440
rect 11072 8022 11100 8434
rect 11060 8016 11112 8022
rect 11060 7958 11112 7964
rect 11152 7880 11204 7886
rect 10980 7840 11152 7868
rect 10876 7822 10928 7828
rect 11348 7868 11376 9846
rect 11426 9840 11482 10300
rect 11532 9846 11652 9874
rect 11532 9840 11560 9846
rect 11440 9812 11560 9840
rect 11520 9648 11572 9654
rect 11520 9590 11572 9596
rect 11532 8616 11560 9590
rect 11440 8588 11560 8616
rect 11440 7970 11468 8588
rect 11520 8492 11572 8498
rect 11520 8434 11572 8440
rect 11532 8090 11560 8434
rect 11520 8084 11572 8090
rect 11520 8026 11572 8032
rect 11440 7942 11560 7970
rect 11428 7880 11480 7886
rect 11348 7840 11428 7868
rect 11152 7822 11204 7828
rect 11428 7822 11480 7828
rect 10324 7404 10376 7410
rect 9600 7364 9674 7392
rect 9324 7274 9536 7290
rect 9312 7268 9548 7274
rect 9364 7262 9496 7268
rect 9312 7210 9364 7216
rect 9496 7210 9548 7216
rect 9646 7206 9674 7364
rect 10324 7346 10376 7352
rect 7380 7200 7432 7206
rect 7380 7142 7432 7148
rect 9036 7200 9088 7206
rect 9036 7142 9088 7148
rect 9634 7200 9686 7206
rect 9634 7142 9686 7148
rect 9747 7100 10055 7109
rect 9747 7098 9753 7100
rect 9809 7098 9833 7100
rect 9889 7098 9913 7100
rect 9969 7098 9993 7100
rect 10049 7098 10055 7100
rect 9809 7046 9811 7098
rect 9991 7046 9993 7098
rect 9747 7044 9753 7046
rect 9809 7044 9833 7046
rect 9889 7044 9913 7046
rect 9969 7044 9993 7046
rect 10049 7044 10055 7046
rect 9747 7035 10055 7044
rect 6552 6996 6604 7002
rect 6552 6938 6604 6944
rect 6814 6556 7122 6565
rect 6814 6554 6820 6556
rect 6876 6554 6900 6556
rect 6956 6554 6980 6556
rect 7036 6554 7060 6556
rect 7116 6554 7122 6556
rect 6876 6502 6878 6554
rect 7058 6502 7060 6554
rect 6814 6500 6820 6502
rect 6876 6500 6900 6502
rect 6956 6500 6980 6502
rect 7036 6500 7060 6502
rect 7116 6500 7122 6502
rect 6814 6491 7122 6500
rect 5448 6384 5500 6390
rect 5448 6326 5500 6332
rect 3882 6012 4190 6021
rect 3882 6010 3888 6012
rect 3944 6010 3968 6012
rect 4024 6010 4048 6012
rect 4104 6010 4128 6012
rect 4184 6010 4190 6012
rect 3944 5958 3946 6010
rect 4126 5958 4128 6010
rect 3882 5956 3888 5958
rect 3944 5956 3968 5958
rect 4024 5956 4048 5958
rect 4104 5956 4128 5958
rect 4184 5956 4190 5958
rect 3882 5947 4190 5956
rect 9747 6012 10055 6021
rect 9747 6010 9753 6012
rect 9809 6010 9833 6012
rect 9889 6010 9913 6012
rect 9969 6010 9993 6012
rect 10049 6010 10055 6012
rect 9809 5958 9811 6010
rect 9991 5958 9993 6010
rect 9747 5956 9753 5958
rect 9809 5956 9833 5958
rect 9889 5956 9913 5958
rect 9969 5956 9993 5958
rect 10049 5956 10055 5958
rect 9747 5947 10055 5956
rect 6814 5468 7122 5477
rect 6814 5466 6820 5468
rect 6876 5466 6900 5468
rect 6956 5466 6980 5468
rect 7036 5466 7060 5468
rect 7116 5466 7122 5468
rect 6876 5414 6878 5466
rect 7058 5414 7060 5466
rect 6814 5412 6820 5414
rect 6876 5412 6900 5414
rect 6956 5412 6980 5414
rect 7036 5412 7060 5414
rect 7116 5412 7122 5414
rect 6814 5403 7122 5412
rect 3882 4924 4190 4933
rect 3882 4922 3888 4924
rect 3944 4922 3968 4924
rect 4024 4922 4048 4924
rect 4104 4922 4128 4924
rect 4184 4922 4190 4924
rect 3944 4870 3946 4922
rect 4126 4870 4128 4922
rect 3882 4868 3888 4870
rect 3944 4868 3968 4870
rect 4024 4868 4048 4870
rect 4104 4868 4128 4870
rect 4184 4868 4190 4870
rect 3882 4859 4190 4868
rect 9747 4924 10055 4933
rect 9747 4922 9753 4924
rect 9809 4922 9833 4924
rect 9889 4922 9913 4924
rect 9969 4922 9993 4924
rect 10049 4922 10055 4924
rect 9809 4870 9811 4922
rect 9991 4870 9993 4922
rect 9747 4868 9753 4870
rect 9809 4868 9833 4870
rect 9889 4868 9913 4870
rect 9969 4868 9993 4870
rect 10049 4868 10055 4870
rect 9747 4859 10055 4868
rect 6814 4380 7122 4389
rect 6814 4378 6820 4380
rect 6876 4378 6900 4380
rect 6956 4378 6980 4380
rect 7036 4378 7060 4380
rect 7116 4378 7122 4380
rect 6876 4326 6878 4378
rect 7058 4326 7060 4378
rect 6814 4324 6820 4326
rect 6876 4324 6900 4326
rect 6956 4324 6980 4326
rect 7036 4324 7060 4326
rect 7116 4324 7122 4326
rect 6814 4315 7122 4324
rect 3882 3836 4190 3845
rect 3882 3834 3888 3836
rect 3944 3834 3968 3836
rect 4024 3834 4048 3836
rect 4104 3834 4128 3836
rect 4184 3834 4190 3836
rect 3944 3782 3946 3834
rect 4126 3782 4128 3834
rect 3882 3780 3888 3782
rect 3944 3780 3968 3782
rect 4024 3780 4048 3782
rect 4104 3780 4128 3782
rect 4184 3780 4190 3782
rect 3882 3771 4190 3780
rect 9747 3836 10055 3845
rect 9747 3834 9753 3836
rect 9809 3834 9833 3836
rect 9889 3834 9913 3836
rect 9969 3834 9993 3836
rect 10049 3834 10055 3836
rect 9809 3782 9811 3834
rect 9991 3782 9993 3834
rect 9747 3780 9753 3782
rect 9809 3780 9833 3782
rect 9889 3780 9913 3782
rect 9969 3780 9993 3782
rect 10049 3780 10055 3782
rect 9747 3771 10055 3780
rect 6814 3292 7122 3301
rect 6814 3290 6820 3292
rect 6876 3290 6900 3292
rect 6956 3290 6980 3292
rect 7036 3290 7060 3292
rect 7116 3290 7122 3292
rect 6876 3238 6878 3290
rect 7058 3238 7060 3290
rect 6814 3236 6820 3238
rect 6876 3236 6900 3238
rect 6956 3236 6980 3238
rect 7036 3236 7060 3238
rect 7116 3236 7122 3238
rect 6814 3227 7122 3236
rect 3882 2748 4190 2757
rect 3882 2746 3888 2748
rect 3944 2746 3968 2748
rect 4024 2746 4048 2748
rect 4104 2746 4128 2748
rect 4184 2746 4190 2748
rect 3944 2694 3946 2746
rect 4126 2694 4128 2746
rect 3882 2692 3888 2694
rect 3944 2692 3968 2694
rect 4024 2692 4048 2694
rect 4104 2692 4128 2694
rect 4184 2692 4190 2694
rect 3882 2683 4190 2692
rect 9747 2748 10055 2757
rect 9747 2746 9753 2748
rect 9809 2746 9833 2748
rect 9889 2746 9913 2748
rect 9969 2746 9993 2748
rect 10049 2746 10055 2748
rect 9809 2694 9811 2746
rect 9991 2694 9993 2746
rect 9747 2692 9753 2694
rect 9809 2692 9833 2694
rect 9889 2692 9913 2694
rect 9969 2692 9993 2694
rect 10049 2692 10055 2694
rect 9747 2683 10055 2692
rect 10690 2408 10746 2417
rect 10690 2343 10746 2352
rect 10416 2304 10468 2310
rect 10416 2246 10468 2252
rect 6814 2204 7122 2213
rect 6814 2202 6820 2204
rect 6876 2202 6900 2204
rect 6956 2202 6980 2204
rect 7036 2202 7060 2204
rect 7116 2202 7122 2204
rect 6876 2150 6878 2202
rect 7058 2150 7060 2202
rect 6814 2148 6820 2150
rect 6876 2148 6900 2150
rect 6956 2148 6980 2150
rect 7036 2148 7060 2150
rect 7116 2148 7122 2150
rect 6814 2139 7122 2148
rect 10428 2106 10456 2246
rect 10704 2106 10732 2343
rect 11532 2106 11560 7942
rect 11624 7868 11652 9846
rect 11702 9840 11758 10300
rect 11796 9988 11848 9994
rect 11796 9930 11848 9936
rect 11888 9988 11940 9994
rect 11888 9930 11940 9936
rect 11716 8498 11744 9840
rect 11808 9178 11836 9930
rect 11900 9518 11928 9930
rect 11978 9840 12034 10300
rect 12254 9840 12310 10300
rect 12530 9840 12586 10300
rect 12806 9840 12862 10300
rect 12912 9846 13032 9874
rect 12912 9840 12940 9846
rect 11888 9512 11940 9518
rect 11888 9454 11940 9460
rect 11796 9172 11848 9178
rect 11796 9114 11848 9120
rect 11704 8492 11756 8498
rect 11704 8434 11756 8440
rect 11796 8288 11848 8294
rect 11796 8230 11848 8236
rect 11704 7880 11756 7886
rect 11624 7840 11704 7868
rect 11704 7822 11756 7828
rect 11612 7744 11664 7750
rect 11612 7686 11664 7692
rect 11624 7342 11652 7686
rect 11808 7478 11836 8230
rect 11992 7886 12020 9840
rect 12072 9376 12124 9382
rect 12072 9318 12124 9324
rect 12084 8294 12112 9318
rect 12072 8288 12124 8294
rect 12072 8230 12124 8236
rect 11980 7880 12032 7886
rect 12268 7868 12296 9840
rect 12348 9036 12400 9042
rect 12348 8978 12400 8984
rect 12360 8362 12388 8978
rect 12544 8514 12572 9840
rect 12820 9812 12940 9840
rect 13004 9738 13032 9846
rect 13082 9840 13138 10300
rect 13188 9846 13308 9874
rect 13188 9840 13216 9846
rect 13096 9812 13216 9840
rect 13004 9710 13124 9738
rect 12679 8732 12987 8741
rect 12679 8730 12685 8732
rect 12741 8730 12765 8732
rect 12821 8730 12845 8732
rect 12901 8730 12925 8732
rect 12981 8730 12987 8732
rect 12741 8678 12743 8730
rect 12923 8678 12925 8730
rect 12679 8676 12685 8678
rect 12741 8676 12765 8678
rect 12821 8676 12845 8678
rect 12901 8676 12925 8678
rect 12981 8676 12987 8678
rect 12679 8667 12987 8676
rect 12900 8628 12952 8634
rect 12900 8570 12952 8576
rect 12544 8486 12664 8514
rect 12440 8424 12492 8430
rect 12440 8366 12492 8372
rect 12348 8356 12400 8362
rect 12348 8298 12400 8304
rect 12452 8090 12480 8366
rect 12440 8084 12492 8090
rect 12440 8026 12492 8032
rect 12532 7880 12584 7886
rect 12268 7840 12532 7868
rect 11980 7822 12032 7828
rect 12636 7868 12664 8486
rect 12912 8090 12940 8570
rect 12900 8084 12952 8090
rect 12900 8026 12952 8032
rect 13096 7886 13124 9710
rect 13176 8424 13228 8430
rect 13176 8366 13228 8372
rect 13188 8090 13216 8366
rect 13176 8084 13228 8090
rect 13176 8026 13228 8032
rect 12808 7880 12860 7886
rect 12636 7840 12808 7868
rect 12532 7822 12584 7828
rect 12808 7822 12860 7828
rect 13084 7880 13136 7886
rect 13280 7868 13308 9846
rect 13358 9840 13414 10300
rect 13634 9840 13690 10300
rect 13910 9840 13966 10300
rect 14186 9840 14242 10300
rect 14280 9920 14332 9926
rect 14280 9862 14332 9868
rect 13372 8498 13400 9840
rect 13452 9240 13504 9246
rect 13452 9182 13504 9188
rect 13360 8492 13412 8498
rect 13360 8434 13412 8440
rect 13464 8362 13492 9182
rect 13648 8498 13676 9840
rect 13636 8492 13688 8498
rect 13924 8480 13952 9840
rect 14200 8566 14228 9840
rect 14188 8560 14240 8566
rect 14188 8502 14240 8508
rect 14004 8492 14056 8498
rect 13924 8452 14004 8480
rect 13636 8434 13688 8440
rect 14004 8434 14056 8440
rect 14292 8362 14320 9862
rect 14462 9840 14518 10300
rect 14648 9852 14700 9858
rect 13452 8356 13504 8362
rect 13452 8298 13504 8304
rect 13636 8356 13688 8362
rect 13636 8298 13688 8304
rect 14280 8356 14332 8362
rect 14280 8298 14332 8304
rect 13648 7993 13676 8298
rect 13634 7984 13690 7993
rect 13634 7919 13690 7928
rect 14476 7886 14504 9840
rect 14738 9840 14794 10300
rect 14844 9846 14964 9874
rect 14844 9840 14872 9846
rect 14752 9812 14872 9840
rect 14648 9794 14700 9800
rect 14556 9172 14608 9178
rect 14556 9114 14608 9120
rect 14568 8634 14596 9114
rect 14660 8650 14688 9794
rect 14832 9716 14884 9722
rect 14832 9658 14884 9664
rect 14556 8628 14608 8634
rect 14660 8622 14780 8650
rect 14844 8634 14872 9658
rect 14556 8570 14608 8576
rect 14752 8498 14780 8622
rect 14832 8628 14884 8634
rect 14832 8570 14884 8576
rect 14648 8492 14700 8498
rect 14648 8434 14700 8440
rect 14740 8492 14792 8498
rect 14740 8434 14792 8440
rect 14660 8090 14688 8434
rect 14648 8084 14700 8090
rect 14648 8026 14700 8032
rect 13360 7880 13412 7886
rect 13280 7840 13360 7868
rect 13084 7822 13136 7828
rect 13360 7822 13412 7828
rect 14464 7880 14516 7886
rect 14936 7868 14964 9846
rect 15014 9840 15070 10300
rect 15290 9840 15346 10300
rect 15396 9846 15516 9874
rect 15396 9840 15424 9846
rect 15028 8922 15056 9840
rect 15304 9812 15424 9840
rect 15384 9308 15436 9314
rect 15384 9250 15436 9256
rect 15028 8894 15148 8922
rect 15016 8628 15068 8634
rect 15016 8570 15068 8576
rect 15028 8537 15056 8570
rect 15014 8528 15070 8537
rect 15014 8463 15070 8472
rect 15016 7880 15068 7886
rect 14936 7840 15016 7868
rect 14464 7822 14516 7828
rect 15120 7868 15148 8894
rect 15396 8566 15424 9250
rect 15384 8560 15436 8566
rect 15384 8502 15436 8508
rect 15200 8492 15252 8498
rect 15200 8434 15252 8440
rect 15292 8492 15344 8498
rect 15292 8434 15344 8440
rect 15212 8090 15240 8434
rect 15304 8090 15332 8434
rect 15384 8424 15436 8430
rect 15384 8366 15436 8372
rect 15396 8090 15424 8366
rect 15200 8084 15252 8090
rect 15200 8026 15252 8032
rect 15292 8084 15344 8090
rect 15292 8026 15344 8032
rect 15384 8084 15436 8090
rect 15384 8026 15436 8032
rect 15292 7880 15344 7886
rect 15120 7840 15292 7868
rect 15016 7822 15068 7828
rect 15488 7868 15516 9846
rect 15566 9840 15622 10300
rect 15672 9846 15792 9874
rect 15672 9840 15700 9846
rect 15580 9812 15700 9840
rect 15764 9738 15792 9846
rect 15842 9840 15898 10300
rect 15948 9846 16068 9874
rect 15948 9840 15976 9846
rect 15856 9812 15976 9840
rect 15764 9710 15976 9738
rect 15842 8392 15898 8401
rect 15842 8327 15898 8336
rect 15856 8294 15884 8327
rect 15844 8288 15896 8294
rect 15844 8230 15896 8236
rect 15612 8188 15920 8197
rect 15612 8186 15618 8188
rect 15674 8186 15698 8188
rect 15754 8186 15778 8188
rect 15834 8186 15858 8188
rect 15914 8186 15920 8188
rect 15674 8134 15676 8186
rect 15856 8134 15858 8186
rect 15612 8132 15618 8134
rect 15674 8132 15698 8134
rect 15754 8132 15778 8134
rect 15834 8132 15858 8134
rect 15914 8132 15920 8134
rect 15612 8123 15920 8132
rect 15568 7880 15620 7886
rect 15488 7840 15568 7868
rect 15292 7822 15344 7828
rect 15568 7822 15620 7828
rect 15844 7880 15896 7886
rect 15948 7868 15976 9710
rect 15896 7840 15976 7868
rect 16040 7868 16068 9846
rect 16118 9840 16174 10300
rect 16224 9846 16344 9874
rect 16224 9840 16252 9846
rect 16132 9812 16252 9840
rect 16212 8968 16264 8974
rect 16212 8910 16264 8916
rect 16120 8492 16172 8498
rect 16120 8434 16172 8440
rect 16132 8090 16160 8434
rect 16224 8362 16252 8910
rect 16212 8356 16264 8362
rect 16212 8298 16264 8304
rect 16120 8084 16172 8090
rect 16120 8026 16172 8032
rect 16212 7948 16264 7954
rect 16212 7890 16264 7896
rect 16120 7880 16172 7886
rect 16040 7840 16120 7868
rect 15844 7822 15896 7828
rect 16120 7822 16172 7828
rect 12679 7644 12987 7653
rect 12679 7642 12685 7644
rect 12741 7642 12765 7644
rect 12821 7642 12845 7644
rect 12901 7642 12925 7644
rect 12981 7642 12987 7644
rect 12741 7590 12743 7642
rect 12923 7590 12925 7642
rect 12679 7588 12685 7590
rect 12741 7588 12765 7590
rect 12821 7588 12845 7590
rect 12901 7588 12925 7590
rect 12981 7588 12987 7590
rect 12679 7579 12987 7588
rect 11796 7472 11848 7478
rect 11796 7414 11848 7420
rect 11612 7336 11664 7342
rect 11612 7278 11664 7284
rect 15612 7100 15920 7109
rect 15612 7098 15618 7100
rect 15674 7098 15698 7100
rect 15754 7098 15778 7100
rect 15834 7098 15858 7100
rect 15914 7098 15920 7100
rect 15674 7046 15676 7098
rect 15856 7046 15858 7098
rect 15612 7044 15618 7046
rect 15674 7044 15698 7046
rect 15754 7044 15778 7046
rect 15834 7044 15858 7046
rect 15914 7044 15920 7046
rect 15612 7035 15920 7044
rect 12679 6556 12987 6565
rect 12679 6554 12685 6556
rect 12741 6554 12765 6556
rect 12821 6554 12845 6556
rect 12901 6554 12925 6556
rect 12981 6554 12987 6556
rect 12741 6502 12743 6554
rect 12923 6502 12925 6554
rect 12679 6500 12685 6502
rect 12741 6500 12765 6502
rect 12821 6500 12845 6502
rect 12901 6500 12925 6502
rect 12981 6500 12987 6502
rect 12679 6491 12987 6500
rect 15612 6012 15920 6021
rect 15612 6010 15618 6012
rect 15674 6010 15698 6012
rect 15754 6010 15778 6012
rect 15834 6010 15858 6012
rect 15914 6010 15920 6012
rect 15674 5958 15676 6010
rect 15856 5958 15858 6010
rect 15612 5956 15618 5958
rect 15674 5956 15698 5958
rect 15754 5956 15778 5958
rect 15834 5956 15858 5958
rect 15914 5956 15920 5958
rect 15612 5947 15920 5956
rect 12679 5468 12987 5477
rect 12679 5466 12685 5468
rect 12741 5466 12765 5468
rect 12821 5466 12845 5468
rect 12901 5466 12925 5468
rect 12981 5466 12987 5468
rect 12741 5414 12743 5466
rect 12923 5414 12925 5466
rect 12679 5412 12685 5414
rect 12741 5412 12765 5414
rect 12821 5412 12845 5414
rect 12901 5412 12925 5414
rect 12981 5412 12987 5414
rect 12679 5403 12987 5412
rect 15612 4924 15920 4933
rect 15612 4922 15618 4924
rect 15674 4922 15698 4924
rect 15754 4922 15778 4924
rect 15834 4922 15858 4924
rect 15914 4922 15920 4924
rect 15674 4870 15676 4922
rect 15856 4870 15858 4922
rect 15612 4868 15618 4870
rect 15674 4868 15698 4870
rect 15754 4868 15778 4870
rect 15834 4868 15858 4870
rect 15914 4868 15920 4870
rect 15612 4859 15920 4868
rect 14832 4616 14884 4622
rect 14832 4558 14884 4564
rect 12679 4380 12987 4389
rect 12679 4378 12685 4380
rect 12741 4378 12765 4380
rect 12821 4378 12845 4380
rect 12901 4378 12925 4380
rect 12981 4378 12987 4380
rect 12741 4326 12743 4378
rect 12923 4326 12925 4378
rect 12679 4324 12685 4326
rect 12741 4324 12765 4326
rect 12821 4324 12845 4326
rect 12901 4324 12925 4326
rect 12981 4324 12987 4326
rect 12679 4315 12987 4324
rect 14844 4282 14872 4558
rect 14832 4276 14884 4282
rect 14832 4218 14884 4224
rect 14464 4140 14516 4146
rect 14464 4082 14516 4088
rect 12679 3292 12987 3301
rect 12679 3290 12685 3292
rect 12741 3290 12765 3292
rect 12821 3290 12845 3292
rect 12901 3290 12925 3292
rect 12981 3290 12987 3292
rect 12741 3238 12743 3290
rect 12923 3238 12925 3290
rect 12679 3236 12685 3238
rect 12741 3236 12765 3238
rect 12821 3236 12845 3238
rect 12901 3236 12925 3238
rect 12981 3236 12987 3238
rect 12679 3227 12987 3236
rect 13820 2372 13872 2378
rect 13820 2314 13872 2320
rect 12679 2204 12987 2213
rect 12679 2202 12685 2204
rect 12741 2202 12765 2204
rect 12821 2202 12845 2204
rect 12901 2202 12925 2204
rect 12981 2202 12987 2204
rect 12741 2150 12743 2202
rect 12923 2150 12925 2202
rect 12679 2148 12685 2150
rect 12741 2148 12765 2150
rect 12821 2148 12845 2150
rect 12901 2148 12925 2150
rect 12981 2148 12987 2150
rect 12679 2139 12987 2148
rect 13832 2106 13860 2314
rect 9036 2100 9088 2106
rect 9036 2042 9088 2048
rect 10416 2100 10468 2106
rect 10416 2042 10468 2048
rect 10692 2100 10744 2106
rect 10692 2042 10744 2048
rect 11520 2100 11572 2106
rect 11520 2042 11572 2048
rect 13820 2100 13872 2106
rect 13820 2042 13872 2048
rect 9048 2009 9076 2042
rect 9034 2000 9090 2009
rect 7656 1964 7708 1970
rect 7656 1906 7708 1912
rect 8852 1964 8904 1970
rect 9034 1935 9090 1944
rect 10232 1964 10284 1970
rect 8852 1906 8904 1912
rect 10232 1906 10284 1912
rect 10508 1964 10560 1970
rect 10508 1906 10560 1912
rect 11520 1964 11572 1970
rect 11520 1906 11572 1912
rect 11796 1964 11848 1970
rect 11796 1906 11848 1912
rect 12440 1964 12492 1970
rect 12440 1906 12492 1912
rect 12808 1964 12860 1970
rect 12808 1906 12860 1912
rect 13636 1964 13688 1970
rect 13636 1906 13688 1912
rect 14096 1964 14148 1970
rect 14096 1906 14148 1912
rect 3882 1660 4190 1669
rect 3882 1658 3888 1660
rect 3944 1658 3968 1660
rect 4024 1658 4048 1660
rect 4104 1658 4128 1660
rect 4184 1658 4190 1660
rect 3944 1606 3946 1658
rect 4126 1606 4128 1658
rect 3882 1604 3888 1606
rect 3944 1604 3968 1606
rect 4024 1604 4048 1606
rect 4104 1604 4128 1606
rect 4184 1604 4190 1606
rect 3882 1595 4190 1604
rect 7668 1562 7696 1906
rect 7838 1864 7894 1873
rect 7838 1799 7840 1808
rect 7892 1799 7894 1808
rect 7840 1770 7892 1776
rect 8864 1562 8892 1906
rect 9747 1660 10055 1669
rect 9747 1658 9753 1660
rect 9809 1658 9833 1660
rect 9889 1658 9913 1660
rect 9969 1658 9993 1660
rect 10049 1658 10055 1660
rect 9809 1606 9811 1658
rect 9991 1606 9993 1658
rect 9747 1604 9753 1606
rect 9809 1604 9833 1606
rect 9889 1604 9913 1606
rect 9969 1604 9993 1606
rect 10049 1604 10055 1606
rect 9747 1595 10055 1604
rect 10244 1562 10272 1906
rect 10520 1562 10548 1906
rect 11532 1562 11560 1906
rect 7656 1556 7708 1562
rect 7656 1498 7708 1504
rect 8852 1556 8904 1562
rect 8852 1498 8904 1504
rect 10232 1556 10284 1562
rect 10232 1498 10284 1504
rect 10508 1556 10560 1562
rect 10508 1498 10560 1504
rect 11520 1556 11572 1562
rect 11520 1498 11572 1504
rect 11808 1358 11836 1906
rect 12452 1358 12480 1906
rect 12820 1562 12848 1906
rect 13648 1562 13676 1906
rect 12808 1556 12860 1562
rect 12808 1498 12860 1504
rect 13636 1556 13688 1562
rect 13636 1498 13688 1504
rect 14108 1358 14136 1906
rect 14476 1358 14504 4082
rect 15612 3836 15920 3845
rect 15612 3834 15618 3836
rect 15674 3834 15698 3836
rect 15754 3834 15778 3836
rect 15834 3834 15858 3836
rect 15914 3834 15920 3836
rect 15674 3782 15676 3834
rect 15856 3782 15858 3834
rect 15612 3780 15618 3782
rect 15674 3780 15698 3782
rect 15754 3780 15778 3782
rect 15834 3780 15858 3782
rect 15914 3780 15920 3782
rect 15612 3771 15920 3780
rect 15612 2748 15920 2757
rect 15612 2746 15618 2748
rect 15674 2746 15698 2748
rect 15754 2746 15778 2748
rect 15834 2746 15858 2748
rect 15914 2746 15920 2748
rect 15674 2694 15676 2746
rect 15856 2694 15858 2746
rect 15612 2692 15618 2694
rect 15674 2692 15698 2694
rect 15754 2692 15778 2694
rect 15834 2692 15858 2694
rect 15914 2692 15920 2694
rect 15612 2683 15920 2692
rect 16224 2038 16252 7890
rect 16316 7868 16344 9846
rect 16394 9840 16450 10300
rect 16500 9846 16620 9874
rect 16500 9840 16528 9846
rect 16408 9812 16528 9840
rect 16488 8492 16540 8498
rect 16488 8434 16540 8440
rect 16500 8022 16528 8434
rect 16592 8430 16620 9846
rect 16670 9840 16726 10300
rect 16946 9840 17002 10300
rect 17052 9846 17172 9874
rect 17052 9840 17080 9846
rect 16580 8424 16632 8430
rect 16580 8366 16632 8372
rect 16488 8016 16540 8022
rect 16488 7958 16540 7964
rect 16684 7886 16712 9840
rect 16960 9812 17080 9840
rect 16948 8900 17000 8906
rect 16948 8842 17000 8848
rect 16960 8634 16988 8842
rect 16948 8628 17000 8634
rect 16948 8570 17000 8576
rect 16856 8492 16908 8498
rect 16856 8434 16908 8440
rect 16868 8090 16896 8434
rect 17144 8362 17172 9846
rect 17222 9840 17278 10300
rect 17498 9840 17554 10300
rect 17774 9840 17830 10300
rect 17868 9988 17920 9994
rect 17868 9930 17920 9936
rect 17132 8356 17184 8362
rect 17132 8298 17184 8304
rect 16856 8084 16908 8090
rect 16856 8026 16908 8032
rect 17236 7886 17264 9840
rect 17316 8832 17368 8838
rect 17316 8774 17368 8780
rect 17328 8634 17356 8774
rect 17316 8628 17368 8634
rect 17316 8570 17368 8576
rect 17512 8430 17540 9840
rect 17500 8424 17552 8430
rect 17500 8366 17552 8372
rect 17788 7886 17816 9840
rect 17880 8634 17908 9930
rect 18050 9840 18106 10300
rect 18156 9846 18276 9874
rect 18156 9840 18184 9846
rect 18064 9812 18184 9840
rect 18144 9716 18196 9722
rect 18144 9658 18196 9664
rect 17868 8628 17920 8634
rect 17868 8570 17920 8576
rect 17868 8492 17920 8498
rect 17868 8434 17920 8440
rect 17880 8362 17908 8434
rect 18156 8362 18184 9658
rect 17868 8356 17920 8362
rect 17868 8298 17920 8304
rect 18144 8356 18196 8362
rect 18144 8298 18196 8304
rect 16396 7880 16448 7886
rect 16316 7840 16396 7868
rect 16396 7822 16448 7828
rect 16672 7880 16724 7886
rect 16672 7822 16724 7828
rect 17224 7880 17276 7886
rect 17224 7822 17276 7828
rect 17776 7880 17828 7886
rect 18248 7868 18276 9846
rect 18326 9840 18382 10300
rect 18602 9840 18658 10300
rect 18878 9840 18934 10300
rect 19154 9840 19210 10300
rect 19430 9840 19486 10300
rect 19706 9840 19762 10300
rect 19982 9840 20038 10300
rect 20258 9840 20314 10300
rect 20534 9840 20590 10300
rect 20810 9840 20866 10300
rect 21086 9840 21142 10300
rect 21362 9840 21418 10300
rect 21638 9840 21694 10300
rect 21914 9840 21970 10300
rect 22190 9840 22246 10300
rect 22466 9840 22522 10300
rect 22572 9846 22692 9874
rect 22572 9840 22600 9846
rect 18340 9194 18368 9840
rect 18340 9166 18460 9194
rect 18432 8634 18460 9166
rect 18616 8838 18644 9840
rect 18892 8906 18920 9840
rect 18972 9580 19024 9586
rect 18972 9522 19024 9528
rect 18880 8900 18932 8906
rect 18880 8842 18932 8848
rect 18604 8832 18656 8838
rect 18604 8774 18656 8780
rect 18544 8732 18852 8741
rect 18544 8730 18550 8732
rect 18606 8730 18630 8732
rect 18686 8730 18710 8732
rect 18766 8730 18790 8732
rect 18846 8730 18852 8732
rect 18606 8678 18608 8730
rect 18788 8678 18790 8730
rect 18544 8676 18550 8678
rect 18606 8676 18630 8678
rect 18686 8676 18710 8678
rect 18766 8676 18790 8678
rect 18846 8676 18852 8678
rect 18544 8667 18852 8676
rect 18420 8628 18472 8634
rect 18420 8570 18472 8576
rect 18604 8492 18656 8498
rect 18604 8434 18656 8440
rect 18616 8090 18644 8434
rect 18984 8430 19012 9522
rect 18972 8424 19024 8430
rect 18972 8366 19024 8372
rect 18604 8084 18656 8090
rect 18604 8026 18656 8032
rect 18328 7880 18380 7886
rect 18248 7840 18328 7868
rect 17776 7822 17828 7828
rect 19168 7868 19196 9840
rect 19340 9104 19392 9110
rect 19340 9046 19392 9052
rect 19352 8498 19380 9046
rect 19340 8492 19392 8498
rect 19340 8434 19392 8440
rect 19340 7880 19392 7886
rect 18328 7822 18380 7828
rect 18602 7848 18658 7857
rect 19168 7840 19340 7868
rect 19444 7868 19472 9840
rect 19616 9648 19668 9654
rect 19616 9590 19668 9596
rect 19524 8832 19576 8838
rect 19524 8774 19576 8780
rect 19536 8498 19564 8774
rect 19628 8634 19656 9590
rect 19616 8628 19668 8634
rect 19616 8570 19668 8576
rect 19524 8492 19576 8498
rect 19524 8434 19576 8440
rect 19524 8288 19576 8294
rect 19524 8230 19576 8236
rect 19536 8090 19564 8230
rect 19524 8084 19576 8090
rect 19524 8026 19576 8032
rect 19524 7880 19576 7886
rect 19444 7840 19524 7868
rect 19340 7822 19392 7828
rect 19720 7868 19748 9840
rect 19800 8900 19852 8906
rect 19800 8842 19852 8848
rect 19812 8498 19840 8842
rect 19996 8634 20024 9840
rect 20272 9058 20300 9840
rect 20272 9030 20392 9058
rect 20364 8634 20392 9030
rect 19984 8628 20036 8634
rect 19984 8570 20036 8576
rect 20352 8628 20404 8634
rect 20352 8570 20404 8576
rect 19800 8492 19852 8498
rect 19800 8434 19852 8440
rect 20076 8492 20128 8498
rect 20076 8434 20128 8440
rect 19800 7880 19852 7886
rect 19720 7840 19800 7868
rect 19524 7822 19576 7828
rect 19800 7822 19852 7828
rect 18602 7783 18658 7792
rect 18616 7750 18644 7783
rect 16764 7744 16816 7750
rect 16764 7686 16816 7692
rect 17316 7744 17368 7750
rect 17316 7686 17368 7692
rect 18604 7744 18656 7750
rect 18604 7686 18656 7692
rect 19064 7744 19116 7750
rect 19064 7686 19116 7692
rect 19708 7744 19760 7750
rect 19708 7686 19760 7692
rect 19984 7744 20036 7750
rect 19984 7686 20036 7692
rect 16776 7546 16804 7686
rect 17328 7546 17356 7686
rect 18544 7644 18852 7653
rect 18544 7642 18550 7644
rect 18606 7642 18630 7644
rect 18686 7642 18710 7644
rect 18766 7642 18790 7644
rect 18846 7642 18852 7644
rect 18606 7590 18608 7642
rect 18788 7590 18790 7642
rect 18544 7588 18550 7590
rect 18606 7588 18630 7590
rect 18686 7588 18710 7590
rect 18766 7588 18790 7590
rect 18846 7588 18852 7590
rect 18544 7579 18852 7588
rect 16764 7540 16816 7546
rect 16764 7482 16816 7488
rect 17316 7540 17368 7546
rect 17316 7482 17368 7488
rect 17408 7404 17460 7410
rect 17408 7346 17460 7352
rect 17420 7002 17448 7346
rect 19076 7002 19104 7686
rect 19720 7313 19748 7686
rect 19996 7449 20024 7686
rect 19982 7440 20038 7449
rect 19982 7375 20038 7384
rect 19706 7304 19762 7313
rect 19706 7239 19762 7248
rect 17408 6996 17460 7002
rect 17408 6938 17460 6944
rect 19064 6996 19116 7002
rect 19064 6938 19116 6944
rect 16856 6792 16908 6798
rect 16856 6734 16908 6740
rect 16868 2774 16896 6734
rect 18544 6556 18852 6565
rect 18544 6554 18550 6556
rect 18606 6554 18630 6556
rect 18686 6554 18710 6556
rect 18766 6554 18790 6556
rect 18846 6554 18852 6556
rect 18606 6502 18608 6554
rect 18788 6502 18790 6554
rect 18544 6500 18550 6502
rect 18606 6500 18630 6502
rect 18686 6500 18710 6502
rect 18766 6500 18790 6502
rect 18846 6500 18852 6502
rect 18544 6491 18852 6500
rect 18544 5468 18852 5477
rect 18544 5466 18550 5468
rect 18606 5466 18630 5468
rect 18686 5466 18710 5468
rect 18766 5466 18790 5468
rect 18846 5466 18852 5468
rect 18606 5414 18608 5466
rect 18788 5414 18790 5466
rect 18544 5412 18550 5414
rect 18606 5412 18630 5414
rect 18686 5412 18710 5414
rect 18766 5412 18790 5414
rect 18846 5412 18852 5414
rect 18544 5403 18852 5412
rect 18544 4380 18852 4389
rect 18544 4378 18550 4380
rect 18606 4378 18630 4380
rect 18686 4378 18710 4380
rect 18766 4378 18790 4380
rect 18846 4378 18852 4380
rect 18606 4326 18608 4378
rect 18788 4326 18790 4378
rect 18544 4324 18550 4326
rect 18606 4324 18630 4326
rect 18686 4324 18710 4326
rect 18766 4324 18790 4326
rect 18846 4324 18852 4326
rect 18544 4315 18852 4324
rect 17776 3528 17828 3534
rect 17776 3470 17828 3476
rect 16776 2746 16896 2774
rect 16212 2032 16264 2038
rect 16212 1974 16264 1980
rect 16120 1964 16172 1970
rect 16120 1906 16172 1912
rect 16304 1964 16356 1970
rect 16304 1906 16356 1912
rect 15612 1660 15920 1669
rect 15612 1658 15618 1660
rect 15674 1658 15698 1660
rect 15754 1658 15778 1660
rect 15834 1658 15858 1660
rect 15914 1658 15920 1660
rect 15674 1606 15676 1658
rect 15856 1606 15858 1658
rect 15612 1604 15618 1606
rect 15674 1604 15698 1606
rect 15754 1604 15778 1606
rect 15834 1604 15858 1606
rect 15914 1604 15920 1606
rect 15612 1595 15920 1604
rect 16132 1562 16160 1906
rect 16316 1766 16344 1906
rect 16304 1760 16356 1766
rect 16304 1702 16356 1708
rect 16120 1556 16172 1562
rect 16120 1498 16172 1504
rect 848 1352 900 1358
rect 848 1294 900 1300
rect 2136 1352 2188 1358
rect 2136 1294 2188 1300
rect 3332 1352 3384 1358
rect 3332 1294 3384 1300
rect 4712 1352 4764 1358
rect 4712 1294 4764 1300
rect 5908 1352 5960 1358
rect 5908 1294 5960 1300
rect 7564 1352 7616 1358
rect 8760 1352 8812 1358
rect 7564 1294 7616 1300
rect 8496 1312 8760 1340
rect 860 160 888 1294
rect 1584 1216 1636 1222
rect 1584 1158 1636 1164
rect 1596 1018 1624 1158
rect 1584 1012 1636 1018
rect 1584 954 1636 960
rect 846 -300 902 160
rect 2042 82 2098 160
rect 2148 82 2176 1294
rect 2320 1216 2372 1222
rect 2320 1158 2372 1164
rect 2332 814 2360 1158
rect 2320 808 2372 814
rect 2320 750 2372 756
rect 2042 54 2176 82
rect 3238 82 3294 160
rect 3344 82 3372 1294
rect 4528 1216 4580 1222
rect 4528 1158 4580 1164
rect 4540 1018 4568 1158
rect 4528 1012 4580 1018
rect 4528 954 4580 960
rect 3238 54 3372 82
rect 4434 82 4490 160
rect 4724 82 4752 1294
rect 5724 1216 5776 1222
rect 5724 1158 5776 1164
rect 5736 1018 5764 1158
rect 5724 1012 5776 1018
rect 5724 954 5776 960
rect 4434 54 4752 82
rect 5630 82 5686 160
rect 5920 82 5948 1294
rect 7288 1216 7340 1222
rect 7288 1158 7340 1164
rect 6814 1116 7122 1125
rect 6814 1114 6820 1116
rect 6876 1114 6900 1116
rect 6956 1114 6980 1116
rect 7036 1114 7060 1116
rect 7116 1114 7122 1116
rect 6876 1062 6878 1114
rect 7058 1062 7060 1114
rect 6814 1060 6820 1062
rect 6876 1060 6900 1062
rect 6956 1060 6980 1062
rect 7036 1060 7060 1062
rect 7116 1060 7122 1062
rect 6814 1051 7122 1060
rect 7300 950 7328 1158
rect 7288 944 7340 950
rect 7288 886 7340 892
rect 7576 610 7604 1294
rect 6920 604 6972 610
rect 6920 546 6972 552
rect 7564 604 7616 610
rect 7564 546 7616 552
rect 5630 54 5948 82
rect 6826 82 6882 160
rect 6932 82 6960 546
rect 6826 54 6960 82
rect 8022 82 8078 160
rect 8496 82 8524 1312
rect 8760 1294 8812 1300
rect 9496 1352 9548 1358
rect 9496 1294 9548 1300
rect 9864 1352 9916 1358
rect 9864 1294 9916 1300
rect 10692 1352 10744 1358
rect 10692 1294 10744 1300
rect 11244 1352 11296 1358
rect 11244 1294 11296 1300
rect 11796 1352 11848 1358
rect 11796 1294 11848 1300
rect 11888 1352 11940 1358
rect 11888 1294 11940 1300
rect 12440 1352 12492 1358
rect 12440 1294 12492 1300
rect 12532 1352 12584 1358
rect 12532 1294 12584 1300
rect 12992 1352 13044 1358
rect 13728 1352 13780 1358
rect 13044 1312 13124 1340
rect 12992 1294 13044 1300
rect 8022 54 8524 82
rect 9218 82 9274 160
rect 9508 82 9536 1294
rect 9876 1018 9904 1294
rect 9864 1012 9916 1018
rect 9864 954 9916 960
rect 9218 54 9536 82
rect 10414 82 10470 160
rect 10704 82 10732 1294
rect 11256 678 11284 1294
rect 11244 672 11296 678
rect 11244 614 11296 620
rect 10414 54 10732 82
rect 11610 82 11666 160
rect 11900 82 11928 1294
rect 12544 882 12572 1294
rect 12679 1116 12987 1125
rect 12679 1114 12685 1116
rect 12741 1114 12765 1116
rect 12821 1114 12845 1116
rect 12901 1114 12925 1116
rect 12981 1114 12987 1116
rect 12741 1062 12743 1114
rect 12923 1062 12925 1114
rect 12679 1060 12685 1062
rect 12741 1060 12765 1062
rect 12821 1060 12845 1062
rect 12901 1060 12925 1062
rect 12981 1060 12987 1062
rect 12679 1051 12987 1060
rect 12532 876 12584 882
rect 12532 818 12584 824
rect 12820 190 12940 218
rect 12820 160 12848 190
rect 11610 54 11928 82
rect 2042 -300 2098 54
rect 3238 -300 3294 54
rect 4434 -300 4490 54
rect 5630 -300 5686 54
rect 6826 -300 6882 54
rect 8022 -300 8078 54
rect 9218 -300 9274 54
rect 10414 -300 10470 54
rect 11610 -300 11666 54
rect 12806 -300 12862 160
rect 12912 82 12940 190
rect 13096 82 13124 1312
rect 13728 1294 13780 1300
rect 14096 1352 14148 1358
rect 14096 1294 14148 1300
rect 14280 1352 14332 1358
rect 14280 1294 14332 1300
rect 14372 1352 14424 1358
rect 14372 1294 14424 1300
rect 14464 1352 14516 1358
rect 14464 1294 14516 1300
rect 15476 1352 15528 1358
rect 16672 1352 16724 1358
rect 15476 1294 15528 1300
rect 16500 1312 16672 1340
rect 13740 1018 13768 1294
rect 13728 1012 13780 1018
rect 13728 954 13780 960
rect 12912 54 13124 82
rect 14002 82 14058 160
rect 14292 82 14320 1294
rect 14384 1018 14412 1294
rect 14556 1216 14608 1222
rect 14556 1158 14608 1164
rect 14568 1018 14596 1158
rect 14372 1012 14424 1018
rect 14372 954 14424 960
rect 14556 1012 14608 1018
rect 14556 954 14608 960
rect 14002 54 14320 82
rect 15198 82 15254 160
rect 15488 82 15516 1294
rect 15198 54 15516 82
rect 16394 82 16450 160
rect 16500 82 16528 1312
rect 16672 1294 16724 1300
rect 16776 1290 16804 2746
rect 17788 1290 17816 3470
rect 18544 3292 18852 3301
rect 18544 3290 18550 3292
rect 18606 3290 18630 3292
rect 18686 3290 18710 3292
rect 18766 3290 18790 3292
rect 18846 3290 18852 3292
rect 18606 3238 18608 3290
rect 18788 3238 18790 3290
rect 18544 3236 18550 3238
rect 18606 3236 18630 3238
rect 18686 3236 18710 3238
rect 18766 3236 18790 3238
rect 18846 3236 18852 3238
rect 18544 3227 18852 3236
rect 20088 2774 20116 8434
rect 20548 8362 20576 9840
rect 20720 8492 20772 8498
rect 20720 8434 20772 8440
rect 20536 8356 20588 8362
rect 20536 8298 20588 8304
rect 19904 2746 20116 2774
rect 18544 2204 18852 2213
rect 18544 2202 18550 2204
rect 18606 2202 18630 2204
rect 18686 2202 18710 2204
rect 18766 2202 18790 2204
rect 18846 2202 18852 2204
rect 18606 2150 18608 2202
rect 18788 2150 18790 2202
rect 18544 2148 18550 2150
rect 18606 2148 18630 2150
rect 18686 2148 18710 2150
rect 18766 2148 18790 2150
rect 18846 2148 18852 2150
rect 18544 2139 18852 2148
rect 17868 1352 17920 1358
rect 17868 1294 17920 1300
rect 19064 1352 19116 1358
rect 19064 1294 19116 1300
rect 16764 1284 16816 1290
rect 16764 1226 16816 1232
rect 17776 1284 17828 1290
rect 17776 1226 17828 1232
rect 16394 54 16528 82
rect 17590 82 17646 160
rect 17880 82 17908 1294
rect 18544 1116 18852 1125
rect 18544 1114 18550 1116
rect 18606 1114 18630 1116
rect 18686 1114 18710 1116
rect 18766 1114 18790 1116
rect 18846 1114 18852 1116
rect 18606 1062 18608 1114
rect 18788 1062 18790 1114
rect 18544 1060 18550 1062
rect 18606 1060 18630 1062
rect 18686 1060 18710 1062
rect 18766 1060 18790 1062
rect 18846 1060 18852 1062
rect 18544 1051 18852 1060
rect 17590 54 17908 82
rect 18786 82 18842 160
rect 19076 82 19104 1294
rect 19904 1018 19932 2746
rect 20732 2106 20760 8434
rect 20824 8090 20852 9840
rect 21100 8634 21128 9840
rect 21088 8628 21140 8634
rect 21088 8570 21140 8576
rect 21376 8566 21404 9840
rect 21364 8560 21416 8566
rect 21364 8502 21416 8508
rect 21180 8492 21232 8498
rect 21180 8434 21232 8440
rect 20812 8084 20864 8090
rect 20812 8026 20864 8032
rect 21192 2310 21220 8434
rect 21652 8362 21680 9840
rect 21640 8356 21692 8362
rect 21640 8298 21692 8304
rect 21477 8188 21785 8197
rect 21477 8186 21483 8188
rect 21539 8186 21563 8188
rect 21619 8186 21643 8188
rect 21699 8186 21723 8188
rect 21779 8186 21785 8188
rect 21539 8134 21541 8186
rect 21721 8134 21723 8186
rect 21477 8132 21483 8134
rect 21539 8132 21563 8134
rect 21619 8132 21643 8134
rect 21699 8132 21723 8134
rect 21779 8132 21785 8134
rect 21477 8123 21785 8132
rect 21928 8090 21956 9840
rect 21916 8084 21968 8090
rect 22204 8072 22232 9840
rect 22480 9812 22600 9840
rect 22468 8492 22520 8498
rect 22468 8434 22520 8440
rect 22480 8401 22508 8434
rect 22466 8392 22522 8401
rect 22466 8327 22522 8336
rect 22284 8084 22336 8090
rect 22204 8044 22284 8072
rect 21916 8026 21968 8032
rect 22664 8072 22692 9846
rect 22742 9840 22798 10300
rect 22848 9846 22968 9874
rect 22848 9840 22876 9846
rect 22756 9812 22876 9840
rect 22836 8084 22888 8090
rect 22664 8044 22836 8072
rect 22284 8026 22336 8032
rect 22836 8026 22888 8032
rect 22940 8004 22968 9846
rect 23018 9840 23074 10300
rect 23124 9846 23244 9874
rect 23124 9840 23152 9846
rect 23032 9812 23152 9840
rect 23216 8634 23244 9846
rect 23294 9840 23350 10300
rect 23570 9840 23626 10300
rect 23676 9846 23796 9874
rect 23676 9840 23704 9846
rect 23204 8628 23256 8634
rect 23204 8570 23256 8576
rect 23020 8492 23072 8498
rect 23020 8434 23072 8440
rect 23032 8401 23060 8434
rect 23018 8392 23074 8401
rect 23018 8327 23074 8336
rect 23204 8016 23256 8022
rect 22940 7976 23204 8004
rect 23204 7958 23256 7964
rect 22100 7812 22152 7818
rect 22100 7754 22152 7760
rect 22652 7812 22704 7818
rect 22652 7754 22704 7760
rect 22744 7812 22796 7818
rect 22744 7754 22796 7760
rect 22112 7313 22140 7754
rect 22468 7404 22520 7410
rect 22468 7346 22520 7352
rect 22098 7304 22154 7313
rect 22098 7239 22154 7248
rect 22100 7200 22152 7206
rect 22100 7142 22152 7148
rect 21477 7100 21785 7109
rect 21477 7098 21483 7100
rect 21539 7098 21563 7100
rect 21619 7098 21643 7100
rect 21699 7098 21723 7100
rect 21779 7098 21785 7100
rect 21539 7046 21541 7098
rect 21721 7046 21723 7098
rect 21477 7044 21483 7046
rect 21539 7044 21563 7046
rect 21619 7044 21643 7046
rect 21699 7044 21723 7046
rect 21779 7044 21785 7046
rect 21477 7035 21785 7044
rect 22112 6390 22140 7142
rect 22100 6384 22152 6390
rect 22100 6326 22152 6332
rect 21477 6012 21785 6021
rect 21477 6010 21483 6012
rect 21539 6010 21563 6012
rect 21619 6010 21643 6012
rect 21699 6010 21723 6012
rect 21779 6010 21785 6012
rect 21539 5958 21541 6010
rect 21721 5958 21723 6010
rect 21477 5956 21483 5958
rect 21539 5956 21563 5958
rect 21619 5956 21643 5958
rect 21699 5956 21723 5958
rect 21779 5956 21785 5958
rect 21477 5947 21785 5956
rect 21477 4924 21785 4933
rect 21477 4922 21483 4924
rect 21539 4922 21563 4924
rect 21619 4922 21643 4924
rect 21699 4922 21723 4924
rect 21779 4922 21785 4924
rect 21539 4870 21541 4922
rect 21721 4870 21723 4922
rect 21477 4868 21483 4870
rect 21539 4868 21563 4870
rect 21619 4868 21643 4870
rect 21699 4868 21723 4870
rect 21779 4868 21785 4870
rect 21477 4859 21785 4868
rect 21477 3836 21785 3845
rect 21477 3834 21483 3836
rect 21539 3834 21563 3836
rect 21619 3834 21643 3836
rect 21699 3834 21723 3836
rect 21779 3834 21785 3836
rect 21539 3782 21541 3834
rect 21721 3782 21723 3834
rect 21477 3780 21483 3782
rect 21539 3780 21563 3782
rect 21619 3780 21643 3782
rect 21699 3780 21723 3782
rect 21779 3780 21785 3782
rect 21477 3771 21785 3780
rect 22480 3194 22508 7346
rect 22468 3188 22520 3194
rect 22468 3130 22520 3136
rect 22468 3052 22520 3058
rect 22468 2994 22520 3000
rect 21477 2748 21785 2757
rect 21477 2746 21483 2748
rect 21539 2746 21563 2748
rect 21619 2746 21643 2748
rect 21699 2746 21723 2748
rect 21779 2746 21785 2748
rect 21539 2694 21541 2746
rect 21721 2694 21723 2746
rect 21477 2692 21483 2694
rect 21539 2692 21563 2694
rect 21619 2692 21643 2694
rect 21699 2692 21723 2694
rect 21779 2692 21785 2694
rect 21477 2683 21785 2692
rect 21180 2304 21232 2310
rect 21180 2246 21232 2252
rect 20720 2100 20772 2106
rect 20720 2042 20772 2048
rect 22192 1964 22244 1970
rect 22192 1906 22244 1912
rect 21477 1660 21785 1669
rect 21477 1658 21483 1660
rect 21539 1658 21563 1660
rect 21619 1658 21643 1660
rect 21699 1658 21723 1660
rect 21779 1658 21785 1660
rect 21539 1606 21541 1658
rect 21721 1606 21723 1658
rect 21477 1604 21483 1606
rect 21539 1604 21563 1606
rect 21619 1604 21643 1606
rect 21699 1604 21723 1606
rect 21779 1604 21785 1606
rect 21477 1595 21785 1604
rect 22204 1562 22232 1906
rect 22192 1556 22244 1562
rect 22192 1498 22244 1504
rect 20260 1352 20312 1358
rect 20260 1294 20312 1300
rect 21456 1352 21508 1358
rect 21456 1294 21508 1300
rect 19984 1216 20036 1222
rect 19984 1158 20036 1164
rect 19996 1018 20024 1158
rect 19892 1012 19944 1018
rect 19892 954 19944 960
rect 19984 1012 20036 1018
rect 19984 954 20036 960
rect 18786 54 19104 82
rect 19982 82 20038 160
rect 20272 82 20300 1294
rect 19982 54 20300 82
rect 21178 82 21234 160
rect 21468 82 21496 1294
rect 22480 1222 22508 2994
rect 22664 1834 22692 7754
rect 22756 1902 22784 7754
rect 22836 7744 22888 7750
rect 22836 7686 22888 7692
rect 22848 3126 22876 7686
rect 23020 7404 23072 7410
rect 23020 7346 23072 7352
rect 22836 3120 22888 3126
rect 22836 3062 22888 3068
rect 23032 2106 23060 7346
rect 23112 6724 23164 6730
rect 23112 6666 23164 6672
rect 23124 3738 23152 6666
rect 23308 6458 23336 9840
rect 23584 9812 23704 9840
rect 23572 8492 23624 8498
rect 23492 8452 23572 8480
rect 23388 6724 23440 6730
rect 23388 6666 23440 6672
rect 23296 6452 23348 6458
rect 23296 6394 23348 6400
rect 23204 6316 23256 6322
rect 23204 6258 23256 6264
rect 23112 3732 23164 3738
rect 23112 3674 23164 3680
rect 23216 2106 23244 6258
rect 23296 2440 23348 2446
rect 23296 2382 23348 2388
rect 23020 2100 23072 2106
rect 23020 2042 23072 2048
rect 23204 2100 23256 2106
rect 23204 2042 23256 2048
rect 22836 1964 22888 1970
rect 22836 1906 22888 1912
rect 22744 1896 22796 1902
rect 22744 1838 22796 1844
rect 22652 1828 22704 1834
rect 22652 1770 22704 1776
rect 22848 1562 22876 1906
rect 23112 1896 23164 1902
rect 23112 1838 23164 1844
rect 23124 1562 23152 1838
rect 23308 1562 23336 2382
rect 23400 2106 23428 6666
rect 23492 4486 23520 8452
rect 23572 8434 23624 8440
rect 23768 8242 23796 9846
rect 23846 9840 23902 10300
rect 24122 9840 24178 10300
rect 24398 9840 24454 10300
rect 24674 9840 24730 10300
rect 24950 9840 25006 10300
rect 25226 9840 25282 10300
rect 25502 9840 25558 10300
rect 23860 8378 23888 9840
rect 23860 8350 23980 8378
rect 23768 8214 23888 8242
rect 23756 7812 23808 7818
rect 23756 7754 23808 7760
rect 23572 7404 23624 7410
rect 23572 7346 23624 7352
rect 23480 4480 23532 4486
rect 23480 4422 23532 4428
rect 23584 2106 23612 7346
rect 23768 2378 23796 7754
rect 23860 6458 23888 8214
rect 23952 6730 23980 8350
rect 24136 7546 24164 9840
rect 24412 8922 24440 9840
rect 24320 8894 24440 8922
rect 24688 8922 24716 9840
rect 24688 8894 24808 8922
rect 24124 7540 24176 7546
rect 24124 7482 24176 7488
rect 24320 6866 24348 8894
rect 24409 8732 24717 8741
rect 24409 8730 24415 8732
rect 24471 8730 24495 8732
rect 24551 8730 24575 8732
rect 24631 8730 24655 8732
rect 24711 8730 24717 8732
rect 24471 8678 24473 8730
rect 24653 8678 24655 8730
rect 24409 8676 24415 8678
rect 24471 8676 24495 8678
rect 24551 8676 24575 8678
rect 24631 8676 24655 8678
rect 24711 8676 24717 8678
rect 24409 8667 24717 8676
rect 24409 7644 24717 7653
rect 24409 7642 24415 7644
rect 24471 7642 24495 7644
rect 24551 7642 24575 7644
rect 24631 7642 24655 7644
rect 24711 7642 24717 7644
rect 24471 7590 24473 7642
rect 24653 7590 24655 7642
rect 24409 7588 24415 7590
rect 24471 7588 24495 7590
rect 24551 7588 24575 7590
rect 24631 7588 24655 7590
rect 24711 7588 24717 7590
rect 24409 7579 24717 7588
rect 24780 7546 24808 8894
rect 24768 7540 24820 7546
rect 24768 7482 24820 7488
rect 24964 7342 24992 9840
rect 24952 7336 25004 7342
rect 24952 7278 25004 7284
rect 24308 6860 24360 6866
rect 24308 6802 24360 6808
rect 23940 6724 23992 6730
rect 23940 6666 23992 6672
rect 24409 6556 24717 6565
rect 24409 6554 24415 6556
rect 24471 6554 24495 6556
rect 24551 6554 24575 6556
rect 24631 6554 24655 6556
rect 24711 6554 24717 6556
rect 24471 6502 24473 6554
rect 24653 6502 24655 6554
rect 24409 6500 24415 6502
rect 24471 6500 24495 6502
rect 24551 6500 24575 6502
rect 24631 6500 24655 6502
rect 24711 6500 24717 6502
rect 24409 6491 24717 6500
rect 23848 6452 23900 6458
rect 23848 6394 23900 6400
rect 25240 5914 25268 9840
rect 25516 7886 25544 9840
rect 25504 7880 25556 7886
rect 25504 7822 25556 7828
rect 25228 5908 25280 5914
rect 25228 5850 25280 5856
rect 23848 5636 23900 5642
rect 23848 5578 23900 5584
rect 23756 2372 23808 2378
rect 23756 2314 23808 2320
rect 23860 2106 23888 5578
rect 24409 5468 24717 5477
rect 24409 5466 24415 5468
rect 24471 5466 24495 5468
rect 24551 5466 24575 5468
rect 24631 5466 24655 5468
rect 24711 5466 24717 5468
rect 24471 5414 24473 5466
rect 24653 5414 24655 5466
rect 24409 5412 24415 5414
rect 24471 5412 24495 5414
rect 24551 5412 24575 5414
rect 24631 5412 24655 5414
rect 24711 5412 24717 5414
rect 24409 5403 24717 5412
rect 24409 4380 24717 4389
rect 24409 4378 24415 4380
rect 24471 4378 24495 4380
rect 24551 4378 24575 4380
rect 24631 4378 24655 4380
rect 24711 4378 24717 4380
rect 24471 4326 24473 4378
rect 24653 4326 24655 4378
rect 24409 4324 24415 4326
rect 24471 4324 24495 4326
rect 24551 4324 24575 4326
rect 24631 4324 24655 4326
rect 24711 4324 24717 4326
rect 24409 4315 24717 4324
rect 24409 3292 24717 3301
rect 24409 3290 24415 3292
rect 24471 3290 24495 3292
rect 24551 3290 24575 3292
rect 24631 3290 24655 3292
rect 24711 3290 24717 3292
rect 24471 3238 24473 3290
rect 24653 3238 24655 3290
rect 24409 3236 24415 3238
rect 24471 3236 24495 3238
rect 24551 3236 24575 3238
rect 24631 3236 24655 3238
rect 24711 3236 24717 3238
rect 24409 3227 24717 3236
rect 24032 3052 24084 3058
rect 24032 2994 24084 3000
rect 24044 2650 24072 2994
rect 24032 2644 24084 2650
rect 24032 2586 24084 2592
rect 24409 2204 24717 2213
rect 24409 2202 24415 2204
rect 24471 2202 24495 2204
rect 24551 2202 24575 2204
rect 24631 2202 24655 2204
rect 24711 2202 24717 2204
rect 24471 2150 24473 2202
rect 24653 2150 24655 2202
rect 24409 2148 24415 2150
rect 24471 2148 24495 2150
rect 24551 2148 24575 2150
rect 24631 2148 24655 2150
rect 24711 2148 24717 2150
rect 24409 2139 24717 2148
rect 23388 2100 23440 2106
rect 23388 2042 23440 2048
rect 23572 2100 23624 2106
rect 23572 2042 23624 2048
rect 23848 2100 23900 2106
rect 23848 2042 23900 2048
rect 24124 1964 24176 1970
rect 24124 1906 24176 1912
rect 24136 1562 24164 1906
rect 22836 1556 22888 1562
rect 22836 1498 22888 1504
rect 23112 1556 23164 1562
rect 23112 1498 23164 1504
rect 23296 1556 23348 1562
rect 23296 1498 23348 1504
rect 24124 1556 24176 1562
rect 24124 1498 24176 1504
rect 22652 1352 22704 1358
rect 22652 1294 22704 1300
rect 23572 1352 23624 1358
rect 24124 1352 24176 1358
rect 23572 1294 23624 1300
rect 23952 1312 24124 1340
rect 22468 1216 22520 1222
rect 22468 1158 22520 1164
rect 22560 1216 22612 1222
rect 22560 1158 22612 1164
rect 22572 1018 22600 1158
rect 22560 1012 22612 1018
rect 22560 954 22612 960
rect 21178 54 21496 82
rect 22374 82 22430 160
rect 22664 82 22692 1294
rect 23584 746 23612 1294
rect 23572 740 23624 746
rect 23572 682 23624 688
rect 23584 190 23704 218
rect 23584 160 23612 190
rect 22374 54 22692 82
rect 14002 -300 14058 54
rect 15198 -300 15254 54
rect 16394 -300 16450 54
rect 17590 -300 17646 54
rect 18786 -300 18842 54
rect 19982 -300 20038 54
rect 21178 -300 21234 54
rect 22374 -300 22430 54
rect 23570 -300 23626 160
rect 23676 82 23704 190
rect 23952 82 23980 1312
rect 24124 1294 24176 1300
rect 24409 1116 24717 1125
rect 24409 1114 24415 1116
rect 24471 1114 24495 1116
rect 24551 1114 24575 1116
rect 24631 1114 24655 1116
rect 24711 1114 24717 1116
rect 24471 1062 24473 1114
rect 24653 1062 24655 1114
rect 24409 1060 24415 1062
rect 24471 1060 24495 1062
rect 24551 1060 24575 1062
rect 24631 1060 24655 1062
rect 24711 1060 24717 1062
rect 24409 1051 24717 1060
rect 24768 740 24820 746
rect 24768 682 24820 688
rect 24780 160 24808 682
rect 23676 54 23980 82
rect 24766 -300 24822 160
<< via2 >>
rect 2594 7828 2596 7848
rect 2596 7828 2648 7848
rect 2648 7828 2650 7848
rect 2594 7792 2650 7828
rect 3888 8186 3944 8188
rect 3968 8186 4024 8188
rect 4048 8186 4104 8188
rect 4128 8186 4184 8188
rect 3888 8134 3934 8186
rect 3934 8134 3944 8186
rect 3968 8134 3998 8186
rect 3998 8134 4010 8186
rect 4010 8134 4024 8186
rect 4048 8134 4062 8186
rect 4062 8134 4074 8186
rect 4074 8134 4104 8186
rect 4128 8134 4138 8186
rect 4138 8134 4184 8186
rect 3888 8132 3944 8134
rect 3968 8132 4024 8134
rect 4048 8132 4104 8134
rect 4128 8132 4184 8134
rect 3888 7098 3944 7100
rect 3968 7098 4024 7100
rect 4048 7098 4104 7100
rect 4128 7098 4184 7100
rect 3888 7046 3934 7098
rect 3934 7046 3944 7098
rect 3968 7046 3998 7098
rect 3998 7046 4010 7098
rect 4010 7046 4024 7098
rect 4048 7046 4062 7098
rect 4062 7046 4074 7098
rect 4074 7046 4104 7098
rect 4128 7046 4138 7098
rect 4138 7046 4184 7098
rect 3888 7044 3944 7046
rect 3968 7044 4024 7046
rect 4048 7044 4104 7046
rect 4128 7044 4184 7046
rect 2686 6724 2742 6760
rect 2686 6704 2688 6724
rect 2688 6704 2740 6724
rect 2740 6704 2742 6724
rect 5630 7404 5686 7440
rect 5630 7384 5632 7404
rect 5632 7384 5684 7404
rect 5684 7384 5686 7404
rect 6820 8730 6876 8732
rect 6900 8730 6956 8732
rect 6980 8730 7036 8732
rect 7060 8730 7116 8732
rect 6820 8678 6866 8730
rect 6866 8678 6876 8730
rect 6900 8678 6930 8730
rect 6930 8678 6942 8730
rect 6942 8678 6956 8730
rect 6980 8678 6994 8730
rect 6994 8678 7006 8730
rect 7006 8678 7036 8730
rect 7060 8678 7070 8730
rect 7070 8678 7116 8730
rect 6820 8676 6876 8678
rect 6900 8676 6956 8678
rect 6980 8676 7036 8678
rect 7060 8676 7116 8678
rect 6734 7812 6790 7848
rect 6734 7792 6736 7812
rect 6736 7792 6788 7812
rect 6788 7792 6790 7812
rect 6182 7248 6238 7304
rect 6820 7642 6876 7644
rect 6900 7642 6956 7644
rect 6980 7642 7036 7644
rect 7060 7642 7116 7644
rect 6820 7590 6866 7642
rect 6866 7590 6876 7642
rect 6900 7590 6930 7642
rect 6930 7590 6942 7642
rect 6942 7590 6956 7642
rect 6980 7590 6994 7642
rect 6994 7590 7006 7642
rect 7006 7590 7036 7642
rect 7060 7590 7070 7642
rect 7070 7590 7116 7642
rect 6820 7588 6876 7590
rect 6900 7588 6956 7590
rect 6980 7588 7036 7590
rect 7060 7588 7116 7590
rect 10230 8472 10286 8528
rect 9753 8186 9809 8188
rect 9833 8186 9889 8188
rect 9913 8186 9969 8188
rect 9993 8186 10049 8188
rect 9753 8134 9799 8186
rect 9799 8134 9809 8186
rect 9833 8134 9863 8186
rect 9863 8134 9875 8186
rect 9875 8134 9889 8186
rect 9913 8134 9927 8186
rect 9927 8134 9939 8186
rect 9939 8134 9969 8186
rect 9993 8134 10003 8186
rect 10003 8134 10049 8186
rect 9753 8132 9809 8134
rect 9833 8132 9889 8134
rect 9913 8132 9969 8134
rect 9993 8132 10049 8134
rect 9753 7098 9809 7100
rect 9833 7098 9889 7100
rect 9913 7098 9969 7100
rect 9993 7098 10049 7100
rect 9753 7046 9799 7098
rect 9799 7046 9809 7098
rect 9833 7046 9863 7098
rect 9863 7046 9875 7098
rect 9875 7046 9889 7098
rect 9913 7046 9927 7098
rect 9927 7046 9939 7098
rect 9939 7046 9969 7098
rect 9993 7046 10003 7098
rect 10003 7046 10049 7098
rect 9753 7044 9809 7046
rect 9833 7044 9889 7046
rect 9913 7044 9969 7046
rect 9993 7044 10049 7046
rect 6820 6554 6876 6556
rect 6900 6554 6956 6556
rect 6980 6554 7036 6556
rect 7060 6554 7116 6556
rect 6820 6502 6866 6554
rect 6866 6502 6876 6554
rect 6900 6502 6930 6554
rect 6930 6502 6942 6554
rect 6942 6502 6956 6554
rect 6980 6502 6994 6554
rect 6994 6502 7006 6554
rect 7006 6502 7036 6554
rect 7060 6502 7070 6554
rect 7070 6502 7116 6554
rect 6820 6500 6876 6502
rect 6900 6500 6956 6502
rect 6980 6500 7036 6502
rect 7060 6500 7116 6502
rect 3888 6010 3944 6012
rect 3968 6010 4024 6012
rect 4048 6010 4104 6012
rect 4128 6010 4184 6012
rect 3888 5958 3934 6010
rect 3934 5958 3944 6010
rect 3968 5958 3998 6010
rect 3998 5958 4010 6010
rect 4010 5958 4024 6010
rect 4048 5958 4062 6010
rect 4062 5958 4074 6010
rect 4074 5958 4104 6010
rect 4128 5958 4138 6010
rect 4138 5958 4184 6010
rect 3888 5956 3944 5958
rect 3968 5956 4024 5958
rect 4048 5956 4104 5958
rect 4128 5956 4184 5958
rect 9753 6010 9809 6012
rect 9833 6010 9889 6012
rect 9913 6010 9969 6012
rect 9993 6010 10049 6012
rect 9753 5958 9799 6010
rect 9799 5958 9809 6010
rect 9833 5958 9863 6010
rect 9863 5958 9875 6010
rect 9875 5958 9889 6010
rect 9913 5958 9927 6010
rect 9927 5958 9939 6010
rect 9939 5958 9969 6010
rect 9993 5958 10003 6010
rect 10003 5958 10049 6010
rect 9753 5956 9809 5958
rect 9833 5956 9889 5958
rect 9913 5956 9969 5958
rect 9993 5956 10049 5958
rect 6820 5466 6876 5468
rect 6900 5466 6956 5468
rect 6980 5466 7036 5468
rect 7060 5466 7116 5468
rect 6820 5414 6866 5466
rect 6866 5414 6876 5466
rect 6900 5414 6930 5466
rect 6930 5414 6942 5466
rect 6942 5414 6956 5466
rect 6980 5414 6994 5466
rect 6994 5414 7006 5466
rect 7006 5414 7036 5466
rect 7060 5414 7070 5466
rect 7070 5414 7116 5466
rect 6820 5412 6876 5414
rect 6900 5412 6956 5414
rect 6980 5412 7036 5414
rect 7060 5412 7116 5414
rect 3888 4922 3944 4924
rect 3968 4922 4024 4924
rect 4048 4922 4104 4924
rect 4128 4922 4184 4924
rect 3888 4870 3934 4922
rect 3934 4870 3944 4922
rect 3968 4870 3998 4922
rect 3998 4870 4010 4922
rect 4010 4870 4024 4922
rect 4048 4870 4062 4922
rect 4062 4870 4074 4922
rect 4074 4870 4104 4922
rect 4128 4870 4138 4922
rect 4138 4870 4184 4922
rect 3888 4868 3944 4870
rect 3968 4868 4024 4870
rect 4048 4868 4104 4870
rect 4128 4868 4184 4870
rect 9753 4922 9809 4924
rect 9833 4922 9889 4924
rect 9913 4922 9969 4924
rect 9993 4922 10049 4924
rect 9753 4870 9799 4922
rect 9799 4870 9809 4922
rect 9833 4870 9863 4922
rect 9863 4870 9875 4922
rect 9875 4870 9889 4922
rect 9913 4870 9927 4922
rect 9927 4870 9939 4922
rect 9939 4870 9969 4922
rect 9993 4870 10003 4922
rect 10003 4870 10049 4922
rect 9753 4868 9809 4870
rect 9833 4868 9889 4870
rect 9913 4868 9969 4870
rect 9993 4868 10049 4870
rect 6820 4378 6876 4380
rect 6900 4378 6956 4380
rect 6980 4378 7036 4380
rect 7060 4378 7116 4380
rect 6820 4326 6866 4378
rect 6866 4326 6876 4378
rect 6900 4326 6930 4378
rect 6930 4326 6942 4378
rect 6942 4326 6956 4378
rect 6980 4326 6994 4378
rect 6994 4326 7006 4378
rect 7006 4326 7036 4378
rect 7060 4326 7070 4378
rect 7070 4326 7116 4378
rect 6820 4324 6876 4326
rect 6900 4324 6956 4326
rect 6980 4324 7036 4326
rect 7060 4324 7116 4326
rect 3888 3834 3944 3836
rect 3968 3834 4024 3836
rect 4048 3834 4104 3836
rect 4128 3834 4184 3836
rect 3888 3782 3934 3834
rect 3934 3782 3944 3834
rect 3968 3782 3998 3834
rect 3998 3782 4010 3834
rect 4010 3782 4024 3834
rect 4048 3782 4062 3834
rect 4062 3782 4074 3834
rect 4074 3782 4104 3834
rect 4128 3782 4138 3834
rect 4138 3782 4184 3834
rect 3888 3780 3944 3782
rect 3968 3780 4024 3782
rect 4048 3780 4104 3782
rect 4128 3780 4184 3782
rect 9753 3834 9809 3836
rect 9833 3834 9889 3836
rect 9913 3834 9969 3836
rect 9993 3834 10049 3836
rect 9753 3782 9799 3834
rect 9799 3782 9809 3834
rect 9833 3782 9863 3834
rect 9863 3782 9875 3834
rect 9875 3782 9889 3834
rect 9913 3782 9927 3834
rect 9927 3782 9939 3834
rect 9939 3782 9969 3834
rect 9993 3782 10003 3834
rect 10003 3782 10049 3834
rect 9753 3780 9809 3782
rect 9833 3780 9889 3782
rect 9913 3780 9969 3782
rect 9993 3780 10049 3782
rect 6820 3290 6876 3292
rect 6900 3290 6956 3292
rect 6980 3290 7036 3292
rect 7060 3290 7116 3292
rect 6820 3238 6866 3290
rect 6866 3238 6876 3290
rect 6900 3238 6930 3290
rect 6930 3238 6942 3290
rect 6942 3238 6956 3290
rect 6980 3238 6994 3290
rect 6994 3238 7006 3290
rect 7006 3238 7036 3290
rect 7060 3238 7070 3290
rect 7070 3238 7116 3290
rect 6820 3236 6876 3238
rect 6900 3236 6956 3238
rect 6980 3236 7036 3238
rect 7060 3236 7116 3238
rect 3888 2746 3944 2748
rect 3968 2746 4024 2748
rect 4048 2746 4104 2748
rect 4128 2746 4184 2748
rect 3888 2694 3934 2746
rect 3934 2694 3944 2746
rect 3968 2694 3998 2746
rect 3998 2694 4010 2746
rect 4010 2694 4024 2746
rect 4048 2694 4062 2746
rect 4062 2694 4074 2746
rect 4074 2694 4104 2746
rect 4128 2694 4138 2746
rect 4138 2694 4184 2746
rect 3888 2692 3944 2694
rect 3968 2692 4024 2694
rect 4048 2692 4104 2694
rect 4128 2692 4184 2694
rect 9753 2746 9809 2748
rect 9833 2746 9889 2748
rect 9913 2746 9969 2748
rect 9993 2746 10049 2748
rect 9753 2694 9799 2746
rect 9799 2694 9809 2746
rect 9833 2694 9863 2746
rect 9863 2694 9875 2746
rect 9875 2694 9889 2746
rect 9913 2694 9927 2746
rect 9927 2694 9939 2746
rect 9939 2694 9969 2746
rect 9993 2694 10003 2746
rect 10003 2694 10049 2746
rect 9753 2692 9809 2694
rect 9833 2692 9889 2694
rect 9913 2692 9969 2694
rect 9993 2692 10049 2694
rect 10690 2352 10746 2408
rect 6820 2202 6876 2204
rect 6900 2202 6956 2204
rect 6980 2202 7036 2204
rect 7060 2202 7116 2204
rect 6820 2150 6866 2202
rect 6866 2150 6876 2202
rect 6900 2150 6930 2202
rect 6930 2150 6942 2202
rect 6942 2150 6956 2202
rect 6980 2150 6994 2202
rect 6994 2150 7006 2202
rect 7006 2150 7036 2202
rect 7060 2150 7070 2202
rect 7070 2150 7116 2202
rect 6820 2148 6876 2150
rect 6900 2148 6956 2150
rect 6980 2148 7036 2150
rect 7060 2148 7116 2150
rect 12685 8730 12741 8732
rect 12765 8730 12821 8732
rect 12845 8730 12901 8732
rect 12925 8730 12981 8732
rect 12685 8678 12731 8730
rect 12731 8678 12741 8730
rect 12765 8678 12795 8730
rect 12795 8678 12807 8730
rect 12807 8678 12821 8730
rect 12845 8678 12859 8730
rect 12859 8678 12871 8730
rect 12871 8678 12901 8730
rect 12925 8678 12935 8730
rect 12935 8678 12981 8730
rect 12685 8676 12741 8678
rect 12765 8676 12821 8678
rect 12845 8676 12901 8678
rect 12925 8676 12981 8678
rect 13634 7928 13690 7984
rect 15014 8472 15070 8528
rect 15842 8336 15898 8392
rect 15618 8186 15674 8188
rect 15698 8186 15754 8188
rect 15778 8186 15834 8188
rect 15858 8186 15914 8188
rect 15618 8134 15664 8186
rect 15664 8134 15674 8186
rect 15698 8134 15728 8186
rect 15728 8134 15740 8186
rect 15740 8134 15754 8186
rect 15778 8134 15792 8186
rect 15792 8134 15804 8186
rect 15804 8134 15834 8186
rect 15858 8134 15868 8186
rect 15868 8134 15914 8186
rect 15618 8132 15674 8134
rect 15698 8132 15754 8134
rect 15778 8132 15834 8134
rect 15858 8132 15914 8134
rect 12685 7642 12741 7644
rect 12765 7642 12821 7644
rect 12845 7642 12901 7644
rect 12925 7642 12981 7644
rect 12685 7590 12731 7642
rect 12731 7590 12741 7642
rect 12765 7590 12795 7642
rect 12795 7590 12807 7642
rect 12807 7590 12821 7642
rect 12845 7590 12859 7642
rect 12859 7590 12871 7642
rect 12871 7590 12901 7642
rect 12925 7590 12935 7642
rect 12935 7590 12981 7642
rect 12685 7588 12741 7590
rect 12765 7588 12821 7590
rect 12845 7588 12901 7590
rect 12925 7588 12981 7590
rect 15618 7098 15674 7100
rect 15698 7098 15754 7100
rect 15778 7098 15834 7100
rect 15858 7098 15914 7100
rect 15618 7046 15664 7098
rect 15664 7046 15674 7098
rect 15698 7046 15728 7098
rect 15728 7046 15740 7098
rect 15740 7046 15754 7098
rect 15778 7046 15792 7098
rect 15792 7046 15804 7098
rect 15804 7046 15834 7098
rect 15858 7046 15868 7098
rect 15868 7046 15914 7098
rect 15618 7044 15674 7046
rect 15698 7044 15754 7046
rect 15778 7044 15834 7046
rect 15858 7044 15914 7046
rect 12685 6554 12741 6556
rect 12765 6554 12821 6556
rect 12845 6554 12901 6556
rect 12925 6554 12981 6556
rect 12685 6502 12731 6554
rect 12731 6502 12741 6554
rect 12765 6502 12795 6554
rect 12795 6502 12807 6554
rect 12807 6502 12821 6554
rect 12845 6502 12859 6554
rect 12859 6502 12871 6554
rect 12871 6502 12901 6554
rect 12925 6502 12935 6554
rect 12935 6502 12981 6554
rect 12685 6500 12741 6502
rect 12765 6500 12821 6502
rect 12845 6500 12901 6502
rect 12925 6500 12981 6502
rect 15618 6010 15674 6012
rect 15698 6010 15754 6012
rect 15778 6010 15834 6012
rect 15858 6010 15914 6012
rect 15618 5958 15664 6010
rect 15664 5958 15674 6010
rect 15698 5958 15728 6010
rect 15728 5958 15740 6010
rect 15740 5958 15754 6010
rect 15778 5958 15792 6010
rect 15792 5958 15804 6010
rect 15804 5958 15834 6010
rect 15858 5958 15868 6010
rect 15868 5958 15914 6010
rect 15618 5956 15674 5958
rect 15698 5956 15754 5958
rect 15778 5956 15834 5958
rect 15858 5956 15914 5958
rect 12685 5466 12741 5468
rect 12765 5466 12821 5468
rect 12845 5466 12901 5468
rect 12925 5466 12981 5468
rect 12685 5414 12731 5466
rect 12731 5414 12741 5466
rect 12765 5414 12795 5466
rect 12795 5414 12807 5466
rect 12807 5414 12821 5466
rect 12845 5414 12859 5466
rect 12859 5414 12871 5466
rect 12871 5414 12901 5466
rect 12925 5414 12935 5466
rect 12935 5414 12981 5466
rect 12685 5412 12741 5414
rect 12765 5412 12821 5414
rect 12845 5412 12901 5414
rect 12925 5412 12981 5414
rect 15618 4922 15674 4924
rect 15698 4922 15754 4924
rect 15778 4922 15834 4924
rect 15858 4922 15914 4924
rect 15618 4870 15664 4922
rect 15664 4870 15674 4922
rect 15698 4870 15728 4922
rect 15728 4870 15740 4922
rect 15740 4870 15754 4922
rect 15778 4870 15792 4922
rect 15792 4870 15804 4922
rect 15804 4870 15834 4922
rect 15858 4870 15868 4922
rect 15868 4870 15914 4922
rect 15618 4868 15674 4870
rect 15698 4868 15754 4870
rect 15778 4868 15834 4870
rect 15858 4868 15914 4870
rect 12685 4378 12741 4380
rect 12765 4378 12821 4380
rect 12845 4378 12901 4380
rect 12925 4378 12981 4380
rect 12685 4326 12731 4378
rect 12731 4326 12741 4378
rect 12765 4326 12795 4378
rect 12795 4326 12807 4378
rect 12807 4326 12821 4378
rect 12845 4326 12859 4378
rect 12859 4326 12871 4378
rect 12871 4326 12901 4378
rect 12925 4326 12935 4378
rect 12935 4326 12981 4378
rect 12685 4324 12741 4326
rect 12765 4324 12821 4326
rect 12845 4324 12901 4326
rect 12925 4324 12981 4326
rect 12685 3290 12741 3292
rect 12765 3290 12821 3292
rect 12845 3290 12901 3292
rect 12925 3290 12981 3292
rect 12685 3238 12731 3290
rect 12731 3238 12741 3290
rect 12765 3238 12795 3290
rect 12795 3238 12807 3290
rect 12807 3238 12821 3290
rect 12845 3238 12859 3290
rect 12859 3238 12871 3290
rect 12871 3238 12901 3290
rect 12925 3238 12935 3290
rect 12935 3238 12981 3290
rect 12685 3236 12741 3238
rect 12765 3236 12821 3238
rect 12845 3236 12901 3238
rect 12925 3236 12981 3238
rect 12685 2202 12741 2204
rect 12765 2202 12821 2204
rect 12845 2202 12901 2204
rect 12925 2202 12981 2204
rect 12685 2150 12731 2202
rect 12731 2150 12741 2202
rect 12765 2150 12795 2202
rect 12795 2150 12807 2202
rect 12807 2150 12821 2202
rect 12845 2150 12859 2202
rect 12859 2150 12871 2202
rect 12871 2150 12901 2202
rect 12925 2150 12935 2202
rect 12935 2150 12981 2202
rect 12685 2148 12741 2150
rect 12765 2148 12821 2150
rect 12845 2148 12901 2150
rect 12925 2148 12981 2150
rect 9034 1944 9090 2000
rect 3888 1658 3944 1660
rect 3968 1658 4024 1660
rect 4048 1658 4104 1660
rect 4128 1658 4184 1660
rect 3888 1606 3934 1658
rect 3934 1606 3944 1658
rect 3968 1606 3998 1658
rect 3998 1606 4010 1658
rect 4010 1606 4024 1658
rect 4048 1606 4062 1658
rect 4062 1606 4074 1658
rect 4074 1606 4104 1658
rect 4128 1606 4138 1658
rect 4138 1606 4184 1658
rect 3888 1604 3944 1606
rect 3968 1604 4024 1606
rect 4048 1604 4104 1606
rect 4128 1604 4184 1606
rect 7838 1828 7894 1864
rect 7838 1808 7840 1828
rect 7840 1808 7892 1828
rect 7892 1808 7894 1828
rect 9753 1658 9809 1660
rect 9833 1658 9889 1660
rect 9913 1658 9969 1660
rect 9993 1658 10049 1660
rect 9753 1606 9799 1658
rect 9799 1606 9809 1658
rect 9833 1606 9863 1658
rect 9863 1606 9875 1658
rect 9875 1606 9889 1658
rect 9913 1606 9927 1658
rect 9927 1606 9939 1658
rect 9939 1606 9969 1658
rect 9993 1606 10003 1658
rect 10003 1606 10049 1658
rect 9753 1604 9809 1606
rect 9833 1604 9889 1606
rect 9913 1604 9969 1606
rect 9993 1604 10049 1606
rect 15618 3834 15674 3836
rect 15698 3834 15754 3836
rect 15778 3834 15834 3836
rect 15858 3834 15914 3836
rect 15618 3782 15664 3834
rect 15664 3782 15674 3834
rect 15698 3782 15728 3834
rect 15728 3782 15740 3834
rect 15740 3782 15754 3834
rect 15778 3782 15792 3834
rect 15792 3782 15804 3834
rect 15804 3782 15834 3834
rect 15858 3782 15868 3834
rect 15868 3782 15914 3834
rect 15618 3780 15674 3782
rect 15698 3780 15754 3782
rect 15778 3780 15834 3782
rect 15858 3780 15914 3782
rect 15618 2746 15674 2748
rect 15698 2746 15754 2748
rect 15778 2746 15834 2748
rect 15858 2746 15914 2748
rect 15618 2694 15664 2746
rect 15664 2694 15674 2746
rect 15698 2694 15728 2746
rect 15728 2694 15740 2746
rect 15740 2694 15754 2746
rect 15778 2694 15792 2746
rect 15792 2694 15804 2746
rect 15804 2694 15834 2746
rect 15858 2694 15868 2746
rect 15868 2694 15914 2746
rect 15618 2692 15674 2694
rect 15698 2692 15754 2694
rect 15778 2692 15834 2694
rect 15858 2692 15914 2694
rect 18550 8730 18606 8732
rect 18630 8730 18686 8732
rect 18710 8730 18766 8732
rect 18790 8730 18846 8732
rect 18550 8678 18596 8730
rect 18596 8678 18606 8730
rect 18630 8678 18660 8730
rect 18660 8678 18672 8730
rect 18672 8678 18686 8730
rect 18710 8678 18724 8730
rect 18724 8678 18736 8730
rect 18736 8678 18766 8730
rect 18790 8678 18800 8730
rect 18800 8678 18846 8730
rect 18550 8676 18606 8678
rect 18630 8676 18686 8678
rect 18710 8676 18766 8678
rect 18790 8676 18846 8678
rect 18602 7792 18658 7848
rect 18550 7642 18606 7644
rect 18630 7642 18686 7644
rect 18710 7642 18766 7644
rect 18790 7642 18846 7644
rect 18550 7590 18596 7642
rect 18596 7590 18606 7642
rect 18630 7590 18660 7642
rect 18660 7590 18672 7642
rect 18672 7590 18686 7642
rect 18710 7590 18724 7642
rect 18724 7590 18736 7642
rect 18736 7590 18766 7642
rect 18790 7590 18800 7642
rect 18800 7590 18846 7642
rect 18550 7588 18606 7590
rect 18630 7588 18686 7590
rect 18710 7588 18766 7590
rect 18790 7588 18846 7590
rect 19982 7384 20038 7440
rect 19706 7248 19762 7304
rect 18550 6554 18606 6556
rect 18630 6554 18686 6556
rect 18710 6554 18766 6556
rect 18790 6554 18846 6556
rect 18550 6502 18596 6554
rect 18596 6502 18606 6554
rect 18630 6502 18660 6554
rect 18660 6502 18672 6554
rect 18672 6502 18686 6554
rect 18710 6502 18724 6554
rect 18724 6502 18736 6554
rect 18736 6502 18766 6554
rect 18790 6502 18800 6554
rect 18800 6502 18846 6554
rect 18550 6500 18606 6502
rect 18630 6500 18686 6502
rect 18710 6500 18766 6502
rect 18790 6500 18846 6502
rect 18550 5466 18606 5468
rect 18630 5466 18686 5468
rect 18710 5466 18766 5468
rect 18790 5466 18846 5468
rect 18550 5414 18596 5466
rect 18596 5414 18606 5466
rect 18630 5414 18660 5466
rect 18660 5414 18672 5466
rect 18672 5414 18686 5466
rect 18710 5414 18724 5466
rect 18724 5414 18736 5466
rect 18736 5414 18766 5466
rect 18790 5414 18800 5466
rect 18800 5414 18846 5466
rect 18550 5412 18606 5414
rect 18630 5412 18686 5414
rect 18710 5412 18766 5414
rect 18790 5412 18846 5414
rect 18550 4378 18606 4380
rect 18630 4378 18686 4380
rect 18710 4378 18766 4380
rect 18790 4378 18846 4380
rect 18550 4326 18596 4378
rect 18596 4326 18606 4378
rect 18630 4326 18660 4378
rect 18660 4326 18672 4378
rect 18672 4326 18686 4378
rect 18710 4326 18724 4378
rect 18724 4326 18736 4378
rect 18736 4326 18766 4378
rect 18790 4326 18800 4378
rect 18800 4326 18846 4378
rect 18550 4324 18606 4326
rect 18630 4324 18686 4326
rect 18710 4324 18766 4326
rect 18790 4324 18846 4326
rect 15618 1658 15674 1660
rect 15698 1658 15754 1660
rect 15778 1658 15834 1660
rect 15858 1658 15914 1660
rect 15618 1606 15664 1658
rect 15664 1606 15674 1658
rect 15698 1606 15728 1658
rect 15728 1606 15740 1658
rect 15740 1606 15754 1658
rect 15778 1606 15792 1658
rect 15792 1606 15804 1658
rect 15804 1606 15834 1658
rect 15858 1606 15868 1658
rect 15868 1606 15914 1658
rect 15618 1604 15674 1606
rect 15698 1604 15754 1606
rect 15778 1604 15834 1606
rect 15858 1604 15914 1606
rect 6820 1114 6876 1116
rect 6900 1114 6956 1116
rect 6980 1114 7036 1116
rect 7060 1114 7116 1116
rect 6820 1062 6866 1114
rect 6866 1062 6876 1114
rect 6900 1062 6930 1114
rect 6930 1062 6942 1114
rect 6942 1062 6956 1114
rect 6980 1062 6994 1114
rect 6994 1062 7006 1114
rect 7006 1062 7036 1114
rect 7060 1062 7070 1114
rect 7070 1062 7116 1114
rect 6820 1060 6876 1062
rect 6900 1060 6956 1062
rect 6980 1060 7036 1062
rect 7060 1060 7116 1062
rect 12685 1114 12741 1116
rect 12765 1114 12821 1116
rect 12845 1114 12901 1116
rect 12925 1114 12981 1116
rect 12685 1062 12731 1114
rect 12731 1062 12741 1114
rect 12765 1062 12795 1114
rect 12795 1062 12807 1114
rect 12807 1062 12821 1114
rect 12845 1062 12859 1114
rect 12859 1062 12871 1114
rect 12871 1062 12901 1114
rect 12925 1062 12935 1114
rect 12935 1062 12981 1114
rect 12685 1060 12741 1062
rect 12765 1060 12821 1062
rect 12845 1060 12901 1062
rect 12925 1060 12981 1062
rect 18550 3290 18606 3292
rect 18630 3290 18686 3292
rect 18710 3290 18766 3292
rect 18790 3290 18846 3292
rect 18550 3238 18596 3290
rect 18596 3238 18606 3290
rect 18630 3238 18660 3290
rect 18660 3238 18672 3290
rect 18672 3238 18686 3290
rect 18710 3238 18724 3290
rect 18724 3238 18736 3290
rect 18736 3238 18766 3290
rect 18790 3238 18800 3290
rect 18800 3238 18846 3290
rect 18550 3236 18606 3238
rect 18630 3236 18686 3238
rect 18710 3236 18766 3238
rect 18790 3236 18846 3238
rect 18550 2202 18606 2204
rect 18630 2202 18686 2204
rect 18710 2202 18766 2204
rect 18790 2202 18846 2204
rect 18550 2150 18596 2202
rect 18596 2150 18606 2202
rect 18630 2150 18660 2202
rect 18660 2150 18672 2202
rect 18672 2150 18686 2202
rect 18710 2150 18724 2202
rect 18724 2150 18736 2202
rect 18736 2150 18766 2202
rect 18790 2150 18800 2202
rect 18800 2150 18846 2202
rect 18550 2148 18606 2150
rect 18630 2148 18686 2150
rect 18710 2148 18766 2150
rect 18790 2148 18846 2150
rect 18550 1114 18606 1116
rect 18630 1114 18686 1116
rect 18710 1114 18766 1116
rect 18790 1114 18846 1116
rect 18550 1062 18596 1114
rect 18596 1062 18606 1114
rect 18630 1062 18660 1114
rect 18660 1062 18672 1114
rect 18672 1062 18686 1114
rect 18710 1062 18724 1114
rect 18724 1062 18736 1114
rect 18736 1062 18766 1114
rect 18790 1062 18800 1114
rect 18800 1062 18846 1114
rect 18550 1060 18606 1062
rect 18630 1060 18686 1062
rect 18710 1060 18766 1062
rect 18790 1060 18846 1062
rect 21483 8186 21539 8188
rect 21563 8186 21619 8188
rect 21643 8186 21699 8188
rect 21723 8186 21779 8188
rect 21483 8134 21529 8186
rect 21529 8134 21539 8186
rect 21563 8134 21593 8186
rect 21593 8134 21605 8186
rect 21605 8134 21619 8186
rect 21643 8134 21657 8186
rect 21657 8134 21669 8186
rect 21669 8134 21699 8186
rect 21723 8134 21733 8186
rect 21733 8134 21779 8186
rect 21483 8132 21539 8134
rect 21563 8132 21619 8134
rect 21643 8132 21699 8134
rect 21723 8132 21779 8134
rect 22466 8336 22522 8392
rect 23018 8336 23074 8392
rect 22098 7248 22154 7304
rect 21483 7098 21539 7100
rect 21563 7098 21619 7100
rect 21643 7098 21699 7100
rect 21723 7098 21779 7100
rect 21483 7046 21529 7098
rect 21529 7046 21539 7098
rect 21563 7046 21593 7098
rect 21593 7046 21605 7098
rect 21605 7046 21619 7098
rect 21643 7046 21657 7098
rect 21657 7046 21669 7098
rect 21669 7046 21699 7098
rect 21723 7046 21733 7098
rect 21733 7046 21779 7098
rect 21483 7044 21539 7046
rect 21563 7044 21619 7046
rect 21643 7044 21699 7046
rect 21723 7044 21779 7046
rect 21483 6010 21539 6012
rect 21563 6010 21619 6012
rect 21643 6010 21699 6012
rect 21723 6010 21779 6012
rect 21483 5958 21529 6010
rect 21529 5958 21539 6010
rect 21563 5958 21593 6010
rect 21593 5958 21605 6010
rect 21605 5958 21619 6010
rect 21643 5958 21657 6010
rect 21657 5958 21669 6010
rect 21669 5958 21699 6010
rect 21723 5958 21733 6010
rect 21733 5958 21779 6010
rect 21483 5956 21539 5958
rect 21563 5956 21619 5958
rect 21643 5956 21699 5958
rect 21723 5956 21779 5958
rect 21483 4922 21539 4924
rect 21563 4922 21619 4924
rect 21643 4922 21699 4924
rect 21723 4922 21779 4924
rect 21483 4870 21529 4922
rect 21529 4870 21539 4922
rect 21563 4870 21593 4922
rect 21593 4870 21605 4922
rect 21605 4870 21619 4922
rect 21643 4870 21657 4922
rect 21657 4870 21669 4922
rect 21669 4870 21699 4922
rect 21723 4870 21733 4922
rect 21733 4870 21779 4922
rect 21483 4868 21539 4870
rect 21563 4868 21619 4870
rect 21643 4868 21699 4870
rect 21723 4868 21779 4870
rect 21483 3834 21539 3836
rect 21563 3834 21619 3836
rect 21643 3834 21699 3836
rect 21723 3834 21779 3836
rect 21483 3782 21529 3834
rect 21529 3782 21539 3834
rect 21563 3782 21593 3834
rect 21593 3782 21605 3834
rect 21605 3782 21619 3834
rect 21643 3782 21657 3834
rect 21657 3782 21669 3834
rect 21669 3782 21699 3834
rect 21723 3782 21733 3834
rect 21733 3782 21779 3834
rect 21483 3780 21539 3782
rect 21563 3780 21619 3782
rect 21643 3780 21699 3782
rect 21723 3780 21779 3782
rect 21483 2746 21539 2748
rect 21563 2746 21619 2748
rect 21643 2746 21699 2748
rect 21723 2746 21779 2748
rect 21483 2694 21529 2746
rect 21529 2694 21539 2746
rect 21563 2694 21593 2746
rect 21593 2694 21605 2746
rect 21605 2694 21619 2746
rect 21643 2694 21657 2746
rect 21657 2694 21669 2746
rect 21669 2694 21699 2746
rect 21723 2694 21733 2746
rect 21733 2694 21779 2746
rect 21483 2692 21539 2694
rect 21563 2692 21619 2694
rect 21643 2692 21699 2694
rect 21723 2692 21779 2694
rect 21483 1658 21539 1660
rect 21563 1658 21619 1660
rect 21643 1658 21699 1660
rect 21723 1658 21779 1660
rect 21483 1606 21529 1658
rect 21529 1606 21539 1658
rect 21563 1606 21593 1658
rect 21593 1606 21605 1658
rect 21605 1606 21619 1658
rect 21643 1606 21657 1658
rect 21657 1606 21669 1658
rect 21669 1606 21699 1658
rect 21723 1606 21733 1658
rect 21733 1606 21779 1658
rect 21483 1604 21539 1606
rect 21563 1604 21619 1606
rect 21643 1604 21699 1606
rect 21723 1604 21779 1606
rect 24415 8730 24471 8732
rect 24495 8730 24551 8732
rect 24575 8730 24631 8732
rect 24655 8730 24711 8732
rect 24415 8678 24461 8730
rect 24461 8678 24471 8730
rect 24495 8678 24525 8730
rect 24525 8678 24537 8730
rect 24537 8678 24551 8730
rect 24575 8678 24589 8730
rect 24589 8678 24601 8730
rect 24601 8678 24631 8730
rect 24655 8678 24665 8730
rect 24665 8678 24711 8730
rect 24415 8676 24471 8678
rect 24495 8676 24551 8678
rect 24575 8676 24631 8678
rect 24655 8676 24711 8678
rect 24415 7642 24471 7644
rect 24495 7642 24551 7644
rect 24575 7642 24631 7644
rect 24655 7642 24711 7644
rect 24415 7590 24461 7642
rect 24461 7590 24471 7642
rect 24495 7590 24525 7642
rect 24525 7590 24537 7642
rect 24537 7590 24551 7642
rect 24575 7590 24589 7642
rect 24589 7590 24601 7642
rect 24601 7590 24631 7642
rect 24655 7590 24665 7642
rect 24665 7590 24711 7642
rect 24415 7588 24471 7590
rect 24495 7588 24551 7590
rect 24575 7588 24631 7590
rect 24655 7588 24711 7590
rect 24415 6554 24471 6556
rect 24495 6554 24551 6556
rect 24575 6554 24631 6556
rect 24655 6554 24711 6556
rect 24415 6502 24461 6554
rect 24461 6502 24471 6554
rect 24495 6502 24525 6554
rect 24525 6502 24537 6554
rect 24537 6502 24551 6554
rect 24575 6502 24589 6554
rect 24589 6502 24601 6554
rect 24601 6502 24631 6554
rect 24655 6502 24665 6554
rect 24665 6502 24711 6554
rect 24415 6500 24471 6502
rect 24495 6500 24551 6502
rect 24575 6500 24631 6502
rect 24655 6500 24711 6502
rect 24415 5466 24471 5468
rect 24495 5466 24551 5468
rect 24575 5466 24631 5468
rect 24655 5466 24711 5468
rect 24415 5414 24461 5466
rect 24461 5414 24471 5466
rect 24495 5414 24525 5466
rect 24525 5414 24537 5466
rect 24537 5414 24551 5466
rect 24575 5414 24589 5466
rect 24589 5414 24601 5466
rect 24601 5414 24631 5466
rect 24655 5414 24665 5466
rect 24665 5414 24711 5466
rect 24415 5412 24471 5414
rect 24495 5412 24551 5414
rect 24575 5412 24631 5414
rect 24655 5412 24711 5414
rect 24415 4378 24471 4380
rect 24495 4378 24551 4380
rect 24575 4378 24631 4380
rect 24655 4378 24711 4380
rect 24415 4326 24461 4378
rect 24461 4326 24471 4378
rect 24495 4326 24525 4378
rect 24525 4326 24537 4378
rect 24537 4326 24551 4378
rect 24575 4326 24589 4378
rect 24589 4326 24601 4378
rect 24601 4326 24631 4378
rect 24655 4326 24665 4378
rect 24665 4326 24711 4378
rect 24415 4324 24471 4326
rect 24495 4324 24551 4326
rect 24575 4324 24631 4326
rect 24655 4324 24711 4326
rect 24415 3290 24471 3292
rect 24495 3290 24551 3292
rect 24575 3290 24631 3292
rect 24655 3290 24711 3292
rect 24415 3238 24461 3290
rect 24461 3238 24471 3290
rect 24495 3238 24525 3290
rect 24525 3238 24537 3290
rect 24537 3238 24551 3290
rect 24575 3238 24589 3290
rect 24589 3238 24601 3290
rect 24601 3238 24631 3290
rect 24655 3238 24665 3290
rect 24665 3238 24711 3290
rect 24415 3236 24471 3238
rect 24495 3236 24551 3238
rect 24575 3236 24631 3238
rect 24655 3236 24711 3238
rect 24415 2202 24471 2204
rect 24495 2202 24551 2204
rect 24575 2202 24631 2204
rect 24655 2202 24711 2204
rect 24415 2150 24461 2202
rect 24461 2150 24471 2202
rect 24495 2150 24525 2202
rect 24525 2150 24537 2202
rect 24537 2150 24551 2202
rect 24575 2150 24589 2202
rect 24589 2150 24601 2202
rect 24601 2150 24631 2202
rect 24655 2150 24665 2202
rect 24665 2150 24711 2202
rect 24415 2148 24471 2150
rect 24495 2148 24551 2150
rect 24575 2148 24631 2150
rect 24655 2148 24711 2150
rect 24415 1114 24471 1116
rect 24495 1114 24551 1116
rect 24575 1114 24631 1116
rect 24655 1114 24711 1116
rect 24415 1062 24461 1114
rect 24461 1062 24471 1114
rect 24495 1062 24525 1114
rect 24525 1062 24537 1114
rect 24537 1062 24551 1114
rect 24575 1062 24589 1114
rect 24589 1062 24601 1114
rect 24601 1062 24631 1114
rect 24655 1062 24665 1114
rect 24665 1062 24711 1114
rect 24415 1060 24471 1062
rect 24495 1060 24551 1062
rect 24575 1060 24631 1062
rect 24655 1060 24711 1062
<< metal3 >>
rect 6810 8736 7126 8737
rect 6810 8672 6816 8736
rect 6880 8672 6896 8736
rect 6960 8672 6976 8736
rect 7040 8672 7056 8736
rect 7120 8672 7126 8736
rect 6810 8671 7126 8672
rect 12675 8736 12991 8737
rect 12675 8672 12681 8736
rect 12745 8672 12761 8736
rect 12825 8672 12841 8736
rect 12905 8672 12921 8736
rect 12985 8672 12991 8736
rect 12675 8671 12991 8672
rect 18540 8736 18856 8737
rect 18540 8672 18546 8736
rect 18610 8672 18626 8736
rect 18690 8672 18706 8736
rect 18770 8672 18786 8736
rect 18850 8672 18856 8736
rect 18540 8671 18856 8672
rect 24405 8736 24721 8737
rect 24405 8672 24411 8736
rect 24475 8672 24491 8736
rect 24555 8672 24571 8736
rect 24635 8672 24651 8736
rect 24715 8672 24721 8736
rect 24405 8671 24721 8672
rect 10225 8530 10291 8533
rect 15009 8530 15075 8533
rect 10225 8528 15075 8530
rect 10225 8472 10230 8528
rect 10286 8472 15014 8528
rect 15070 8472 15075 8528
rect 10225 8470 15075 8472
rect 10225 8467 10291 8470
rect 15009 8467 15075 8470
rect 15142 8332 15148 8396
rect 15212 8394 15218 8396
rect 15837 8394 15903 8397
rect 15212 8392 15903 8394
rect 15212 8336 15842 8392
rect 15898 8336 15903 8392
rect 15212 8334 15903 8336
rect 15212 8332 15218 8334
rect 15837 8331 15903 8334
rect 22318 8332 22324 8396
rect 22388 8394 22394 8396
rect 22461 8394 22527 8397
rect 22388 8392 22527 8394
rect 22388 8336 22466 8392
rect 22522 8336 22527 8392
rect 22388 8334 22527 8336
rect 22388 8332 22394 8334
rect 22461 8331 22527 8334
rect 22686 8332 22692 8396
rect 22756 8394 22762 8396
rect 23013 8394 23079 8397
rect 22756 8392 23079 8394
rect 22756 8336 23018 8392
rect 23074 8336 23079 8392
rect 22756 8334 23079 8336
rect 22756 8332 22762 8334
rect 23013 8331 23079 8334
rect 3878 8192 4194 8193
rect 3878 8128 3884 8192
rect 3948 8128 3964 8192
rect 4028 8128 4044 8192
rect 4108 8128 4124 8192
rect 4188 8128 4194 8192
rect 3878 8127 4194 8128
rect 9743 8192 10059 8193
rect 9743 8128 9749 8192
rect 9813 8128 9829 8192
rect 9893 8128 9909 8192
rect 9973 8128 9989 8192
rect 10053 8128 10059 8192
rect 9743 8127 10059 8128
rect 15608 8192 15924 8193
rect 15608 8128 15614 8192
rect 15678 8128 15694 8192
rect 15758 8128 15774 8192
rect 15838 8128 15854 8192
rect 15918 8128 15924 8192
rect 15608 8127 15924 8128
rect 21473 8192 21789 8193
rect 21473 8128 21479 8192
rect 21543 8128 21559 8192
rect 21623 8128 21639 8192
rect 21703 8128 21719 8192
rect 21783 8128 21789 8192
rect 21473 8127 21789 8128
rect 13629 7986 13695 7989
rect 2730 7984 13695 7986
rect 2730 7928 13634 7984
rect 13690 7928 13695 7984
rect 2730 7926 13695 7928
rect 2589 7850 2655 7853
rect 2730 7850 2790 7926
rect 13629 7923 13695 7926
rect 2589 7848 2790 7850
rect 2589 7792 2594 7848
rect 2650 7792 2790 7848
rect 2589 7790 2790 7792
rect 6729 7850 6795 7853
rect 18597 7850 18663 7853
rect 6729 7848 18663 7850
rect 6729 7792 6734 7848
rect 6790 7792 18602 7848
rect 18658 7792 18663 7848
rect 6729 7790 18663 7792
rect 2589 7787 2655 7790
rect 6729 7787 6795 7790
rect 18597 7787 18663 7790
rect 6810 7648 7126 7649
rect 6810 7584 6816 7648
rect 6880 7584 6896 7648
rect 6960 7584 6976 7648
rect 7040 7584 7056 7648
rect 7120 7584 7126 7648
rect 6810 7583 7126 7584
rect 12675 7648 12991 7649
rect 12675 7584 12681 7648
rect 12745 7584 12761 7648
rect 12825 7584 12841 7648
rect 12905 7584 12921 7648
rect 12985 7584 12991 7648
rect 12675 7583 12991 7584
rect 18540 7648 18856 7649
rect 18540 7584 18546 7648
rect 18610 7584 18626 7648
rect 18690 7584 18706 7648
rect 18770 7584 18786 7648
rect 18850 7584 18856 7648
rect 18540 7583 18856 7584
rect 24405 7648 24721 7649
rect 24405 7584 24411 7648
rect 24475 7584 24491 7648
rect 24555 7584 24571 7648
rect 24635 7584 24651 7648
rect 24715 7584 24721 7648
rect 24405 7583 24721 7584
rect 5625 7442 5691 7445
rect 19977 7442 20043 7445
rect 5625 7440 20043 7442
rect 5625 7384 5630 7440
rect 5686 7384 19982 7440
rect 20038 7384 20043 7440
rect 5625 7382 20043 7384
rect 5625 7379 5691 7382
rect 19977 7379 20043 7382
rect 6177 7306 6243 7309
rect 19701 7306 19767 7309
rect 6177 7304 19767 7306
rect 6177 7248 6182 7304
rect 6238 7248 19706 7304
rect 19762 7248 19767 7304
rect 6177 7246 19767 7248
rect 6177 7243 6243 7246
rect 19701 7243 19767 7246
rect 22093 7308 22159 7309
rect 22093 7304 22140 7308
rect 22204 7306 22210 7308
rect 22093 7248 22098 7304
rect 22093 7244 22140 7248
rect 22204 7246 22250 7306
rect 22204 7244 22210 7246
rect 22093 7243 22159 7244
rect 3878 7104 4194 7105
rect 3878 7040 3884 7104
rect 3948 7040 3964 7104
rect 4028 7040 4044 7104
rect 4108 7040 4124 7104
rect 4188 7040 4194 7104
rect 3878 7039 4194 7040
rect 9743 7104 10059 7105
rect 9743 7040 9749 7104
rect 9813 7040 9829 7104
rect 9893 7040 9909 7104
rect 9973 7040 9989 7104
rect 10053 7040 10059 7104
rect 9743 7039 10059 7040
rect 15608 7104 15924 7105
rect 15608 7040 15614 7104
rect 15678 7040 15694 7104
rect 15758 7040 15774 7104
rect 15838 7040 15854 7104
rect 15918 7040 15924 7104
rect 15608 7039 15924 7040
rect 21473 7104 21789 7105
rect 21473 7040 21479 7104
rect 21543 7040 21559 7104
rect 21623 7040 21639 7104
rect 21703 7040 21719 7104
rect 21783 7040 21789 7104
rect 21473 7039 21789 7040
rect 2681 6762 2747 6765
rect 15142 6762 15148 6764
rect 2681 6760 15148 6762
rect 2681 6704 2686 6760
rect 2742 6704 15148 6760
rect 2681 6702 15148 6704
rect 2681 6699 2747 6702
rect 15142 6700 15148 6702
rect 15212 6700 15218 6764
rect 6810 6560 7126 6561
rect 6810 6496 6816 6560
rect 6880 6496 6896 6560
rect 6960 6496 6976 6560
rect 7040 6496 7056 6560
rect 7120 6496 7126 6560
rect 6810 6495 7126 6496
rect 12675 6560 12991 6561
rect 12675 6496 12681 6560
rect 12745 6496 12761 6560
rect 12825 6496 12841 6560
rect 12905 6496 12921 6560
rect 12985 6496 12991 6560
rect 12675 6495 12991 6496
rect 18540 6560 18856 6561
rect 18540 6496 18546 6560
rect 18610 6496 18626 6560
rect 18690 6496 18706 6560
rect 18770 6496 18786 6560
rect 18850 6496 18856 6560
rect 18540 6495 18856 6496
rect 24405 6560 24721 6561
rect 24405 6496 24411 6560
rect 24475 6496 24491 6560
rect 24555 6496 24571 6560
rect 24635 6496 24651 6560
rect 24715 6496 24721 6560
rect 24405 6495 24721 6496
rect 3878 6016 4194 6017
rect 3878 5952 3884 6016
rect 3948 5952 3964 6016
rect 4028 5952 4044 6016
rect 4108 5952 4124 6016
rect 4188 5952 4194 6016
rect 3878 5951 4194 5952
rect 9743 6016 10059 6017
rect 9743 5952 9749 6016
rect 9813 5952 9829 6016
rect 9893 5952 9909 6016
rect 9973 5952 9989 6016
rect 10053 5952 10059 6016
rect 9743 5951 10059 5952
rect 15608 6016 15924 6017
rect 15608 5952 15614 6016
rect 15678 5952 15694 6016
rect 15758 5952 15774 6016
rect 15838 5952 15854 6016
rect 15918 5952 15924 6016
rect 15608 5951 15924 5952
rect 21473 6016 21789 6017
rect 21473 5952 21479 6016
rect 21543 5952 21559 6016
rect 21623 5952 21639 6016
rect 21703 5952 21719 6016
rect 21783 5952 21789 6016
rect 21473 5951 21789 5952
rect 6810 5472 7126 5473
rect 6810 5408 6816 5472
rect 6880 5408 6896 5472
rect 6960 5408 6976 5472
rect 7040 5408 7056 5472
rect 7120 5408 7126 5472
rect 6810 5407 7126 5408
rect 12675 5472 12991 5473
rect 12675 5408 12681 5472
rect 12745 5408 12761 5472
rect 12825 5408 12841 5472
rect 12905 5408 12921 5472
rect 12985 5408 12991 5472
rect 12675 5407 12991 5408
rect 18540 5472 18856 5473
rect 18540 5408 18546 5472
rect 18610 5408 18626 5472
rect 18690 5408 18706 5472
rect 18770 5408 18786 5472
rect 18850 5408 18856 5472
rect 18540 5407 18856 5408
rect 24405 5472 24721 5473
rect 24405 5408 24411 5472
rect 24475 5408 24491 5472
rect 24555 5408 24571 5472
rect 24635 5408 24651 5472
rect 24715 5408 24721 5472
rect 24405 5407 24721 5408
rect 3878 4928 4194 4929
rect 3878 4864 3884 4928
rect 3948 4864 3964 4928
rect 4028 4864 4044 4928
rect 4108 4864 4124 4928
rect 4188 4864 4194 4928
rect 3878 4863 4194 4864
rect 9743 4928 10059 4929
rect 9743 4864 9749 4928
rect 9813 4864 9829 4928
rect 9893 4864 9909 4928
rect 9973 4864 9989 4928
rect 10053 4864 10059 4928
rect 9743 4863 10059 4864
rect 15608 4928 15924 4929
rect 15608 4864 15614 4928
rect 15678 4864 15694 4928
rect 15758 4864 15774 4928
rect 15838 4864 15854 4928
rect 15918 4864 15924 4928
rect 15608 4863 15924 4864
rect 21473 4928 21789 4929
rect 21473 4864 21479 4928
rect 21543 4864 21559 4928
rect 21623 4864 21639 4928
rect 21703 4864 21719 4928
rect 21783 4864 21789 4928
rect 21473 4863 21789 4864
rect 6810 4384 7126 4385
rect 6810 4320 6816 4384
rect 6880 4320 6896 4384
rect 6960 4320 6976 4384
rect 7040 4320 7056 4384
rect 7120 4320 7126 4384
rect 6810 4319 7126 4320
rect 12675 4384 12991 4385
rect 12675 4320 12681 4384
rect 12745 4320 12761 4384
rect 12825 4320 12841 4384
rect 12905 4320 12921 4384
rect 12985 4320 12991 4384
rect 12675 4319 12991 4320
rect 18540 4384 18856 4385
rect 18540 4320 18546 4384
rect 18610 4320 18626 4384
rect 18690 4320 18706 4384
rect 18770 4320 18786 4384
rect 18850 4320 18856 4384
rect 18540 4319 18856 4320
rect 24405 4384 24721 4385
rect 24405 4320 24411 4384
rect 24475 4320 24491 4384
rect 24555 4320 24571 4384
rect 24635 4320 24651 4384
rect 24715 4320 24721 4384
rect 24405 4319 24721 4320
rect 3878 3840 4194 3841
rect 3878 3776 3884 3840
rect 3948 3776 3964 3840
rect 4028 3776 4044 3840
rect 4108 3776 4124 3840
rect 4188 3776 4194 3840
rect 3878 3775 4194 3776
rect 9743 3840 10059 3841
rect 9743 3776 9749 3840
rect 9813 3776 9829 3840
rect 9893 3776 9909 3840
rect 9973 3776 9989 3840
rect 10053 3776 10059 3840
rect 9743 3775 10059 3776
rect 15608 3840 15924 3841
rect 15608 3776 15614 3840
rect 15678 3776 15694 3840
rect 15758 3776 15774 3840
rect 15838 3776 15854 3840
rect 15918 3776 15924 3840
rect 15608 3775 15924 3776
rect 21473 3840 21789 3841
rect 21473 3776 21479 3840
rect 21543 3776 21559 3840
rect 21623 3776 21639 3840
rect 21703 3776 21719 3840
rect 21783 3776 21789 3840
rect 21473 3775 21789 3776
rect 6810 3296 7126 3297
rect 6810 3232 6816 3296
rect 6880 3232 6896 3296
rect 6960 3232 6976 3296
rect 7040 3232 7056 3296
rect 7120 3232 7126 3296
rect 6810 3231 7126 3232
rect 12675 3296 12991 3297
rect 12675 3232 12681 3296
rect 12745 3232 12761 3296
rect 12825 3232 12841 3296
rect 12905 3232 12921 3296
rect 12985 3232 12991 3296
rect 12675 3231 12991 3232
rect 18540 3296 18856 3297
rect 18540 3232 18546 3296
rect 18610 3232 18626 3296
rect 18690 3232 18706 3296
rect 18770 3232 18786 3296
rect 18850 3232 18856 3296
rect 18540 3231 18856 3232
rect 24405 3296 24721 3297
rect 24405 3232 24411 3296
rect 24475 3232 24491 3296
rect 24555 3232 24571 3296
rect 24635 3232 24651 3296
rect 24715 3232 24721 3296
rect 24405 3231 24721 3232
rect 3878 2752 4194 2753
rect 3878 2688 3884 2752
rect 3948 2688 3964 2752
rect 4028 2688 4044 2752
rect 4108 2688 4124 2752
rect 4188 2688 4194 2752
rect 3878 2687 4194 2688
rect 9743 2752 10059 2753
rect 9743 2688 9749 2752
rect 9813 2688 9829 2752
rect 9893 2688 9909 2752
rect 9973 2688 9989 2752
rect 10053 2688 10059 2752
rect 9743 2687 10059 2688
rect 15608 2752 15924 2753
rect 15608 2688 15614 2752
rect 15678 2688 15694 2752
rect 15758 2688 15774 2752
rect 15838 2688 15854 2752
rect 15918 2688 15924 2752
rect 15608 2687 15924 2688
rect 21473 2752 21789 2753
rect 21473 2688 21479 2752
rect 21543 2688 21559 2752
rect 21623 2688 21639 2752
rect 21703 2688 21719 2752
rect 21783 2688 21789 2752
rect 21473 2687 21789 2688
rect 10685 2410 10751 2413
rect 22134 2410 22140 2412
rect 10685 2408 22140 2410
rect 10685 2352 10690 2408
rect 10746 2352 22140 2408
rect 10685 2350 22140 2352
rect 10685 2347 10751 2350
rect 22134 2348 22140 2350
rect 22204 2348 22210 2412
rect 6810 2208 7126 2209
rect 6810 2144 6816 2208
rect 6880 2144 6896 2208
rect 6960 2144 6976 2208
rect 7040 2144 7056 2208
rect 7120 2144 7126 2208
rect 6810 2143 7126 2144
rect 12675 2208 12991 2209
rect 12675 2144 12681 2208
rect 12745 2144 12761 2208
rect 12825 2144 12841 2208
rect 12905 2144 12921 2208
rect 12985 2144 12991 2208
rect 12675 2143 12991 2144
rect 18540 2208 18856 2209
rect 18540 2144 18546 2208
rect 18610 2144 18626 2208
rect 18690 2144 18706 2208
rect 18770 2144 18786 2208
rect 18850 2144 18856 2208
rect 18540 2143 18856 2144
rect 24405 2208 24721 2209
rect 24405 2144 24411 2208
rect 24475 2144 24491 2208
rect 24555 2144 24571 2208
rect 24635 2144 24651 2208
rect 24715 2144 24721 2208
rect 24405 2143 24721 2144
rect 9029 2002 9095 2005
rect 22502 2002 22508 2004
rect 9029 2000 22508 2002
rect 9029 1944 9034 2000
rect 9090 1944 22508 2000
rect 9029 1942 22508 1944
rect 9029 1939 9095 1942
rect 22502 1940 22508 1942
rect 22572 1940 22578 2004
rect 7833 1866 7899 1869
rect 22318 1866 22324 1868
rect 7833 1864 22324 1866
rect 7833 1808 7838 1864
rect 7894 1808 22324 1864
rect 7833 1806 22324 1808
rect 7833 1803 7899 1806
rect 22318 1804 22324 1806
rect 22388 1804 22394 1868
rect 3878 1664 4194 1665
rect 3878 1600 3884 1664
rect 3948 1600 3964 1664
rect 4028 1600 4044 1664
rect 4108 1600 4124 1664
rect 4188 1600 4194 1664
rect 3878 1599 4194 1600
rect 9743 1664 10059 1665
rect 9743 1600 9749 1664
rect 9813 1600 9829 1664
rect 9893 1600 9909 1664
rect 9973 1600 9989 1664
rect 10053 1600 10059 1664
rect 9743 1599 10059 1600
rect 15608 1664 15924 1665
rect 15608 1600 15614 1664
rect 15678 1600 15694 1664
rect 15758 1600 15774 1664
rect 15838 1600 15854 1664
rect 15918 1600 15924 1664
rect 15608 1599 15924 1600
rect 21473 1664 21789 1665
rect 21473 1600 21479 1664
rect 21543 1600 21559 1664
rect 21623 1600 21639 1664
rect 21703 1600 21719 1664
rect 21783 1600 21789 1664
rect 21473 1599 21789 1600
rect 6810 1120 7126 1121
rect 6810 1056 6816 1120
rect 6880 1056 6896 1120
rect 6960 1056 6976 1120
rect 7040 1056 7056 1120
rect 7120 1056 7126 1120
rect 6810 1055 7126 1056
rect 12675 1120 12991 1121
rect 12675 1056 12681 1120
rect 12745 1056 12761 1120
rect 12825 1056 12841 1120
rect 12905 1056 12921 1120
rect 12985 1056 12991 1120
rect 12675 1055 12991 1056
rect 18540 1120 18856 1121
rect 18540 1056 18546 1120
rect 18610 1056 18626 1120
rect 18690 1056 18706 1120
rect 18770 1056 18786 1120
rect 18850 1056 18856 1120
rect 18540 1055 18856 1056
rect 24405 1120 24721 1121
rect 24405 1056 24411 1120
rect 24475 1056 24491 1120
rect 24555 1056 24571 1120
rect 24635 1056 24651 1120
rect 24715 1056 24721 1120
rect 24405 1055 24721 1056
<< via3 >>
rect 6816 8732 6880 8736
rect 6816 8676 6820 8732
rect 6820 8676 6876 8732
rect 6876 8676 6880 8732
rect 6816 8672 6880 8676
rect 6896 8732 6960 8736
rect 6896 8676 6900 8732
rect 6900 8676 6956 8732
rect 6956 8676 6960 8732
rect 6896 8672 6960 8676
rect 6976 8732 7040 8736
rect 6976 8676 6980 8732
rect 6980 8676 7036 8732
rect 7036 8676 7040 8732
rect 6976 8672 7040 8676
rect 7056 8732 7120 8736
rect 7056 8676 7060 8732
rect 7060 8676 7116 8732
rect 7116 8676 7120 8732
rect 7056 8672 7120 8676
rect 12681 8732 12745 8736
rect 12681 8676 12685 8732
rect 12685 8676 12741 8732
rect 12741 8676 12745 8732
rect 12681 8672 12745 8676
rect 12761 8732 12825 8736
rect 12761 8676 12765 8732
rect 12765 8676 12821 8732
rect 12821 8676 12825 8732
rect 12761 8672 12825 8676
rect 12841 8732 12905 8736
rect 12841 8676 12845 8732
rect 12845 8676 12901 8732
rect 12901 8676 12905 8732
rect 12841 8672 12905 8676
rect 12921 8732 12985 8736
rect 12921 8676 12925 8732
rect 12925 8676 12981 8732
rect 12981 8676 12985 8732
rect 12921 8672 12985 8676
rect 18546 8732 18610 8736
rect 18546 8676 18550 8732
rect 18550 8676 18606 8732
rect 18606 8676 18610 8732
rect 18546 8672 18610 8676
rect 18626 8732 18690 8736
rect 18626 8676 18630 8732
rect 18630 8676 18686 8732
rect 18686 8676 18690 8732
rect 18626 8672 18690 8676
rect 18706 8732 18770 8736
rect 18706 8676 18710 8732
rect 18710 8676 18766 8732
rect 18766 8676 18770 8732
rect 18706 8672 18770 8676
rect 18786 8732 18850 8736
rect 18786 8676 18790 8732
rect 18790 8676 18846 8732
rect 18846 8676 18850 8732
rect 18786 8672 18850 8676
rect 24411 8732 24475 8736
rect 24411 8676 24415 8732
rect 24415 8676 24471 8732
rect 24471 8676 24475 8732
rect 24411 8672 24475 8676
rect 24491 8732 24555 8736
rect 24491 8676 24495 8732
rect 24495 8676 24551 8732
rect 24551 8676 24555 8732
rect 24491 8672 24555 8676
rect 24571 8732 24635 8736
rect 24571 8676 24575 8732
rect 24575 8676 24631 8732
rect 24631 8676 24635 8732
rect 24571 8672 24635 8676
rect 24651 8732 24715 8736
rect 24651 8676 24655 8732
rect 24655 8676 24711 8732
rect 24711 8676 24715 8732
rect 24651 8672 24715 8676
rect 15148 8332 15212 8396
rect 22324 8332 22388 8396
rect 22692 8332 22756 8396
rect 3884 8188 3948 8192
rect 3884 8132 3888 8188
rect 3888 8132 3944 8188
rect 3944 8132 3948 8188
rect 3884 8128 3948 8132
rect 3964 8188 4028 8192
rect 3964 8132 3968 8188
rect 3968 8132 4024 8188
rect 4024 8132 4028 8188
rect 3964 8128 4028 8132
rect 4044 8188 4108 8192
rect 4044 8132 4048 8188
rect 4048 8132 4104 8188
rect 4104 8132 4108 8188
rect 4044 8128 4108 8132
rect 4124 8188 4188 8192
rect 4124 8132 4128 8188
rect 4128 8132 4184 8188
rect 4184 8132 4188 8188
rect 4124 8128 4188 8132
rect 9749 8188 9813 8192
rect 9749 8132 9753 8188
rect 9753 8132 9809 8188
rect 9809 8132 9813 8188
rect 9749 8128 9813 8132
rect 9829 8188 9893 8192
rect 9829 8132 9833 8188
rect 9833 8132 9889 8188
rect 9889 8132 9893 8188
rect 9829 8128 9893 8132
rect 9909 8188 9973 8192
rect 9909 8132 9913 8188
rect 9913 8132 9969 8188
rect 9969 8132 9973 8188
rect 9909 8128 9973 8132
rect 9989 8188 10053 8192
rect 9989 8132 9993 8188
rect 9993 8132 10049 8188
rect 10049 8132 10053 8188
rect 9989 8128 10053 8132
rect 15614 8188 15678 8192
rect 15614 8132 15618 8188
rect 15618 8132 15674 8188
rect 15674 8132 15678 8188
rect 15614 8128 15678 8132
rect 15694 8188 15758 8192
rect 15694 8132 15698 8188
rect 15698 8132 15754 8188
rect 15754 8132 15758 8188
rect 15694 8128 15758 8132
rect 15774 8188 15838 8192
rect 15774 8132 15778 8188
rect 15778 8132 15834 8188
rect 15834 8132 15838 8188
rect 15774 8128 15838 8132
rect 15854 8188 15918 8192
rect 15854 8132 15858 8188
rect 15858 8132 15914 8188
rect 15914 8132 15918 8188
rect 15854 8128 15918 8132
rect 21479 8188 21543 8192
rect 21479 8132 21483 8188
rect 21483 8132 21539 8188
rect 21539 8132 21543 8188
rect 21479 8128 21543 8132
rect 21559 8188 21623 8192
rect 21559 8132 21563 8188
rect 21563 8132 21619 8188
rect 21619 8132 21623 8188
rect 21559 8128 21623 8132
rect 21639 8188 21703 8192
rect 21639 8132 21643 8188
rect 21643 8132 21699 8188
rect 21699 8132 21703 8188
rect 21639 8128 21703 8132
rect 21719 8188 21783 8192
rect 21719 8132 21723 8188
rect 21723 8132 21779 8188
rect 21779 8132 21783 8188
rect 21719 8128 21783 8132
rect 6816 7644 6880 7648
rect 6816 7588 6820 7644
rect 6820 7588 6876 7644
rect 6876 7588 6880 7644
rect 6816 7584 6880 7588
rect 6896 7644 6960 7648
rect 6896 7588 6900 7644
rect 6900 7588 6956 7644
rect 6956 7588 6960 7644
rect 6896 7584 6960 7588
rect 6976 7644 7040 7648
rect 6976 7588 6980 7644
rect 6980 7588 7036 7644
rect 7036 7588 7040 7644
rect 6976 7584 7040 7588
rect 7056 7644 7120 7648
rect 7056 7588 7060 7644
rect 7060 7588 7116 7644
rect 7116 7588 7120 7644
rect 7056 7584 7120 7588
rect 12681 7644 12745 7648
rect 12681 7588 12685 7644
rect 12685 7588 12741 7644
rect 12741 7588 12745 7644
rect 12681 7584 12745 7588
rect 12761 7644 12825 7648
rect 12761 7588 12765 7644
rect 12765 7588 12821 7644
rect 12821 7588 12825 7644
rect 12761 7584 12825 7588
rect 12841 7644 12905 7648
rect 12841 7588 12845 7644
rect 12845 7588 12901 7644
rect 12901 7588 12905 7644
rect 12841 7584 12905 7588
rect 12921 7644 12985 7648
rect 12921 7588 12925 7644
rect 12925 7588 12981 7644
rect 12981 7588 12985 7644
rect 12921 7584 12985 7588
rect 18546 7644 18610 7648
rect 18546 7588 18550 7644
rect 18550 7588 18606 7644
rect 18606 7588 18610 7644
rect 18546 7584 18610 7588
rect 18626 7644 18690 7648
rect 18626 7588 18630 7644
rect 18630 7588 18686 7644
rect 18686 7588 18690 7644
rect 18626 7584 18690 7588
rect 18706 7644 18770 7648
rect 18706 7588 18710 7644
rect 18710 7588 18766 7644
rect 18766 7588 18770 7644
rect 18706 7584 18770 7588
rect 18786 7644 18850 7648
rect 18786 7588 18790 7644
rect 18790 7588 18846 7644
rect 18846 7588 18850 7644
rect 18786 7584 18850 7588
rect 24411 7644 24475 7648
rect 24411 7588 24415 7644
rect 24415 7588 24471 7644
rect 24471 7588 24475 7644
rect 24411 7584 24475 7588
rect 24491 7644 24555 7648
rect 24491 7588 24495 7644
rect 24495 7588 24551 7644
rect 24551 7588 24555 7644
rect 24491 7584 24555 7588
rect 24571 7644 24635 7648
rect 24571 7588 24575 7644
rect 24575 7588 24631 7644
rect 24631 7588 24635 7644
rect 24571 7584 24635 7588
rect 24651 7644 24715 7648
rect 24651 7588 24655 7644
rect 24655 7588 24711 7644
rect 24711 7588 24715 7644
rect 24651 7584 24715 7588
rect 22140 7304 22204 7308
rect 22140 7248 22154 7304
rect 22154 7248 22204 7304
rect 22140 7244 22204 7248
rect 3884 7100 3948 7104
rect 3884 7044 3888 7100
rect 3888 7044 3944 7100
rect 3944 7044 3948 7100
rect 3884 7040 3948 7044
rect 3964 7100 4028 7104
rect 3964 7044 3968 7100
rect 3968 7044 4024 7100
rect 4024 7044 4028 7100
rect 3964 7040 4028 7044
rect 4044 7100 4108 7104
rect 4044 7044 4048 7100
rect 4048 7044 4104 7100
rect 4104 7044 4108 7100
rect 4044 7040 4108 7044
rect 4124 7100 4188 7104
rect 4124 7044 4128 7100
rect 4128 7044 4184 7100
rect 4184 7044 4188 7100
rect 4124 7040 4188 7044
rect 9749 7100 9813 7104
rect 9749 7044 9753 7100
rect 9753 7044 9809 7100
rect 9809 7044 9813 7100
rect 9749 7040 9813 7044
rect 9829 7100 9893 7104
rect 9829 7044 9833 7100
rect 9833 7044 9889 7100
rect 9889 7044 9893 7100
rect 9829 7040 9893 7044
rect 9909 7100 9973 7104
rect 9909 7044 9913 7100
rect 9913 7044 9969 7100
rect 9969 7044 9973 7100
rect 9909 7040 9973 7044
rect 9989 7100 10053 7104
rect 9989 7044 9993 7100
rect 9993 7044 10049 7100
rect 10049 7044 10053 7100
rect 9989 7040 10053 7044
rect 15614 7100 15678 7104
rect 15614 7044 15618 7100
rect 15618 7044 15674 7100
rect 15674 7044 15678 7100
rect 15614 7040 15678 7044
rect 15694 7100 15758 7104
rect 15694 7044 15698 7100
rect 15698 7044 15754 7100
rect 15754 7044 15758 7100
rect 15694 7040 15758 7044
rect 15774 7100 15838 7104
rect 15774 7044 15778 7100
rect 15778 7044 15834 7100
rect 15834 7044 15838 7100
rect 15774 7040 15838 7044
rect 15854 7100 15918 7104
rect 15854 7044 15858 7100
rect 15858 7044 15914 7100
rect 15914 7044 15918 7100
rect 15854 7040 15918 7044
rect 21479 7100 21543 7104
rect 21479 7044 21483 7100
rect 21483 7044 21539 7100
rect 21539 7044 21543 7100
rect 21479 7040 21543 7044
rect 21559 7100 21623 7104
rect 21559 7044 21563 7100
rect 21563 7044 21619 7100
rect 21619 7044 21623 7100
rect 21559 7040 21623 7044
rect 21639 7100 21703 7104
rect 21639 7044 21643 7100
rect 21643 7044 21699 7100
rect 21699 7044 21703 7100
rect 21639 7040 21703 7044
rect 21719 7100 21783 7104
rect 21719 7044 21723 7100
rect 21723 7044 21779 7100
rect 21779 7044 21783 7100
rect 21719 7040 21783 7044
rect 15148 6700 15212 6764
rect 6816 6556 6880 6560
rect 6816 6500 6820 6556
rect 6820 6500 6876 6556
rect 6876 6500 6880 6556
rect 6816 6496 6880 6500
rect 6896 6556 6960 6560
rect 6896 6500 6900 6556
rect 6900 6500 6956 6556
rect 6956 6500 6960 6556
rect 6896 6496 6960 6500
rect 6976 6556 7040 6560
rect 6976 6500 6980 6556
rect 6980 6500 7036 6556
rect 7036 6500 7040 6556
rect 6976 6496 7040 6500
rect 7056 6556 7120 6560
rect 7056 6500 7060 6556
rect 7060 6500 7116 6556
rect 7116 6500 7120 6556
rect 7056 6496 7120 6500
rect 12681 6556 12745 6560
rect 12681 6500 12685 6556
rect 12685 6500 12741 6556
rect 12741 6500 12745 6556
rect 12681 6496 12745 6500
rect 12761 6556 12825 6560
rect 12761 6500 12765 6556
rect 12765 6500 12821 6556
rect 12821 6500 12825 6556
rect 12761 6496 12825 6500
rect 12841 6556 12905 6560
rect 12841 6500 12845 6556
rect 12845 6500 12901 6556
rect 12901 6500 12905 6556
rect 12841 6496 12905 6500
rect 12921 6556 12985 6560
rect 12921 6500 12925 6556
rect 12925 6500 12981 6556
rect 12981 6500 12985 6556
rect 12921 6496 12985 6500
rect 18546 6556 18610 6560
rect 18546 6500 18550 6556
rect 18550 6500 18606 6556
rect 18606 6500 18610 6556
rect 18546 6496 18610 6500
rect 18626 6556 18690 6560
rect 18626 6500 18630 6556
rect 18630 6500 18686 6556
rect 18686 6500 18690 6556
rect 18626 6496 18690 6500
rect 18706 6556 18770 6560
rect 18706 6500 18710 6556
rect 18710 6500 18766 6556
rect 18766 6500 18770 6556
rect 18706 6496 18770 6500
rect 18786 6556 18850 6560
rect 18786 6500 18790 6556
rect 18790 6500 18846 6556
rect 18846 6500 18850 6556
rect 18786 6496 18850 6500
rect 24411 6556 24475 6560
rect 24411 6500 24415 6556
rect 24415 6500 24471 6556
rect 24471 6500 24475 6556
rect 24411 6496 24475 6500
rect 24491 6556 24555 6560
rect 24491 6500 24495 6556
rect 24495 6500 24551 6556
rect 24551 6500 24555 6556
rect 24491 6496 24555 6500
rect 24571 6556 24635 6560
rect 24571 6500 24575 6556
rect 24575 6500 24631 6556
rect 24631 6500 24635 6556
rect 24571 6496 24635 6500
rect 24651 6556 24715 6560
rect 24651 6500 24655 6556
rect 24655 6500 24711 6556
rect 24711 6500 24715 6556
rect 24651 6496 24715 6500
rect 3884 6012 3948 6016
rect 3884 5956 3888 6012
rect 3888 5956 3944 6012
rect 3944 5956 3948 6012
rect 3884 5952 3948 5956
rect 3964 6012 4028 6016
rect 3964 5956 3968 6012
rect 3968 5956 4024 6012
rect 4024 5956 4028 6012
rect 3964 5952 4028 5956
rect 4044 6012 4108 6016
rect 4044 5956 4048 6012
rect 4048 5956 4104 6012
rect 4104 5956 4108 6012
rect 4044 5952 4108 5956
rect 4124 6012 4188 6016
rect 4124 5956 4128 6012
rect 4128 5956 4184 6012
rect 4184 5956 4188 6012
rect 4124 5952 4188 5956
rect 9749 6012 9813 6016
rect 9749 5956 9753 6012
rect 9753 5956 9809 6012
rect 9809 5956 9813 6012
rect 9749 5952 9813 5956
rect 9829 6012 9893 6016
rect 9829 5956 9833 6012
rect 9833 5956 9889 6012
rect 9889 5956 9893 6012
rect 9829 5952 9893 5956
rect 9909 6012 9973 6016
rect 9909 5956 9913 6012
rect 9913 5956 9969 6012
rect 9969 5956 9973 6012
rect 9909 5952 9973 5956
rect 9989 6012 10053 6016
rect 9989 5956 9993 6012
rect 9993 5956 10049 6012
rect 10049 5956 10053 6012
rect 9989 5952 10053 5956
rect 15614 6012 15678 6016
rect 15614 5956 15618 6012
rect 15618 5956 15674 6012
rect 15674 5956 15678 6012
rect 15614 5952 15678 5956
rect 15694 6012 15758 6016
rect 15694 5956 15698 6012
rect 15698 5956 15754 6012
rect 15754 5956 15758 6012
rect 15694 5952 15758 5956
rect 15774 6012 15838 6016
rect 15774 5956 15778 6012
rect 15778 5956 15834 6012
rect 15834 5956 15838 6012
rect 15774 5952 15838 5956
rect 15854 6012 15918 6016
rect 15854 5956 15858 6012
rect 15858 5956 15914 6012
rect 15914 5956 15918 6012
rect 15854 5952 15918 5956
rect 21479 6012 21543 6016
rect 21479 5956 21483 6012
rect 21483 5956 21539 6012
rect 21539 5956 21543 6012
rect 21479 5952 21543 5956
rect 21559 6012 21623 6016
rect 21559 5956 21563 6012
rect 21563 5956 21619 6012
rect 21619 5956 21623 6012
rect 21559 5952 21623 5956
rect 21639 6012 21703 6016
rect 21639 5956 21643 6012
rect 21643 5956 21699 6012
rect 21699 5956 21703 6012
rect 21639 5952 21703 5956
rect 21719 6012 21783 6016
rect 21719 5956 21723 6012
rect 21723 5956 21779 6012
rect 21779 5956 21783 6012
rect 21719 5952 21783 5956
rect 6816 5468 6880 5472
rect 6816 5412 6820 5468
rect 6820 5412 6876 5468
rect 6876 5412 6880 5468
rect 6816 5408 6880 5412
rect 6896 5468 6960 5472
rect 6896 5412 6900 5468
rect 6900 5412 6956 5468
rect 6956 5412 6960 5468
rect 6896 5408 6960 5412
rect 6976 5468 7040 5472
rect 6976 5412 6980 5468
rect 6980 5412 7036 5468
rect 7036 5412 7040 5468
rect 6976 5408 7040 5412
rect 7056 5468 7120 5472
rect 7056 5412 7060 5468
rect 7060 5412 7116 5468
rect 7116 5412 7120 5468
rect 7056 5408 7120 5412
rect 12681 5468 12745 5472
rect 12681 5412 12685 5468
rect 12685 5412 12741 5468
rect 12741 5412 12745 5468
rect 12681 5408 12745 5412
rect 12761 5468 12825 5472
rect 12761 5412 12765 5468
rect 12765 5412 12821 5468
rect 12821 5412 12825 5468
rect 12761 5408 12825 5412
rect 12841 5468 12905 5472
rect 12841 5412 12845 5468
rect 12845 5412 12901 5468
rect 12901 5412 12905 5468
rect 12841 5408 12905 5412
rect 12921 5468 12985 5472
rect 12921 5412 12925 5468
rect 12925 5412 12981 5468
rect 12981 5412 12985 5468
rect 12921 5408 12985 5412
rect 18546 5468 18610 5472
rect 18546 5412 18550 5468
rect 18550 5412 18606 5468
rect 18606 5412 18610 5468
rect 18546 5408 18610 5412
rect 18626 5468 18690 5472
rect 18626 5412 18630 5468
rect 18630 5412 18686 5468
rect 18686 5412 18690 5468
rect 18626 5408 18690 5412
rect 18706 5468 18770 5472
rect 18706 5412 18710 5468
rect 18710 5412 18766 5468
rect 18766 5412 18770 5468
rect 18706 5408 18770 5412
rect 18786 5468 18850 5472
rect 18786 5412 18790 5468
rect 18790 5412 18846 5468
rect 18846 5412 18850 5468
rect 18786 5408 18850 5412
rect 24411 5468 24475 5472
rect 24411 5412 24415 5468
rect 24415 5412 24471 5468
rect 24471 5412 24475 5468
rect 24411 5408 24475 5412
rect 24491 5468 24555 5472
rect 24491 5412 24495 5468
rect 24495 5412 24551 5468
rect 24551 5412 24555 5468
rect 24491 5408 24555 5412
rect 24571 5468 24635 5472
rect 24571 5412 24575 5468
rect 24575 5412 24631 5468
rect 24631 5412 24635 5468
rect 24571 5408 24635 5412
rect 24651 5468 24715 5472
rect 24651 5412 24655 5468
rect 24655 5412 24711 5468
rect 24711 5412 24715 5468
rect 24651 5408 24715 5412
rect 3884 4924 3948 4928
rect 3884 4868 3888 4924
rect 3888 4868 3944 4924
rect 3944 4868 3948 4924
rect 3884 4864 3948 4868
rect 3964 4924 4028 4928
rect 3964 4868 3968 4924
rect 3968 4868 4024 4924
rect 4024 4868 4028 4924
rect 3964 4864 4028 4868
rect 4044 4924 4108 4928
rect 4044 4868 4048 4924
rect 4048 4868 4104 4924
rect 4104 4868 4108 4924
rect 4044 4864 4108 4868
rect 4124 4924 4188 4928
rect 4124 4868 4128 4924
rect 4128 4868 4184 4924
rect 4184 4868 4188 4924
rect 4124 4864 4188 4868
rect 9749 4924 9813 4928
rect 9749 4868 9753 4924
rect 9753 4868 9809 4924
rect 9809 4868 9813 4924
rect 9749 4864 9813 4868
rect 9829 4924 9893 4928
rect 9829 4868 9833 4924
rect 9833 4868 9889 4924
rect 9889 4868 9893 4924
rect 9829 4864 9893 4868
rect 9909 4924 9973 4928
rect 9909 4868 9913 4924
rect 9913 4868 9969 4924
rect 9969 4868 9973 4924
rect 9909 4864 9973 4868
rect 9989 4924 10053 4928
rect 9989 4868 9993 4924
rect 9993 4868 10049 4924
rect 10049 4868 10053 4924
rect 9989 4864 10053 4868
rect 15614 4924 15678 4928
rect 15614 4868 15618 4924
rect 15618 4868 15674 4924
rect 15674 4868 15678 4924
rect 15614 4864 15678 4868
rect 15694 4924 15758 4928
rect 15694 4868 15698 4924
rect 15698 4868 15754 4924
rect 15754 4868 15758 4924
rect 15694 4864 15758 4868
rect 15774 4924 15838 4928
rect 15774 4868 15778 4924
rect 15778 4868 15834 4924
rect 15834 4868 15838 4924
rect 15774 4864 15838 4868
rect 15854 4924 15918 4928
rect 15854 4868 15858 4924
rect 15858 4868 15914 4924
rect 15914 4868 15918 4924
rect 15854 4864 15918 4868
rect 21479 4924 21543 4928
rect 21479 4868 21483 4924
rect 21483 4868 21539 4924
rect 21539 4868 21543 4924
rect 21479 4864 21543 4868
rect 21559 4924 21623 4928
rect 21559 4868 21563 4924
rect 21563 4868 21619 4924
rect 21619 4868 21623 4924
rect 21559 4864 21623 4868
rect 21639 4924 21703 4928
rect 21639 4868 21643 4924
rect 21643 4868 21699 4924
rect 21699 4868 21703 4924
rect 21639 4864 21703 4868
rect 21719 4924 21783 4928
rect 21719 4868 21723 4924
rect 21723 4868 21779 4924
rect 21779 4868 21783 4924
rect 21719 4864 21783 4868
rect 6816 4380 6880 4384
rect 6816 4324 6820 4380
rect 6820 4324 6876 4380
rect 6876 4324 6880 4380
rect 6816 4320 6880 4324
rect 6896 4380 6960 4384
rect 6896 4324 6900 4380
rect 6900 4324 6956 4380
rect 6956 4324 6960 4380
rect 6896 4320 6960 4324
rect 6976 4380 7040 4384
rect 6976 4324 6980 4380
rect 6980 4324 7036 4380
rect 7036 4324 7040 4380
rect 6976 4320 7040 4324
rect 7056 4380 7120 4384
rect 7056 4324 7060 4380
rect 7060 4324 7116 4380
rect 7116 4324 7120 4380
rect 7056 4320 7120 4324
rect 12681 4380 12745 4384
rect 12681 4324 12685 4380
rect 12685 4324 12741 4380
rect 12741 4324 12745 4380
rect 12681 4320 12745 4324
rect 12761 4380 12825 4384
rect 12761 4324 12765 4380
rect 12765 4324 12821 4380
rect 12821 4324 12825 4380
rect 12761 4320 12825 4324
rect 12841 4380 12905 4384
rect 12841 4324 12845 4380
rect 12845 4324 12901 4380
rect 12901 4324 12905 4380
rect 12841 4320 12905 4324
rect 12921 4380 12985 4384
rect 12921 4324 12925 4380
rect 12925 4324 12981 4380
rect 12981 4324 12985 4380
rect 12921 4320 12985 4324
rect 18546 4380 18610 4384
rect 18546 4324 18550 4380
rect 18550 4324 18606 4380
rect 18606 4324 18610 4380
rect 18546 4320 18610 4324
rect 18626 4380 18690 4384
rect 18626 4324 18630 4380
rect 18630 4324 18686 4380
rect 18686 4324 18690 4380
rect 18626 4320 18690 4324
rect 18706 4380 18770 4384
rect 18706 4324 18710 4380
rect 18710 4324 18766 4380
rect 18766 4324 18770 4380
rect 18706 4320 18770 4324
rect 18786 4380 18850 4384
rect 18786 4324 18790 4380
rect 18790 4324 18846 4380
rect 18846 4324 18850 4380
rect 18786 4320 18850 4324
rect 24411 4380 24475 4384
rect 24411 4324 24415 4380
rect 24415 4324 24471 4380
rect 24471 4324 24475 4380
rect 24411 4320 24475 4324
rect 24491 4380 24555 4384
rect 24491 4324 24495 4380
rect 24495 4324 24551 4380
rect 24551 4324 24555 4380
rect 24491 4320 24555 4324
rect 24571 4380 24635 4384
rect 24571 4324 24575 4380
rect 24575 4324 24631 4380
rect 24631 4324 24635 4380
rect 24571 4320 24635 4324
rect 24651 4380 24715 4384
rect 24651 4324 24655 4380
rect 24655 4324 24711 4380
rect 24711 4324 24715 4380
rect 24651 4320 24715 4324
rect 3884 3836 3948 3840
rect 3884 3780 3888 3836
rect 3888 3780 3944 3836
rect 3944 3780 3948 3836
rect 3884 3776 3948 3780
rect 3964 3836 4028 3840
rect 3964 3780 3968 3836
rect 3968 3780 4024 3836
rect 4024 3780 4028 3836
rect 3964 3776 4028 3780
rect 4044 3836 4108 3840
rect 4044 3780 4048 3836
rect 4048 3780 4104 3836
rect 4104 3780 4108 3836
rect 4044 3776 4108 3780
rect 4124 3836 4188 3840
rect 4124 3780 4128 3836
rect 4128 3780 4184 3836
rect 4184 3780 4188 3836
rect 4124 3776 4188 3780
rect 9749 3836 9813 3840
rect 9749 3780 9753 3836
rect 9753 3780 9809 3836
rect 9809 3780 9813 3836
rect 9749 3776 9813 3780
rect 9829 3836 9893 3840
rect 9829 3780 9833 3836
rect 9833 3780 9889 3836
rect 9889 3780 9893 3836
rect 9829 3776 9893 3780
rect 9909 3836 9973 3840
rect 9909 3780 9913 3836
rect 9913 3780 9969 3836
rect 9969 3780 9973 3836
rect 9909 3776 9973 3780
rect 9989 3836 10053 3840
rect 9989 3780 9993 3836
rect 9993 3780 10049 3836
rect 10049 3780 10053 3836
rect 9989 3776 10053 3780
rect 15614 3836 15678 3840
rect 15614 3780 15618 3836
rect 15618 3780 15674 3836
rect 15674 3780 15678 3836
rect 15614 3776 15678 3780
rect 15694 3836 15758 3840
rect 15694 3780 15698 3836
rect 15698 3780 15754 3836
rect 15754 3780 15758 3836
rect 15694 3776 15758 3780
rect 15774 3836 15838 3840
rect 15774 3780 15778 3836
rect 15778 3780 15834 3836
rect 15834 3780 15838 3836
rect 15774 3776 15838 3780
rect 15854 3836 15918 3840
rect 15854 3780 15858 3836
rect 15858 3780 15914 3836
rect 15914 3780 15918 3836
rect 15854 3776 15918 3780
rect 21479 3836 21543 3840
rect 21479 3780 21483 3836
rect 21483 3780 21539 3836
rect 21539 3780 21543 3836
rect 21479 3776 21543 3780
rect 21559 3836 21623 3840
rect 21559 3780 21563 3836
rect 21563 3780 21619 3836
rect 21619 3780 21623 3836
rect 21559 3776 21623 3780
rect 21639 3836 21703 3840
rect 21639 3780 21643 3836
rect 21643 3780 21699 3836
rect 21699 3780 21703 3836
rect 21639 3776 21703 3780
rect 21719 3836 21783 3840
rect 21719 3780 21723 3836
rect 21723 3780 21779 3836
rect 21779 3780 21783 3836
rect 21719 3776 21783 3780
rect 6816 3292 6880 3296
rect 6816 3236 6820 3292
rect 6820 3236 6876 3292
rect 6876 3236 6880 3292
rect 6816 3232 6880 3236
rect 6896 3292 6960 3296
rect 6896 3236 6900 3292
rect 6900 3236 6956 3292
rect 6956 3236 6960 3292
rect 6896 3232 6960 3236
rect 6976 3292 7040 3296
rect 6976 3236 6980 3292
rect 6980 3236 7036 3292
rect 7036 3236 7040 3292
rect 6976 3232 7040 3236
rect 7056 3292 7120 3296
rect 7056 3236 7060 3292
rect 7060 3236 7116 3292
rect 7116 3236 7120 3292
rect 7056 3232 7120 3236
rect 12681 3292 12745 3296
rect 12681 3236 12685 3292
rect 12685 3236 12741 3292
rect 12741 3236 12745 3292
rect 12681 3232 12745 3236
rect 12761 3292 12825 3296
rect 12761 3236 12765 3292
rect 12765 3236 12821 3292
rect 12821 3236 12825 3292
rect 12761 3232 12825 3236
rect 12841 3292 12905 3296
rect 12841 3236 12845 3292
rect 12845 3236 12901 3292
rect 12901 3236 12905 3292
rect 12841 3232 12905 3236
rect 12921 3292 12985 3296
rect 12921 3236 12925 3292
rect 12925 3236 12981 3292
rect 12981 3236 12985 3292
rect 12921 3232 12985 3236
rect 18546 3292 18610 3296
rect 18546 3236 18550 3292
rect 18550 3236 18606 3292
rect 18606 3236 18610 3292
rect 18546 3232 18610 3236
rect 18626 3292 18690 3296
rect 18626 3236 18630 3292
rect 18630 3236 18686 3292
rect 18686 3236 18690 3292
rect 18626 3232 18690 3236
rect 18706 3292 18770 3296
rect 18706 3236 18710 3292
rect 18710 3236 18766 3292
rect 18766 3236 18770 3292
rect 18706 3232 18770 3236
rect 18786 3292 18850 3296
rect 18786 3236 18790 3292
rect 18790 3236 18846 3292
rect 18846 3236 18850 3292
rect 18786 3232 18850 3236
rect 24411 3292 24475 3296
rect 24411 3236 24415 3292
rect 24415 3236 24471 3292
rect 24471 3236 24475 3292
rect 24411 3232 24475 3236
rect 24491 3292 24555 3296
rect 24491 3236 24495 3292
rect 24495 3236 24551 3292
rect 24551 3236 24555 3292
rect 24491 3232 24555 3236
rect 24571 3292 24635 3296
rect 24571 3236 24575 3292
rect 24575 3236 24631 3292
rect 24631 3236 24635 3292
rect 24571 3232 24635 3236
rect 24651 3292 24715 3296
rect 24651 3236 24655 3292
rect 24655 3236 24711 3292
rect 24711 3236 24715 3292
rect 24651 3232 24715 3236
rect 3884 2748 3948 2752
rect 3884 2692 3888 2748
rect 3888 2692 3944 2748
rect 3944 2692 3948 2748
rect 3884 2688 3948 2692
rect 3964 2748 4028 2752
rect 3964 2692 3968 2748
rect 3968 2692 4024 2748
rect 4024 2692 4028 2748
rect 3964 2688 4028 2692
rect 4044 2748 4108 2752
rect 4044 2692 4048 2748
rect 4048 2692 4104 2748
rect 4104 2692 4108 2748
rect 4044 2688 4108 2692
rect 4124 2748 4188 2752
rect 4124 2692 4128 2748
rect 4128 2692 4184 2748
rect 4184 2692 4188 2748
rect 4124 2688 4188 2692
rect 9749 2748 9813 2752
rect 9749 2692 9753 2748
rect 9753 2692 9809 2748
rect 9809 2692 9813 2748
rect 9749 2688 9813 2692
rect 9829 2748 9893 2752
rect 9829 2692 9833 2748
rect 9833 2692 9889 2748
rect 9889 2692 9893 2748
rect 9829 2688 9893 2692
rect 9909 2748 9973 2752
rect 9909 2692 9913 2748
rect 9913 2692 9969 2748
rect 9969 2692 9973 2748
rect 9909 2688 9973 2692
rect 9989 2748 10053 2752
rect 9989 2692 9993 2748
rect 9993 2692 10049 2748
rect 10049 2692 10053 2748
rect 9989 2688 10053 2692
rect 15614 2748 15678 2752
rect 15614 2692 15618 2748
rect 15618 2692 15674 2748
rect 15674 2692 15678 2748
rect 15614 2688 15678 2692
rect 15694 2748 15758 2752
rect 15694 2692 15698 2748
rect 15698 2692 15754 2748
rect 15754 2692 15758 2748
rect 15694 2688 15758 2692
rect 15774 2748 15838 2752
rect 15774 2692 15778 2748
rect 15778 2692 15834 2748
rect 15834 2692 15838 2748
rect 15774 2688 15838 2692
rect 15854 2748 15918 2752
rect 15854 2692 15858 2748
rect 15858 2692 15914 2748
rect 15914 2692 15918 2748
rect 15854 2688 15918 2692
rect 21479 2748 21543 2752
rect 21479 2692 21483 2748
rect 21483 2692 21539 2748
rect 21539 2692 21543 2748
rect 21479 2688 21543 2692
rect 21559 2748 21623 2752
rect 21559 2692 21563 2748
rect 21563 2692 21619 2748
rect 21619 2692 21623 2748
rect 21559 2688 21623 2692
rect 21639 2748 21703 2752
rect 21639 2692 21643 2748
rect 21643 2692 21699 2748
rect 21699 2692 21703 2748
rect 21639 2688 21703 2692
rect 21719 2748 21783 2752
rect 21719 2692 21723 2748
rect 21723 2692 21779 2748
rect 21779 2692 21783 2748
rect 21719 2688 21783 2692
rect 22140 2348 22204 2412
rect 6816 2204 6880 2208
rect 6816 2148 6820 2204
rect 6820 2148 6876 2204
rect 6876 2148 6880 2204
rect 6816 2144 6880 2148
rect 6896 2204 6960 2208
rect 6896 2148 6900 2204
rect 6900 2148 6956 2204
rect 6956 2148 6960 2204
rect 6896 2144 6960 2148
rect 6976 2204 7040 2208
rect 6976 2148 6980 2204
rect 6980 2148 7036 2204
rect 7036 2148 7040 2204
rect 6976 2144 7040 2148
rect 7056 2204 7120 2208
rect 7056 2148 7060 2204
rect 7060 2148 7116 2204
rect 7116 2148 7120 2204
rect 7056 2144 7120 2148
rect 12681 2204 12745 2208
rect 12681 2148 12685 2204
rect 12685 2148 12741 2204
rect 12741 2148 12745 2204
rect 12681 2144 12745 2148
rect 12761 2204 12825 2208
rect 12761 2148 12765 2204
rect 12765 2148 12821 2204
rect 12821 2148 12825 2204
rect 12761 2144 12825 2148
rect 12841 2204 12905 2208
rect 12841 2148 12845 2204
rect 12845 2148 12901 2204
rect 12901 2148 12905 2204
rect 12841 2144 12905 2148
rect 12921 2204 12985 2208
rect 12921 2148 12925 2204
rect 12925 2148 12981 2204
rect 12981 2148 12985 2204
rect 12921 2144 12985 2148
rect 18546 2204 18610 2208
rect 18546 2148 18550 2204
rect 18550 2148 18606 2204
rect 18606 2148 18610 2204
rect 18546 2144 18610 2148
rect 18626 2204 18690 2208
rect 18626 2148 18630 2204
rect 18630 2148 18686 2204
rect 18686 2148 18690 2204
rect 18626 2144 18690 2148
rect 18706 2204 18770 2208
rect 18706 2148 18710 2204
rect 18710 2148 18766 2204
rect 18766 2148 18770 2204
rect 18706 2144 18770 2148
rect 18786 2204 18850 2208
rect 18786 2148 18790 2204
rect 18790 2148 18846 2204
rect 18846 2148 18850 2204
rect 18786 2144 18850 2148
rect 24411 2204 24475 2208
rect 24411 2148 24415 2204
rect 24415 2148 24471 2204
rect 24471 2148 24475 2204
rect 24411 2144 24475 2148
rect 24491 2204 24555 2208
rect 24491 2148 24495 2204
rect 24495 2148 24551 2204
rect 24551 2148 24555 2204
rect 24491 2144 24555 2148
rect 24571 2204 24635 2208
rect 24571 2148 24575 2204
rect 24575 2148 24631 2204
rect 24631 2148 24635 2204
rect 24571 2144 24635 2148
rect 24651 2204 24715 2208
rect 24651 2148 24655 2204
rect 24655 2148 24711 2204
rect 24711 2148 24715 2204
rect 24651 2144 24715 2148
rect 22508 1940 22572 2004
rect 22324 1804 22388 1868
rect 3884 1660 3948 1664
rect 3884 1604 3888 1660
rect 3888 1604 3944 1660
rect 3944 1604 3948 1660
rect 3884 1600 3948 1604
rect 3964 1660 4028 1664
rect 3964 1604 3968 1660
rect 3968 1604 4024 1660
rect 4024 1604 4028 1660
rect 3964 1600 4028 1604
rect 4044 1660 4108 1664
rect 4044 1604 4048 1660
rect 4048 1604 4104 1660
rect 4104 1604 4108 1660
rect 4044 1600 4108 1604
rect 4124 1660 4188 1664
rect 4124 1604 4128 1660
rect 4128 1604 4184 1660
rect 4184 1604 4188 1660
rect 4124 1600 4188 1604
rect 9749 1660 9813 1664
rect 9749 1604 9753 1660
rect 9753 1604 9809 1660
rect 9809 1604 9813 1660
rect 9749 1600 9813 1604
rect 9829 1660 9893 1664
rect 9829 1604 9833 1660
rect 9833 1604 9889 1660
rect 9889 1604 9893 1660
rect 9829 1600 9893 1604
rect 9909 1660 9973 1664
rect 9909 1604 9913 1660
rect 9913 1604 9969 1660
rect 9969 1604 9973 1660
rect 9909 1600 9973 1604
rect 9989 1660 10053 1664
rect 9989 1604 9993 1660
rect 9993 1604 10049 1660
rect 10049 1604 10053 1660
rect 9989 1600 10053 1604
rect 15614 1660 15678 1664
rect 15614 1604 15618 1660
rect 15618 1604 15674 1660
rect 15674 1604 15678 1660
rect 15614 1600 15678 1604
rect 15694 1660 15758 1664
rect 15694 1604 15698 1660
rect 15698 1604 15754 1660
rect 15754 1604 15758 1660
rect 15694 1600 15758 1604
rect 15774 1660 15838 1664
rect 15774 1604 15778 1660
rect 15778 1604 15834 1660
rect 15834 1604 15838 1660
rect 15774 1600 15838 1604
rect 15854 1660 15918 1664
rect 15854 1604 15858 1660
rect 15858 1604 15914 1660
rect 15914 1604 15918 1660
rect 15854 1600 15918 1604
rect 21479 1660 21543 1664
rect 21479 1604 21483 1660
rect 21483 1604 21539 1660
rect 21539 1604 21543 1660
rect 21479 1600 21543 1604
rect 21559 1660 21623 1664
rect 21559 1604 21563 1660
rect 21563 1604 21619 1660
rect 21619 1604 21623 1660
rect 21559 1600 21623 1604
rect 21639 1660 21703 1664
rect 21639 1604 21643 1660
rect 21643 1604 21699 1660
rect 21699 1604 21703 1660
rect 21639 1600 21703 1604
rect 21719 1660 21783 1664
rect 21719 1604 21723 1660
rect 21723 1604 21779 1660
rect 21779 1604 21783 1660
rect 21719 1600 21783 1604
rect 6816 1116 6880 1120
rect 6816 1060 6820 1116
rect 6820 1060 6876 1116
rect 6876 1060 6880 1116
rect 6816 1056 6880 1060
rect 6896 1116 6960 1120
rect 6896 1060 6900 1116
rect 6900 1060 6956 1116
rect 6956 1060 6960 1116
rect 6896 1056 6960 1060
rect 6976 1116 7040 1120
rect 6976 1060 6980 1116
rect 6980 1060 7036 1116
rect 7036 1060 7040 1116
rect 6976 1056 7040 1060
rect 7056 1116 7120 1120
rect 7056 1060 7060 1116
rect 7060 1060 7116 1116
rect 7116 1060 7120 1116
rect 7056 1056 7120 1060
rect 12681 1116 12745 1120
rect 12681 1060 12685 1116
rect 12685 1060 12741 1116
rect 12741 1060 12745 1116
rect 12681 1056 12745 1060
rect 12761 1116 12825 1120
rect 12761 1060 12765 1116
rect 12765 1060 12821 1116
rect 12821 1060 12825 1116
rect 12761 1056 12825 1060
rect 12841 1116 12905 1120
rect 12841 1060 12845 1116
rect 12845 1060 12901 1116
rect 12901 1060 12905 1116
rect 12841 1056 12905 1060
rect 12921 1116 12985 1120
rect 12921 1060 12925 1116
rect 12925 1060 12981 1116
rect 12981 1060 12985 1116
rect 12921 1056 12985 1060
rect 18546 1116 18610 1120
rect 18546 1060 18550 1116
rect 18550 1060 18606 1116
rect 18606 1060 18610 1116
rect 18546 1056 18610 1060
rect 18626 1116 18690 1120
rect 18626 1060 18630 1116
rect 18630 1060 18686 1116
rect 18686 1060 18690 1116
rect 18626 1056 18690 1060
rect 18706 1116 18770 1120
rect 18706 1060 18710 1116
rect 18710 1060 18766 1116
rect 18766 1060 18770 1116
rect 18706 1056 18770 1060
rect 18786 1116 18850 1120
rect 18786 1060 18790 1116
rect 18790 1060 18846 1116
rect 18846 1060 18850 1116
rect 18786 1056 18850 1060
rect 24411 1116 24475 1120
rect 24411 1060 24415 1116
rect 24415 1060 24471 1116
rect 24471 1060 24475 1116
rect 24411 1056 24475 1060
rect 24491 1116 24555 1120
rect 24491 1060 24495 1116
rect 24495 1060 24551 1116
rect 24551 1060 24555 1116
rect 24491 1056 24555 1060
rect 24571 1116 24635 1120
rect 24571 1060 24575 1116
rect 24575 1060 24631 1116
rect 24631 1060 24635 1116
rect 24571 1056 24635 1060
rect 24651 1116 24715 1120
rect 24651 1060 24655 1116
rect 24655 1060 24711 1116
rect 24711 1060 24715 1116
rect 24651 1056 24715 1060
<< metal4 >>
rect 3876 8192 4196 8752
rect 3876 8128 3884 8192
rect 3948 8128 3964 8192
rect 4028 8128 4044 8192
rect 4108 8128 4124 8192
rect 4188 8128 4196 8192
rect 3876 7104 4196 8128
rect 3876 7040 3884 7104
rect 3948 7040 3964 7104
rect 4028 7040 4044 7104
rect 4108 7040 4124 7104
rect 4188 7040 4196 7104
rect 3876 6016 4196 7040
rect 3876 5952 3884 6016
rect 3948 5952 3964 6016
rect 4028 5952 4044 6016
rect 4108 5952 4124 6016
rect 4188 5952 4196 6016
rect 3876 4928 4196 5952
rect 3876 4864 3884 4928
rect 3948 4864 3964 4928
rect 4028 4864 4044 4928
rect 4108 4864 4124 4928
rect 4188 4864 4196 4928
rect 3876 3840 4196 4864
rect 3876 3776 3884 3840
rect 3948 3776 3964 3840
rect 4028 3776 4044 3840
rect 4108 3776 4124 3840
rect 4188 3776 4196 3840
rect 3876 2752 4196 3776
rect 3876 2688 3884 2752
rect 3948 2688 3964 2752
rect 4028 2688 4044 2752
rect 4108 2688 4124 2752
rect 4188 2688 4196 2752
rect 3876 1664 4196 2688
rect 3876 1600 3884 1664
rect 3948 1600 3964 1664
rect 4028 1600 4044 1664
rect 4108 1600 4124 1664
rect 4188 1600 4196 1664
rect 3876 1040 4196 1600
rect 6808 8736 7128 8752
rect 6808 8672 6816 8736
rect 6880 8672 6896 8736
rect 6960 8672 6976 8736
rect 7040 8672 7056 8736
rect 7120 8672 7128 8736
rect 6808 7648 7128 8672
rect 6808 7584 6816 7648
rect 6880 7584 6896 7648
rect 6960 7584 6976 7648
rect 7040 7584 7056 7648
rect 7120 7584 7128 7648
rect 6808 6560 7128 7584
rect 6808 6496 6816 6560
rect 6880 6496 6896 6560
rect 6960 6496 6976 6560
rect 7040 6496 7056 6560
rect 7120 6496 7128 6560
rect 6808 5472 7128 6496
rect 6808 5408 6816 5472
rect 6880 5408 6896 5472
rect 6960 5408 6976 5472
rect 7040 5408 7056 5472
rect 7120 5408 7128 5472
rect 6808 4384 7128 5408
rect 6808 4320 6816 4384
rect 6880 4320 6896 4384
rect 6960 4320 6976 4384
rect 7040 4320 7056 4384
rect 7120 4320 7128 4384
rect 6808 3296 7128 4320
rect 6808 3232 6816 3296
rect 6880 3232 6896 3296
rect 6960 3232 6976 3296
rect 7040 3232 7056 3296
rect 7120 3232 7128 3296
rect 6808 2208 7128 3232
rect 6808 2144 6816 2208
rect 6880 2144 6896 2208
rect 6960 2144 6976 2208
rect 7040 2144 7056 2208
rect 7120 2144 7128 2208
rect 6808 1120 7128 2144
rect 6808 1056 6816 1120
rect 6880 1056 6896 1120
rect 6960 1056 6976 1120
rect 7040 1056 7056 1120
rect 7120 1056 7128 1120
rect 6808 1040 7128 1056
rect 9741 8192 10061 8752
rect 9741 8128 9749 8192
rect 9813 8128 9829 8192
rect 9893 8128 9909 8192
rect 9973 8128 9989 8192
rect 10053 8128 10061 8192
rect 9741 7104 10061 8128
rect 9741 7040 9749 7104
rect 9813 7040 9829 7104
rect 9893 7040 9909 7104
rect 9973 7040 9989 7104
rect 10053 7040 10061 7104
rect 9741 6016 10061 7040
rect 9741 5952 9749 6016
rect 9813 5952 9829 6016
rect 9893 5952 9909 6016
rect 9973 5952 9989 6016
rect 10053 5952 10061 6016
rect 9741 4928 10061 5952
rect 9741 4864 9749 4928
rect 9813 4864 9829 4928
rect 9893 4864 9909 4928
rect 9973 4864 9989 4928
rect 10053 4864 10061 4928
rect 9741 3840 10061 4864
rect 9741 3776 9749 3840
rect 9813 3776 9829 3840
rect 9893 3776 9909 3840
rect 9973 3776 9989 3840
rect 10053 3776 10061 3840
rect 9741 2752 10061 3776
rect 9741 2688 9749 2752
rect 9813 2688 9829 2752
rect 9893 2688 9909 2752
rect 9973 2688 9989 2752
rect 10053 2688 10061 2752
rect 9741 1664 10061 2688
rect 9741 1600 9749 1664
rect 9813 1600 9829 1664
rect 9893 1600 9909 1664
rect 9973 1600 9989 1664
rect 10053 1600 10061 1664
rect 9741 1040 10061 1600
rect 12673 8736 12993 8752
rect 12673 8672 12681 8736
rect 12745 8672 12761 8736
rect 12825 8672 12841 8736
rect 12905 8672 12921 8736
rect 12985 8672 12993 8736
rect 12673 7648 12993 8672
rect 15147 8396 15213 8397
rect 15147 8332 15148 8396
rect 15212 8332 15213 8396
rect 15147 8331 15213 8332
rect 12673 7584 12681 7648
rect 12745 7584 12761 7648
rect 12825 7584 12841 7648
rect 12905 7584 12921 7648
rect 12985 7584 12993 7648
rect 12673 6560 12993 7584
rect 15150 6765 15210 8331
rect 15606 8192 15926 8752
rect 15606 8128 15614 8192
rect 15678 8128 15694 8192
rect 15758 8128 15774 8192
rect 15838 8128 15854 8192
rect 15918 8128 15926 8192
rect 15606 7104 15926 8128
rect 15606 7040 15614 7104
rect 15678 7040 15694 7104
rect 15758 7040 15774 7104
rect 15838 7040 15854 7104
rect 15918 7040 15926 7104
rect 15147 6764 15213 6765
rect 15147 6700 15148 6764
rect 15212 6700 15213 6764
rect 15147 6699 15213 6700
rect 12673 6496 12681 6560
rect 12745 6496 12761 6560
rect 12825 6496 12841 6560
rect 12905 6496 12921 6560
rect 12985 6496 12993 6560
rect 12673 5472 12993 6496
rect 12673 5408 12681 5472
rect 12745 5408 12761 5472
rect 12825 5408 12841 5472
rect 12905 5408 12921 5472
rect 12985 5408 12993 5472
rect 12673 4384 12993 5408
rect 12673 4320 12681 4384
rect 12745 4320 12761 4384
rect 12825 4320 12841 4384
rect 12905 4320 12921 4384
rect 12985 4320 12993 4384
rect 12673 3296 12993 4320
rect 12673 3232 12681 3296
rect 12745 3232 12761 3296
rect 12825 3232 12841 3296
rect 12905 3232 12921 3296
rect 12985 3232 12993 3296
rect 12673 2208 12993 3232
rect 12673 2144 12681 2208
rect 12745 2144 12761 2208
rect 12825 2144 12841 2208
rect 12905 2144 12921 2208
rect 12985 2144 12993 2208
rect 12673 1120 12993 2144
rect 12673 1056 12681 1120
rect 12745 1056 12761 1120
rect 12825 1056 12841 1120
rect 12905 1056 12921 1120
rect 12985 1056 12993 1120
rect 12673 1040 12993 1056
rect 15606 6016 15926 7040
rect 15606 5952 15614 6016
rect 15678 5952 15694 6016
rect 15758 5952 15774 6016
rect 15838 5952 15854 6016
rect 15918 5952 15926 6016
rect 15606 4928 15926 5952
rect 15606 4864 15614 4928
rect 15678 4864 15694 4928
rect 15758 4864 15774 4928
rect 15838 4864 15854 4928
rect 15918 4864 15926 4928
rect 15606 3840 15926 4864
rect 15606 3776 15614 3840
rect 15678 3776 15694 3840
rect 15758 3776 15774 3840
rect 15838 3776 15854 3840
rect 15918 3776 15926 3840
rect 15606 2752 15926 3776
rect 15606 2688 15614 2752
rect 15678 2688 15694 2752
rect 15758 2688 15774 2752
rect 15838 2688 15854 2752
rect 15918 2688 15926 2752
rect 15606 1664 15926 2688
rect 15606 1600 15614 1664
rect 15678 1600 15694 1664
rect 15758 1600 15774 1664
rect 15838 1600 15854 1664
rect 15918 1600 15926 1664
rect 15606 1040 15926 1600
rect 18538 8736 18858 8752
rect 18538 8672 18546 8736
rect 18610 8672 18626 8736
rect 18690 8672 18706 8736
rect 18770 8672 18786 8736
rect 18850 8672 18858 8736
rect 18538 7648 18858 8672
rect 18538 7584 18546 7648
rect 18610 7584 18626 7648
rect 18690 7584 18706 7648
rect 18770 7584 18786 7648
rect 18850 7584 18858 7648
rect 18538 6560 18858 7584
rect 18538 6496 18546 6560
rect 18610 6496 18626 6560
rect 18690 6496 18706 6560
rect 18770 6496 18786 6560
rect 18850 6496 18858 6560
rect 18538 5472 18858 6496
rect 18538 5408 18546 5472
rect 18610 5408 18626 5472
rect 18690 5408 18706 5472
rect 18770 5408 18786 5472
rect 18850 5408 18858 5472
rect 18538 4384 18858 5408
rect 18538 4320 18546 4384
rect 18610 4320 18626 4384
rect 18690 4320 18706 4384
rect 18770 4320 18786 4384
rect 18850 4320 18858 4384
rect 18538 3296 18858 4320
rect 18538 3232 18546 3296
rect 18610 3232 18626 3296
rect 18690 3232 18706 3296
rect 18770 3232 18786 3296
rect 18850 3232 18858 3296
rect 18538 2208 18858 3232
rect 18538 2144 18546 2208
rect 18610 2144 18626 2208
rect 18690 2144 18706 2208
rect 18770 2144 18786 2208
rect 18850 2144 18858 2208
rect 18538 1120 18858 2144
rect 18538 1056 18546 1120
rect 18610 1056 18626 1120
rect 18690 1056 18706 1120
rect 18770 1056 18786 1120
rect 18850 1056 18858 1120
rect 18538 1040 18858 1056
rect 21471 8192 21791 8752
rect 24403 8736 24723 8752
rect 24403 8672 24411 8736
rect 24475 8672 24491 8736
rect 24555 8672 24571 8736
rect 24635 8672 24651 8736
rect 24715 8672 24723 8736
rect 22323 8396 22389 8397
rect 22323 8332 22324 8396
rect 22388 8332 22389 8396
rect 22323 8331 22389 8332
rect 22691 8396 22757 8397
rect 22691 8332 22692 8396
rect 22756 8332 22757 8396
rect 22691 8331 22757 8332
rect 21471 8128 21479 8192
rect 21543 8128 21559 8192
rect 21623 8128 21639 8192
rect 21703 8128 21719 8192
rect 21783 8128 21791 8192
rect 21471 7104 21791 8128
rect 22139 7308 22205 7309
rect 22139 7244 22140 7308
rect 22204 7244 22205 7308
rect 22139 7243 22205 7244
rect 21471 7040 21479 7104
rect 21543 7040 21559 7104
rect 21623 7040 21639 7104
rect 21703 7040 21719 7104
rect 21783 7040 21791 7104
rect 21471 6016 21791 7040
rect 21471 5952 21479 6016
rect 21543 5952 21559 6016
rect 21623 5952 21639 6016
rect 21703 5952 21719 6016
rect 21783 5952 21791 6016
rect 21471 4928 21791 5952
rect 21471 4864 21479 4928
rect 21543 4864 21559 4928
rect 21623 4864 21639 4928
rect 21703 4864 21719 4928
rect 21783 4864 21791 4928
rect 21471 3840 21791 4864
rect 21471 3776 21479 3840
rect 21543 3776 21559 3840
rect 21623 3776 21639 3840
rect 21703 3776 21719 3840
rect 21783 3776 21791 3840
rect 21471 2752 21791 3776
rect 21471 2688 21479 2752
rect 21543 2688 21559 2752
rect 21623 2688 21639 2752
rect 21703 2688 21719 2752
rect 21783 2688 21791 2752
rect 21471 1664 21791 2688
rect 22142 2413 22202 7243
rect 22139 2412 22205 2413
rect 22139 2348 22140 2412
rect 22204 2348 22205 2412
rect 22139 2347 22205 2348
rect 22326 1869 22386 8331
rect 22694 6930 22754 8331
rect 22510 6870 22754 6930
rect 24403 7648 24723 8672
rect 24403 7584 24411 7648
rect 24475 7584 24491 7648
rect 24555 7584 24571 7648
rect 24635 7584 24651 7648
rect 24715 7584 24723 7648
rect 22510 2005 22570 6870
rect 24403 6560 24723 7584
rect 24403 6496 24411 6560
rect 24475 6496 24491 6560
rect 24555 6496 24571 6560
rect 24635 6496 24651 6560
rect 24715 6496 24723 6560
rect 24403 5472 24723 6496
rect 24403 5408 24411 5472
rect 24475 5408 24491 5472
rect 24555 5408 24571 5472
rect 24635 5408 24651 5472
rect 24715 5408 24723 5472
rect 24403 4384 24723 5408
rect 24403 4320 24411 4384
rect 24475 4320 24491 4384
rect 24555 4320 24571 4384
rect 24635 4320 24651 4384
rect 24715 4320 24723 4384
rect 24403 3296 24723 4320
rect 24403 3232 24411 3296
rect 24475 3232 24491 3296
rect 24555 3232 24571 3296
rect 24635 3232 24651 3296
rect 24715 3232 24723 3296
rect 24403 2208 24723 3232
rect 24403 2144 24411 2208
rect 24475 2144 24491 2208
rect 24555 2144 24571 2208
rect 24635 2144 24651 2208
rect 24715 2144 24723 2208
rect 22507 2004 22573 2005
rect 22507 1940 22508 2004
rect 22572 1940 22573 2004
rect 22507 1939 22573 1940
rect 22323 1868 22389 1869
rect 22323 1804 22324 1868
rect 22388 1804 22389 1868
rect 22323 1803 22389 1804
rect 21471 1600 21479 1664
rect 21543 1600 21559 1664
rect 21623 1600 21639 1664
rect 21703 1600 21719 1664
rect 21783 1600 21791 1664
rect 21471 1040 21791 1600
rect 24403 1120 24723 2144
rect 24403 1056 24411 1120
rect 24475 1056 24491 1120
rect 24555 1056 24571 1120
rect 24635 1056 24651 1120
rect 24715 1056 24723 1120
rect 24403 1040 24723 1056
use sky130_fd_sc_hd__diode_2  ANTENNA_1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 1748 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_6 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1656 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_10 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2024 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_14 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2392 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_22 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3128 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27
timestamp 1688980957
transform 1 0 3588 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_29
timestamp 1688980957
transform 1 0 3772 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_40
timestamp 1688980957
transform 1 0 4784 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_48
timestamp 1688980957
transform 1 0 5520 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_53 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5980 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_57
timestamp 1688980957
transform 1 0 6348 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_71 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 7636 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_77
timestamp 1688980957
transform 1 0 8188 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_85
timestamp 1688980957
transform 1 0 8924 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_92
timestamp 1688980957
transform 1 0 9568 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_99
timestamp 1688980957
transform 1 0 10212 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_111
timestamp 1688980957
transform 1 0 11316 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_113
timestamp 1688980957
transform 1 0 11500 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_121
timestamp 1688980957
transform 1 0 12236 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_125
timestamp 1688980957
transform 1 0 12604 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_133
timestamp 1688980957
transform 1 0 13340 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_138
timestamp 1688980957
transform 1 0 13800 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_147
timestamp 1688980957
transform 1 0 14628 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_153
timestamp 1688980957
transform 1 0 15180 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_160
timestamp 1688980957
transform 1 0 15824 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_172
timestamp 1688980957
transform 1 0 16928 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_183
timestamp 1688980957
transform 1 0 17940 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_191
timestamp 1688980957
transform 1 0 18676 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_197
timestamp 1688980957
transform 1 0 19228 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_205
timestamp 1688980957
transform 1 0 19964 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_209
timestamp 1688980957
transform 1 0 20332 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_217
timestamp 1688980957
transform 1 0 21068 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_222
timestamp 1688980957
transform 1 0 21528 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_228
timestamp 1688980957
transform 1 0 22080 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_235
timestamp 1688980957
transform 1 0 22724 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_251
timestamp 1688980957
transform 1 0 24196 0 1 1088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1380 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 1688980957
transform 1 0 2484 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_27
timestamp 1688980957
transform 1 0 3588 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_39
timestamp 1688980957
transform 1 0 4692 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_51
timestamp 1688980957
transform 1 0 5796 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 1688980957
transform 1 0 6164 0 -1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_57
timestamp 1688980957
transform 1 0 6348 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_69
timestamp 1688980957
transform 1 0 7452 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_74
timestamp 1688980957
transform 1 0 7912 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_82
timestamp 1688980957
transform 1 0 8648 0 -1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_87
timestamp 1688980957
transform 1 0 9108 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_105
timestamp 1688980957
transform 1 0 10764 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_111
timestamp 1688980957
transform 1 0 11316 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_119
timestamp 1688980957
transform 1 0 12052 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_126
timestamp 1688980957
transform 1 0 12696 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_130
timestamp 1688980957
transform 1 0 13064 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_139
timestamp 1688980957
transform 1 0 13892 0 -1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_144
timestamp 1688980957
transform 1 0 14352 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_156
timestamp 1688980957
transform 1 0 15456 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_162
timestamp 1688980957
transform 1 0 16008 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_166
timestamp 1688980957
transform 1 0 16376 0 -1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_169
timestamp 1688980957
transform 1 0 16652 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_181
timestamp 1688980957
transform 1 0 17756 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_193
timestamp 1688980957
transform 1 0 18860 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_205
timestamp 1688980957
transform 1 0 19964 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_217
timestamp 1688980957
transform 1 0 21068 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_223
timestamp 1688980957
transform 1 0 21620 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_225
timestamp 1688980957
transform 1 0 21804 0 -1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_230
timestamp 1688980957
transform 1 0 22264 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_251
timestamp 1688980957
transform 1 0 24196 0 -1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1688980957
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 1688980957
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1688980957
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 1688980957
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 1688980957
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_53
timestamp 1688980957
transform 1 0 5980 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_65
timestamp 1688980957
transform 1 0 7084 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_77
timestamp 1688980957
transform 1 0 8188 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 1688980957
transform 1 0 8740 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_85
timestamp 1688980957
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_97
timestamp 1688980957
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_109
timestamp 1688980957
transform 1 0 11132 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_121
timestamp 1688980957
transform 1 0 12236 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_133
timestamp 1688980957
transform 1 0 13340 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_139
timestamp 1688980957
transform 1 0 13892 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_141
timestamp 1688980957
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_153
timestamp 1688980957
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_165
timestamp 1688980957
transform 1 0 16284 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_177
timestamp 1688980957
transform 1 0 17388 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_189
timestamp 1688980957
transform 1 0 18492 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_195
timestamp 1688980957
transform 1 0 19044 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_197
timestamp 1688980957
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_209
timestamp 1688980957
transform 1 0 20332 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_221
timestamp 1688980957
transform 1 0 21436 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_233
timestamp 1688980957
transform 1 0 22540 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_245
timestamp 1688980957
transform 1 0 23644 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_250
timestamp 1688980957
transform 1 0 24104 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1688980957
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1688980957
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 1688980957
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 1688980957
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 1688980957
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1688980957
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 1688980957
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_69
timestamp 1688980957
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_81
timestamp 1688980957
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_93
timestamp 1688980957
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_105
timestamp 1688980957
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_111
timestamp 1688980957
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_113
timestamp 1688980957
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_125
timestamp 1688980957
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_137
timestamp 1688980957
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_149
timestamp 1688980957
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_161
timestamp 1688980957
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_167
timestamp 1688980957
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_169
timestamp 1688980957
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_181
timestamp 1688980957
transform 1 0 17756 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_193
timestamp 1688980957
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_205
timestamp 1688980957
transform 1 0 19964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_217
timestamp 1688980957
transform 1 0 21068 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_223
timestamp 1688980957
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_225
timestamp 1688980957
transform 1 0 21804 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_233
timestamp 1688980957
transform 1 0 22540 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_238
timestamp 1688980957
transform 1 0 23000 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_244
timestamp 1688980957
transform 1 0 23552 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_250
timestamp 1688980957
transform 1 0 24104 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1688980957
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 1688980957
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1688980957
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 1688980957
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 1688980957
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_53
timestamp 1688980957
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_65
timestamp 1688980957
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_77
timestamp 1688980957
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp 1688980957
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_85
timestamp 1688980957
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_97
timestamp 1688980957
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_109
timestamp 1688980957
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_121
timestamp 1688980957
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_133
timestamp 1688980957
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_139
timestamp 1688980957
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_141
timestamp 1688980957
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_153
timestamp 1688980957
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_165
timestamp 1688980957
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_177
timestamp 1688980957
transform 1 0 17388 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_181
timestamp 1688980957
transform 1 0 17756 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_185
timestamp 1688980957
transform 1 0 18124 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_193
timestamp 1688980957
transform 1 0 18860 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_197
timestamp 1688980957
transform 1 0 19228 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_209
timestamp 1688980957
transform 1 0 20332 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_221
timestamp 1688980957
transform 1 0 21436 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_233
timestamp 1688980957
transform 1 0 22540 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_244
timestamp 1688980957
transform 1 0 23552 0 1 3264
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 1688980957
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 1688980957
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_27
timestamp 1688980957
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_39
timestamp 1688980957
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_51
timestamp 1688980957
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 1688980957
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_57
timestamp 1688980957
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_69
timestamp 1688980957
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_81
timestamp 1688980957
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_93
timestamp 1688980957
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_105
timestamp 1688980957
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_111
timestamp 1688980957
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_113
timestamp 1688980957
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_125
timestamp 1688980957
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_137
timestamp 1688980957
transform 1 0 13708 0 -1 4352
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_146
timestamp 1688980957
transform 1 0 14536 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_158
timestamp 1688980957
transform 1 0 15640 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_166
timestamp 1688980957
transform 1 0 16376 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_169
timestamp 1688980957
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_181
timestamp 1688980957
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_193
timestamp 1688980957
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_205
timestamp 1688980957
transform 1 0 19964 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_217
timestamp 1688980957
transform 1 0 21068 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_223
timestamp 1688980957
transform 1 0 21620 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_225
timestamp 1688980957
transform 1 0 21804 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_237
timestamp 1688980957
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_249
timestamp 1688980957
transform 1 0 24012 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 1688980957
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_15
timestamp 1688980957
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1688980957
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 1688980957
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_41
timestamp 1688980957
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_53
timestamp 1688980957
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_65
timestamp 1688980957
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_77
timestamp 1688980957
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_83
timestamp 1688980957
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_85
timestamp 1688980957
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_97
timestamp 1688980957
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_109
timestamp 1688980957
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_121
timestamp 1688980957
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_133
timestamp 1688980957
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_139
timestamp 1688980957
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_141
timestamp 1688980957
transform 1 0 14076 0 1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_152
timestamp 1688980957
transform 1 0 15088 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_164
timestamp 1688980957
transform 1 0 16192 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_176
timestamp 1688980957
transform 1 0 17296 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_188
timestamp 1688980957
transform 1 0 18400 0 1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_197
timestamp 1688980957
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_209
timestamp 1688980957
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_221
timestamp 1688980957
transform 1 0 21436 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_233
timestamp 1688980957
transform 1 0 22540 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_245
timestamp 1688980957
transform 1 0 23644 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_251
timestamp 1688980957
transform 1 0 24196 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 1688980957
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 1688980957
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_27
timestamp 1688980957
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_39
timestamp 1688980957
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_51
timestamp 1688980957
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 1688980957
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_57
timestamp 1688980957
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_69
timestamp 1688980957
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_81
timestamp 1688980957
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_93
timestamp 1688980957
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_105
timestamp 1688980957
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_111
timestamp 1688980957
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_113
timestamp 1688980957
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_125
timestamp 1688980957
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_137
timestamp 1688980957
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_149
timestamp 1688980957
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_161
timestamp 1688980957
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_167
timestamp 1688980957
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_169
timestamp 1688980957
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_181
timestamp 1688980957
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_193
timestamp 1688980957
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_205
timestamp 1688980957
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_217
timestamp 1688980957
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_223
timestamp 1688980957
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_225
timestamp 1688980957
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_237
timestamp 1688980957
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_249
timestamp 1688980957
transform 1 0 24012 0 -1 5440
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 1688980957
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 1688980957
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1688980957
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 1688980957
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_41
timestamp 1688980957
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_53
timestamp 1688980957
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_65
timestamp 1688980957
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_77
timestamp 1688980957
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_83
timestamp 1688980957
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_85
timestamp 1688980957
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_97
timestamp 1688980957
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_109
timestamp 1688980957
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_121
timestamp 1688980957
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_133
timestamp 1688980957
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_139
timestamp 1688980957
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_141
timestamp 1688980957
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_153
timestamp 1688980957
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_165
timestamp 1688980957
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_177
timestamp 1688980957
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_189
timestamp 1688980957
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_195
timestamp 1688980957
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_197
timestamp 1688980957
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_209
timestamp 1688980957
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_221
timestamp 1688980957
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_233
timestamp 1688980957
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_245
timestamp 1688980957
transform 1 0 23644 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_9
timestamp 1688980957
transform 1 0 1932 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_21
timestamp 1688980957
transform 1 0 3036 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_33
timestamp 1688980957
transform 1 0 4140 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_45
timestamp 1688980957
transform 1 0 5244 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_53
timestamp 1688980957
transform 1 0 5980 0 -1 6528
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_57
timestamp 1688980957
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_69
timestamp 1688980957
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_81
timestamp 1688980957
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_93
timestamp 1688980957
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_105
timestamp 1688980957
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_111
timestamp 1688980957
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_113
timestamp 1688980957
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_125
timestamp 1688980957
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_137
timestamp 1688980957
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_149
timestamp 1688980957
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_161
timestamp 1688980957
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_167
timestamp 1688980957
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_169
timestamp 1688980957
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_181
timestamp 1688980957
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_193
timestamp 1688980957
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_205
timestamp 1688980957
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_217
timestamp 1688980957
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_223
timestamp 1688980957
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_225
timestamp 1688980957
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_237
timestamp 1688980957
transform 1 0 22908 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_251
timestamp 1688980957
transform 1 0 24196 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_3
timestamp 1688980957
transform 1 0 1380 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_7
timestamp 1688980957
transform 1 0 1748 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_15
timestamp 1688980957
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 1688980957
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_29
timestamp 1688980957
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_41
timestamp 1688980957
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_53
timestamp 1688980957
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_65
timestamp 1688980957
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_77
timestamp 1688980957
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_83
timestamp 1688980957
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_85
timestamp 1688980957
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_97
timestamp 1688980957
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_109
timestamp 1688980957
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_121
timestamp 1688980957
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_133
timestamp 1688980957
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_139
timestamp 1688980957
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_141
timestamp 1688980957
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_153
timestamp 1688980957
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_165
timestamp 1688980957
transform 1 0 16284 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_172
timestamp 1688980957
transform 1 0 16928 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_184
timestamp 1688980957
transform 1 0 18032 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_197
timestamp 1688980957
transform 1 0 19228 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_209
timestamp 1688980957
transform 1 0 20332 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_221
timestamp 1688980957
transform 1 0 21436 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_233
timestamp 1688980957
transform 1 0 22540 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_237
timestamp 1688980957
transform 1 0 22908 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_250
timestamp 1688980957
transform 1 0 24104 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_3
timestamp 1688980957
transform 1 0 1380 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_22
timestamp 1688980957
transform 1 0 3128 0 -1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_28
timestamp 1688980957
transform 1 0 3680 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_40
timestamp 1688980957
transform 1 0 4784 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_46
timestamp 1688980957
transform 1 0 5336 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_50
timestamp 1688980957
transform 1 0 5704 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_60
timestamp 1688980957
transform 1 0 6624 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_69
timestamp 1688980957
transform 1 0 7452 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_74
timestamp 1688980957
transform 1 0 7912 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_84
timestamp 1688980957
transform 1 0 8832 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_96
timestamp 1688980957
transform 1 0 9936 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_101
timestamp 1688980957
transform 1 0 10396 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_109
timestamp 1688980957
transform 1 0 11132 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_113
timestamp 1688980957
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_125
timestamp 1688980957
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_137
timestamp 1688980957
transform 1 0 13708 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_149
timestamp 1688980957
transform 1 0 14812 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_161
timestamp 1688980957
transform 1 0 15916 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_167
timestamp 1688980957
transform 1 0 16468 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_169
timestamp 1688980957
transform 1 0 16652 0 -1 7616
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_178
timestamp 1688980957
transform 1 0 17480 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_190
timestamp 1688980957
transform 1 0 18584 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_202
timestamp 1688980957
transform 1 0 19688 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_214
timestamp 1688980957
transform 1 0 20792 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_222
timestamp 1688980957
transform 1 0 21528 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_225
timestamp 1688980957
transform 1 0 21804 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_249
timestamp 1688980957
transform 1 0 24012 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 1688980957
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_29
timestamp 1688980957
transform 1 0 3772 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_46
timestamp 1688980957
transform 1 0 5336 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_70
timestamp 1688980957
transform 1 0 7544 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_78
timestamp 1688980957
transform 1 0 8280 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_85
timestamp 1688980957
transform 1 0 8924 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_116
timestamp 1688980957
transform 1 0 11776 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_134
timestamp 1688980957
transform 1 0 13432 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_141
timestamp 1688980957
transform 1 0 14076 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_145
timestamp 1688980957
transform 1 0 14444 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_167
timestamp 1688980957
transform 1 0 16468 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_173
timestamp 1688980957
transform 1 0 17020 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_179
timestamp 1688980957
transform 1 0 17572 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_191
timestamp 1688980957
transform 1 0 18676 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_206
timestamp 1688980957
transform 1 0 20056 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_214
timestamp 1688980957
transform 1 0 20792 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_251
timestamp 1688980957
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_3
timestamp 1688980957
transform 1 0 1380 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_26
timestamp 1688980957
transform 1 0 3496 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_29
timestamp 1688980957
transform 1 0 3772 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_57
timestamp 1688980957
transform 1 0 6348 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_64
timestamp 1688980957
transform 1 0 6992 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_85
timestamp 1688980957
transform 1 0 8924 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_222
timestamp 1688980957
transform 1 0 21528 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_249
timestamp 1688980957
transform 1 0 24012 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2116 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14076 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1688980957
transform 1 0 15272 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1688980957
transform 1 0 16652 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1688980957
transform 1 0 17664 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1688980957
transform 1 0 18860 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1688980957
transform 1 0 20056 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1688980957
transform 1 0 21252 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1688980957
transform 1 0 22448 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1688980957
transform 1 0 23920 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1688980957
transform 1 0 23368 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input12
timestamp 1688980957
transform 1 0 3312 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input13
timestamp 1688980957
transform 1 0 4508 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input14
timestamp 1688980957
transform 1 0 5704 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input15
timestamp 1688980957
transform 1 0 7360 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1688980957
transform 1 0 8556 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1688980957
transform 1 0 9292 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1688980957
transform 1 0 10488 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1688980957
transform 1 0 11684 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1688980957
transform 1 0 12788 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1688980957
transform 1 0 10120 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1688980957
transform 1 0 10396 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1688980957
transform 1 0 10672 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 1688980957
transform 1 0 10948 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1688980957
transform 1 0 11224 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 1688980957
transform 1 0 11500 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1688980957
transform 1 0 11500 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1688980957
transform 1 0 12052 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1688980957
transform 1 0 12328 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1688980957
transform 1 0 12604 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1688980957
transform 1 0 12880 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 1688980957
transform 1 0 13156 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1688980957
transform 1 0 13156 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input34
timestamp 1688980957
transform 1 0 13708 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input35
timestamp 1688980957
transform 1 0 14076 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input36
timestamp 1688980957
transform 1 0 14904 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 1688980957
transform 1 0 14536 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input38
timestamp 1688980957
transform 1 0 14812 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input39
timestamp 1688980957
transform 1 0 15088 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input40
timestamp 1688980957
transform 1 0 15364 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input41
timestamp 1688980957
transform 1 0 15640 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input42
timestamp 1688980957
transform 1 0 19228 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input43
timestamp 1688980957
transform 1 0 19504 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input44
timestamp 1688980957
transform 1 0 19780 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input45
timestamp 1688980957
transform 1 0 19228 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input46
timestamp 1688980957
transform 1 0 19504 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input47
timestamp 1688980957
transform 1 0 19780 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input48
timestamp 1688980957
transform 1 0 15916 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input49
timestamp 1688980957
transform 1 0 16192 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input50
timestamp 1688980957
transform 1 0 17204 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input51
timestamp 1688980957
transform 1 0 16744 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input52
timestamp 1688980957
transform 1 0 17756 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input53
timestamp 1688980957
transform 1 0 17296 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input54
timestamp 1688980957
transform 1 0 18308 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input55
timestamp 1688980957
transform 1 0 17848 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input56
timestamp 1688980957
transform 1 0 18124 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input57
timestamp 1688980957
transform 1 0 1380 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  inst_clk_buf
timestamp 1688980957
transform 1 0 14352 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_RAM_IO_switch_matrix__00_
timestamp 1688980957
transform 1 0 9844 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_RAM_IO_switch_matrix__01_
timestamp 1688980957
transform 1 0 9016 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_RAM_IO_switch_matrix__02_
timestamp 1688980957
transform 1 0 7176 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_RAM_IO_switch_matrix__03_
timestamp 1688980957
transform 1 0 9292 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_RAM_IO_switch_matrix__04_
timestamp 1688980957
transform 1 0 15732 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_RAM_IO_switch_matrix__05_
timestamp 1688980957
transform 1 0 15456 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_RAM_IO_switch_matrix__06_
timestamp 1688980957
transform 1 0 15180 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_RAM_IO_switch_matrix__07_
timestamp 1688980957
transform 1 0 14628 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_RAM_IO_switch_matrix__08_
timestamp 1688980957
transform 1 0 14352 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_RAM_IO_switch_matrix__09_
timestamp 1688980957
transform 1 0 13432 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_RAM_IO_switch_matrix__10_
timestamp 1688980957
transform 1 0 12880 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_RAM_IO_switch_matrix__11_
timestamp 1688980957
transform 1 0 12604 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_RAM_IO_switch_matrix__12_
timestamp 1688980957
transform 1 0 12328 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_RAM_IO_switch_matrix__13_
timestamp 1688980957
transform 1 0 12052 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_RAM_IO_switch_matrix__14_
timestamp 1688980957
transform 1 0 11776 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_RAM_IO_switch_matrix__15_
timestamp 1688980957
transform 1 0 11132 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_RAM_IO_switch_matrix__16_
timestamp 1688980957
transform 1 0 10856 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_RAM_IO_switch_matrix__17_
timestamp 1688980957
transform 1 0 10580 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_RAM_IO_switch_matrix__18_
timestamp 1688980957
transform 1 0 10120 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_RAM_IO_switch_matrix__19_
timestamp 1688980957
transform 1 0 9568 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_RAM_IO_switch_matrix__20_
timestamp 1688980957
transform 1 0 5428 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_RAM_IO_switch_matrix__21_
timestamp 1688980957
transform 1 0 5980 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_RAM_IO_switch_matrix__22_
timestamp 1688980957
transform 1 0 17480 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_RAM_IO_switch_matrix__23_
timestamp 1688980957
transform 1 0 8556 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_RAM_IO_switch_matrix__24_
timestamp 1688980957
transform 1 0 16928 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_RAM_IO_switch_matrix__25_
timestamp 1688980957
transform 1 0 16652 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_RAM_IO_switch_matrix__26_
timestamp 1688980957
transform 1 0 16284 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_RAM_IO_switch_matrix__27_
timestamp 1688980957
transform 1 0 16008 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_RAM_IO_switch_matrix__28_
timestamp 1688980957
transform 1 0 18860 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_RAM_IO_switch_matrix__29_
timestamp 1688980957
transform 1 0 6348 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_RAM_IO_switch_matrix__30_
timestamp 1688980957
transform 1 0 18400 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_RAM_IO_switch_matrix__31_
timestamp 1688980957
transform 1 0 18860 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_RAM_IO_switch_matrix__32_
timestamp 1688980957
transform 1 0 18584 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_RAM_IO_switch_matrix__33_
timestamp 1688980957
transform 1 0 7636 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_RAM_IO_switch_matrix__34_
timestamp 1688980957
transform 1 0 18032 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_RAM_IO_switch_matrix__35_
timestamp 1688980957
transform 1 0 8280 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  output58 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 20424 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output59
timestamp 1688980957
transform 1 0 23460 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output60
timestamp 1688980957
transform 1 0 23092 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output61
timestamp 1688980957
transform 1 0 23644 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output62
timestamp 1688980957
transform 1 0 23000 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output63
timestamp 1688980957
transform 1 0 23460 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output64
timestamp 1688980957
transform 1 0 23552 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output65
timestamp 1688980957
transform 1 0 22908 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output66
timestamp 1688980957
transform 1 0 22356 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output67
timestamp 1688980957
transform 1 0 23736 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output68
timestamp 1688980957
transform 1 0 21436 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output69
timestamp 1688980957
transform 1 0 20976 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output70 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 21068 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output71
timestamp 1688980957
transform 1 0 21804 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output72
timestamp 1688980957
transform 1 0 22356 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output73
timestamp 1688980957
transform 1 0 22908 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output74
timestamp 1688980957
transform 1 0 21988 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output75
timestamp 1688980957
transform 1 0 22540 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output76
timestamp 1688980957
transform 1 0 23092 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output77
timestamp 1688980957
transform 1 0 23644 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output78
timestamp 1688980957
transform 1 0 2944 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output79
timestamp 1688980957
transform 1 0 1840 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output80
timestamp 1688980957
transform 1 0 2576 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output81
timestamp 1688980957
transform 1 0 1380 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output82
timestamp 1688980957
transform -1 0 2484 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output83
timestamp 1688980957
transform 1 0 2024 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output84
timestamp 1688980957
transform 1 0 1472 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output85
timestamp 1688980957
transform 1 0 1380 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output86
timestamp 1688980957
transform 1 0 1932 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output87
timestamp 1688980957
transform 1 0 2484 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output88
timestamp 1688980957
transform 1 0 2392 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output89
timestamp 1688980957
transform 1 0 3036 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output90
timestamp 1688980957
transform 1 0 1472 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output91
timestamp 1688980957
transform 1 0 3312 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output92
timestamp 1688980957
transform 1 0 3864 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output93
timestamp 1688980957
transform 1 0 3864 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output94
timestamp 1688980957
transform 1 0 4416 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output95
timestamp 1688980957
transform 1 0 4968 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output96
timestamp 1688980957
transform 1 0 4416 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output97
timestamp 1688980957
transform 1 0 4784 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output98
timestamp 1688980957
transform 1 0 5520 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output99
timestamp 1688980957
transform 1 0 7912 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output100
timestamp 1688980957
transform 1 0 8464 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output101
timestamp 1688980957
transform 1 0 8464 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output102
timestamp 1688980957
transform 1 0 9108 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output103
timestamp 1688980957
transform 1 0 10028 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output104
timestamp 1688980957
transform 1 0 9476 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output105
timestamp 1688980957
transform 1 0 5336 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output106
timestamp 1688980957
transform 1 0 6072 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output107
timestamp 1688980957
transform 1 0 5888 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output108
timestamp 1688980957
transform 1 0 6624 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output109
timestamp 1688980957
transform 1 0 6440 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output110
timestamp 1688980957
transform 1 0 7176 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output111
timestamp 1688980957
transform 1 0 7176 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output112
timestamp 1688980957
transform 1 0 7728 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output113
timestamp 1688980957
transform 1 0 7544 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output114
timestamp 1688980957
transform 1 0 20056 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1688980957
transform 1 0 1104 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1688980957
transform -1 0 24564 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1688980957
transform 1 0 1104 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1688980957
transform -1 0 24564 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1688980957
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1688980957
transform -1 0 24564 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1688980957
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1688980957
transform -1 0 24564 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1688980957
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1688980957
transform -1 0 24564 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1688980957
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1688980957
transform -1 0 24564 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1688980957
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1688980957
transform -1 0 24564 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1688980957
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1688980957
transform -1 0 24564 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1688980957
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1688980957
transform -1 0 24564 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1688980957
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1688980957
transform -1 0 24564 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1688980957
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1688980957
transform -1 0 24564 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1688980957
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1688980957
transform -1 0 24564 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1688980957
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1688980957
transform -1 0 24564 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1688980957
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1688980957
transform -1 0 24564 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_0__0_
timestamp 1688980957
transform 1 0 11040 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_1__0_
timestamp 1688980957
transform 1 0 13524 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_2__0_
timestamp 1688980957
transform 1 0 12328 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_3__0_
timestamp 1688980957
transform 1 0 9660 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_4__0_
timestamp 1688980957
transform 1 0 7084 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_5__0_
timestamp 1688980957
transform 1 0 8280 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_6__0_
timestamp 1688980957
transform 1 0 9936 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_7__0_
timestamp 1688980957
transform 1 0 10764 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_8__0_
timestamp 1688980957
transform 1 0 11960 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_9__0_
timestamp 1688980957
transform 1 0 13064 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_10__0_
timestamp 1688980957
transform 1 0 14260 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_11__0_
timestamp 1688980957
transform 1 0 15548 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_12__0_
timestamp 1688980957
transform 1 0 16652 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_13__0_
timestamp 1688980957
transform 1 0 17848 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_14__0_
timestamp 1688980957
transform 1 0 23092 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_15__0_
timestamp 1688980957
transform 1 0 22816 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_16__0_
timestamp 1688980957
transform 1 0 21804 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_17__0_
timestamp 1688980957
transform 1 0 22724 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_18__0_
timestamp 1688980957
transform 1 0 23644 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_19__0_
timestamp 1688980957
transform 1 0 23828 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  strobe_outbuf_0__0_
timestamp 1688980957
transform 1 0 11500 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  strobe_outbuf_1__0_
timestamp 1688980957
transform 1 0 14076 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  strobe_outbuf_2__0_
timestamp 1688980957
transform 1 0 12788 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  strobe_outbuf_3__0_
timestamp 1688980957
transform 1 0 10212 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  strobe_outbuf_4__0_
timestamp 1688980957
transform 1 0 7636 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  strobe_outbuf_5__0_
timestamp 1688980957
transform 1 0 8832 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  strobe_outbuf_6__0_
timestamp 1688980957
transform 1 0 10488 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  strobe_outbuf_7__0_
timestamp 1688980957
transform 1 0 11776 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  strobe_outbuf_8__0_
timestamp 1688980957
transform 1 0 12420 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  strobe_outbuf_9__0_
timestamp 1688980957
transform 1 0 13616 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  strobe_outbuf_10__0_
timestamp 1688980957
transform 1 0 14812 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  strobe_outbuf_11__0_
timestamp 1688980957
transform 1 0 16100 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_12__0_
timestamp 1688980957
transform 1 0 17204 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_13__0_
timestamp 1688980957
transform 1 0 23276 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_14__0_
timestamp 1688980957
transform 1 0 23644 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_15__0_
timestamp 1688980957
transform 1 0 23368 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_16__0_
timestamp 1688980957
transform 1 0 21988 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_17__0_
timestamp 1688980957
transform 1 0 23276 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_18__0_
timestamp 1688980957
transform 1 0 23920 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_19__0_
timestamp 1688980957
transform 1 0 23828 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_28 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3680 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_29
timestamp 1688980957
transform 1 0 6256 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_30
timestamp 1688980957
transform 1 0 8832 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_31
timestamp 1688980957
transform 1 0 11408 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_32
timestamp 1688980957
transform 1 0 13984 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_33
timestamp 1688980957
transform 1 0 16560 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_34
timestamp 1688980957
transform 1 0 19136 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_35
timestamp 1688980957
transform 1 0 21712 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_36
timestamp 1688980957
transform 1 0 6256 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_37
timestamp 1688980957
transform 1 0 11408 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_38
timestamp 1688980957
transform 1 0 16560 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_39
timestamp 1688980957
transform 1 0 21712 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_40
timestamp 1688980957
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_41
timestamp 1688980957
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_42
timestamp 1688980957
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_43
timestamp 1688980957
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_44
timestamp 1688980957
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_45
timestamp 1688980957
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_46
timestamp 1688980957
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_47
timestamp 1688980957
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_48
timestamp 1688980957
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_49
timestamp 1688980957
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_50
timestamp 1688980957
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_51
timestamp 1688980957
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_52
timestamp 1688980957
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_53
timestamp 1688980957
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_54
timestamp 1688980957
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_55
timestamp 1688980957
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56
timestamp 1688980957
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1688980957
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1688980957
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1688980957
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1688980957
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1688980957
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1688980957
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1688980957
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1688980957
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1688980957
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 1688980957
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 1688980957
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 1688980957
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1688980957
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1688980957
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1688980957
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1688980957
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1688980957
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1688980957
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1688980957
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1688980957
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1688980957
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1688980957
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1688980957
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1688980957
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1688980957
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1688980957
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1688980957
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1688980957
transform 1 0 3680 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1688980957
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1688980957
transform 1 0 8832 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1688980957
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1688980957
transform 1 0 13984 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1688980957
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1688980957
transform 1 0 19136 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1688980957
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
<< labels >>
flabel metal2 s 2042 -300 2098 160 0 FreeSans 224 90 0 0 FrameStrobe[0]
port 0 nsew signal input
flabel metal2 s 14002 -300 14058 160 0 FreeSans 224 90 0 0 FrameStrobe[10]
port 1 nsew signal input
flabel metal2 s 15198 -300 15254 160 0 FreeSans 224 90 0 0 FrameStrobe[11]
port 2 nsew signal input
flabel metal2 s 16394 -300 16450 160 0 FreeSans 224 90 0 0 FrameStrobe[12]
port 3 nsew signal input
flabel metal2 s 17590 -300 17646 160 0 FreeSans 224 90 0 0 FrameStrobe[13]
port 4 nsew signal input
flabel metal2 s 18786 -300 18842 160 0 FreeSans 224 90 0 0 FrameStrobe[14]
port 5 nsew signal input
flabel metal2 s 19982 -300 20038 160 0 FreeSans 224 90 0 0 FrameStrobe[15]
port 6 nsew signal input
flabel metal2 s 21178 -300 21234 160 0 FreeSans 224 90 0 0 FrameStrobe[16]
port 7 nsew signal input
flabel metal2 s 22374 -300 22430 160 0 FreeSans 224 90 0 0 FrameStrobe[17]
port 8 nsew signal input
flabel metal2 s 23570 -300 23626 160 0 FreeSans 224 90 0 0 FrameStrobe[18]
port 9 nsew signal input
flabel metal2 s 24766 -300 24822 160 0 FreeSans 224 90 0 0 FrameStrobe[19]
port 10 nsew signal input
flabel metal2 s 3238 -300 3294 160 0 FreeSans 224 90 0 0 FrameStrobe[1]
port 11 nsew signal input
flabel metal2 s 4434 -300 4490 160 0 FreeSans 224 90 0 0 FrameStrobe[2]
port 12 nsew signal input
flabel metal2 s 5630 -300 5686 160 0 FreeSans 224 90 0 0 FrameStrobe[3]
port 13 nsew signal input
flabel metal2 s 6826 -300 6882 160 0 FreeSans 224 90 0 0 FrameStrobe[4]
port 14 nsew signal input
flabel metal2 s 8022 -300 8078 160 0 FreeSans 224 90 0 0 FrameStrobe[5]
port 15 nsew signal input
flabel metal2 s 9218 -300 9274 160 0 FreeSans 224 90 0 0 FrameStrobe[6]
port 16 nsew signal input
flabel metal2 s 10414 -300 10470 160 0 FreeSans 224 90 0 0 FrameStrobe[7]
port 17 nsew signal input
flabel metal2 s 11610 -300 11666 160 0 FreeSans 224 90 0 0 FrameStrobe[8]
port 18 nsew signal input
flabel metal2 s 12806 -300 12862 160 0 FreeSans 224 90 0 0 FrameStrobe[9]
port 19 nsew signal input
flabel metal2 s 20258 9840 20314 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[0]
port 20 nsew signal tristate
flabel metal2 s 23018 9840 23074 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[10]
port 21 nsew signal tristate
flabel metal2 s 23294 9840 23350 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[11]
port 22 nsew signal tristate
flabel metal2 s 23570 9840 23626 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[12]
port 23 nsew signal tristate
flabel metal2 s 23846 9840 23902 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[13]
port 24 nsew signal tristate
flabel metal2 s 24122 9840 24178 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[14]
port 25 nsew signal tristate
flabel metal2 s 24398 9840 24454 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[15]
port 26 nsew signal tristate
flabel metal2 s 24674 9840 24730 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[16]
port 27 nsew signal tristate
flabel metal2 s 24950 9840 25006 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[17]
port 28 nsew signal tristate
flabel metal2 s 25226 9840 25282 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[18]
port 29 nsew signal tristate
flabel metal2 s 25502 9840 25558 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[19]
port 30 nsew signal tristate
flabel metal2 s 20534 9840 20590 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[1]
port 31 nsew signal tristate
flabel metal2 s 20810 9840 20866 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[2]
port 32 nsew signal tristate
flabel metal2 s 21086 9840 21142 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[3]
port 33 nsew signal tristate
flabel metal2 s 21362 9840 21418 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[4]
port 34 nsew signal tristate
flabel metal2 s 21638 9840 21694 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[5]
port 35 nsew signal tristate
flabel metal2 s 21914 9840 21970 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[6]
port 36 nsew signal tristate
flabel metal2 s 22190 9840 22246 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[7]
port 37 nsew signal tristate
flabel metal2 s 22466 9840 22522 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[8]
port 38 nsew signal tristate
flabel metal2 s 22742 9840 22798 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[9]
port 39 nsew signal tristate
flabel metal2 s 110 9840 166 10300 0 FreeSans 224 90 0 0 N1BEG[0]
port 40 nsew signal tristate
flabel metal2 s 386 9840 442 10300 0 FreeSans 224 90 0 0 N1BEG[1]
port 41 nsew signal tristate
flabel metal2 s 662 9840 718 10300 0 FreeSans 224 90 0 0 N1BEG[2]
port 42 nsew signal tristate
flabel metal2 s 938 9840 994 10300 0 FreeSans 224 90 0 0 N1BEG[3]
port 43 nsew signal tristate
flabel metal2 s 1214 9840 1270 10300 0 FreeSans 224 90 0 0 N2BEG[0]
port 44 nsew signal tristate
flabel metal2 s 1490 9840 1546 10300 0 FreeSans 224 90 0 0 N2BEG[1]
port 45 nsew signal tristate
flabel metal2 s 1766 9840 1822 10300 0 FreeSans 224 90 0 0 N2BEG[2]
port 46 nsew signal tristate
flabel metal2 s 2042 9840 2098 10300 0 FreeSans 224 90 0 0 N2BEG[3]
port 47 nsew signal tristate
flabel metal2 s 2318 9840 2374 10300 0 FreeSans 224 90 0 0 N2BEG[4]
port 48 nsew signal tristate
flabel metal2 s 2594 9840 2650 10300 0 FreeSans 224 90 0 0 N2BEG[5]
port 49 nsew signal tristate
flabel metal2 s 2870 9840 2926 10300 0 FreeSans 224 90 0 0 N2BEG[6]
port 50 nsew signal tristate
flabel metal2 s 3146 9840 3202 10300 0 FreeSans 224 90 0 0 N2BEG[7]
port 51 nsew signal tristate
flabel metal2 s 3422 9840 3478 10300 0 FreeSans 224 90 0 0 N2BEGb[0]
port 52 nsew signal tristate
flabel metal2 s 3698 9840 3754 10300 0 FreeSans 224 90 0 0 N2BEGb[1]
port 53 nsew signal tristate
flabel metal2 s 3974 9840 4030 10300 0 FreeSans 224 90 0 0 N2BEGb[2]
port 54 nsew signal tristate
flabel metal2 s 4250 9840 4306 10300 0 FreeSans 224 90 0 0 N2BEGb[3]
port 55 nsew signal tristate
flabel metal2 s 4526 9840 4582 10300 0 FreeSans 224 90 0 0 N2BEGb[4]
port 56 nsew signal tristate
flabel metal2 s 4802 9840 4858 10300 0 FreeSans 224 90 0 0 N2BEGb[5]
port 57 nsew signal tristate
flabel metal2 s 5078 9840 5134 10300 0 FreeSans 224 90 0 0 N2BEGb[6]
port 58 nsew signal tristate
flabel metal2 s 5354 9840 5410 10300 0 FreeSans 224 90 0 0 N2BEGb[7]
port 59 nsew signal tristate
flabel metal2 s 5630 9840 5686 10300 0 FreeSans 224 90 0 0 N4BEG[0]
port 60 nsew signal tristate
flabel metal2 s 8390 9840 8446 10300 0 FreeSans 224 90 0 0 N4BEG[10]
port 61 nsew signal tristate
flabel metal2 s 8666 9840 8722 10300 0 FreeSans 224 90 0 0 N4BEG[11]
port 62 nsew signal tristate
flabel metal2 s 8942 9840 8998 10300 0 FreeSans 224 90 0 0 N4BEG[12]
port 63 nsew signal tristate
flabel metal2 s 9218 9840 9274 10300 0 FreeSans 224 90 0 0 N4BEG[13]
port 64 nsew signal tristate
flabel metal2 s 9494 9840 9550 10300 0 FreeSans 224 90 0 0 N4BEG[14]
port 65 nsew signal tristate
flabel metal2 s 9770 9840 9826 10300 0 FreeSans 224 90 0 0 N4BEG[15]
port 66 nsew signal tristate
flabel metal2 s 5906 9840 5962 10300 0 FreeSans 224 90 0 0 N4BEG[1]
port 67 nsew signal tristate
flabel metal2 s 6182 9840 6238 10300 0 FreeSans 224 90 0 0 N4BEG[2]
port 68 nsew signal tristate
flabel metal2 s 6458 9840 6514 10300 0 FreeSans 224 90 0 0 N4BEG[3]
port 69 nsew signal tristate
flabel metal2 s 6734 9840 6790 10300 0 FreeSans 224 90 0 0 N4BEG[4]
port 70 nsew signal tristate
flabel metal2 s 7010 9840 7066 10300 0 FreeSans 224 90 0 0 N4BEG[5]
port 71 nsew signal tristate
flabel metal2 s 7286 9840 7342 10300 0 FreeSans 224 90 0 0 N4BEG[6]
port 72 nsew signal tristate
flabel metal2 s 7562 9840 7618 10300 0 FreeSans 224 90 0 0 N4BEG[7]
port 73 nsew signal tristate
flabel metal2 s 7838 9840 7894 10300 0 FreeSans 224 90 0 0 N4BEG[8]
port 74 nsew signal tristate
flabel metal2 s 8114 9840 8170 10300 0 FreeSans 224 90 0 0 N4BEG[9]
port 75 nsew signal tristate
flabel metal2 s 10046 9840 10102 10300 0 FreeSans 224 90 0 0 S1END[0]
port 76 nsew signal input
flabel metal2 s 10322 9840 10378 10300 0 FreeSans 224 90 0 0 S1END[1]
port 77 nsew signal input
flabel metal2 s 10598 9840 10654 10300 0 FreeSans 224 90 0 0 S1END[2]
port 78 nsew signal input
flabel metal2 s 10874 9840 10930 10300 0 FreeSans 224 90 0 0 S1END[3]
port 79 nsew signal input
flabel metal2 s 11150 9840 11206 10300 0 FreeSans 224 90 0 0 S2END[0]
port 80 nsew signal input
flabel metal2 s 11426 9840 11482 10300 0 FreeSans 224 90 0 0 S2END[1]
port 81 nsew signal input
flabel metal2 s 11702 9840 11758 10300 0 FreeSans 224 90 0 0 S2END[2]
port 82 nsew signal input
flabel metal2 s 11978 9840 12034 10300 0 FreeSans 224 90 0 0 S2END[3]
port 83 nsew signal input
flabel metal2 s 12254 9840 12310 10300 0 FreeSans 224 90 0 0 S2END[4]
port 84 nsew signal input
flabel metal2 s 12530 9840 12586 10300 0 FreeSans 224 90 0 0 S2END[5]
port 85 nsew signal input
flabel metal2 s 12806 9840 12862 10300 0 FreeSans 224 90 0 0 S2END[6]
port 86 nsew signal input
flabel metal2 s 13082 9840 13138 10300 0 FreeSans 224 90 0 0 S2END[7]
port 87 nsew signal input
flabel metal2 s 13358 9840 13414 10300 0 FreeSans 224 90 0 0 S2MID[0]
port 88 nsew signal input
flabel metal2 s 13634 9840 13690 10300 0 FreeSans 224 90 0 0 S2MID[1]
port 89 nsew signal input
flabel metal2 s 13910 9840 13966 10300 0 FreeSans 224 90 0 0 S2MID[2]
port 90 nsew signal input
flabel metal2 s 14186 9840 14242 10300 0 FreeSans 224 90 0 0 S2MID[3]
port 91 nsew signal input
flabel metal2 s 14462 9840 14518 10300 0 FreeSans 224 90 0 0 S2MID[4]
port 92 nsew signal input
flabel metal2 s 14738 9840 14794 10300 0 FreeSans 224 90 0 0 S2MID[5]
port 93 nsew signal input
flabel metal2 s 15014 9840 15070 10300 0 FreeSans 224 90 0 0 S2MID[6]
port 94 nsew signal input
flabel metal2 s 15290 9840 15346 10300 0 FreeSans 224 90 0 0 S2MID[7]
port 95 nsew signal input
flabel metal2 s 15566 9840 15622 10300 0 FreeSans 224 90 0 0 S4END[0]
port 96 nsew signal input
flabel metal2 s 18326 9840 18382 10300 0 FreeSans 224 90 0 0 S4END[10]
port 97 nsew signal input
flabel metal2 s 18602 9840 18658 10300 0 FreeSans 224 90 0 0 S4END[11]
port 98 nsew signal input
flabel metal2 s 18878 9840 18934 10300 0 FreeSans 224 90 0 0 S4END[12]
port 99 nsew signal input
flabel metal2 s 19154 9840 19210 10300 0 FreeSans 224 90 0 0 S4END[13]
port 100 nsew signal input
flabel metal2 s 19430 9840 19486 10300 0 FreeSans 224 90 0 0 S4END[14]
port 101 nsew signal input
flabel metal2 s 19706 9840 19762 10300 0 FreeSans 224 90 0 0 S4END[15]
port 102 nsew signal input
flabel metal2 s 15842 9840 15898 10300 0 FreeSans 224 90 0 0 S4END[1]
port 103 nsew signal input
flabel metal2 s 16118 9840 16174 10300 0 FreeSans 224 90 0 0 S4END[2]
port 104 nsew signal input
flabel metal2 s 16394 9840 16450 10300 0 FreeSans 224 90 0 0 S4END[3]
port 105 nsew signal input
flabel metal2 s 16670 9840 16726 10300 0 FreeSans 224 90 0 0 S4END[4]
port 106 nsew signal input
flabel metal2 s 16946 9840 17002 10300 0 FreeSans 224 90 0 0 S4END[5]
port 107 nsew signal input
flabel metal2 s 17222 9840 17278 10300 0 FreeSans 224 90 0 0 S4END[6]
port 108 nsew signal input
flabel metal2 s 17498 9840 17554 10300 0 FreeSans 224 90 0 0 S4END[7]
port 109 nsew signal input
flabel metal2 s 17774 9840 17830 10300 0 FreeSans 224 90 0 0 S4END[8]
port 110 nsew signal input
flabel metal2 s 18050 9840 18106 10300 0 FreeSans 224 90 0 0 S4END[9]
port 111 nsew signal input
flabel metal2 s 846 -300 902 160 0 FreeSans 224 90 0 0 UserCLK
port 112 nsew signal input
flabel metal2 s 19982 9840 20038 10300 0 FreeSans 224 90 0 0 UserCLKo
port 113 nsew signal tristate
flabel metal4 s 6808 1040 7128 8752 0 FreeSans 1920 90 0 0 VGND
port 114 nsew ground bidirectional
flabel metal4 s 12673 1040 12993 8752 0 FreeSans 1920 90 0 0 VGND
port 114 nsew ground bidirectional
flabel metal4 s 18538 1040 18858 8752 0 FreeSans 1920 90 0 0 VGND
port 114 nsew ground bidirectional
flabel metal4 s 24403 1040 24723 8752 0 FreeSans 1920 90 0 0 VGND
port 114 nsew ground bidirectional
flabel metal4 s 3876 1040 4196 8752 0 FreeSans 1920 90 0 0 VPWR
port 115 nsew power bidirectional
flabel metal4 s 9741 1040 10061 8752 0 FreeSans 1920 90 0 0 VPWR
port 115 nsew power bidirectional
flabel metal4 s 15606 1040 15926 8752 0 FreeSans 1920 90 0 0 VPWR
port 115 nsew power bidirectional
flabel metal4 s 21471 1040 21791 8752 0 FreeSans 1920 90 0 0 VPWR
port 115 nsew power bidirectional
rlabel via1 12913 8704 12913 8704 0 VGND
rlabel metal1 12834 8160 12834 8160 0 VPWR
rlabel metal2 2123 68 2123 68 0 FrameStrobe[0]
rlabel metal2 14175 68 14175 68 0 FrameStrobe[10]
rlabel metal2 15371 68 15371 68 0 FrameStrobe[11]
rlabel metal1 16790 1326 16790 1326 0 FrameStrobe[12]
rlabel metal2 17763 68 17763 68 0 FrameStrobe[13]
rlabel metal2 18959 68 18959 68 0 FrameStrobe[14]
rlabel metal2 20155 68 20155 68 0 FrameStrobe[15]
rlabel metal2 21351 68 21351 68 0 FrameStrobe[16]
rlabel metal2 22547 68 22547 68 0 FrameStrobe[17]
rlabel metal2 23598 143 23598 143 0 FrameStrobe[18]
rlabel metal2 24794 398 24794 398 0 FrameStrobe[19]
rlabel metal2 3319 68 3319 68 0 FrameStrobe[1]
rlabel metal2 4607 68 4607 68 0 FrameStrobe[2]
rlabel metal2 5803 68 5803 68 0 FrameStrobe[3]
rlabel metal2 6946 323 6946 323 0 FrameStrobe[4]
rlabel metal2 8287 68 8287 68 0 FrameStrobe[5]
rlabel metal2 9391 68 9391 68 0 FrameStrobe[6]
rlabel metal2 10587 68 10587 68 0 FrameStrobe[7]
rlabel metal2 11783 68 11783 68 0 FrameStrobe[8]
rlabel metal2 12834 143 12834 143 0 FrameStrobe[9]
rlabel metal2 20286 9445 20286 9445 0 FrameStrobe_O[0]
rlabel metal2 23046 9836 23046 9836 0 FrameStrobe_O[10]
rlabel metal2 23322 8136 23322 8136 0 FrameStrobe_O[11]
rlabel metal2 23598 9836 23598 9836 0 FrameStrobe_O[12]
rlabel metal1 23736 6766 23736 6766 0 FrameStrobe_O[13]
rlabel metal1 24012 7514 24012 7514 0 FrameStrobe_O[14]
rlabel metal1 24150 6834 24150 6834 0 FrameStrobe_O[15]
rlabel metal1 24104 7446 24104 7446 0 FrameStrobe_O[16]
rlabel metal1 23874 7310 23874 7310 0 FrameStrobe_O[17]
rlabel metal1 24702 5882 24702 5882 0 FrameStrobe_O[18]
rlabel metal2 25530 8850 25530 8850 0 FrameStrobe_O[19]
rlabel metal2 20562 9088 20562 9088 0 FrameStrobe_O[1]
rlabel metal1 21068 8058 21068 8058 0 FrameStrobe_O[2]
rlabel metal1 21574 8602 21574 8602 0 FrameStrobe_O[3]
rlabel metal1 22586 8568 22586 8568 0 FrameStrobe_O[4]
rlabel metal2 21666 9088 21666 9088 0 FrameStrobe_O[5]
rlabel metal2 21942 8952 21942 8952 0 FrameStrobe_O[6]
rlabel metal2 22218 8952 22218 8952 0 FrameStrobe_O[7]
rlabel metal2 22494 9836 22494 9836 0 FrameStrobe_O[8]
rlabel metal2 22770 9836 22770 9836 0 FrameStrobe_O[9]
rlabel metal1 11316 1530 11316 1530 0 FrameStrobe_O_i\[0\]
rlabel metal1 14582 4250 14582 4250 0 FrameStrobe_O_i\[10\]
rlabel metal1 15870 1530 15870 1530 0 FrameStrobe_O_i\[11\]
rlabel metal1 17066 6970 17066 6970 0 FrameStrobe_O_i\[12\]
rlabel metal1 23506 3468 23506 3468 0 FrameStrobe_O_i\[13\]
rlabel metal2 23138 1700 23138 1700 0 FrameStrobe_O_i\[14\]
rlabel metal2 22862 1734 22862 1734 0 FrameStrobe_O_i\[15\]
rlabel metal1 22034 1530 22034 1530 0 FrameStrobe_O_i\[16\]
rlabel metal1 23506 2992 23506 2992 0 FrameStrobe_O_i\[17\]
rlabel metal1 23920 1530 23920 1530 0 FrameStrobe_O_i\[18\]
rlabel metal1 23966 2618 23966 2618 0 FrameStrobe_O_i\[19\]
rlabel metal1 13570 1224 13570 1224 0 FrameStrobe_O_i\[1\]
rlabel metal1 12604 1530 12604 1530 0 FrameStrobe_O_i\[2\]
rlabel metal1 9982 1530 9982 1530 0 FrameStrobe_O_i\[3\]
rlabel metal1 7406 1530 7406 1530 0 FrameStrobe_O_i\[4\]
rlabel metal1 8602 1530 8602 1530 0 FrameStrobe_O_i\[5\]
rlabel metal1 10258 1462 10258 1462 0 FrameStrobe_O_i\[6\]
rlabel metal1 11086 1190 11086 1190 0 FrameStrobe_O_i\[7\]
rlabel metal1 12144 1190 12144 1190 0 FrameStrobe_O_i\[8\]
rlabel metal1 13386 1530 13386 1530 0 FrameStrobe_O_i\[9\]
rlabel metal2 138 9326 138 9326 0 N1BEG[0]
rlabel metal2 414 9224 414 9224 0 N1BEG[1]
rlabel metal2 690 8340 690 8340 0 N1BEG[2]
rlabel metal1 1288 6426 1288 6426 0 N1BEG[3]
rlabel metal1 1610 6766 1610 6766 0 N2BEG[0]
rlabel metal2 1518 8646 1518 8646 0 N2BEG[1]
rlabel metal2 1794 8680 1794 8680 0 N2BEG[2]
rlabel metal1 1932 8058 1932 8058 0 N2BEG[3]
rlabel metal2 2346 8952 2346 8952 0 N2BEG[4]
rlabel metal2 2622 8918 2622 8918 0 N2BEG[5]
rlabel metal1 2852 8602 2852 8602 0 N2BEG[6]
rlabel metal2 3174 8952 3174 8952 0 N2BEG[7]
rlabel metal2 3450 9088 3450 9088 0 N2BEGb[0]
rlabel metal1 3634 7514 3634 7514 0 N2BEGb[1]
rlabel metal2 4002 9105 4002 9105 0 N2BEGb[2]
rlabel metal2 4278 9224 4278 9224 0 N2BEGb[3]
rlabel metal2 4554 8952 4554 8952 0 N2BEGb[4]
rlabel metal1 5014 8058 5014 8058 0 N2BEGb[5]
rlabel metal1 4876 8602 4876 8602 0 N2BEGb[6]
rlabel metal1 5290 8602 5290 8602 0 N2BEGb[7]
rlabel metal2 5658 8952 5658 8952 0 N4BEG[0]
rlabel metal1 8372 8602 8372 8602 0 N4BEG[10]
rlabel metal2 8694 8952 8694 8952 0 N4BEG[11]
rlabel metal1 8832 8602 8832 8602 0 N4BEG[12]
rlabel metal1 9292 8602 9292 8602 0 N4BEG[13]
rlabel metal2 9522 9734 9522 9734 0 N4BEG[14]
rlabel metal2 9798 9224 9798 9224 0 N4BEG[15]
rlabel metal1 5842 8602 5842 8602 0 N4BEG[1]
rlabel metal2 6210 8952 6210 8952 0 N4BEG[2]
rlabel metal1 6302 8602 6302 8602 0 N4BEG[3]
rlabel metal2 6762 8918 6762 8918 0 N4BEG[4]
rlabel metal1 7038 8602 7038 8602 0 N4BEG[5]
rlabel metal1 7360 8058 7360 8058 0 N4BEG[6]
rlabel metal1 7498 8602 7498 8602 0 N4BEG[7]
rlabel metal2 7866 8952 7866 8952 0 N4BEG[8]
rlabel metal1 7958 8602 7958 8602 0 N4BEG[9]
rlabel metal2 10074 9836 10074 9836 0 S1END[0]
rlabel metal2 10350 9836 10350 9836 0 S1END[1]
rlabel metal2 10626 9836 10626 9836 0 S1END[2]
rlabel metal2 10902 9581 10902 9581 0 S1END[3]
rlabel metal2 11178 9836 11178 9836 0 S2END[0]
rlabel metal2 11454 9836 11454 9836 0 S2END[1]
rlabel metal2 11730 9156 11730 9156 0 S2END[2]
rlabel metal2 12006 8850 12006 8850 0 S2END[3]
rlabel metal2 12282 8850 12282 8850 0 S2END[4]
rlabel metal2 12558 9173 12558 9173 0 S2END[5]
rlabel metal2 12834 9836 12834 9836 0 S2END[6]
rlabel metal2 13110 9836 13110 9836 0 S2END[7]
rlabel metal2 13386 9156 13386 9156 0 S2MID[0]
rlabel metal2 13662 9156 13662 9156 0 S2MID[1]
rlabel metal2 13938 9156 13938 9156 0 S2MID[2]
rlabel metal2 14214 9190 14214 9190 0 S2MID[3]
rlabel metal2 14490 8850 14490 8850 0 S2MID[4]
rlabel metal2 14766 9836 14766 9836 0 S2MID[5]
rlabel metal2 15042 9377 15042 9377 0 S2MID[6]
rlabel metal2 15318 9836 15318 9836 0 S2MID[7]
rlabel metal2 15594 9836 15594 9836 0 S4END[0]
rlabel metal2 18354 9513 18354 9513 0 S4END[10]
rlabel metal2 18630 9326 18630 9326 0 S4END[11]
rlabel metal2 18906 9360 18906 9360 0 S4END[12]
rlabel metal2 19182 8850 19182 8850 0 S4END[13]
rlabel metal2 19458 8850 19458 8850 0 S4END[14]
rlabel metal2 19734 8850 19734 8850 0 S4END[15]
rlabel metal2 15870 9836 15870 9836 0 S4END[1]
rlabel metal2 16146 9836 16146 9836 0 S4END[2]
rlabel metal2 16422 9836 16422 9836 0 S4END[3]
rlabel metal2 16698 8850 16698 8850 0 S4END[4]
rlabel metal2 16974 9836 16974 9836 0 S4END[5]
rlabel metal2 17250 8850 17250 8850 0 S4END[6]
rlabel metal2 17526 9122 17526 9122 0 S4END[7]
rlabel metal2 17802 8850 17802 8850 0 S4END[8]
rlabel metal2 18078 9836 18078 9836 0 S4END[9]
rlabel metal2 874 704 874 704 0 UserCLK
rlabel metal1 20148 8602 20148 8602 0 UserCLKo
rlabel metal2 2346 986 2346 986 0 net1
rlabel metal1 23920 1326 23920 1326 0 net10
rlabel metal1 8556 7514 8556 7514 0 net100
rlabel metal2 16974 8738 16974 8738 0 net101
rlabel metal1 9154 8432 9154 8432 0 net102
rlabel metal1 16284 8330 16284 8330 0 net103
rlabel metal1 16100 8262 16100 8262 0 net104
rlabel metal1 5934 7174 5934 7174 0 net105
rlabel metal1 19090 6936 19090 6936 0 net106
rlabel metal1 6164 7514 6164 7514 0 net107
rlabel metal2 18630 7769 18630 7769 0 net108
rlabel metal1 19044 8330 19044 8330 0 net109
rlabel metal1 23368 1530 23368 1530 0 net11
rlabel metal1 18492 8330 18492 8330 0 net110
rlabel metal1 7452 7514 7452 7514 0 net111
rlabel metal1 18078 8602 18078 8602 0 net112
rlabel metal2 8326 7956 8326 7956 0 net113
rlabel metal2 14582 1088 14582 1088 0 net114
rlabel metal1 3542 1224 3542 1224 0 net12
rlabel metal1 4554 952 4554 952 0 net13
rlabel metal2 5750 1088 5750 1088 0 net14
rlabel metal1 7360 1326 7360 1326 0 net15
rlabel metal1 8556 1326 8556 1326 0 net16
rlabel metal1 10166 1292 10166 1292 0 net17
rlabel metal1 10994 1292 10994 1292 0 net18
rlabel metal1 12190 1292 12190 1292 0 net19
rlabel metal1 14306 1190 14306 1190 0 net2
rlabel metal1 13294 1292 13294 1292 0 net20
rlabel metal1 9913 7174 9913 7174 0 net21
rlabel metal1 10258 7752 10258 7752 0 net22
rlabel metal1 9246 7888 9246 7888 0 net23
rlabel metal1 9890 7888 9890 7888 0 net24
rlabel metal2 9798 7956 9798 7956 0 net25
rlabel metal1 10350 7820 10350 7820 0 net26
rlabel metal1 10810 8432 10810 8432 0 net27
rlabel metal1 11592 7990 11592 7990 0 net28
rlabel metal1 11960 8058 11960 8058 0 net29
rlabel metal1 15778 1292 15778 1292 0 net3
rlabel metal1 12558 8058 12558 8058 0 net30
rlabel metal2 12926 8330 12926 8330 0 net31
rlabel metal2 13202 8228 13202 8228 0 net32
rlabel metal1 12650 8500 12650 8500 0 net33
rlabel metal1 13110 8466 13110 8466 0 net34
rlabel metal1 13478 8432 13478 8432 0 net35
rlabel metal1 14398 8432 14398 8432 0 net36
rlabel metal1 14628 8058 14628 8058 0 net37
rlabel metal1 15042 8058 15042 8058 0 net38
rlabel metal1 15226 7990 15226 7990 0 net39
rlabel metal1 16744 1190 16744 1190 0 net4
rlabel metal2 15410 8228 15410 8228 0 net40
rlabel metal1 15916 8058 15916 8058 0 net41
rlabel metal1 19090 8466 19090 8466 0 net42
rlabel metal1 18630 7854 18630 7854 0 net43
rlabel metal1 19688 8330 19688 8330 0 net44
rlabel metal1 19090 7854 19090 7854 0 net45
rlabel metal2 19734 7497 19734 7497 0 net46
rlabel metal2 20010 7565 20010 7565 0 net47
rlabel metal1 16238 7990 16238 7990 0 net48
rlabel metal1 16560 8058 16560 8058 0 net49
rlabel metal1 17756 1190 17756 1190 0 net5
rlabel metal1 17204 8466 17204 8466 0 net50
rlabel metal2 16790 7616 16790 7616 0 net51
rlabel metal1 17756 8466 17756 8466 0 net52
rlabel metal1 17342 7378 17342 7378 0 net53
rlabel metal1 18216 8466 18216 8466 0 net54
rlabel metal1 17894 7752 17894 7752 0 net55
rlabel metal1 18400 8058 18400 8058 0 net56
rlabel metal1 1610 918 1610 918 0 net57
rlabel metal1 11638 2074 11638 2074 0 net58
rlabel metal2 23552 8466 23552 8466 0 net59
rlabel metal1 23322 1258 23322 1258 0 net6
rlabel metal1 23230 2040 23230 2040 0 net60
rlabel metal1 22954 6358 22954 6358 0 net61
rlabel metal1 23230 3706 23230 3706 0 net62
rlabel metal1 23644 2074 23644 2074 0 net63
rlabel metal2 23414 4386 23414 4386 0 net64
rlabel metal1 22540 2074 22540 2074 0 net65
rlabel metal1 22908 3162 22908 3162 0 net66
rlabel metal1 23920 2074 23920 2074 0 net67
rlabel metal1 23874 3128 23874 3128 0 net68
rlabel metal1 17526 2074 17526 2074 0 net69
rlabel metal1 23046 1292 23046 1292 0 net7
rlabel metal1 13018 2040 13018 2040 0 net70
rlabel metal2 10442 2176 10442 2176 0 net71
rlabel metal3 22425 8364 22425 8364 0 net72
rlabel metal4 22540 4436 22540 4436 0 net73
rlabel via3 22149 7276 22149 7276 0 net74
rlabel metal2 22678 4794 22678 4794 0 net75
rlabel metal1 23000 7786 23000 7786 0 net76
rlabel metal2 23782 5066 23782 5066 0 net77
rlabel metal1 9522 7718 9522 7718 0 net78
rlabel metal1 1978 9248 1978 9248 0 net79
rlabel metal1 22034 1292 22034 1292 0 net8
rlabel metal1 2714 7344 2714 7344 0 net80
rlabel metal2 5474 7140 5474 7140 0 net81
rlabel metal1 2530 6698 2530 6698 0 net82
rlabel metal1 15686 8296 15686 8296 0 net83
rlabel metal2 1610 8602 1610 8602 0 net84
rlabel metal2 14858 9146 14858 9146 0 net85
rlabel metal2 2254 8874 2254 8874 0 net86
rlabel via2 2622 7837 2622 7837 0 net87
rlabel metal2 2530 8840 2530 8840 0 net88
rlabel metal1 12466 8296 12466 8296 0 net89
rlabel metal2 22494 2108 22494 2108 0 net9
rlabel metal1 1518 8500 1518 8500 0 net90
rlabel metal1 3358 7344 3358 7344 0 net91
rlabel metal1 4002 7752 4002 7752 0 net92
rlabel metal1 5244 8534 5244 8534 0 net93
rlabel metal1 5060 7786 5060 7786 0 net94
rlabel metal1 5842 7854 5842 7854 0 net95
rlabel metal2 10166 8041 10166 8041 0 net96
rlabel metal1 9522 8058 9522 8058 0 net97
rlabel metal1 5566 7514 5566 7514 0 net98
rlabel metal1 17434 8602 17434 8602 0 net99
<< properties >>
string FIXED_BBOX 0 0 25700 10000
<< end >>
