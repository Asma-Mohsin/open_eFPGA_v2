magic
tech sky130A
magscale 1 2
timestamp 1734828903
<< obsli1 >>
rect 1104 1071 21896 43537
<< obsm1 >>
rect 14 620 22986 43920
<< metal2 >>
rect 2962 44540 3018 45000
rect 3146 44540 3202 45000
rect 3330 44540 3386 45000
rect 3514 44540 3570 45000
rect 3698 44540 3754 45000
rect 3882 44540 3938 45000
rect 4066 44540 4122 45000
rect 4250 44540 4306 45000
rect 4434 44540 4490 45000
rect 4618 44540 4674 45000
rect 4802 44540 4858 45000
rect 4986 44540 5042 45000
rect 5170 44540 5226 45000
rect 5354 44540 5410 45000
rect 5538 44540 5594 45000
rect 5722 44540 5778 45000
rect 5906 44540 5962 45000
rect 6090 44540 6146 45000
rect 6274 44540 6330 45000
rect 6458 44540 6514 45000
rect 6642 44540 6698 45000
rect 6826 44540 6882 45000
rect 7010 44540 7066 45000
rect 7194 44540 7250 45000
rect 7378 44540 7434 45000
rect 7562 44540 7618 45000
rect 7746 44540 7802 45000
rect 7930 44540 7986 45000
rect 8114 44540 8170 45000
rect 8298 44540 8354 45000
rect 8482 44540 8538 45000
rect 8666 44540 8722 45000
rect 8850 44540 8906 45000
rect 9034 44540 9090 45000
rect 9218 44540 9274 45000
rect 9402 44540 9458 45000
rect 9586 44540 9642 45000
rect 9770 44540 9826 45000
rect 9954 44540 10010 45000
rect 10138 44540 10194 45000
rect 10322 44540 10378 45000
rect 10506 44540 10562 45000
rect 10690 44540 10746 45000
rect 10874 44540 10930 45000
rect 11058 44540 11114 45000
rect 11242 44540 11298 45000
rect 11426 44540 11482 45000
rect 11610 44540 11666 45000
rect 11794 44540 11850 45000
rect 11978 44540 12034 45000
rect 12162 44540 12218 45000
rect 12346 44540 12402 45000
rect 12530 44540 12586 45000
rect 12714 44540 12770 45000
rect 12898 44540 12954 45000
rect 13082 44540 13138 45000
rect 13266 44540 13322 45000
rect 13450 44540 13506 45000
rect 13634 44540 13690 45000
rect 13818 44540 13874 45000
rect 14002 44540 14058 45000
rect 14186 44540 14242 45000
rect 14370 44540 14426 45000
rect 14554 44540 14610 45000
rect 14738 44540 14794 45000
rect 14922 44540 14978 45000
rect 15106 44540 15162 45000
rect 15290 44540 15346 45000
rect 15474 44540 15530 45000
rect 15658 44540 15714 45000
rect 15842 44540 15898 45000
rect 16026 44540 16082 45000
rect 16210 44540 16266 45000
rect 16394 44540 16450 45000
rect 16578 44540 16634 45000
rect 16762 44540 16818 45000
rect 16946 44540 17002 45000
rect 17130 44540 17186 45000
rect 17314 44540 17370 45000
rect 17498 44540 17554 45000
rect 17682 44540 17738 45000
rect 17866 44540 17922 45000
rect 18050 44540 18106 45000
rect 18234 44540 18290 45000
rect 18418 44540 18474 45000
rect 18602 44540 18658 45000
rect 18786 44540 18842 45000
rect 18970 44540 19026 45000
rect 19154 44540 19210 45000
rect 19338 44540 19394 45000
rect 19522 44540 19578 45000
rect 19706 44540 19762 45000
rect 19890 44540 19946 45000
rect 2962 -300 3018 160
rect 3146 -300 3202 160
rect 3330 -300 3386 160
rect 3514 -300 3570 160
rect 3698 -300 3754 160
rect 3882 -300 3938 160
rect 4066 -300 4122 160
rect 4250 -300 4306 160
rect 4434 -300 4490 160
rect 4618 -300 4674 160
rect 4802 -300 4858 160
rect 4986 -300 5042 160
rect 5170 -300 5226 160
rect 5354 -300 5410 160
rect 5538 -300 5594 160
rect 5722 -300 5778 160
rect 5906 -300 5962 160
rect 6090 -300 6146 160
rect 6274 -300 6330 160
rect 6458 -300 6514 160
rect 6642 -300 6698 160
rect 6826 -300 6882 160
rect 7010 -300 7066 160
rect 7194 -300 7250 160
rect 7378 -300 7434 160
rect 7562 -300 7618 160
rect 7746 -300 7802 160
rect 7930 -300 7986 160
rect 8114 -300 8170 160
rect 8298 -300 8354 160
rect 8482 -300 8538 160
rect 8666 -300 8722 160
rect 8850 -300 8906 160
rect 9034 -300 9090 160
rect 9218 -300 9274 160
rect 9402 -300 9458 160
rect 9586 -300 9642 160
rect 9770 -300 9826 160
rect 9954 -300 10010 160
rect 10138 -300 10194 160
rect 10322 -300 10378 160
rect 10506 -300 10562 160
rect 10690 -300 10746 160
rect 10874 -300 10930 160
rect 11058 -300 11114 160
rect 11242 -300 11298 160
rect 11426 -300 11482 160
rect 11610 -300 11666 160
rect 11794 -300 11850 160
rect 11978 -300 12034 160
rect 12162 -300 12218 160
rect 12346 -300 12402 160
rect 12530 -300 12586 160
rect 12714 -300 12770 160
rect 12898 -300 12954 160
rect 13082 -300 13138 160
rect 13266 -300 13322 160
rect 13450 -300 13506 160
rect 13634 -300 13690 160
rect 13818 -300 13874 160
rect 14002 -300 14058 160
rect 14186 -300 14242 160
rect 14370 -300 14426 160
rect 14554 -300 14610 160
rect 14738 -300 14794 160
rect 14922 -300 14978 160
rect 15106 -300 15162 160
rect 15290 -300 15346 160
rect 15474 -300 15530 160
rect 15658 -300 15714 160
rect 15842 -300 15898 160
rect 16026 -300 16082 160
rect 16210 -300 16266 160
rect 16394 -300 16450 160
rect 16578 -300 16634 160
rect 16762 -300 16818 160
rect 16946 -300 17002 160
rect 17130 -300 17186 160
rect 17314 -300 17370 160
rect 17498 -300 17554 160
rect 17682 -300 17738 160
rect 17866 -300 17922 160
rect 18050 -300 18106 160
rect 18234 -300 18290 160
rect 18418 -300 18474 160
rect 18602 -300 18658 160
rect 18786 -300 18842 160
rect 18970 -300 19026 160
rect 19154 -300 19210 160
rect 19338 -300 19394 160
rect 19522 -300 19578 160
rect 19706 -300 19762 160
rect 19890 -300 19946 160
<< obsm2 >>
rect 18 44484 2906 44540
rect 3074 44484 3090 44540
rect 3258 44484 3274 44540
rect 3442 44484 3458 44540
rect 3626 44484 3642 44540
rect 3810 44484 3826 44540
rect 3994 44484 4010 44540
rect 4178 44484 4194 44540
rect 4362 44484 4378 44540
rect 4546 44484 4562 44540
rect 4730 44484 4746 44540
rect 4914 44484 4930 44540
rect 5098 44484 5114 44540
rect 5282 44484 5298 44540
rect 5466 44484 5482 44540
rect 5650 44484 5666 44540
rect 5834 44484 5850 44540
rect 6018 44484 6034 44540
rect 6202 44484 6218 44540
rect 6386 44484 6402 44540
rect 6570 44484 6586 44540
rect 6754 44484 6770 44540
rect 6938 44484 6954 44540
rect 7122 44484 7138 44540
rect 7306 44484 7322 44540
rect 7490 44484 7506 44540
rect 7674 44484 7690 44540
rect 7858 44484 7874 44540
rect 8042 44484 8058 44540
rect 8226 44484 8242 44540
rect 8410 44484 8426 44540
rect 8594 44484 8610 44540
rect 8778 44484 8794 44540
rect 8962 44484 8978 44540
rect 9146 44484 9162 44540
rect 9330 44484 9346 44540
rect 9514 44484 9530 44540
rect 9698 44484 9714 44540
rect 9882 44484 9898 44540
rect 10066 44484 10082 44540
rect 10250 44484 10266 44540
rect 10434 44484 10450 44540
rect 10618 44484 10634 44540
rect 10802 44484 10818 44540
rect 10986 44484 11002 44540
rect 11170 44484 11186 44540
rect 11354 44484 11370 44540
rect 11538 44484 11554 44540
rect 11722 44484 11738 44540
rect 11906 44484 11922 44540
rect 12090 44484 12106 44540
rect 12274 44484 12290 44540
rect 12458 44484 12474 44540
rect 12642 44484 12658 44540
rect 12826 44484 12842 44540
rect 13010 44484 13026 44540
rect 13194 44484 13210 44540
rect 13378 44484 13394 44540
rect 13562 44484 13578 44540
rect 13746 44484 13762 44540
rect 13930 44484 13946 44540
rect 14114 44484 14130 44540
rect 14298 44484 14314 44540
rect 14482 44484 14498 44540
rect 14666 44484 14682 44540
rect 14850 44484 14866 44540
rect 15034 44484 15050 44540
rect 15218 44484 15234 44540
rect 15402 44484 15418 44540
rect 15586 44484 15602 44540
rect 15770 44484 15786 44540
rect 15954 44484 15970 44540
rect 16138 44484 16154 44540
rect 16322 44484 16338 44540
rect 16506 44484 16522 44540
rect 16690 44484 16706 44540
rect 16874 44484 16890 44540
rect 17058 44484 17074 44540
rect 17242 44484 17258 44540
rect 17426 44484 17442 44540
rect 17610 44484 17626 44540
rect 17794 44484 17810 44540
rect 17978 44484 17994 44540
rect 18162 44484 18178 44540
rect 18346 44484 18362 44540
rect 18530 44484 18546 44540
rect 18714 44484 18730 44540
rect 18898 44484 18914 44540
rect 19082 44484 19098 44540
rect 19266 44484 19282 44540
rect 19450 44484 19466 44540
rect 19634 44484 19650 44540
rect 19818 44484 19834 44540
rect 20002 44484 22980 44540
rect 18 216 22980 44484
rect 18 31 2906 216
rect 3074 31 3090 216
rect 3258 31 3274 216
rect 3442 31 3458 216
rect 3626 31 3642 216
rect 3810 31 3826 216
rect 3994 31 4010 216
rect 4178 31 4194 216
rect 4362 31 4378 216
rect 4546 31 4562 216
rect 4730 31 4746 216
rect 4914 31 4930 216
rect 5098 31 5114 216
rect 5282 31 5298 216
rect 5466 31 5482 216
rect 5650 31 5666 216
rect 5834 31 5850 216
rect 6018 31 6034 216
rect 6202 31 6218 216
rect 6386 31 6402 216
rect 6570 31 6586 216
rect 6754 31 6770 216
rect 6938 31 6954 216
rect 7122 31 7138 216
rect 7306 31 7322 216
rect 7490 31 7506 216
rect 7674 31 7690 216
rect 7858 31 7874 216
rect 8042 31 8058 216
rect 8226 31 8242 216
rect 8410 31 8426 216
rect 8594 31 8610 216
rect 8778 31 8794 216
rect 8962 31 8978 216
rect 9146 31 9162 216
rect 9330 31 9346 216
rect 9514 31 9530 216
rect 9698 31 9714 216
rect 9882 31 9898 216
rect 10066 31 10082 216
rect 10250 31 10266 216
rect 10434 31 10450 216
rect 10618 31 10634 216
rect 10802 31 10818 216
rect 10986 31 11002 216
rect 11170 31 11186 216
rect 11354 31 11370 216
rect 11538 31 11554 216
rect 11722 31 11738 216
rect 11906 31 11922 216
rect 12090 31 12106 216
rect 12274 31 12290 216
rect 12458 31 12474 216
rect 12642 31 12658 216
rect 12826 31 12842 216
rect 13010 31 13026 216
rect 13194 31 13210 216
rect 13378 31 13394 216
rect 13562 31 13578 216
rect 13746 31 13762 216
rect 13930 31 13946 216
rect 14114 31 14130 216
rect 14298 31 14314 216
rect 14482 31 14498 216
rect 14666 31 14682 216
rect 14850 31 14866 216
rect 15034 31 15050 216
rect 15218 31 15234 216
rect 15402 31 15418 216
rect 15586 31 15602 216
rect 15770 31 15786 216
rect 15954 31 15970 216
rect 16138 31 16154 216
rect 16322 31 16338 216
rect 16506 31 16522 216
rect 16690 31 16706 216
rect 16874 31 16890 216
rect 17058 31 17074 216
rect 17242 31 17258 216
rect 17426 31 17442 216
rect 17610 31 17626 216
rect 17794 31 17810 216
rect 17978 31 17994 216
rect 18162 31 18178 216
rect 18346 31 18362 216
rect 18530 31 18546 216
rect 18714 31 18730 216
rect 18898 31 18914 216
rect 19082 31 19098 216
rect 19266 31 19282 216
rect 19450 31 19466 216
rect 19634 31 19650 216
rect 19818 31 19834 216
rect 20002 31 22980 216
<< metal3 >>
rect 22840 43528 23300 43648
rect 22840 42984 23300 43104
rect 22840 42440 23300 42560
rect 22840 41896 23300 42016
rect 22840 41352 23300 41472
rect 22840 40808 23300 40928
rect 22840 40264 23300 40384
rect 22840 39720 23300 39840
rect -300 39448 160 39568
rect -300 39176 160 39296
rect 22840 39176 23300 39296
rect -300 38904 160 39024
rect -300 38632 160 38752
rect 22840 38632 23300 38752
rect -300 38360 160 38480
rect -300 38088 160 38208
rect 22840 38088 23300 38208
rect -300 37816 160 37936
rect -300 37544 160 37664
rect 22840 37544 23300 37664
rect -300 37272 160 37392
rect -300 37000 160 37120
rect 22840 37000 23300 37120
rect -300 36728 160 36848
rect -300 36456 160 36576
rect 22840 36456 23300 36576
rect -300 36184 160 36304
rect -300 35912 160 36032
rect 22840 35912 23300 36032
rect -300 35640 160 35760
rect -300 35368 160 35488
rect 22840 35368 23300 35488
rect -300 35096 160 35216
rect -300 34824 160 34944
rect 22840 34824 23300 34944
rect -300 34552 160 34672
rect -300 34280 160 34400
rect 22840 34280 23300 34400
rect -300 34008 160 34128
rect -300 33736 160 33856
rect 22840 33736 23300 33856
rect -300 33464 160 33584
rect -300 33192 160 33312
rect 22840 33192 23300 33312
rect -300 32920 160 33040
rect -300 32648 160 32768
rect 22840 32648 23300 32768
rect -300 32376 160 32496
rect -300 32104 160 32224
rect 22840 32104 23300 32224
rect -300 31832 160 31952
rect -300 31560 160 31680
rect 22840 31560 23300 31680
rect -300 31288 160 31408
rect -300 31016 160 31136
rect 22840 31016 23300 31136
rect -300 30744 160 30864
rect -300 30472 160 30592
rect 22840 30472 23300 30592
rect -300 30200 160 30320
rect -300 29928 160 30048
rect 22840 29928 23300 30048
rect -300 29656 160 29776
rect -300 29384 160 29504
rect 22840 29384 23300 29504
rect -300 29112 160 29232
rect -300 28840 160 28960
rect 22840 28840 23300 28960
rect -300 28568 160 28688
rect -300 28296 160 28416
rect 22840 28296 23300 28416
rect -300 28024 160 28144
rect -300 27752 160 27872
rect 22840 27752 23300 27872
rect -300 27480 160 27600
rect -300 27208 160 27328
rect 22840 27208 23300 27328
rect -300 26936 160 27056
rect -300 26664 160 26784
rect 22840 26664 23300 26784
rect -300 26392 160 26512
rect -300 26120 160 26240
rect 22840 26120 23300 26240
rect -300 25848 160 25968
rect -300 25576 160 25696
rect 22840 25576 23300 25696
rect -300 25304 160 25424
rect -300 25032 160 25152
rect 22840 25032 23300 25152
rect -300 24760 160 24880
rect -300 24488 160 24608
rect 22840 24488 23300 24608
rect -300 24216 160 24336
rect -300 23944 160 24064
rect 22840 23944 23300 24064
rect -300 23672 160 23792
rect -300 23400 160 23520
rect 22840 23400 23300 23520
rect -300 23128 160 23248
rect -300 22856 160 22976
rect 22840 22856 23300 22976
rect -300 22584 160 22704
rect -300 22312 160 22432
rect 22840 22312 23300 22432
rect -300 22040 160 22160
rect -300 21768 160 21888
rect 22840 21768 23300 21888
rect -300 21496 160 21616
rect -300 21224 160 21344
rect 22840 21224 23300 21344
rect -300 20952 160 21072
rect -300 20680 160 20800
rect 22840 20680 23300 20800
rect -300 20408 160 20528
rect -300 20136 160 20256
rect 22840 20136 23300 20256
rect -300 19864 160 19984
rect -300 19592 160 19712
rect 22840 19592 23300 19712
rect -300 19320 160 19440
rect -300 19048 160 19168
rect 22840 19048 23300 19168
rect -300 18776 160 18896
rect -300 18504 160 18624
rect 22840 18504 23300 18624
rect -300 18232 160 18352
rect -300 17960 160 18080
rect 22840 17960 23300 18080
rect -300 17688 160 17808
rect -300 17416 160 17536
rect 22840 17416 23300 17536
rect -300 17144 160 17264
rect -300 16872 160 16992
rect 22840 16872 23300 16992
rect -300 16600 160 16720
rect -300 16328 160 16448
rect 22840 16328 23300 16448
rect -300 16056 160 16176
rect -300 15784 160 15904
rect 22840 15784 23300 15904
rect -300 15512 160 15632
rect -300 15240 160 15360
rect 22840 15240 23300 15360
rect -300 14968 160 15088
rect -300 14696 160 14816
rect 22840 14696 23300 14816
rect -300 14424 160 14544
rect -300 14152 160 14272
rect 22840 14152 23300 14272
rect -300 13880 160 14000
rect -300 13608 160 13728
rect 22840 13608 23300 13728
rect -300 13336 160 13456
rect -300 13064 160 13184
rect 22840 13064 23300 13184
rect -300 12792 160 12912
rect -300 12520 160 12640
rect 22840 12520 23300 12640
rect -300 12248 160 12368
rect -300 11976 160 12096
rect 22840 11976 23300 12096
rect -300 11704 160 11824
rect -300 11432 160 11552
rect 22840 11432 23300 11552
rect -300 11160 160 11280
rect -300 10888 160 11008
rect 22840 10888 23300 11008
rect -300 10616 160 10736
rect -300 10344 160 10464
rect 22840 10344 23300 10464
rect -300 10072 160 10192
rect -300 9800 160 9920
rect 22840 9800 23300 9920
rect -300 9528 160 9648
rect -300 9256 160 9376
rect 22840 9256 23300 9376
rect -300 8984 160 9104
rect -300 8712 160 8832
rect 22840 8712 23300 8832
rect -300 8440 160 8560
rect -300 8168 160 8288
rect 22840 8168 23300 8288
rect -300 7896 160 8016
rect -300 7624 160 7744
rect 22840 7624 23300 7744
rect -300 7352 160 7472
rect -300 7080 160 7200
rect 22840 7080 23300 7200
rect -300 6808 160 6928
rect -300 6536 160 6656
rect 22840 6536 23300 6656
rect -300 6264 160 6384
rect -300 5992 160 6112
rect 22840 5992 23300 6112
rect -300 5720 160 5840
rect -300 5448 160 5568
rect 22840 5448 23300 5568
rect -300 5176 160 5296
rect -300 4904 160 5024
rect 22840 4904 23300 5024
rect 22840 4360 23300 4480
rect 22840 3816 23300 3936
rect 22840 3272 23300 3392
rect 22840 2728 23300 2848
rect 22840 2184 23300 2304
rect 22840 1640 23300 1760
rect 22840 1096 23300 1216
rect 22840 552 23300 672
<< obsm3 >>
rect 13 43728 22895 43893
rect 13 43448 22760 43728
rect 13 43184 22895 43448
rect 13 42904 22760 43184
rect 13 42640 22895 42904
rect 13 42360 22760 42640
rect 13 42096 22895 42360
rect 13 41816 22760 42096
rect 13 41552 22895 41816
rect 13 41272 22760 41552
rect 13 41008 22895 41272
rect 13 40728 22760 41008
rect 13 40464 22895 40728
rect 13 40184 22760 40464
rect 13 39920 22895 40184
rect 13 39648 22760 39920
rect 240 39640 22760 39648
rect 240 39376 22895 39640
rect 240 39096 22760 39376
rect 240 38832 22895 39096
rect 240 38552 22760 38832
rect 240 38288 22895 38552
rect 240 38008 22760 38288
rect 240 37744 22895 38008
rect 240 37464 22760 37744
rect 240 37200 22895 37464
rect 240 36920 22760 37200
rect 240 36656 22895 36920
rect 240 36376 22760 36656
rect 240 36112 22895 36376
rect 240 35832 22760 36112
rect 240 35568 22895 35832
rect 240 35288 22760 35568
rect 240 35024 22895 35288
rect 240 34744 22760 35024
rect 240 34480 22895 34744
rect 240 34200 22760 34480
rect 240 33936 22895 34200
rect 240 33656 22760 33936
rect 240 33392 22895 33656
rect 240 33112 22760 33392
rect 240 32848 22895 33112
rect 240 32568 22760 32848
rect 240 32304 22895 32568
rect 240 32024 22760 32304
rect 240 31760 22895 32024
rect 240 31480 22760 31760
rect 240 31216 22895 31480
rect 240 30936 22760 31216
rect 240 30672 22895 30936
rect 240 30392 22760 30672
rect 240 30128 22895 30392
rect 240 29848 22760 30128
rect 240 29584 22895 29848
rect 240 29304 22760 29584
rect 240 29040 22895 29304
rect 240 28760 22760 29040
rect 240 28496 22895 28760
rect 240 28216 22760 28496
rect 240 27952 22895 28216
rect 240 27672 22760 27952
rect 240 27408 22895 27672
rect 240 27128 22760 27408
rect 240 26864 22895 27128
rect 240 26584 22760 26864
rect 240 26320 22895 26584
rect 240 26040 22760 26320
rect 240 25776 22895 26040
rect 240 25496 22760 25776
rect 240 25232 22895 25496
rect 240 24952 22760 25232
rect 240 24688 22895 24952
rect 240 24408 22760 24688
rect 240 24144 22895 24408
rect 240 23864 22760 24144
rect 240 23600 22895 23864
rect 240 23320 22760 23600
rect 240 23056 22895 23320
rect 240 22776 22760 23056
rect 240 22512 22895 22776
rect 240 22232 22760 22512
rect 240 21968 22895 22232
rect 240 21688 22760 21968
rect 240 21424 22895 21688
rect 240 21144 22760 21424
rect 240 20880 22895 21144
rect 240 20600 22760 20880
rect 240 20336 22895 20600
rect 240 20056 22760 20336
rect 240 19792 22895 20056
rect 240 19512 22760 19792
rect 240 19248 22895 19512
rect 240 18968 22760 19248
rect 240 18704 22895 18968
rect 240 18424 22760 18704
rect 240 18160 22895 18424
rect 240 17880 22760 18160
rect 240 17616 22895 17880
rect 240 17336 22760 17616
rect 240 17072 22895 17336
rect 240 16792 22760 17072
rect 240 16528 22895 16792
rect 240 16248 22760 16528
rect 240 15984 22895 16248
rect 240 15704 22760 15984
rect 240 15440 22895 15704
rect 240 15160 22760 15440
rect 240 14896 22895 15160
rect 240 14616 22760 14896
rect 240 14352 22895 14616
rect 240 14072 22760 14352
rect 240 13808 22895 14072
rect 240 13528 22760 13808
rect 240 13264 22895 13528
rect 240 12984 22760 13264
rect 240 12720 22895 12984
rect 240 12440 22760 12720
rect 240 12176 22895 12440
rect 240 11896 22760 12176
rect 240 11632 22895 11896
rect 240 11352 22760 11632
rect 240 11088 22895 11352
rect 240 10808 22760 11088
rect 240 10544 22895 10808
rect 240 10264 22760 10544
rect 240 10000 22895 10264
rect 240 9720 22760 10000
rect 240 9456 22895 9720
rect 240 9176 22760 9456
rect 240 8912 22895 9176
rect 240 8632 22760 8912
rect 240 8368 22895 8632
rect 240 8088 22760 8368
rect 240 7824 22895 8088
rect 240 7544 22760 7824
rect 240 7280 22895 7544
rect 240 7000 22760 7280
rect 240 6736 22895 7000
rect 240 6456 22760 6736
rect 240 6192 22895 6456
rect 240 5912 22760 6192
rect 240 5648 22895 5912
rect 240 5368 22760 5648
rect 240 5104 22895 5368
rect 240 4824 22760 5104
rect 13 4560 22895 4824
rect 13 4280 22760 4560
rect 13 4016 22895 4280
rect 13 3736 22760 4016
rect 13 3472 22895 3736
rect 13 3192 22760 3472
rect 13 2928 22895 3192
rect 13 2648 22760 2928
rect 13 2384 22895 2648
rect 13 2104 22760 2384
rect 13 1840 22895 2104
rect 13 1560 22760 1840
rect 13 1296 22895 1560
rect 13 1016 22760 1296
rect 13 752 22895 1016
rect 13 472 22760 752
rect 13 35 22895 472
<< metal4 >>
rect 3543 1040 3863 43568
rect 6142 1040 6462 43568
rect 8741 1040 9061 43568
rect 11340 1040 11660 43568
rect 13939 1040 14259 43568
rect 16538 1040 16858 43568
rect 19137 1040 19457 43568
rect 21736 1040 22056 43568
<< obsm4 >>
rect 243 960 3463 43213
rect 3943 960 6062 43213
rect 6542 960 8661 43213
rect 9141 960 11260 43213
rect 11740 960 13859 43213
rect 14339 960 16458 43213
rect 16938 960 19057 43213
rect 19537 960 21469 43213
rect 243 35 21469 960
<< labels >>
rlabel metal3 s 22840 9256 23300 9376 6 Config_accessC_bit0
port 1 nsew signal output
rlabel metal3 s 22840 9800 23300 9920 6 Config_accessC_bit1
port 2 nsew signal output
rlabel metal3 s 22840 10344 23300 10464 6 Config_accessC_bit2
port 3 nsew signal output
rlabel metal3 s 22840 10888 23300 11008 6 Config_accessC_bit3
port 4 nsew signal output
rlabel metal3 s -300 17960 160 18080 4 E1END[0]
port 5 nsew signal input
rlabel metal3 s -300 18232 160 18352 4 E1END[1]
port 6 nsew signal input
rlabel metal3 s -300 18504 160 18624 4 E1END[2]
port 7 nsew signal input
rlabel metal3 s -300 18776 160 18896 4 E1END[3]
port 8 nsew signal input
rlabel metal3 s -300 21224 160 21344 4 E2END[0]
port 9 nsew signal input
rlabel metal3 s -300 21496 160 21616 4 E2END[1]
port 10 nsew signal input
rlabel metal3 s -300 21768 160 21888 4 E2END[2]
port 11 nsew signal input
rlabel metal3 s -300 22040 160 22160 4 E2END[3]
port 12 nsew signal input
rlabel metal3 s -300 22312 160 22432 4 E2END[4]
port 13 nsew signal input
rlabel metal3 s -300 22584 160 22704 4 E2END[5]
port 14 nsew signal input
rlabel metal3 s -300 22856 160 22976 4 E2END[6]
port 15 nsew signal input
rlabel metal3 s -300 23128 160 23248 4 E2END[7]
port 16 nsew signal input
rlabel metal3 s -300 19048 160 19168 4 E2MID[0]
port 17 nsew signal input
rlabel metal3 s -300 19320 160 19440 4 E2MID[1]
port 18 nsew signal input
rlabel metal3 s -300 19592 160 19712 4 E2MID[2]
port 19 nsew signal input
rlabel metal3 s -300 19864 160 19984 4 E2MID[3]
port 20 nsew signal input
rlabel metal3 s -300 20136 160 20256 4 E2MID[4]
port 21 nsew signal input
rlabel metal3 s -300 20408 160 20528 4 E2MID[5]
port 22 nsew signal input
rlabel metal3 s -300 20680 160 20800 4 E2MID[6]
port 23 nsew signal input
rlabel metal3 s -300 20952 160 21072 4 E2MID[7]
port 24 nsew signal input
rlabel metal3 s -300 27752 160 27872 4 E6END[0]
port 25 nsew signal input
rlabel metal3 s -300 30472 160 30592 4 E6END[10]
port 26 nsew signal input
rlabel metal3 s -300 30744 160 30864 4 E6END[11]
port 27 nsew signal input
rlabel metal3 s -300 28024 160 28144 4 E6END[1]
port 28 nsew signal input
rlabel metal3 s -300 28296 160 28416 4 E6END[2]
port 29 nsew signal input
rlabel metal3 s -300 28568 160 28688 4 E6END[3]
port 30 nsew signal input
rlabel metal3 s -300 28840 160 28960 4 E6END[4]
port 31 nsew signal input
rlabel metal3 s -300 29112 160 29232 4 E6END[5]
port 32 nsew signal input
rlabel metal3 s -300 29384 160 29504 4 E6END[6]
port 33 nsew signal input
rlabel metal3 s -300 29656 160 29776 4 E6END[7]
port 34 nsew signal input
rlabel metal3 s -300 29928 160 30048 4 E6END[8]
port 35 nsew signal input
rlabel metal3 s -300 30200 160 30320 4 E6END[9]
port 36 nsew signal input
rlabel metal3 s -300 23400 160 23520 4 EE4END[0]
port 37 nsew signal input
rlabel metal3 s -300 26120 160 26240 4 EE4END[10]
port 38 nsew signal input
rlabel metal3 s -300 26392 160 26512 4 EE4END[11]
port 39 nsew signal input
rlabel metal3 s -300 26664 160 26784 4 EE4END[12]
port 40 nsew signal input
rlabel metal3 s -300 26936 160 27056 4 EE4END[13]
port 41 nsew signal input
rlabel metal3 s -300 27208 160 27328 4 EE4END[14]
port 42 nsew signal input
rlabel metal3 s -300 27480 160 27600 4 EE4END[15]
port 43 nsew signal input
rlabel metal3 s -300 23672 160 23792 4 EE4END[1]
port 44 nsew signal input
rlabel metal3 s -300 23944 160 24064 4 EE4END[2]
port 45 nsew signal input
rlabel metal3 s -300 24216 160 24336 4 EE4END[3]
port 46 nsew signal input
rlabel metal3 s -300 24488 160 24608 4 EE4END[4]
port 47 nsew signal input
rlabel metal3 s -300 24760 160 24880 4 EE4END[5]
port 48 nsew signal input
rlabel metal3 s -300 25032 160 25152 4 EE4END[6]
port 49 nsew signal input
rlabel metal3 s -300 25304 160 25424 4 EE4END[7]
port 50 nsew signal input
rlabel metal3 s -300 25576 160 25696 4 EE4END[8]
port 51 nsew signal input
rlabel metal3 s -300 25848 160 25968 4 EE4END[9]
port 52 nsew signal input
rlabel metal3 s 22840 15784 23300 15904 6 FAB2RAM_A0_O0
port 53 nsew signal output
rlabel metal3 s 22840 16328 23300 16448 6 FAB2RAM_A0_O1
port 54 nsew signal output
rlabel metal3 s 22840 16872 23300 16992 6 FAB2RAM_A0_O2
port 55 nsew signal output
rlabel metal3 s 22840 17416 23300 17536 6 FAB2RAM_A0_O3
port 56 nsew signal output
rlabel metal3 s 22840 13608 23300 13728 6 FAB2RAM_A1_O0
port 57 nsew signal output
rlabel metal3 s 22840 14152 23300 14272 6 FAB2RAM_A1_O1
port 58 nsew signal output
rlabel metal3 s 22840 14696 23300 14816 6 FAB2RAM_A1_O2
port 59 nsew signal output
rlabel metal3 s 22840 15240 23300 15360 6 FAB2RAM_A1_O3
port 60 nsew signal output
rlabel metal3 s 22840 11432 23300 11552 6 FAB2RAM_C_O0
port 61 nsew signal output
rlabel metal3 s 22840 11976 23300 12096 6 FAB2RAM_C_O1
port 62 nsew signal output
rlabel metal3 s 22840 12520 23300 12640 6 FAB2RAM_C_O2
port 63 nsew signal output
rlabel metal3 s 22840 13064 23300 13184 6 FAB2RAM_C_O3
port 64 nsew signal output
rlabel metal3 s 22840 24488 23300 24608 6 FAB2RAM_D0_O0
port 65 nsew signal output
rlabel metal3 s 22840 25032 23300 25152 6 FAB2RAM_D0_O1
port 66 nsew signal output
rlabel metal3 s 22840 25576 23300 25696 6 FAB2RAM_D0_O2
port 67 nsew signal output
rlabel metal3 s 22840 26120 23300 26240 6 FAB2RAM_D0_O3
port 68 nsew signal output
rlabel metal3 s 22840 22312 23300 22432 6 FAB2RAM_D1_O0
port 69 nsew signal output
rlabel metal3 s 22840 22856 23300 22976 6 FAB2RAM_D1_O1
port 70 nsew signal output
rlabel metal3 s 22840 23400 23300 23520 6 FAB2RAM_D1_O2
port 71 nsew signal output
rlabel metal3 s 22840 23944 23300 24064 6 FAB2RAM_D1_O3
port 72 nsew signal output
rlabel metal3 s 22840 20136 23300 20256 6 FAB2RAM_D2_O0
port 73 nsew signal output
rlabel metal3 s 22840 20680 23300 20800 6 FAB2RAM_D2_O1
port 74 nsew signal output
rlabel metal3 s 22840 21224 23300 21344 6 FAB2RAM_D2_O2
port 75 nsew signal output
rlabel metal3 s 22840 21768 23300 21888 6 FAB2RAM_D2_O3
port 76 nsew signal output
rlabel metal3 s 22840 17960 23300 18080 6 FAB2RAM_D3_O0
port 77 nsew signal output
rlabel metal3 s 22840 18504 23300 18624 6 FAB2RAM_D3_O1
port 78 nsew signal output
rlabel metal3 s 22840 19048 23300 19168 6 FAB2RAM_D3_O2
port 79 nsew signal output
rlabel metal3 s 22840 19592 23300 19712 6 FAB2RAM_D3_O3
port 80 nsew signal output
rlabel metal3 s -300 31016 160 31136 4 FrameData[0]
port 81 nsew signal input
rlabel metal3 s -300 33736 160 33856 4 FrameData[10]
port 82 nsew signal input
rlabel metal3 s -300 34008 160 34128 4 FrameData[11]
port 83 nsew signal input
rlabel metal3 s -300 34280 160 34400 4 FrameData[12]
port 84 nsew signal input
rlabel metal3 s -300 34552 160 34672 4 FrameData[13]
port 85 nsew signal input
rlabel metal3 s -300 34824 160 34944 4 FrameData[14]
port 86 nsew signal input
rlabel metal3 s -300 35096 160 35216 4 FrameData[15]
port 87 nsew signal input
rlabel metal3 s -300 35368 160 35488 4 FrameData[16]
port 88 nsew signal input
rlabel metal3 s -300 35640 160 35760 4 FrameData[17]
port 89 nsew signal input
rlabel metal3 s -300 35912 160 36032 4 FrameData[18]
port 90 nsew signal input
rlabel metal3 s -300 36184 160 36304 4 FrameData[19]
port 91 nsew signal input
rlabel metal3 s -300 31288 160 31408 4 FrameData[1]
port 92 nsew signal input
rlabel metal3 s -300 36456 160 36576 4 FrameData[20]
port 93 nsew signal input
rlabel metal3 s -300 36728 160 36848 4 FrameData[21]
port 94 nsew signal input
rlabel metal3 s -300 37000 160 37120 4 FrameData[22]
port 95 nsew signal input
rlabel metal3 s -300 37272 160 37392 4 FrameData[23]
port 96 nsew signal input
rlabel metal3 s -300 37544 160 37664 4 FrameData[24]
port 97 nsew signal input
rlabel metal3 s -300 37816 160 37936 4 FrameData[25]
port 98 nsew signal input
rlabel metal3 s -300 38088 160 38208 4 FrameData[26]
port 99 nsew signal input
rlabel metal3 s -300 38360 160 38480 4 FrameData[27]
port 100 nsew signal input
rlabel metal3 s -300 38632 160 38752 4 FrameData[28]
port 101 nsew signal input
rlabel metal3 s -300 38904 160 39024 4 FrameData[29]
port 102 nsew signal input
rlabel metal3 s -300 31560 160 31680 4 FrameData[2]
port 103 nsew signal input
rlabel metal3 s -300 39176 160 39296 4 FrameData[30]
port 104 nsew signal input
rlabel metal3 s -300 39448 160 39568 4 FrameData[31]
port 105 nsew signal input
rlabel metal3 s -300 31832 160 31952 4 FrameData[3]
port 106 nsew signal input
rlabel metal3 s -300 32104 160 32224 4 FrameData[4]
port 107 nsew signal input
rlabel metal3 s -300 32376 160 32496 4 FrameData[5]
port 108 nsew signal input
rlabel metal3 s -300 32648 160 32768 4 FrameData[6]
port 109 nsew signal input
rlabel metal3 s -300 32920 160 33040 4 FrameData[7]
port 110 nsew signal input
rlabel metal3 s -300 33192 160 33312 4 FrameData[8]
port 111 nsew signal input
rlabel metal3 s -300 33464 160 33584 4 FrameData[9]
port 112 nsew signal input
rlabel metal3 s 22840 26664 23300 26784 6 FrameData_O[0]
port 113 nsew signal output
rlabel metal3 s 22840 32104 23300 32224 6 FrameData_O[10]
port 114 nsew signal output
rlabel metal3 s 22840 32648 23300 32768 6 FrameData_O[11]
port 115 nsew signal output
rlabel metal3 s 22840 33192 23300 33312 6 FrameData_O[12]
port 116 nsew signal output
rlabel metal3 s 22840 33736 23300 33856 6 FrameData_O[13]
port 117 nsew signal output
rlabel metal3 s 22840 34280 23300 34400 6 FrameData_O[14]
port 118 nsew signal output
rlabel metal3 s 22840 34824 23300 34944 6 FrameData_O[15]
port 119 nsew signal output
rlabel metal3 s 22840 35368 23300 35488 6 FrameData_O[16]
port 120 nsew signal output
rlabel metal3 s 22840 35912 23300 36032 6 FrameData_O[17]
port 121 nsew signal output
rlabel metal3 s 22840 36456 23300 36576 6 FrameData_O[18]
port 122 nsew signal output
rlabel metal3 s 22840 37000 23300 37120 6 FrameData_O[19]
port 123 nsew signal output
rlabel metal3 s 22840 27208 23300 27328 6 FrameData_O[1]
port 124 nsew signal output
rlabel metal3 s 22840 37544 23300 37664 6 FrameData_O[20]
port 125 nsew signal output
rlabel metal3 s 22840 38088 23300 38208 6 FrameData_O[21]
port 126 nsew signal output
rlabel metal3 s 22840 38632 23300 38752 6 FrameData_O[22]
port 127 nsew signal output
rlabel metal3 s 22840 39176 23300 39296 6 FrameData_O[23]
port 128 nsew signal output
rlabel metal3 s 22840 39720 23300 39840 6 FrameData_O[24]
port 129 nsew signal output
rlabel metal3 s 22840 40264 23300 40384 6 FrameData_O[25]
port 130 nsew signal output
rlabel metal3 s 22840 40808 23300 40928 6 FrameData_O[26]
port 131 nsew signal output
rlabel metal3 s 22840 41352 23300 41472 6 FrameData_O[27]
port 132 nsew signal output
rlabel metal3 s 22840 41896 23300 42016 6 FrameData_O[28]
port 133 nsew signal output
rlabel metal3 s 22840 42440 23300 42560 6 FrameData_O[29]
port 134 nsew signal output
rlabel metal3 s 22840 27752 23300 27872 6 FrameData_O[2]
port 135 nsew signal output
rlabel metal3 s 22840 42984 23300 43104 6 FrameData_O[30]
port 136 nsew signal output
rlabel metal3 s 22840 43528 23300 43648 6 FrameData_O[31]
port 137 nsew signal output
rlabel metal3 s 22840 28296 23300 28416 6 FrameData_O[3]
port 138 nsew signal output
rlabel metal3 s 22840 28840 23300 28960 6 FrameData_O[4]
port 139 nsew signal output
rlabel metal3 s 22840 29384 23300 29504 6 FrameData_O[5]
port 140 nsew signal output
rlabel metal3 s 22840 29928 23300 30048 6 FrameData_O[6]
port 141 nsew signal output
rlabel metal3 s 22840 30472 23300 30592 6 FrameData_O[7]
port 142 nsew signal output
rlabel metal3 s 22840 31016 23300 31136 6 FrameData_O[8]
port 143 nsew signal output
rlabel metal3 s 22840 31560 23300 31680 6 FrameData_O[9]
port 144 nsew signal output
rlabel metal2 s 16394 -300 16450 160 8 FrameStrobe[0]
port 145 nsew signal input
rlabel metal2 s 18234 -300 18290 160 8 FrameStrobe[10]
port 146 nsew signal input
rlabel metal2 s 18418 -300 18474 160 8 FrameStrobe[11]
port 147 nsew signal input
rlabel metal2 s 18602 -300 18658 160 8 FrameStrobe[12]
port 148 nsew signal input
rlabel metal2 s 18786 -300 18842 160 8 FrameStrobe[13]
port 149 nsew signal input
rlabel metal2 s 18970 -300 19026 160 8 FrameStrobe[14]
port 150 nsew signal input
rlabel metal2 s 19154 -300 19210 160 8 FrameStrobe[15]
port 151 nsew signal input
rlabel metal2 s 19338 -300 19394 160 8 FrameStrobe[16]
port 152 nsew signal input
rlabel metal2 s 19522 -300 19578 160 8 FrameStrobe[17]
port 153 nsew signal input
rlabel metal2 s 19706 -300 19762 160 8 FrameStrobe[18]
port 154 nsew signal input
rlabel metal2 s 19890 -300 19946 160 8 FrameStrobe[19]
port 155 nsew signal input
rlabel metal2 s 16578 -300 16634 160 8 FrameStrobe[1]
port 156 nsew signal input
rlabel metal2 s 16762 -300 16818 160 8 FrameStrobe[2]
port 157 nsew signal input
rlabel metal2 s 16946 -300 17002 160 8 FrameStrobe[3]
port 158 nsew signal input
rlabel metal2 s 17130 -300 17186 160 8 FrameStrobe[4]
port 159 nsew signal input
rlabel metal2 s 17314 -300 17370 160 8 FrameStrobe[5]
port 160 nsew signal input
rlabel metal2 s 17498 -300 17554 160 8 FrameStrobe[6]
port 161 nsew signal input
rlabel metal2 s 17682 -300 17738 160 8 FrameStrobe[7]
port 162 nsew signal input
rlabel metal2 s 17866 -300 17922 160 8 FrameStrobe[8]
port 163 nsew signal input
rlabel metal2 s 18050 -300 18106 160 8 FrameStrobe[9]
port 164 nsew signal input
rlabel metal2 s 16394 44540 16450 45000 6 FrameStrobe_O[0]
port 165 nsew signal output
rlabel metal2 s 18234 44540 18290 45000 6 FrameStrobe_O[10]
port 166 nsew signal output
rlabel metal2 s 18418 44540 18474 45000 6 FrameStrobe_O[11]
port 167 nsew signal output
rlabel metal2 s 18602 44540 18658 45000 6 FrameStrobe_O[12]
port 168 nsew signal output
rlabel metal2 s 18786 44540 18842 45000 6 FrameStrobe_O[13]
port 169 nsew signal output
rlabel metal2 s 18970 44540 19026 45000 6 FrameStrobe_O[14]
port 170 nsew signal output
rlabel metal2 s 19154 44540 19210 45000 6 FrameStrobe_O[15]
port 171 nsew signal output
rlabel metal2 s 19338 44540 19394 45000 6 FrameStrobe_O[16]
port 172 nsew signal output
rlabel metal2 s 19522 44540 19578 45000 6 FrameStrobe_O[17]
port 173 nsew signal output
rlabel metal2 s 19706 44540 19762 45000 6 FrameStrobe_O[18]
port 174 nsew signal output
rlabel metal2 s 19890 44540 19946 45000 6 FrameStrobe_O[19]
port 175 nsew signal output
rlabel metal2 s 16578 44540 16634 45000 6 FrameStrobe_O[1]
port 176 nsew signal output
rlabel metal2 s 16762 44540 16818 45000 6 FrameStrobe_O[2]
port 177 nsew signal output
rlabel metal2 s 16946 44540 17002 45000 6 FrameStrobe_O[3]
port 178 nsew signal output
rlabel metal2 s 17130 44540 17186 45000 6 FrameStrobe_O[4]
port 179 nsew signal output
rlabel metal2 s 17314 44540 17370 45000 6 FrameStrobe_O[5]
port 180 nsew signal output
rlabel metal2 s 17498 44540 17554 45000 6 FrameStrobe_O[6]
port 181 nsew signal output
rlabel metal2 s 17682 44540 17738 45000 6 FrameStrobe_O[7]
port 182 nsew signal output
rlabel metal2 s 17866 44540 17922 45000 6 FrameStrobe_O[8]
port 183 nsew signal output
rlabel metal2 s 18050 44540 18106 45000 6 FrameStrobe_O[9]
port 184 nsew signal output
rlabel metal2 s 2962 44540 3018 45000 6 N1BEG[0]
port 185 nsew signal output
rlabel metal2 s 3146 44540 3202 45000 6 N1BEG[1]
port 186 nsew signal output
rlabel metal2 s 3330 44540 3386 45000 6 N1BEG[2]
port 187 nsew signal output
rlabel metal2 s 3514 44540 3570 45000 6 N1BEG[3]
port 188 nsew signal output
rlabel metal2 s 2962 -300 3018 160 8 N1END[0]
port 189 nsew signal input
rlabel metal2 s 3146 -300 3202 160 8 N1END[1]
port 190 nsew signal input
rlabel metal2 s 3330 -300 3386 160 8 N1END[2]
port 191 nsew signal input
rlabel metal2 s 3514 -300 3570 160 8 N1END[3]
port 192 nsew signal input
rlabel metal2 s 3698 44540 3754 45000 6 N2BEG[0]
port 193 nsew signal output
rlabel metal2 s 3882 44540 3938 45000 6 N2BEG[1]
port 194 nsew signal output
rlabel metal2 s 4066 44540 4122 45000 6 N2BEG[2]
port 195 nsew signal output
rlabel metal2 s 4250 44540 4306 45000 6 N2BEG[3]
port 196 nsew signal output
rlabel metal2 s 4434 44540 4490 45000 6 N2BEG[4]
port 197 nsew signal output
rlabel metal2 s 4618 44540 4674 45000 6 N2BEG[5]
port 198 nsew signal output
rlabel metal2 s 4802 44540 4858 45000 6 N2BEG[6]
port 199 nsew signal output
rlabel metal2 s 4986 44540 5042 45000 6 N2BEG[7]
port 200 nsew signal output
rlabel metal2 s 5170 44540 5226 45000 6 N2BEGb[0]
port 201 nsew signal output
rlabel metal2 s 5354 44540 5410 45000 6 N2BEGb[1]
port 202 nsew signal output
rlabel metal2 s 5538 44540 5594 45000 6 N2BEGb[2]
port 203 nsew signal output
rlabel metal2 s 5722 44540 5778 45000 6 N2BEGb[3]
port 204 nsew signal output
rlabel metal2 s 5906 44540 5962 45000 6 N2BEGb[4]
port 205 nsew signal output
rlabel metal2 s 6090 44540 6146 45000 6 N2BEGb[5]
port 206 nsew signal output
rlabel metal2 s 6274 44540 6330 45000 6 N2BEGb[6]
port 207 nsew signal output
rlabel metal2 s 6458 44540 6514 45000 6 N2BEGb[7]
port 208 nsew signal output
rlabel metal2 s 5170 -300 5226 160 8 N2END[0]
port 209 nsew signal input
rlabel metal2 s 5354 -300 5410 160 8 N2END[1]
port 210 nsew signal input
rlabel metal2 s 5538 -300 5594 160 8 N2END[2]
port 211 nsew signal input
rlabel metal2 s 5722 -300 5778 160 8 N2END[3]
port 212 nsew signal input
rlabel metal2 s 5906 -300 5962 160 8 N2END[4]
port 213 nsew signal input
rlabel metal2 s 6090 -300 6146 160 8 N2END[5]
port 214 nsew signal input
rlabel metal2 s 6274 -300 6330 160 8 N2END[6]
port 215 nsew signal input
rlabel metal2 s 6458 -300 6514 160 8 N2END[7]
port 216 nsew signal input
rlabel metal2 s 3698 -300 3754 160 8 N2MID[0]
port 217 nsew signal input
rlabel metal2 s 3882 -300 3938 160 8 N2MID[1]
port 218 nsew signal input
rlabel metal2 s 4066 -300 4122 160 8 N2MID[2]
port 219 nsew signal input
rlabel metal2 s 4250 -300 4306 160 8 N2MID[3]
port 220 nsew signal input
rlabel metal2 s 4434 -300 4490 160 8 N2MID[4]
port 221 nsew signal input
rlabel metal2 s 4618 -300 4674 160 8 N2MID[5]
port 222 nsew signal input
rlabel metal2 s 4802 -300 4858 160 8 N2MID[6]
port 223 nsew signal input
rlabel metal2 s 4986 -300 5042 160 8 N2MID[7]
port 224 nsew signal input
rlabel metal2 s 6642 44540 6698 45000 6 N4BEG[0]
port 225 nsew signal output
rlabel metal2 s 8482 44540 8538 45000 6 N4BEG[10]
port 226 nsew signal output
rlabel metal2 s 8666 44540 8722 45000 6 N4BEG[11]
port 227 nsew signal output
rlabel metal2 s 8850 44540 8906 45000 6 N4BEG[12]
port 228 nsew signal output
rlabel metal2 s 9034 44540 9090 45000 6 N4BEG[13]
port 229 nsew signal output
rlabel metal2 s 9218 44540 9274 45000 6 N4BEG[14]
port 230 nsew signal output
rlabel metal2 s 9402 44540 9458 45000 6 N4BEG[15]
port 231 nsew signal output
rlabel metal2 s 6826 44540 6882 45000 6 N4BEG[1]
port 232 nsew signal output
rlabel metal2 s 7010 44540 7066 45000 6 N4BEG[2]
port 233 nsew signal output
rlabel metal2 s 7194 44540 7250 45000 6 N4BEG[3]
port 234 nsew signal output
rlabel metal2 s 7378 44540 7434 45000 6 N4BEG[4]
port 235 nsew signal output
rlabel metal2 s 7562 44540 7618 45000 6 N4BEG[5]
port 236 nsew signal output
rlabel metal2 s 7746 44540 7802 45000 6 N4BEG[6]
port 237 nsew signal output
rlabel metal2 s 7930 44540 7986 45000 6 N4BEG[7]
port 238 nsew signal output
rlabel metal2 s 8114 44540 8170 45000 6 N4BEG[8]
port 239 nsew signal output
rlabel metal2 s 8298 44540 8354 45000 6 N4BEG[9]
port 240 nsew signal output
rlabel metal2 s 6642 -300 6698 160 8 N4END[0]
port 241 nsew signal input
rlabel metal2 s 8482 -300 8538 160 8 N4END[10]
port 242 nsew signal input
rlabel metal2 s 8666 -300 8722 160 8 N4END[11]
port 243 nsew signal input
rlabel metal2 s 8850 -300 8906 160 8 N4END[12]
port 244 nsew signal input
rlabel metal2 s 9034 -300 9090 160 8 N4END[13]
port 245 nsew signal input
rlabel metal2 s 9218 -300 9274 160 8 N4END[14]
port 246 nsew signal input
rlabel metal2 s 9402 -300 9458 160 8 N4END[15]
port 247 nsew signal input
rlabel metal2 s 6826 -300 6882 160 8 N4END[1]
port 248 nsew signal input
rlabel metal2 s 7010 -300 7066 160 8 N4END[2]
port 249 nsew signal input
rlabel metal2 s 7194 -300 7250 160 8 N4END[3]
port 250 nsew signal input
rlabel metal2 s 7378 -300 7434 160 8 N4END[4]
port 251 nsew signal input
rlabel metal2 s 7562 -300 7618 160 8 N4END[5]
port 252 nsew signal input
rlabel metal2 s 7746 -300 7802 160 8 N4END[6]
port 253 nsew signal input
rlabel metal2 s 7930 -300 7986 160 8 N4END[7]
port 254 nsew signal input
rlabel metal2 s 8114 -300 8170 160 8 N4END[8]
port 255 nsew signal input
rlabel metal2 s 8298 -300 8354 160 8 N4END[9]
port 256 nsew signal input
rlabel metal3 s 22840 7080 23300 7200 6 RAM2FAB_D0_I0
port 257 nsew signal input
rlabel metal3 s 22840 7624 23300 7744 6 RAM2FAB_D0_I1
port 258 nsew signal input
rlabel metal3 s 22840 8168 23300 8288 6 RAM2FAB_D0_I2
port 259 nsew signal input
rlabel metal3 s 22840 8712 23300 8832 6 RAM2FAB_D0_I3
port 260 nsew signal input
rlabel metal3 s 22840 4904 23300 5024 6 RAM2FAB_D1_I0
port 261 nsew signal input
rlabel metal3 s 22840 5448 23300 5568 6 RAM2FAB_D1_I1
port 262 nsew signal input
rlabel metal3 s 22840 5992 23300 6112 6 RAM2FAB_D1_I2
port 263 nsew signal input
rlabel metal3 s 22840 6536 23300 6656 6 RAM2FAB_D1_I3
port 264 nsew signal input
rlabel metal3 s 22840 2728 23300 2848 6 RAM2FAB_D2_I0
port 265 nsew signal input
rlabel metal3 s 22840 3272 23300 3392 6 RAM2FAB_D2_I1
port 266 nsew signal input
rlabel metal3 s 22840 3816 23300 3936 6 RAM2FAB_D2_I2
port 267 nsew signal input
rlabel metal3 s 22840 4360 23300 4480 6 RAM2FAB_D2_I3
port 268 nsew signal input
rlabel metal3 s 22840 552 23300 672 6 RAM2FAB_D3_I0
port 269 nsew signal input
rlabel metal3 s 22840 1096 23300 1216 6 RAM2FAB_D3_I1
port 270 nsew signal input
rlabel metal3 s 22840 1640 23300 1760 6 RAM2FAB_D3_I2
port 271 nsew signal input
rlabel metal3 s 22840 2184 23300 2304 6 RAM2FAB_D3_I3
port 272 nsew signal input
rlabel metal2 s 9586 -300 9642 160 8 S1BEG[0]
port 273 nsew signal output
rlabel metal2 s 9770 -300 9826 160 8 S1BEG[1]
port 274 nsew signal output
rlabel metal2 s 9954 -300 10010 160 8 S1BEG[2]
port 275 nsew signal output
rlabel metal2 s 10138 -300 10194 160 8 S1BEG[3]
port 276 nsew signal output
rlabel metal2 s 9586 44540 9642 45000 6 S1END[0]
port 277 nsew signal input
rlabel metal2 s 9770 44540 9826 45000 6 S1END[1]
port 278 nsew signal input
rlabel metal2 s 9954 44540 10010 45000 6 S1END[2]
port 279 nsew signal input
rlabel metal2 s 10138 44540 10194 45000 6 S1END[3]
port 280 nsew signal input
rlabel metal2 s 11794 -300 11850 160 8 S2BEG[0]
port 281 nsew signal output
rlabel metal2 s 11978 -300 12034 160 8 S2BEG[1]
port 282 nsew signal output
rlabel metal2 s 12162 -300 12218 160 8 S2BEG[2]
port 283 nsew signal output
rlabel metal2 s 12346 -300 12402 160 8 S2BEG[3]
port 284 nsew signal output
rlabel metal2 s 12530 -300 12586 160 8 S2BEG[4]
port 285 nsew signal output
rlabel metal2 s 12714 -300 12770 160 8 S2BEG[5]
port 286 nsew signal output
rlabel metal2 s 12898 -300 12954 160 8 S2BEG[6]
port 287 nsew signal output
rlabel metal2 s 13082 -300 13138 160 8 S2BEG[7]
port 288 nsew signal output
rlabel metal2 s 10322 -300 10378 160 8 S2BEGb[0]
port 289 nsew signal output
rlabel metal2 s 10506 -300 10562 160 8 S2BEGb[1]
port 290 nsew signal output
rlabel metal2 s 10690 -300 10746 160 8 S2BEGb[2]
port 291 nsew signal output
rlabel metal2 s 10874 -300 10930 160 8 S2BEGb[3]
port 292 nsew signal output
rlabel metal2 s 11058 -300 11114 160 8 S2BEGb[4]
port 293 nsew signal output
rlabel metal2 s 11242 -300 11298 160 8 S2BEGb[5]
port 294 nsew signal output
rlabel metal2 s 11426 -300 11482 160 8 S2BEGb[6]
port 295 nsew signal output
rlabel metal2 s 11610 -300 11666 160 8 S2BEGb[7]
port 296 nsew signal output
rlabel metal2 s 10322 44540 10378 45000 6 S2END[0]
port 297 nsew signal input
rlabel metal2 s 10506 44540 10562 45000 6 S2END[1]
port 298 nsew signal input
rlabel metal2 s 10690 44540 10746 45000 6 S2END[2]
port 299 nsew signal input
rlabel metal2 s 10874 44540 10930 45000 6 S2END[3]
port 300 nsew signal input
rlabel metal2 s 11058 44540 11114 45000 6 S2END[4]
port 301 nsew signal input
rlabel metal2 s 11242 44540 11298 45000 6 S2END[5]
port 302 nsew signal input
rlabel metal2 s 11426 44540 11482 45000 6 S2END[6]
port 303 nsew signal input
rlabel metal2 s 11610 44540 11666 45000 6 S2END[7]
port 304 nsew signal input
rlabel metal2 s 11794 44540 11850 45000 6 S2MID[0]
port 305 nsew signal input
rlabel metal2 s 11978 44540 12034 45000 6 S2MID[1]
port 306 nsew signal input
rlabel metal2 s 12162 44540 12218 45000 6 S2MID[2]
port 307 nsew signal input
rlabel metal2 s 12346 44540 12402 45000 6 S2MID[3]
port 308 nsew signal input
rlabel metal2 s 12530 44540 12586 45000 6 S2MID[4]
port 309 nsew signal input
rlabel metal2 s 12714 44540 12770 45000 6 S2MID[5]
port 310 nsew signal input
rlabel metal2 s 12898 44540 12954 45000 6 S2MID[6]
port 311 nsew signal input
rlabel metal2 s 13082 44540 13138 45000 6 S2MID[7]
port 312 nsew signal input
rlabel metal2 s 13266 -300 13322 160 8 S4BEG[0]
port 313 nsew signal output
rlabel metal2 s 15106 -300 15162 160 8 S4BEG[10]
port 314 nsew signal output
rlabel metal2 s 15290 -300 15346 160 8 S4BEG[11]
port 315 nsew signal output
rlabel metal2 s 15474 -300 15530 160 8 S4BEG[12]
port 316 nsew signal output
rlabel metal2 s 15658 -300 15714 160 8 S4BEG[13]
port 317 nsew signal output
rlabel metal2 s 15842 -300 15898 160 8 S4BEG[14]
port 318 nsew signal output
rlabel metal2 s 16026 -300 16082 160 8 S4BEG[15]
port 319 nsew signal output
rlabel metal2 s 13450 -300 13506 160 8 S4BEG[1]
port 320 nsew signal output
rlabel metal2 s 13634 -300 13690 160 8 S4BEG[2]
port 321 nsew signal output
rlabel metal2 s 13818 -300 13874 160 8 S4BEG[3]
port 322 nsew signal output
rlabel metal2 s 14002 -300 14058 160 8 S4BEG[4]
port 323 nsew signal output
rlabel metal2 s 14186 -300 14242 160 8 S4BEG[5]
port 324 nsew signal output
rlabel metal2 s 14370 -300 14426 160 8 S4BEG[6]
port 325 nsew signal output
rlabel metal2 s 14554 -300 14610 160 8 S4BEG[7]
port 326 nsew signal output
rlabel metal2 s 14738 -300 14794 160 8 S4BEG[8]
port 327 nsew signal output
rlabel metal2 s 14922 -300 14978 160 8 S4BEG[9]
port 328 nsew signal output
rlabel metal2 s 13266 44540 13322 45000 6 S4END[0]
port 329 nsew signal input
rlabel metal2 s 15106 44540 15162 45000 6 S4END[10]
port 330 nsew signal input
rlabel metal2 s 15290 44540 15346 45000 6 S4END[11]
port 331 nsew signal input
rlabel metal2 s 15474 44540 15530 45000 6 S4END[12]
port 332 nsew signal input
rlabel metal2 s 15658 44540 15714 45000 6 S4END[13]
port 333 nsew signal input
rlabel metal2 s 15842 44540 15898 45000 6 S4END[14]
port 334 nsew signal input
rlabel metal2 s 16026 44540 16082 45000 6 S4END[15]
port 335 nsew signal input
rlabel metal2 s 13450 44540 13506 45000 6 S4END[1]
port 336 nsew signal input
rlabel metal2 s 13634 44540 13690 45000 6 S4END[2]
port 337 nsew signal input
rlabel metal2 s 13818 44540 13874 45000 6 S4END[3]
port 338 nsew signal input
rlabel metal2 s 14002 44540 14058 45000 6 S4END[4]
port 339 nsew signal input
rlabel metal2 s 14186 44540 14242 45000 6 S4END[5]
port 340 nsew signal input
rlabel metal2 s 14370 44540 14426 45000 6 S4END[6]
port 341 nsew signal input
rlabel metal2 s 14554 44540 14610 45000 6 S4END[7]
port 342 nsew signal input
rlabel metal2 s 14738 44540 14794 45000 6 S4END[8]
port 343 nsew signal input
rlabel metal2 s 14922 44540 14978 45000 6 S4END[9]
port 344 nsew signal input
rlabel metal2 s 16210 -300 16266 160 8 UserCLK
port 345 nsew signal input
rlabel metal2 s 16210 44540 16266 45000 6 UserCLKo
port 346 nsew signal output
rlabel metal4 s 6142 1040 6462 43568 6 VGND
port 347 nsew ground bidirectional
rlabel metal4 s 11340 1040 11660 43568 6 VGND
port 347 nsew ground bidirectional
rlabel metal4 s 16538 1040 16858 43568 6 VGND
port 347 nsew ground bidirectional
rlabel metal4 s 21736 1040 22056 43568 6 VGND
port 347 nsew ground bidirectional
rlabel metal4 s 3543 1040 3863 43568 6 VPWR
port 348 nsew power bidirectional
rlabel metal4 s 8741 1040 9061 43568 6 VPWR
port 348 nsew power bidirectional
rlabel metal4 s 13939 1040 14259 43568 6 VPWR
port 348 nsew power bidirectional
rlabel metal4 s 19137 1040 19457 43568 6 VPWR
port 348 nsew power bidirectional
rlabel metal3 s -300 4904 160 5024 4 W1BEG[0]
port 349 nsew signal output
rlabel metal3 s -300 5176 160 5296 4 W1BEG[1]
port 350 nsew signal output
rlabel metal3 s -300 5448 160 5568 4 W1BEG[2]
port 351 nsew signal output
rlabel metal3 s -300 5720 160 5840 4 W1BEG[3]
port 352 nsew signal output
rlabel metal3 s -300 5992 160 6112 4 W2BEG[0]
port 353 nsew signal output
rlabel metal3 s -300 6264 160 6384 4 W2BEG[1]
port 354 nsew signal output
rlabel metal3 s -300 6536 160 6656 4 W2BEG[2]
port 355 nsew signal output
rlabel metal3 s -300 6808 160 6928 4 W2BEG[3]
port 356 nsew signal output
rlabel metal3 s -300 7080 160 7200 4 W2BEG[4]
port 357 nsew signal output
rlabel metal3 s -300 7352 160 7472 4 W2BEG[5]
port 358 nsew signal output
rlabel metal3 s -300 7624 160 7744 4 W2BEG[6]
port 359 nsew signal output
rlabel metal3 s -300 7896 160 8016 4 W2BEG[7]
port 360 nsew signal output
rlabel metal3 s -300 8168 160 8288 4 W2BEGb[0]
port 361 nsew signal output
rlabel metal3 s -300 8440 160 8560 4 W2BEGb[1]
port 362 nsew signal output
rlabel metal3 s -300 8712 160 8832 4 W2BEGb[2]
port 363 nsew signal output
rlabel metal3 s -300 8984 160 9104 4 W2BEGb[3]
port 364 nsew signal output
rlabel metal3 s -300 9256 160 9376 4 W2BEGb[4]
port 365 nsew signal output
rlabel metal3 s -300 9528 160 9648 4 W2BEGb[5]
port 366 nsew signal output
rlabel metal3 s -300 9800 160 9920 4 W2BEGb[6]
port 367 nsew signal output
rlabel metal3 s -300 10072 160 10192 4 W2BEGb[7]
port 368 nsew signal output
rlabel metal3 s -300 14696 160 14816 4 W6BEG[0]
port 369 nsew signal output
rlabel metal3 s -300 17416 160 17536 4 W6BEG[10]
port 370 nsew signal output
rlabel metal3 s -300 17688 160 17808 4 W6BEG[11]
port 371 nsew signal output
rlabel metal3 s -300 14968 160 15088 4 W6BEG[1]
port 372 nsew signal output
rlabel metal3 s -300 15240 160 15360 4 W6BEG[2]
port 373 nsew signal output
rlabel metal3 s -300 15512 160 15632 4 W6BEG[3]
port 374 nsew signal output
rlabel metal3 s -300 15784 160 15904 4 W6BEG[4]
port 375 nsew signal output
rlabel metal3 s -300 16056 160 16176 4 W6BEG[5]
port 376 nsew signal output
rlabel metal3 s -300 16328 160 16448 4 W6BEG[6]
port 377 nsew signal output
rlabel metal3 s -300 16600 160 16720 4 W6BEG[7]
port 378 nsew signal output
rlabel metal3 s -300 16872 160 16992 4 W6BEG[8]
port 379 nsew signal output
rlabel metal3 s -300 17144 160 17264 4 W6BEG[9]
port 380 nsew signal output
rlabel metal3 s -300 10344 160 10464 4 WW4BEG[0]
port 381 nsew signal output
rlabel metal3 s -300 13064 160 13184 4 WW4BEG[10]
port 382 nsew signal output
rlabel metal3 s -300 13336 160 13456 4 WW4BEG[11]
port 383 nsew signal output
rlabel metal3 s -300 13608 160 13728 4 WW4BEG[12]
port 384 nsew signal output
rlabel metal3 s -300 13880 160 14000 4 WW4BEG[13]
port 385 nsew signal output
rlabel metal3 s -300 14152 160 14272 4 WW4BEG[14]
port 386 nsew signal output
rlabel metal3 s -300 14424 160 14544 4 WW4BEG[15]
port 387 nsew signal output
rlabel metal3 s -300 10616 160 10736 4 WW4BEG[1]
port 388 nsew signal output
rlabel metal3 s -300 10888 160 11008 4 WW4BEG[2]
port 389 nsew signal output
rlabel metal3 s -300 11160 160 11280 4 WW4BEG[3]
port 390 nsew signal output
rlabel metal3 s -300 11432 160 11552 4 WW4BEG[4]
port 391 nsew signal output
rlabel metal3 s -300 11704 160 11824 4 WW4BEG[5]
port 392 nsew signal output
rlabel metal3 s -300 11976 160 12096 4 WW4BEG[6]
port 393 nsew signal output
rlabel metal3 s -300 12248 160 12368 4 WW4BEG[7]
port 394 nsew signal output
rlabel metal3 s -300 12520 160 12640 4 WW4BEG[8]
port 395 nsew signal output
rlabel metal3 s -300 12792 160 12912 4 WW4BEG[9]
port 396 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 23000 44700
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 4639224
string GDS_FILE /home/asma/open_eFPGA_v2/openlane/RAM_IO/runs/24_12_22_00_50/results/signoff/RAM_IO.magic.gds
string GDS_START 165798
<< end >>

