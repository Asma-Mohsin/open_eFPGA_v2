magic
tech sky130A
magscale 1 2
timestamp 1733618897
<< nwell >>
rect 1066 6789 43554 7355
rect 1066 5701 43554 6267
rect 1066 4613 43554 5179
rect 1066 3525 43554 4091
rect 1066 2437 43554 3003
<< obsli1 >>
rect 1104 2159 43516 7633
<< obsm1 >>
rect 1104 892 43675 7664
<< metal2 >>
rect 1122 9840 1178 10300
rect 3238 9840 3294 10300
rect 5354 9840 5410 10300
rect 7470 9840 7526 10300
rect 9586 9840 9642 10300
rect 11702 9840 11758 10300
rect 13818 9840 13874 10300
rect 15934 9840 15990 10300
rect 18050 9840 18106 10300
rect 20166 9840 20222 10300
rect 22282 9840 22338 10300
rect 24398 9840 24454 10300
rect 26514 9840 26570 10300
rect 28630 9840 28686 10300
rect 30746 9840 30802 10300
rect 32862 9840 32918 10300
rect 34978 9840 35034 10300
rect 37094 9840 37150 10300
rect 39210 9840 39266 10300
rect 41326 9840 41382 10300
rect 43442 9840 43498 10300
rect 5078 -300 5134 160
rect 5354 -300 5410 160
rect 5630 -300 5686 160
rect 5906 -300 5962 160
rect 6182 -300 6238 160
rect 6458 -300 6514 160
rect 6734 -300 6790 160
rect 7010 -300 7066 160
rect 7286 -300 7342 160
rect 7562 -300 7618 160
rect 7838 -300 7894 160
rect 8114 -300 8170 160
rect 8390 -300 8446 160
rect 8666 -300 8722 160
rect 8942 -300 8998 160
rect 9218 -300 9274 160
rect 9494 -300 9550 160
rect 9770 -300 9826 160
rect 10046 -300 10102 160
rect 10322 -300 10378 160
rect 10598 -300 10654 160
rect 10874 -300 10930 160
rect 11150 -300 11206 160
rect 11426 -300 11482 160
rect 11702 -300 11758 160
rect 11978 -300 12034 160
rect 12254 -300 12310 160
rect 12530 -300 12586 160
rect 12806 -300 12862 160
rect 13082 -300 13138 160
rect 13358 -300 13414 160
rect 13634 -300 13690 160
rect 13910 -300 13966 160
rect 14186 -300 14242 160
rect 14462 -300 14518 160
rect 14738 -300 14794 160
rect 15014 -300 15070 160
rect 15290 -300 15346 160
rect 15566 -300 15622 160
rect 15842 -300 15898 160
rect 16118 -300 16174 160
rect 16394 -300 16450 160
rect 16670 -300 16726 160
rect 16946 -300 17002 160
rect 17222 -300 17278 160
rect 17498 -300 17554 160
rect 17774 -300 17830 160
rect 18050 -300 18106 160
rect 18326 -300 18382 160
rect 18602 -300 18658 160
rect 18878 -300 18934 160
rect 19154 -300 19210 160
rect 19430 -300 19486 160
rect 19706 -300 19762 160
rect 19982 -300 20038 160
rect 20258 -300 20314 160
rect 20534 -300 20590 160
rect 20810 -300 20866 160
rect 21086 -300 21142 160
rect 21362 -300 21418 160
rect 21638 -300 21694 160
rect 21914 -300 21970 160
rect 22190 -300 22246 160
rect 22466 -300 22522 160
rect 22742 -300 22798 160
rect 23018 -300 23074 160
rect 23294 -300 23350 160
rect 23570 -300 23626 160
rect 23846 -300 23902 160
rect 24122 -300 24178 160
rect 24398 -300 24454 160
rect 24674 -300 24730 160
rect 24950 -300 25006 160
rect 25226 -300 25282 160
rect 25502 -300 25558 160
rect 25778 -300 25834 160
rect 26054 -300 26110 160
rect 26330 -300 26386 160
rect 26606 -300 26662 160
rect 26882 -300 26938 160
rect 27158 -300 27214 160
rect 27434 -300 27490 160
rect 27710 -300 27766 160
rect 27986 -300 28042 160
rect 28262 -300 28318 160
rect 28538 -300 28594 160
rect 28814 -300 28870 160
rect 29090 -300 29146 160
rect 29366 -300 29422 160
rect 29642 -300 29698 160
rect 29918 -300 29974 160
rect 30194 -300 30250 160
rect 30470 -300 30526 160
rect 30746 -300 30802 160
rect 31022 -300 31078 160
rect 31298 -300 31354 160
rect 31574 -300 31630 160
rect 31850 -300 31906 160
rect 32126 -300 32182 160
rect 32402 -300 32458 160
rect 32678 -300 32734 160
rect 32954 -300 33010 160
rect 33230 -300 33286 160
rect 33506 -300 33562 160
rect 33782 -300 33838 160
rect 34058 -300 34114 160
rect 34334 -300 34390 160
rect 34610 -300 34666 160
rect 34886 -300 34942 160
rect 35162 -300 35218 160
rect 35438 -300 35494 160
rect 35714 -300 35770 160
rect 35990 -300 36046 160
rect 36266 -300 36322 160
rect 36542 -300 36598 160
rect 36818 -300 36874 160
rect 37094 -300 37150 160
rect 37370 -300 37426 160
rect 37646 -300 37702 160
rect 37922 -300 37978 160
rect 38198 -300 38254 160
rect 38474 -300 38530 160
rect 38750 -300 38806 160
rect 39026 -300 39082 160
rect 39302 -300 39358 160
rect 39578 -300 39634 160
<< obsm2 >>
rect 1234 9784 3182 9874
rect 3350 9784 5298 9874
rect 5466 9784 7414 9874
rect 7582 9784 9530 9874
rect 9698 9784 11646 9874
rect 11814 9784 13762 9874
rect 13930 9784 15878 9874
rect 16046 9784 17994 9874
rect 18162 9784 20110 9874
rect 20278 9784 22226 9874
rect 22394 9784 24342 9874
rect 24510 9784 26458 9874
rect 26626 9784 28574 9874
rect 28742 9784 30690 9874
rect 30858 9784 32806 9874
rect 32974 9784 34922 9874
rect 35090 9784 37038 9874
rect 37206 9784 39154 9874
rect 39322 9784 41270 9874
rect 41438 9784 43386 9874
rect 43554 9784 43669 9874
rect 1124 216 43669 9784
rect 1124 54 5022 216
rect 5190 54 5298 216
rect 5466 54 5574 216
rect 5742 54 5850 216
rect 6018 54 6126 216
rect 6294 54 6402 216
rect 6570 54 6678 216
rect 6846 54 6954 216
rect 7122 54 7230 216
rect 7398 54 7506 216
rect 7674 54 7782 216
rect 7950 54 8058 216
rect 8226 54 8334 216
rect 8502 54 8610 216
rect 8778 54 8886 216
rect 9054 54 9162 216
rect 9330 54 9438 216
rect 9606 54 9714 216
rect 9882 54 9990 216
rect 10158 54 10266 216
rect 10434 54 10542 216
rect 10710 54 10818 216
rect 10986 54 11094 216
rect 11262 54 11370 216
rect 11538 54 11646 216
rect 11814 54 11922 216
rect 12090 54 12198 216
rect 12366 54 12474 216
rect 12642 54 12750 216
rect 12918 54 13026 216
rect 13194 54 13302 216
rect 13470 54 13578 216
rect 13746 54 13854 216
rect 14022 54 14130 216
rect 14298 54 14406 216
rect 14574 54 14682 216
rect 14850 54 14958 216
rect 15126 54 15234 216
rect 15402 54 15510 216
rect 15678 54 15786 216
rect 15954 54 16062 216
rect 16230 54 16338 216
rect 16506 54 16614 216
rect 16782 54 16890 216
rect 17058 54 17166 216
rect 17334 54 17442 216
rect 17610 54 17718 216
rect 17886 54 17994 216
rect 18162 54 18270 216
rect 18438 54 18546 216
rect 18714 54 18822 216
rect 18990 54 19098 216
rect 19266 54 19374 216
rect 19542 54 19650 216
rect 19818 54 19926 216
rect 20094 54 20202 216
rect 20370 54 20478 216
rect 20646 54 20754 216
rect 20922 54 21030 216
rect 21198 54 21306 216
rect 21474 54 21582 216
rect 21750 54 21858 216
rect 22026 54 22134 216
rect 22302 54 22410 216
rect 22578 54 22686 216
rect 22854 54 22962 216
rect 23130 54 23238 216
rect 23406 54 23514 216
rect 23682 54 23790 216
rect 23958 54 24066 216
rect 24234 54 24342 216
rect 24510 54 24618 216
rect 24786 54 24894 216
rect 25062 54 25170 216
rect 25338 54 25446 216
rect 25614 54 25722 216
rect 25890 54 25998 216
rect 26166 54 26274 216
rect 26442 54 26550 216
rect 26718 54 26826 216
rect 26994 54 27102 216
rect 27270 54 27378 216
rect 27546 54 27654 216
rect 27822 54 27930 216
rect 28098 54 28206 216
rect 28374 54 28482 216
rect 28650 54 28758 216
rect 28926 54 29034 216
rect 29202 54 29310 216
rect 29478 54 29586 216
rect 29754 54 29862 216
rect 30030 54 30138 216
rect 30306 54 30414 216
rect 30582 54 30690 216
rect 30858 54 30966 216
rect 31134 54 31242 216
rect 31410 54 31518 216
rect 31686 54 31794 216
rect 31962 54 32070 216
rect 32238 54 32346 216
rect 32514 54 32622 216
rect 32790 54 32898 216
rect 33066 54 33174 216
rect 33342 54 33450 216
rect 33618 54 33726 216
rect 33894 54 34002 216
rect 34170 54 34278 216
rect 34446 54 34554 216
rect 34722 54 34830 216
rect 34998 54 35106 216
rect 35274 54 35382 216
rect 35550 54 35658 216
rect 35826 54 35934 216
rect 36102 54 36210 216
rect 36378 54 36486 216
rect 36654 54 36762 216
rect 36930 54 37038 216
rect 37206 54 37314 216
rect 37482 54 37590 216
rect 37758 54 37866 216
rect 38034 54 38142 216
rect 38310 54 38418 216
rect 38586 54 38694 216
rect 38862 54 38970 216
rect 39138 54 39246 216
rect 39414 54 39522 216
rect 39690 54 43669 216
<< obsm3 >>
rect 5073 851 43673 7649
<< metal4 >>
rect 6245 2128 6565 7664
rect 11546 2128 11866 7664
rect 16848 2128 17168 7664
rect 22149 2128 22469 7664
rect 27451 2128 27771 7664
rect 32752 2128 33072 7664
rect 38054 2128 38374 7664
rect 43355 2128 43675 7664
<< obsm4 >>
rect 30419 2048 32672 5133
rect 33152 2048 36557 5133
rect 30419 1123 36557 2048
<< labels >>
rlabel metal2 s 34058 -300 34114 160 8 Ci
port 1 nsew signal input
rlabel metal2 s 34334 -300 34390 160 8 FrameStrobe[0]
port 2 nsew signal input
rlabel metal2 s 37094 -300 37150 160 8 FrameStrobe[10]
port 3 nsew signal input
rlabel metal2 s 37370 -300 37426 160 8 FrameStrobe[11]
port 4 nsew signal input
rlabel metal2 s 37646 -300 37702 160 8 FrameStrobe[12]
port 5 nsew signal input
rlabel metal2 s 37922 -300 37978 160 8 FrameStrobe[13]
port 6 nsew signal input
rlabel metal2 s 38198 -300 38254 160 8 FrameStrobe[14]
port 7 nsew signal input
rlabel metal2 s 38474 -300 38530 160 8 FrameStrobe[15]
port 8 nsew signal input
rlabel metal2 s 38750 -300 38806 160 8 FrameStrobe[16]
port 9 nsew signal input
rlabel metal2 s 39026 -300 39082 160 8 FrameStrobe[17]
port 10 nsew signal input
rlabel metal2 s 39302 -300 39358 160 8 FrameStrobe[18]
port 11 nsew signal input
rlabel metal2 s 39578 -300 39634 160 8 FrameStrobe[19]
port 12 nsew signal input
rlabel metal2 s 34610 -300 34666 160 8 FrameStrobe[1]
port 13 nsew signal input
rlabel metal2 s 34886 -300 34942 160 8 FrameStrobe[2]
port 14 nsew signal input
rlabel metal2 s 35162 -300 35218 160 8 FrameStrobe[3]
port 15 nsew signal input
rlabel metal2 s 35438 -300 35494 160 8 FrameStrobe[4]
port 16 nsew signal input
rlabel metal2 s 35714 -300 35770 160 8 FrameStrobe[5]
port 17 nsew signal input
rlabel metal2 s 35990 -300 36046 160 8 FrameStrobe[6]
port 18 nsew signal input
rlabel metal2 s 36266 -300 36322 160 8 FrameStrobe[7]
port 19 nsew signal input
rlabel metal2 s 36542 -300 36598 160 8 FrameStrobe[8]
port 20 nsew signal input
rlabel metal2 s 36818 -300 36874 160 8 FrameStrobe[9]
port 21 nsew signal input
rlabel metal2 s 3238 9840 3294 10300 6 FrameStrobe_O[0]
port 22 nsew signal output
rlabel metal2 s 24398 9840 24454 10300 6 FrameStrobe_O[10]
port 23 nsew signal output
rlabel metal2 s 26514 9840 26570 10300 6 FrameStrobe_O[11]
port 24 nsew signal output
rlabel metal2 s 28630 9840 28686 10300 6 FrameStrobe_O[12]
port 25 nsew signal output
rlabel metal2 s 30746 9840 30802 10300 6 FrameStrobe_O[13]
port 26 nsew signal output
rlabel metal2 s 32862 9840 32918 10300 6 FrameStrobe_O[14]
port 27 nsew signal output
rlabel metal2 s 34978 9840 35034 10300 6 FrameStrobe_O[15]
port 28 nsew signal output
rlabel metal2 s 37094 9840 37150 10300 6 FrameStrobe_O[16]
port 29 nsew signal output
rlabel metal2 s 39210 9840 39266 10300 6 FrameStrobe_O[17]
port 30 nsew signal output
rlabel metal2 s 41326 9840 41382 10300 6 FrameStrobe_O[18]
port 31 nsew signal output
rlabel metal2 s 43442 9840 43498 10300 6 FrameStrobe_O[19]
port 32 nsew signal output
rlabel metal2 s 5354 9840 5410 10300 6 FrameStrobe_O[1]
port 33 nsew signal output
rlabel metal2 s 7470 9840 7526 10300 6 FrameStrobe_O[2]
port 34 nsew signal output
rlabel metal2 s 9586 9840 9642 10300 6 FrameStrobe_O[3]
port 35 nsew signal output
rlabel metal2 s 11702 9840 11758 10300 6 FrameStrobe_O[4]
port 36 nsew signal output
rlabel metal2 s 13818 9840 13874 10300 6 FrameStrobe_O[5]
port 37 nsew signal output
rlabel metal2 s 15934 9840 15990 10300 6 FrameStrobe_O[6]
port 38 nsew signal output
rlabel metal2 s 18050 9840 18106 10300 6 FrameStrobe_O[7]
port 39 nsew signal output
rlabel metal2 s 20166 9840 20222 10300 6 FrameStrobe_O[8]
port 40 nsew signal output
rlabel metal2 s 22282 9840 22338 10300 6 FrameStrobe_O[9]
port 41 nsew signal output
rlabel metal2 s 5078 -300 5134 160 8 N1END[0]
port 42 nsew signal input
rlabel metal2 s 5354 -300 5410 160 8 N1END[1]
port 43 nsew signal input
rlabel metal2 s 5630 -300 5686 160 8 N1END[2]
port 44 nsew signal input
rlabel metal2 s 5906 -300 5962 160 8 N1END[3]
port 45 nsew signal input
rlabel metal2 s 8390 -300 8446 160 8 N2END[0]
port 46 nsew signal input
rlabel metal2 s 8666 -300 8722 160 8 N2END[1]
port 47 nsew signal input
rlabel metal2 s 8942 -300 8998 160 8 N2END[2]
port 48 nsew signal input
rlabel metal2 s 9218 -300 9274 160 8 N2END[3]
port 49 nsew signal input
rlabel metal2 s 9494 -300 9550 160 8 N2END[4]
port 50 nsew signal input
rlabel metal2 s 9770 -300 9826 160 8 N2END[5]
port 51 nsew signal input
rlabel metal2 s 10046 -300 10102 160 8 N2END[6]
port 52 nsew signal input
rlabel metal2 s 10322 -300 10378 160 8 N2END[7]
port 53 nsew signal input
rlabel metal2 s 6182 -300 6238 160 8 N2MID[0]
port 54 nsew signal input
rlabel metal2 s 6458 -300 6514 160 8 N2MID[1]
port 55 nsew signal input
rlabel metal2 s 6734 -300 6790 160 8 N2MID[2]
port 56 nsew signal input
rlabel metal2 s 7010 -300 7066 160 8 N2MID[3]
port 57 nsew signal input
rlabel metal2 s 7286 -300 7342 160 8 N2MID[4]
port 58 nsew signal input
rlabel metal2 s 7562 -300 7618 160 8 N2MID[5]
port 59 nsew signal input
rlabel metal2 s 7838 -300 7894 160 8 N2MID[6]
port 60 nsew signal input
rlabel metal2 s 8114 -300 8170 160 8 N2MID[7]
port 61 nsew signal input
rlabel metal2 s 10598 -300 10654 160 8 N4END[0]
port 62 nsew signal input
rlabel metal2 s 13358 -300 13414 160 8 N4END[10]
port 63 nsew signal input
rlabel metal2 s 13634 -300 13690 160 8 N4END[11]
port 64 nsew signal input
rlabel metal2 s 13910 -300 13966 160 8 N4END[12]
port 65 nsew signal input
rlabel metal2 s 14186 -300 14242 160 8 N4END[13]
port 66 nsew signal input
rlabel metal2 s 14462 -300 14518 160 8 N4END[14]
port 67 nsew signal input
rlabel metal2 s 14738 -300 14794 160 8 N4END[15]
port 68 nsew signal input
rlabel metal2 s 10874 -300 10930 160 8 N4END[1]
port 69 nsew signal input
rlabel metal2 s 11150 -300 11206 160 8 N4END[2]
port 70 nsew signal input
rlabel metal2 s 11426 -300 11482 160 8 N4END[3]
port 71 nsew signal input
rlabel metal2 s 11702 -300 11758 160 8 N4END[4]
port 72 nsew signal input
rlabel metal2 s 11978 -300 12034 160 8 N4END[5]
port 73 nsew signal input
rlabel metal2 s 12254 -300 12310 160 8 N4END[6]
port 74 nsew signal input
rlabel metal2 s 12530 -300 12586 160 8 N4END[7]
port 75 nsew signal input
rlabel metal2 s 12806 -300 12862 160 8 N4END[8]
port 76 nsew signal input
rlabel metal2 s 13082 -300 13138 160 8 N4END[9]
port 77 nsew signal input
rlabel metal2 s 15014 -300 15070 160 8 NN4END[0]
port 78 nsew signal input
rlabel metal2 s 17774 -300 17830 160 8 NN4END[10]
port 79 nsew signal input
rlabel metal2 s 18050 -300 18106 160 8 NN4END[11]
port 80 nsew signal input
rlabel metal2 s 18326 -300 18382 160 8 NN4END[12]
port 81 nsew signal input
rlabel metal2 s 18602 -300 18658 160 8 NN4END[13]
port 82 nsew signal input
rlabel metal2 s 18878 -300 18934 160 8 NN4END[14]
port 83 nsew signal input
rlabel metal2 s 19154 -300 19210 160 8 NN4END[15]
port 84 nsew signal input
rlabel metal2 s 15290 -300 15346 160 8 NN4END[1]
port 85 nsew signal input
rlabel metal2 s 15566 -300 15622 160 8 NN4END[2]
port 86 nsew signal input
rlabel metal2 s 15842 -300 15898 160 8 NN4END[3]
port 87 nsew signal input
rlabel metal2 s 16118 -300 16174 160 8 NN4END[4]
port 88 nsew signal input
rlabel metal2 s 16394 -300 16450 160 8 NN4END[5]
port 89 nsew signal input
rlabel metal2 s 16670 -300 16726 160 8 NN4END[6]
port 90 nsew signal input
rlabel metal2 s 16946 -300 17002 160 8 NN4END[7]
port 91 nsew signal input
rlabel metal2 s 17222 -300 17278 160 8 NN4END[8]
port 92 nsew signal input
rlabel metal2 s 17498 -300 17554 160 8 NN4END[9]
port 93 nsew signal input
rlabel metal2 s 19430 -300 19486 160 8 S1BEG[0]
port 94 nsew signal output
rlabel metal2 s 19706 -300 19762 160 8 S1BEG[1]
port 95 nsew signal output
rlabel metal2 s 19982 -300 20038 160 8 S1BEG[2]
port 96 nsew signal output
rlabel metal2 s 20258 -300 20314 160 8 S1BEG[3]
port 97 nsew signal output
rlabel metal2 s 22742 -300 22798 160 8 S2BEG[0]
port 98 nsew signal output
rlabel metal2 s 23018 -300 23074 160 8 S2BEG[1]
port 99 nsew signal output
rlabel metal2 s 23294 -300 23350 160 8 S2BEG[2]
port 100 nsew signal output
rlabel metal2 s 23570 -300 23626 160 8 S2BEG[3]
port 101 nsew signal output
rlabel metal2 s 23846 -300 23902 160 8 S2BEG[4]
port 102 nsew signal output
rlabel metal2 s 24122 -300 24178 160 8 S2BEG[5]
port 103 nsew signal output
rlabel metal2 s 24398 -300 24454 160 8 S2BEG[6]
port 104 nsew signal output
rlabel metal2 s 24674 -300 24730 160 8 S2BEG[7]
port 105 nsew signal output
rlabel metal2 s 20534 -300 20590 160 8 S2BEGb[0]
port 106 nsew signal output
rlabel metal2 s 20810 -300 20866 160 8 S2BEGb[1]
port 107 nsew signal output
rlabel metal2 s 21086 -300 21142 160 8 S2BEGb[2]
port 108 nsew signal output
rlabel metal2 s 21362 -300 21418 160 8 S2BEGb[3]
port 109 nsew signal output
rlabel metal2 s 21638 -300 21694 160 8 S2BEGb[4]
port 110 nsew signal output
rlabel metal2 s 21914 -300 21970 160 8 S2BEGb[5]
port 111 nsew signal output
rlabel metal2 s 22190 -300 22246 160 8 S2BEGb[6]
port 112 nsew signal output
rlabel metal2 s 22466 -300 22522 160 8 S2BEGb[7]
port 113 nsew signal output
rlabel metal2 s 24950 -300 25006 160 8 S4BEG[0]
port 114 nsew signal output
rlabel metal2 s 27710 -300 27766 160 8 S4BEG[10]
port 115 nsew signal output
rlabel metal2 s 27986 -300 28042 160 8 S4BEG[11]
port 116 nsew signal output
rlabel metal2 s 28262 -300 28318 160 8 S4BEG[12]
port 117 nsew signal output
rlabel metal2 s 28538 -300 28594 160 8 S4BEG[13]
port 118 nsew signal output
rlabel metal2 s 28814 -300 28870 160 8 S4BEG[14]
port 119 nsew signal output
rlabel metal2 s 29090 -300 29146 160 8 S4BEG[15]
port 120 nsew signal output
rlabel metal2 s 25226 -300 25282 160 8 S4BEG[1]
port 121 nsew signal output
rlabel metal2 s 25502 -300 25558 160 8 S4BEG[2]
port 122 nsew signal output
rlabel metal2 s 25778 -300 25834 160 8 S4BEG[3]
port 123 nsew signal output
rlabel metal2 s 26054 -300 26110 160 8 S4BEG[4]
port 124 nsew signal output
rlabel metal2 s 26330 -300 26386 160 8 S4BEG[5]
port 125 nsew signal output
rlabel metal2 s 26606 -300 26662 160 8 S4BEG[6]
port 126 nsew signal output
rlabel metal2 s 26882 -300 26938 160 8 S4BEG[7]
port 127 nsew signal output
rlabel metal2 s 27158 -300 27214 160 8 S4BEG[8]
port 128 nsew signal output
rlabel metal2 s 27434 -300 27490 160 8 S4BEG[9]
port 129 nsew signal output
rlabel metal2 s 29366 -300 29422 160 8 SS4BEG[0]
port 130 nsew signal output
rlabel metal2 s 32126 -300 32182 160 8 SS4BEG[10]
port 131 nsew signal output
rlabel metal2 s 32402 -300 32458 160 8 SS4BEG[11]
port 132 nsew signal output
rlabel metal2 s 32678 -300 32734 160 8 SS4BEG[12]
port 133 nsew signal output
rlabel metal2 s 32954 -300 33010 160 8 SS4BEG[13]
port 134 nsew signal output
rlabel metal2 s 33230 -300 33286 160 8 SS4BEG[14]
port 135 nsew signal output
rlabel metal2 s 33506 -300 33562 160 8 SS4BEG[15]
port 136 nsew signal output
rlabel metal2 s 29642 -300 29698 160 8 SS4BEG[1]
port 137 nsew signal output
rlabel metal2 s 29918 -300 29974 160 8 SS4BEG[2]
port 138 nsew signal output
rlabel metal2 s 30194 -300 30250 160 8 SS4BEG[3]
port 139 nsew signal output
rlabel metal2 s 30470 -300 30526 160 8 SS4BEG[4]
port 140 nsew signal output
rlabel metal2 s 30746 -300 30802 160 8 SS4BEG[5]
port 141 nsew signal output
rlabel metal2 s 31022 -300 31078 160 8 SS4BEG[6]
port 142 nsew signal output
rlabel metal2 s 31298 -300 31354 160 8 SS4BEG[7]
port 143 nsew signal output
rlabel metal2 s 31574 -300 31630 160 8 SS4BEG[8]
port 144 nsew signal output
rlabel metal2 s 31850 -300 31906 160 8 SS4BEG[9]
port 145 nsew signal output
rlabel metal2 s 33782 -300 33838 160 8 UserCLK
port 146 nsew signal input
rlabel metal2 s 1122 9840 1178 10300 6 UserCLKo
port 147 nsew signal output
rlabel metal4 s 6245 2128 6565 7664 6 vccd1
port 148 nsew power bidirectional
rlabel metal4 s 16848 2128 17168 7664 6 vccd1
port 148 nsew power bidirectional
rlabel metal4 s 27451 2128 27771 7664 6 vccd1
port 148 nsew power bidirectional
rlabel metal4 s 38054 2128 38374 7664 6 vccd1
port 148 nsew power bidirectional
rlabel metal4 s 11546 2128 11866 7664 6 vssd1
port 149 nsew ground bidirectional
rlabel metal4 s 22149 2128 22469 7664 6 vssd1
port 149 nsew ground bidirectional
rlabel metal4 s 32752 2128 33072 7664 6 vssd1
port 149 nsew ground bidirectional
rlabel metal4 s 43355 2128 43675 7664 6 vssd1
port 149 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 44700 10000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 495066
string GDS_FILE /home/asma/Desktop/open_eFPGA/openlane/N_term_single/runs/24_12_08_00_47/results/signoff/N_term_single.magic.gds
string GDS_START 41474
<< end >>

