magic
tech sky130A
magscale 1 2
timestamp 1733618459
<< viali >>
rect 5089 8585 5123 8619
rect 5641 8585 5675 8619
rect 6009 8585 6043 8619
rect 6745 8585 6779 8619
rect 7481 8585 7515 8619
rect 8033 8585 8067 8619
rect 8585 8585 8619 8619
rect 9505 8585 9539 8619
rect 10241 8585 10275 8619
rect 10793 8585 10827 8619
rect 11161 8585 11195 8619
rect 12265 8585 12299 8619
rect 12817 8585 12851 8619
rect 13185 8585 13219 8619
rect 13737 8585 13771 8619
rect 14657 8585 14691 8619
rect 15025 8585 15059 8619
rect 15761 8585 15795 8619
rect 16313 8585 16347 8619
rect 16865 8585 16899 8619
rect 17233 8585 17267 8619
rect 17785 8585 17819 8619
rect 18245 8585 18279 8619
rect 18889 8585 18923 8619
rect 19901 8585 19935 8619
rect 29561 8585 29595 8619
rect 30665 8585 30699 8619
rect 31493 8585 31527 8619
rect 32137 8585 32171 8619
rect 32413 8585 32447 8619
rect 33517 8585 33551 8619
rect 34161 8585 34195 8619
rect 34897 8585 34931 8619
rect 36185 8585 36219 8619
rect 36553 8585 36587 8619
rect 39313 8585 39347 8619
rect 41153 8585 41187 8619
rect 5181 8517 5215 8551
rect 8125 8517 8159 8551
rect 13829 8517 13863 8551
rect 15301 8517 15335 8551
rect 37933 8517 37967 8551
rect 38485 8517 38519 8551
rect 39037 8517 39071 8551
rect 40877 8517 40911 8551
rect 4721 8449 4755 8483
rect 5733 8449 5767 8483
rect 6193 8449 6227 8483
rect 6837 8449 6871 8483
rect 7297 8449 7331 8483
rect 7665 8449 7699 8483
rect 8677 8449 8711 8483
rect 9321 8449 9355 8483
rect 9781 8449 9815 8483
rect 10425 8449 10459 8483
rect 10885 8449 10919 8483
rect 11345 8449 11379 8483
rect 11897 8449 11931 8483
rect 12357 8449 12391 8483
rect 13001 8449 13035 8483
rect 13369 8449 13403 8483
rect 14749 8449 14783 8483
rect 15945 8449 15979 8483
rect 16405 8449 16439 8483
rect 17049 8449 17083 8483
rect 17417 8449 17451 8483
rect 17877 8449 17911 8483
rect 18153 8449 18187 8483
rect 18981 8449 19015 8483
rect 19263 8449 19297 8483
rect 19809 8449 19843 8483
rect 20453 8449 20487 8483
rect 20729 8449 20763 8483
rect 21005 8449 21039 8483
rect 21281 8449 21315 8483
rect 21557 8449 21591 8483
rect 22017 8449 22051 8483
rect 22293 8449 22327 8483
rect 22569 8449 22603 8483
rect 22845 8449 22879 8483
rect 23121 8449 23155 8483
rect 23397 8449 23431 8483
rect 23673 8449 23707 8483
rect 23949 8449 23983 8483
rect 24225 8449 24259 8483
rect 24409 8449 24443 8483
rect 24685 8449 24719 8483
rect 24961 8449 24995 8483
rect 25237 8449 25271 8483
rect 25697 8449 25731 8483
rect 25789 8449 25823 8483
rect 26065 8449 26099 8483
rect 26341 8449 26375 8483
rect 26617 8449 26651 8483
rect 27169 8449 27203 8483
rect 27261 8449 27295 8483
rect 27537 8449 27571 8483
rect 27813 8449 27847 8483
rect 28273 8449 28307 8483
rect 28549 8449 28583 8483
rect 28825 8449 28859 8483
rect 29101 8449 29135 8483
rect 29377 8449 29411 8483
rect 29745 8449 29779 8483
rect 30021 8449 30055 8483
rect 30297 8449 30331 8483
rect 30573 8449 30607 8483
rect 30849 8449 30883 8483
rect 31125 8449 31159 8483
rect 31401 8449 31435 8483
rect 31677 8449 31711 8483
rect 31953 8449 31987 8483
rect 32321 8449 32355 8483
rect 32597 8449 32631 8483
rect 32873 8449 32907 8483
rect 33149 8449 33183 8483
rect 33425 8449 33459 8483
rect 33701 8449 33735 8483
rect 33977 8449 34011 8483
rect 34529 8449 34563 8483
rect 34805 8449 34839 8483
rect 35357 8449 35391 8483
rect 35909 8449 35943 8483
rect 36461 8449 36495 8483
rect 37381 8449 37415 8483
rect 39957 8449 39991 8483
rect 40509 8449 40543 8483
rect 41061 8449 41095 8483
rect 4537 8313 4571 8347
rect 7113 8313 7147 8347
rect 9137 8313 9171 8347
rect 11713 8313 11747 8347
rect 19441 8313 19475 8347
rect 21373 8313 21407 8347
rect 28365 8313 28399 8347
rect 28917 8313 28951 8347
rect 30941 8313 30975 8347
rect 31217 8313 31251 8347
rect 34345 8313 34379 8347
rect 35541 8313 35575 8347
rect 37565 8313 37599 8347
rect 38117 8313 38151 8347
rect 38669 8313 38703 8347
rect 40141 8313 40175 8347
rect 20269 8245 20303 8279
rect 20545 8245 20579 8279
rect 20821 8245 20855 8279
rect 21097 8245 21131 8279
rect 21833 8245 21867 8279
rect 22109 8245 22143 8279
rect 22385 8245 22419 8279
rect 22661 8245 22695 8279
rect 22937 8245 22971 8279
rect 23213 8245 23247 8279
rect 23489 8245 23523 8279
rect 23765 8245 23799 8279
rect 24041 8245 24075 8279
rect 24593 8245 24627 8279
rect 24869 8245 24903 8279
rect 25145 8245 25179 8279
rect 25421 8245 25455 8279
rect 25513 8245 25547 8279
rect 25973 8245 26007 8279
rect 26249 8245 26283 8279
rect 26525 8245 26559 8279
rect 26801 8245 26835 8279
rect 26985 8245 27019 8279
rect 27445 8245 27479 8279
rect 27721 8245 27755 8279
rect 27997 8245 28031 8279
rect 28089 8245 28123 8279
rect 28641 8245 28675 8279
rect 29193 8245 29227 8279
rect 29837 8245 29871 8279
rect 30113 8245 30147 8279
rect 30389 8245 30423 8279
rect 31769 8245 31803 8279
rect 32689 8245 32723 8279
rect 32965 8245 32999 8279
rect 33241 8245 33275 8279
rect 6009 8041 6043 8075
rect 6561 8041 6595 8075
rect 7113 8041 7147 8075
rect 8033 8041 8067 8075
rect 8585 8041 8619 8075
rect 9321 8041 9355 8075
rect 10425 8041 10459 8075
rect 11253 8041 11287 8075
rect 11805 8041 11839 8075
rect 12633 8041 12667 8075
rect 13461 8041 13495 8075
rect 14289 8041 14323 8075
rect 14841 8041 14875 8075
rect 15577 8041 15611 8075
rect 15945 8041 15979 8075
rect 16497 8041 16531 8075
rect 17785 8041 17819 8075
rect 18153 8041 18187 8075
rect 18521 8041 18555 8075
rect 20637 8041 20671 8075
rect 25513 8041 25547 8075
rect 25789 8041 25823 8075
rect 26065 8041 26099 8075
rect 36369 8041 36403 8075
rect 37473 8041 37507 8075
rect 38025 8041 38059 8075
rect 40049 8041 40083 8075
rect 40601 8041 40635 8075
rect 10057 7973 10091 8007
rect 17141 7973 17175 8007
rect 18889 7973 18923 8007
rect 19257 7973 19291 8007
rect 19533 7973 19567 8007
rect 20913 7973 20947 8007
rect 21189 7973 21223 8007
rect 21741 7973 21775 8007
rect 35909 7973 35943 8007
rect 10241 7837 10275 7871
rect 10701 7837 10735 7871
rect 11529 7837 11563 7871
rect 13737 7837 13771 7871
rect 14565 7837 14599 7871
rect 15761 7837 15795 7871
rect 16221 7837 16255 7871
rect 16773 7837 16807 7871
rect 17609 7833 17643 7867
rect 18061 7837 18095 7871
rect 18337 7837 18371 7871
rect 18705 7837 18739 7871
rect 19073 7837 19107 7871
rect 19441 7837 19475 7871
rect 19717 7837 19751 7871
rect 19993 7837 20027 7871
rect 20269 7837 20303 7871
rect 20545 7837 20579 7871
rect 20821 7837 20855 7871
rect 21097 7837 21131 7871
rect 21373 7837 21407 7871
rect 21649 7837 21683 7871
rect 21925 7837 21959 7871
rect 22201 7837 22235 7871
rect 22477 7837 22511 7871
rect 22753 7837 22787 7871
rect 23029 7837 23063 7871
rect 23305 7837 23339 7871
rect 23581 7837 23615 7871
rect 23857 7837 23891 7871
rect 24133 7837 24167 7871
rect 24593 7837 24627 7871
rect 24869 7837 24903 7871
rect 25145 7837 25179 7871
rect 25421 7837 25455 7871
rect 25697 7837 25731 7871
rect 25973 7837 26007 7871
rect 26249 7837 26283 7871
rect 26525 7837 26559 7871
rect 26801 7837 26835 7871
rect 27077 7837 27111 7871
rect 27353 7837 27387 7871
rect 27629 7837 27663 7871
rect 27905 7837 27939 7871
rect 33609 7837 33643 7871
rect 37381 7837 37415 7871
rect 38485 7837 38519 7871
rect 6285 7769 6319 7803
rect 6837 7769 6871 7803
rect 7389 7769 7423 7803
rect 8125 7769 8159 7803
rect 8677 7769 8711 7803
rect 9597 7769 9631 7803
rect 12081 7769 12115 7803
rect 12909 7769 12943 7803
rect 15117 7769 15151 7803
rect 17325 7769 17359 7803
rect 35725 7769 35759 7803
rect 36277 7769 36311 7803
rect 36829 7769 36863 7803
rect 37933 7769 37967 7803
rect 39037 7769 39071 7803
rect 39957 7769 39991 7803
rect 40509 7769 40543 7803
rect 17877 7701 17911 7735
rect 19809 7701 19843 7735
rect 20085 7701 20119 7735
rect 20361 7701 20395 7735
rect 21465 7701 21499 7735
rect 22017 7701 22051 7735
rect 22293 7701 22327 7735
rect 22569 7701 22603 7735
rect 22845 7701 22879 7735
rect 23121 7701 23155 7735
rect 23397 7701 23431 7735
rect 23673 7701 23707 7735
rect 23949 7701 23983 7735
rect 24409 7701 24443 7735
rect 24685 7701 24719 7735
rect 24961 7701 24995 7735
rect 25237 7701 25271 7735
rect 26341 7701 26375 7735
rect 26617 7701 26651 7735
rect 26893 7701 26927 7735
rect 27169 7701 27203 7735
rect 27445 7701 27479 7735
rect 27721 7701 27755 7735
rect 33425 7701 33459 7735
rect 36921 7701 36955 7735
rect 38761 7701 38795 7735
rect 39129 7701 39163 7735
rect 14473 7497 14507 7531
rect 17693 7497 17727 7531
rect 18245 7497 18279 7531
rect 18797 7497 18831 7531
rect 19257 7497 19291 7531
rect 19533 7497 19567 7531
rect 20269 7497 20303 7531
rect 21465 7497 21499 7531
rect 22569 7497 22603 7531
rect 7297 7361 7331 7395
rect 8769 7361 8803 7395
rect 14657 7361 14691 7395
rect 17601 7361 17635 7395
rect 17877 7361 17911 7395
rect 18153 7361 18187 7395
rect 18429 7361 18463 7395
rect 18981 7361 19015 7395
rect 19073 7361 19107 7395
rect 19349 7361 19383 7395
rect 19809 7361 19843 7395
rect 20177 7361 20211 7395
rect 20453 7361 20487 7395
rect 20821 7361 20855 7395
rect 21097 7361 21131 7395
rect 21373 7361 21407 7395
rect 21649 7361 21683 7395
rect 22017 7361 22051 7395
rect 22753 7361 22787 7395
rect 24961 7361 24995 7395
rect 26341 7361 26375 7395
rect 7113 7225 7147 7259
rect 8585 7225 8619 7259
rect 17969 7225 18003 7259
rect 21189 7225 21223 7259
rect 17417 7157 17451 7191
rect 19625 7157 19659 7191
rect 19993 7157 20027 7191
rect 20637 7157 20671 7191
rect 20913 7157 20947 7191
rect 21833 7157 21867 7191
rect 24777 7157 24811 7191
rect 26157 7157 26191 7191
rect 19809 6749 19843 6783
rect 20085 6749 20119 6783
rect 19625 6613 19659 6647
rect 19901 6613 19935 6647
rect 37565 5321 37599 5355
rect 37381 5185 37415 5219
rect 23029 4777 23063 4811
rect 23857 4777 23891 4811
rect 25973 4777 26007 4811
rect 28089 4777 28123 4811
rect 36921 4777 36955 4811
rect 38209 4777 38243 4811
rect 22753 4709 22787 4743
rect 23305 4709 23339 4743
rect 32321 4709 32355 4743
rect 21557 4573 21591 4607
rect 22569 4573 22603 4607
rect 22845 4573 22879 4607
rect 23121 4573 23155 4607
rect 23673 4573 23707 4607
rect 25789 4573 25823 4607
rect 27905 4573 27939 4607
rect 32137 4573 32171 4607
rect 36737 4573 36771 4607
rect 38025 4573 38059 4607
rect 21741 4437 21775 4471
rect 20913 4233 20947 4267
rect 22017 4233 22051 4267
rect 25145 4233 25179 4267
rect 37657 4233 37691 4267
rect 20729 4097 20763 4131
rect 21833 4097 21867 4131
rect 22109 4097 22143 4131
rect 22385 4097 22419 4131
rect 22661 4097 22695 4131
rect 24961 4097 24995 4131
rect 27077 4097 27111 4131
rect 31309 4097 31343 4131
rect 37473 4097 37507 4131
rect 39773 4097 39807 4131
rect 27261 3961 27295 3995
rect 31493 3961 31527 3995
rect 22293 3893 22327 3927
rect 22569 3893 22603 3927
rect 22845 3893 22879 3927
rect 39957 3893 39991 3927
rect 22109 3689 22143 3723
rect 23029 3689 23063 3723
rect 30205 3689 30239 3723
rect 37289 3689 37323 3723
rect 40509 3689 40543 3723
rect 19625 3621 19659 3655
rect 19441 3485 19475 3519
rect 21925 3485 21959 3519
rect 22201 3485 22235 3519
rect 22477 3485 22511 3519
rect 22845 3485 22879 3519
rect 30021 3485 30055 3519
rect 37105 3485 37139 3519
rect 40693 3485 40727 3519
rect 22385 3349 22419 3383
rect 22661 3349 22695 3383
rect 18797 3145 18831 3179
rect 21281 3145 21315 3179
rect 21557 3145 21591 3179
rect 29377 3145 29411 3179
rect 36185 3145 36219 3179
rect 39957 3145 39991 3179
rect 18613 3009 18647 3043
rect 21097 3009 21131 3043
rect 21373 3009 21407 3043
rect 22661 3009 22695 3043
rect 29193 3009 29227 3043
rect 36001 3009 36035 3043
rect 39773 3009 39807 3043
rect 22845 2873 22879 2907
rect 22109 2601 22143 2635
rect 39221 2601 39255 2635
rect 40233 2601 40267 2635
rect 21925 2397 21959 2431
rect 39037 2397 39071 2431
rect 40417 2397 40451 2431
rect 39037 2057 39071 2091
rect 21373 1921 21407 1955
rect 38853 1921 38887 1955
rect 21557 1717 21591 1751
rect 1593 1513 1627 1547
rect 3525 1513 3559 1547
rect 39313 1513 39347 1547
rect 42993 1513 43027 1547
rect 14289 1445 14323 1479
rect 1409 1309 1443 1343
rect 3341 1309 3375 1343
rect 5457 1309 5491 1343
rect 7573 1309 7607 1343
rect 9689 1309 9723 1343
rect 11805 1309 11839 1343
rect 14105 1309 14139 1343
rect 16037 1309 16071 1343
rect 18153 1309 18187 1343
rect 20269 1309 20303 1343
rect 22385 1309 22419 1343
rect 24501 1309 24535 1343
rect 26617 1309 26651 1343
rect 28733 1309 28767 1343
rect 30849 1309 30883 1343
rect 32965 1309 32999 1343
rect 35081 1309 35115 1343
rect 37289 1309 37323 1343
rect 39497 1309 39531 1343
rect 41613 1309 41647 1343
rect 43177 1309 43211 1343
rect 5641 1173 5675 1207
rect 7757 1173 7791 1207
rect 9873 1173 9907 1207
rect 11989 1173 12023 1207
rect 16221 1173 16255 1207
rect 18337 1173 18371 1207
rect 20453 1173 20487 1207
rect 22569 1173 22603 1207
rect 24685 1173 24719 1207
rect 26801 1173 26835 1207
rect 28917 1173 28951 1207
rect 31033 1173 31067 1207
rect 33149 1173 33183 1207
rect 35265 1173 35299 1207
rect 37473 1173 37507 1207
rect 41429 1173 41463 1207
<< metal1 >>
rect 11146 9936 11152 9988
rect 11204 9976 11210 9988
rect 23014 9976 23020 9988
rect 11204 9948 23020 9976
rect 11204 9936 11210 9948
rect 23014 9936 23020 9948
rect 23072 9936 23078 9988
rect 23198 9936 23204 9988
rect 23256 9976 23262 9988
rect 27154 9976 27160 9988
rect 23256 9948 27160 9976
rect 23256 9936 23262 9948
rect 27154 9936 27160 9948
rect 27212 9936 27218 9988
rect 19978 9908 19984 9920
rect 12406 9880 19984 9908
rect 12406 9840 12434 9880
rect 19978 9868 19984 9880
rect 20036 9868 20042 9920
rect 20162 9868 20168 9920
rect 20220 9908 20226 9920
rect 23566 9908 23572 9920
rect 20220 9880 23572 9908
rect 20220 9868 20226 9880
rect 23566 9868 23572 9880
rect 23624 9868 23630 9920
rect 29270 9868 29276 9920
rect 29328 9908 29334 9920
rect 29328 9880 35894 9908
rect 29328 9868 29334 9880
rect 8588 9812 12434 9840
rect 8588 9648 8616 9812
rect 17218 9800 17224 9852
rect 17276 9840 17282 9852
rect 22094 9840 22100 9852
rect 17276 9812 22100 9840
rect 17276 9800 17282 9812
rect 22094 9800 22100 9812
rect 22152 9800 22158 9852
rect 22186 9800 22192 9852
rect 22244 9840 22250 9852
rect 28166 9840 28172 9852
rect 22244 9812 28172 9840
rect 22244 9800 22250 9812
rect 28166 9800 28172 9812
rect 28224 9800 28230 9852
rect 33410 9840 33416 9852
rect 31726 9812 33416 9840
rect 17788 9744 21036 9772
rect 17788 9716 17816 9744
rect 12452 9676 17080 9704
rect 8570 9596 8576 9648
rect 8628 9596 8634 9648
rect 10778 9596 10784 9648
rect 10836 9636 10842 9648
rect 12452 9636 12480 9676
rect 16850 9636 16856 9648
rect 10836 9608 12480 9636
rect 14568 9608 16856 9636
rect 10836 9596 10842 9608
rect 14568 9568 14596 9608
rect 16850 9596 16856 9608
rect 16908 9596 16914 9648
rect 17052 9636 17080 9676
rect 17770 9664 17776 9716
rect 17828 9664 17834 9716
rect 18322 9664 18328 9716
rect 18380 9704 18386 9716
rect 18380 9676 20944 9704
rect 18380 9664 18386 9676
rect 20162 9636 20168 9648
rect 17052 9608 20168 9636
rect 20162 9596 20168 9608
rect 20220 9596 20226 9648
rect 4724 9540 14596 9568
rect 4724 9240 4752 9540
rect 17494 9528 17500 9580
rect 17552 9568 17558 9580
rect 20714 9568 20720 9580
rect 17552 9540 20720 9568
rect 17552 9528 17558 9540
rect 20714 9528 20720 9540
rect 20772 9528 20778 9580
rect 20916 9568 20944 9676
rect 21008 9636 21036 9744
rect 21082 9732 21088 9784
rect 21140 9772 21146 9784
rect 26786 9772 26792 9784
rect 21140 9744 26792 9772
rect 21140 9732 21146 9744
rect 26786 9732 26792 9744
rect 26844 9732 26850 9784
rect 31726 9772 31754 9812
rect 33410 9800 33416 9812
rect 33468 9800 33474 9852
rect 28966 9744 31754 9772
rect 21542 9664 21548 9716
rect 21600 9704 21606 9716
rect 28966 9704 28994 9744
rect 21600 9676 28994 9704
rect 21600 9664 21606 9676
rect 30466 9664 30472 9716
rect 30524 9704 30530 9716
rect 30524 9676 31984 9704
rect 30524 9664 30530 9676
rect 21910 9636 21916 9648
rect 21008 9608 21916 9636
rect 21910 9596 21916 9608
rect 21968 9596 21974 9648
rect 22922 9596 22928 9648
rect 22980 9636 22986 9648
rect 26878 9636 26884 9648
rect 22980 9608 26884 9636
rect 22980 9596 22986 9608
rect 26878 9596 26884 9608
rect 26936 9596 26942 9648
rect 20990 9568 20996 9580
rect 20916 9540 20996 9568
rect 20990 9528 20996 9540
rect 21048 9528 21054 9580
rect 21818 9528 21824 9580
rect 21876 9568 21882 9580
rect 31478 9568 31484 9580
rect 21876 9540 31484 9568
rect 21876 9528 21882 9540
rect 31478 9528 31484 9540
rect 31536 9528 31542 9580
rect 5534 9460 5540 9512
rect 5592 9500 5598 9512
rect 14642 9500 14648 9512
rect 5592 9472 14648 9500
rect 5592 9460 5598 9472
rect 14642 9460 14648 9472
rect 14700 9460 14706 9512
rect 14734 9460 14740 9512
rect 14792 9500 14798 9512
rect 21358 9500 21364 9512
rect 14792 9472 21364 9500
rect 14792 9460 14798 9472
rect 21358 9460 21364 9472
rect 21416 9460 21422 9512
rect 31018 9500 31024 9512
rect 21836 9472 31024 9500
rect 7282 9392 7288 9444
rect 7340 9432 7346 9444
rect 17954 9432 17960 9444
rect 7340 9404 17960 9432
rect 7340 9392 7346 9404
rect 17954 9392 17960 9404
rect 18012 9392 18018 9444
rect 18598 9392 18604 9444
rect 18656 9432 18662 9444
rect 21836 9432 21864 9472
rect 31018 9460 31024 9472
rect 31076 9460 31082 9512
rect 18656 9404 21864 9432
rect 18656 9392 18662 9404
rect 22186 9392 22192 9444
rect 22244 9432 22250 9444
rect 31846 9432 31852 9444
rect 22244 9404 31852 9432
rect 22244 9392 22250 9404
rect 31846 9392 31852 9404
rect 31904 9392 31910 9444
rect 22922 9364 22928 9376
rect 11348 9336 22928 9364
rect 4706 9188 4712 9240
rect 4764 9188 4770 9240
rect 11348 9172 11376 9336
rect 22922 9324 22928 9336
rect 22980 9324 22986 9376
rect 26786 9324 26792 9376
rect 26844 9364 26850 9376
rect 31956 9364 31984 9676
rect 35866 9432 35894 9880
rect 37550 9432 37556 9444
rect 35866 9404 37556 9432
rect 37550 9392 37556 9404
rect 37608 9392 37614 9444
rect 38010 9364 38016 9376
rect 26844 9336 31892 9364
rect 31956 9336 38016 9364
rect 26844 9324 26850 9336
rect 17218 9296 17224 9308
rect 12268 9268 17224 9296
rect 12268 9172 12296 9268
rect 17218 9256 17224 9268
rect 17276 9256 17282 9308
rect 18874 9256 18880 9308
rect 18932 9296 18938 9308
rect 20990 9296 20996 9308
rect 18932 9268 20996 9296
rect 18932 9256 18938 9268
rect 20990 9256 20996 9268
rect 21048 9256 21054 9308
rect 23290 9256 23296 9308
rect 23348 9296 23354 9308
rect 29914 9296 29920 9308
rect 23348 9268 29920 9296
rect 23348 9256 23354 9268
rect 29914 9256 29920 9268
rect 29972 9256 29978 9308
rect 31864 9296 31892 9336
rect 38010 9324 38016 9336
rect 38068 9324 38074 9376
rect 32122 9296 32128 9308
rect 31864 9268 32128 9296
rect 32122 9256 32128 9268
rect 32180 9256 32186 9308
rect 12526 9188 12532 9240
rect 12584 9228 12590 9240
rect 13814 9228 13820 9240
rect 12584 9200 13820 9228
rect 12584 9188 12590 9200
rect 13814 9188 13820 9200
rect 13872 9188 13878 9240
rect 13906 9188 13912 9240
rect 13964 9228 13970 9240
rect 21634 9228 21640 9240
rect 13964 9200 21640 9228
rect 13964 9188 13970 9200
rect 21634 9188 21640 9200
rect 21692 9188 21698 9240
rect 24578 9188 24584 9240
rect 24636 9228 24642 9240
rect 30742 9228 30748 9240
rect 24636 9200 30748 9228
rect 24636 9188 24642 9200
rect 30742 9188 30748 9200
rect 30800 9188 30806 9240
rect 34698 9188 34704 9240
rect 34756 9228 34762 9240
rect 35066 9228 35072 9240
rect 34756 9200 35072 9228
rect 34756 9188 34762 9200
rect 35066 9188 35072 9200
rect 35124 9188 35130 9240
rect 11330 9120 11336 9172
rect 11388 9120 11394 9172
rect 12250 9120 12256 9172
rect 12308 9120 12314 9172
rect 12986 9120 12992 9172
rect 13044 9160 13050 9172
rect 21818 9160 21824 9172
rect 13044 9132 21824 9160
rect 13044 9120 13050 9132
rect 21818 9120 21824 9132
rect 21876 9120 21882 9172
rect 21910 9120 21916 9172
rect 21968 9160 21974 9172
rect 21968 9132 25084 9160
rect 21968 9120 21974 9132
rect 6886 9064 13768 9092
rect 6178 8780 6184 8832
rect 6236 8820 6242 8832
rect 6886 8820 6914 9064
rect 8386 8984 8392 9036
rect 8444 9024 8450 9036
rect 13630 9024 13636 9036
rect 8444 8996 13636 9024
rect 8444 8984 8450 8996
rect 13630 8984 13636 8996
rect 13688 8984 13694 9036
rect 13740 9024 13768 9064
rect 13814 9052 13820 9104
rect 13872 9092 13878 9104
rect 22094 9092 22100 9104
rect 13872 9064 22100 9092
rect 13872 9052 13878 9064
rect 22094 9052 22100 9064
rect 22152 9052 22158 9104
rect 22186 9052 22192 9104
rect 22244 9092 22250 9104
rect 24946 9092 24952 9104
rect 22244 9064 24952 9092
rect 22244 9052 22250 9064
rect 24946 9052 24952 9064
rect 25004 9052 25010 9104
rect 25056 9092 25084 9132
rect 25406 9120 25412 9172
rect 25464 9160 25470 9172
rect 29362 9160 29368 9172
rect 25464 9132 29368 9160
rect 25464 9120 25470 9132
rect 29362 9120 29368 9132
rect 29420 9120 29426 9172
rect 25056 9064 31064 9092
rect 24118 9024 24124 9036
rect 13740 8996 24124 9024
rect 24118 8984 24124 8996
rect 24176 8984 24182 9036
rect 30926 9024 30932 9036
rect 24596 8996 30932 9024
rect 16114 8956 16120 8968
rect 12406 8928 16120 8956
rect 8662 8848 8668 8900
rect 8720 8888 8726 8900
rect 12406 8888 12434 8928
rect 16114 8916 16120 8928
rect 16172 8916 16178 8968
rect 16298 8916 16304 8968
rect 16356 8956 16362 8968
rect 17494 8956 17500 8968
rect 16356 8928 17500 8956
rect 16356 8916 16362 8928
rect 17494 8916 17500 8928
rect 17552 8916 17558 8968
rect 18506 8916 18512 8968
rect 18564 8956 18570 8968
rect 24596 8956 24624 8996
rect 30926 8984 30932 8996
rect 30984 8984 30990 9036
rect 31036 9024 31064 9064
rect 31570 9024 31576 9036
rect 31036 8996 31576 9024
rect 31570 8984 31576 8996
rect 31628 8984 31634 9036
rect 34606 8984 34612 9036
rect 34664 9024 34670 9036
rect 37458 9024 37464 9036
rect 34664 8996 37464 9024
rect 34664 8984 34670 8996
rect 37458 8984 37464 8996
rect 37516 8984 37522 9036
rect 29822 8956 29828 8968
rect 18564 8928 24624 8956
rect 24780 8928 29828 8956
rect 18564 8916 18570 8928
rect 15194 8888 15200 8900
rect 8720 8860 12434 8888
rect 13280 8860 15200 8888
rect 8720 8848 8726 8860
rect 6236 8792 6914 8820
rect 6236 8780 6242 8792
rect 9674 8780 9680 8832
rect 9732 8820 9738 8832
rect 13280 8820 13308 8860
rect 15194 8848 15200 8860
rect 15252 8848 15258 8900
rect 15286 8848 15292 8900
rect 15344 8888 15350 8900
rect 20806 8888 20812 8900
rect 15344 8860 20812 8888
rect 15344 8848 15350 8860
rect 20806 8848 20812 8860
rect 20864 8848 20870 8900
rect 20990 8848 20996 8900
rect 21048 8888 21054 8900
rect 21048 8860 21772 8888
rect 21048 8848 21054 8860
rect 9732 8792 13308 8820
rect 9732 8780 9738 8792
rect 13354 8780 13360 8832
rect 13412 8820 13418 8832
rect 21634 8820 21640 8832
rect 13412 8792 21640 8820
rect 13412 8780 13418 8792
rect 21634 8780 21640 8792
rect 21692 8780 21698 8832
rect 21744 8820 21772 8860
rect 23106 8848 23112 8900
rect 23164 8888 23170 8900
rect 24578 8888 24584 8900
rect 23164 8860 24584 8888
rect 23164 8848 23170 8860
rect 24578 8848 24584 8860
rect 24636 8848 24642 8900
rect 24780 8820 24808 8928
rect 29822 8916 29828 8928
rect 29880 8916 29886 8968
rect 31110 8916 31116 8968
rect 31168 8956 31174 8968
rect 35894 8956 35900 8968
rect 31168 8928 35900 8956
rect 31168 8916 31174 8928
rect 35894 8916 35900 8928
rect 35952 8916 35958 8968
rect 27062 8848 27068 8900
rect 27120 8888 27126 8900
rect 30374 8888 30380 8900
rect 27120 8860 30380 8888
rect 27120 8848 27126 8860
rect 30374 8848 30380 8860
rect 30432 8848 30438 8900
rect 21744 8792 24808 8820
rect 37642 8780 37648 8832
rect 37700 8820 37706 8832
rect 39298 8820 39304 8832
rect 37700 8792 39304 8820
rect 37700 8780 37706 8792
rect 39298 8780 39304 8792
rect 39356 8780 39362 8832
rect 1104 8730 43675 8752
rect 1104 8678 11552 8730
rect 11604 8678 11616 8730
rect 11668 8678 11680 8730
rect 11732 8678 11744 8730
rect 11796 8678 11808 8730
rect 11860 8678 22155 8730
rect 22207 8678 22219 8730
rect 22271 8678 22283 8730
rect 22335 8678 22347 8730
rect 22399 8678 22411 8730
rect 22463 8678 32758 8730
rect 32810 8678 32822 8730
rect 32874 8678 32886 8730
rect 32938 8678 32950 8730
rect 33002 8678 33014 8730
rect 33066 8678 43361 8730
rect 43413 8678 43425 8730
rect 43477 8678 43489 8730
rect 43541 8678 43553 8730
rect 43605 8678 43617 8730
rect 43669 8678 43675 8730
rect 1104 8656 43675 8678
rect 5077 8619 5135 8625
rect 5077 8585 5089 8619
rect 5123 8616 5135 8619
rect 5442 8616 5448 8628
rect 5123 8588 5448 8616
rect 5123 8585 5135 8588
rect 5077 8579 5135 8585
rect 5442 8576 5448 8588
rect 5500 8576 5506 8628
rect 5534 8576 5540 8628
rect 5592 8576 5598 8628
rect 5629 8619 5687 8625
rect 5629 8585 5641 8619
rect 5675 8616 5687 8619
rect 5718 8616 5724 8628
rect 5675 8588 5724 8616
rect 5675 8585 5687 8588
rect 5629 8579 5687 8585
rect 5718 8576 5724 8588
rect 5776 8576 5782 8628
rect 5997 8619 6055 8625
rect 5997 8585 6009 8619
rect 6043 8616 6055 8619
rect 6270 8616 6276 8628
rect 6043 8588 6276 8616
rect 6043 8585 6055 8588
rect 5997 8579 6055 8585
rect 6270 8576 6276 8588
rect 6328 8576 6334 8628
rect 6733 8619 6791 8625
rect 6733 8585 6745 8619
rect 6779 8616 6791 8619
rect 6822 8616 6828 8628
rect 6779 8588 6828 8616
rect 6779 8585 6791 8588
rect 6733 8579 6791 8585
rect 6822 8576 6828 8588
rect 6880 8576 6886 8628
rect 7282 8576 7288 8628
rect 7340 8576 7346 8628
rect 7469 8619 7527 8625
rect 7469 8585 7481 8619
rect 7515 8616 7527 8619
rect 7926 8616 7932 8628
rect 7515 8588 7932 8616
rect 7515 8585 7527 8588
rect 7469 8579 7527 8585
rect 7926 8576 7932 8588
rect 7984 8576 7990 8628
rect 8021 8619 8079 8625
rect 8021 8585 8033 8619
rect 8067 8616 8079 8619
rect 8478 8616 8484 8628
rect 8067 8588 8484 8616
rect 8067 8585 8079 8588
rect 8021 8579 8079 8585
rect 8478 8576 8484 8588
rect 8536 8576 8542 8628
rect 8573 8619 8631 8625
rect 8573 8585 8585 8619
rect 8619 8585 8631 8619
rect 8573 8579 8631 8585
rect 9493 8619 9551 8625
rect 9493 8585 9505 8619
rect 9539 8616 9551 8619
rect 9858 8616 9864 8628
rect 9539 8588 9864 8616
rect 9539 8585 9551 8588
rect 9493 8579 9551 8585
rect 5169 8551 5227 8557
rect 5169 8517 5181 8551
rect 5215 8548 5227 8551
rect 5552 8548 5580 8576
rect 7300 8548 7328 8576
rect 5215 8520 5580 8548
rect 5736 8520 7328 8548
rect 8113 8551 8171 8557
rect 5215 8517 5227 8520
rect 5169 8511 5227 8517
rect 4706 8440 4712 8492
rect 4764 8440 4770 8492
rect 5736 8489 5764 8520
rect 8113 8517 8125 8551
rect 8159 8548 8171 8551
rect 8386 8548 8392 8560
rect 8159 8520 8392 8548
rect 8159 8517 8171 8520
rect 8113 8511 8171 8517
rect 8386 8508 8392 8520
rect 8444 8508 8450 8560
rect 8588 8548 8616 8579
rect 9858 8576 9864 8588
rect 9916 8576 9922 8628
rect 10229 8619 10287 8625
rect 10229 8585 10241 8619
rect 10275 8585 10287 8619
rect 10229 8579 10287 8585
rect 10781 8619 10839 8625
rect 10781 8585 10793 8619
rect 10827 8616 10839 8619
rect 10962 8616 10968 8628
rect 10827 8588 10968 8616
rect 10827 8585 10839 8588
rect 10781 8579 10839 8585
rect 9582 8548 9588 8560
rect 8588 8520 9588 8548
rect 9582 8508 9588 8520
rect 9640 8508 9646 8560
rect 10244 8548 10272 8579
rect 10962 8576 10968 8588
rect 11020 8576 11026 8628
rect 11149 8619 11207 8625
rect 11149 8585 11161 8619
rect 11195 8616 11207 8619
rect 12066 8616 12072 8628
rect 11195 8588 12072 8616
rect 11195 8585 11207 8588
rect 11149 8579 11207 8585
rect 12066 8576 12072 8588
rect 12124 8576 12130 8628
rect 12253 8619 12311 8625
rect 12253 8585 12265 8619
rect 12299 8616 12311 8619
rect 12342 8616 12348 8628
rect 12299 8588 12348 8616
rect 12299 8585 12311 8588
rect 12253 8579 12311 8585
rect 12342 8576 12348 8588
rect 12400 8576 12406 8628
rect 12805 8619 12863 8625
rect 12805 8585 12817 8619
rect 12851 8616 12863 8619
rect 13078 8616 13084 8628
rect 12851 8588 13084 8616
rect 12851 8585 12863 8588
rect 12805 8579 12863 8585
rect 13078 8576 13084 8588
rect 13136 8576 13142 8628
rect 13173 8619 13231 8625
rect 13173 8585 13185 8619
rect 13219 8616 13231 8619
rect 13538 8616 13544 8628
rect 13219 8588 13544 8616
rect 13219 8585 13231 8588
rect 13173 8579 13231 8585
rect 13538 8576 13544 8588
rect 13596 8576 13602 8628
rect 13630 8576 13636 8628
rect 13688 8576 13694 8628
rect 13725 8619 13783 8625
rect 13725 8585 13737 8619
rect 13771 8616 13783 8619
rect 13998 8616 14004 8628
rect 13771 8588 14004 8616
rect 13771 8585 13783 8588
rect 13725 8579 13783 8585
rect 13998 8576 14004 8588
rect 14056 8576 14062 8628
rect 14645 8619 14703 8625
rect 14645 8585 14657 8619
rect 14691 8585 14703 8619
rect 14645 8579 14703 8585
rect 15013 8619 15071 8625
rect 15013 8585 15025 8619
rect 15059 8616 15071 8619
rect 15378 8616 15384 8628
rect 15059 8588 15384 8616
rect 15059 8585 15071 8588
rect 15013 8579 15071 8585
rect 11422 8548 11428 8560
rect 10244 8520 11428 8548
rect 11422 8508 11428 8520
rect 11480 8508 11486 8560
rect 11624 8520 13492 8548
rect 5721 8483 5779 8489
rect 5721 8449 5733 8483
rect 5767 8449 5779 8483
rect 5721 8443 5779 8449
rect 6178 8440 6184 8492
rect 6236 8440 6242 8492
rect 6825 8483 6883 8489
rect 6825 8449 6837 8483
rect 6871 8480 6883 8483
rect 7190 8480 7196 8492
rect 6871 8452 7196 8480
rect 6871 8449 6883 8452
rect 6825 8443 6883 8449
rect 7190 8440 7196 8452
rect 7248 8440 7254 8492
rect 7285 8483 7343 8489
rect 7285 8449 7297 8483
rect 7331 8449 7343 8483
rect 7285 8443 7343 8449
rect 7653 8483 7711 8489
rect 7653 8449 7665 8483
rect 7699 8480 7711 8483
rect 8570 8480 8576 8492
rect 7699 8452 8576 8480
rect 7699 8449 7711 8452
rect 7653 8443 7711 8449
rect 7300 8412 7328 8443
rect 8570 8440 8576 8452
rect 8628 8440 8634 8492
rect 8662 8440 8668 8492
rect 8720 8440 8726 8492
rect 9309 8483 9367 8489
rect 9309 8449 9321 8483
rect 9355 8480 9367 8483
rect 9674 8480 9680 8492
rect 9355 8452 9680 8480
rect 9355 8449 9367 8452
rect 9309 8443 9367 8449
rect 9674 8440 9680 8452
rect 9732 8440 9738 8492
rect 9769 8483 9827 8489
rect 9769 8449 9781 8483
rect 9815 8449 9827 8483
rect 9769 8443 9827 8449
rect 10413 8483 10471 8489
rect 10413 8449 10425 8483
rect 10459 8480 10471 8483
rect 10778 8480 10784 8492
rect 10459 8452 10784 8480
rect 10459 8449 10471 8452
rect 10413 8443 10471 8449
rect 9784 8412 9812 8443
rect 10778 8440 10784 8452
rect 10836 8440 10842 8492
rect 10873 8483 10931 8489
rect 10873 8449 10885 8483
rect 10919 8480 10931 8483
rect 11146 8480 11152 8492
rect 10919 8452 11152 8480
rect 10919 8449 10931 8452
rect 10873 8443 10931 8449
rect 11146 8440 11152 8452
rect 11204 8440 11210 8492
rect 11330 8440 11336 8492
rect 11388 8440 11394 8492
rect 11624 8412 11652 8520
rect 11885 8483 11943 8489
rect 11885 8449 11897 8483
rect 11931 8480 11943 8483
rect 12250 8480 12256 8492
rect 11931 8452 12256 8480
rect 11931 8449 11943 8452
rect 11885 8443 11943 8449
rect 12250 8440 12256 8452
rect 12308 8440 12314 8492
rect 12345 8483 12403 8489
rect 12345 8449 12357 8483
rect 12391 8480 12403 8483
rect 12526 8480 12532 8492
rect 12391 8452 12532 8480
rect 12391 8449 12403 8452
rect 12345 8443 12403 8449
rect 12526 8440 12532 8452
rect 12584 8440 12590 8492
rect 12986 8440 12992 8492
rect 13044 8440 13050 8492
rect 13354 8440 13360 8492
rect 13412 8440 13418 8492
rect 12710 8412 12716 8424
rect 7300 8384 9720 8412
rect 9784 8384 11652 8412
rect 11716 8384 12716 8412
rect 4525 8347 4583 8353
rect 4525 8313 4537 8347
rect 4571 8344 4583 8347
rect 5166 8344 5172 8356
rect 4571 8316 5172 8344
rect 4571 8313 4583 8316
rect 4525 8307 4583 8313
rect 5166 8304 5172 8316
rect 5224 8304 5230 8356
rect 7101 8347 7159 8353
rect 7101 8313 7113 8347
rect 7147 8344 7159 8347
rect 7650 8344 7656 8356
rect 7147 8316 7656 8344
rect 7147 8313 7159 8316
rect 7101 8307 7159 8313
rect 7650 8304 7656 8316
rect 7708 8304 7714 8356
rect 9122 8304 9128 8356
rect 9180 8304 9186 8356
rect 9692 8344 9720 8384
rect 11716 8353 11744 8384
rect 12710 8372 12716 8384
rect 12768 8372 12774 8424
rect 13464 8412 13492 8520
rect 13648 8412 13676 8576
rect 13814 8508 13820 8560
rect 13872 8508 13878 8560
rect 14660 8548 14688 8579
rect 15378 8576 15384 8588
rect 15436 8576 15442 8628
rect 15749 8619 15807 8625
rect 15749 8585 15761 8619
rect 15795 8616 15807 8619
rect 16206 8616 16212 8628
rect 15795 8588 16212 8616
rect 15795 8585 15807 8588
rect 15749 8579 15807 8585
rect 16206 8576 16212 8588
rect 16264 8576 16270 8628
rect 16301 8619 16359 8625
rect 16301 8585 16313 8619
rect 16347 8616 16359 8619
rect 16758 8616 16764 8628
rect 16347 8588 16764 8616
rect 16347 8585 16359 8588
rect 16301 8579 16359 8585
rect 16758 8576 16764 8588
rect 16816 8576 16822 8628
rect 16853 8619 16911 8625
rect 16853 8585 16865 8619
rect 16899 8585 16911 8619
rect 16853 8579 16911 8585
rect 17221 8619 17279 8625
rect 17221 8585 17233 8619
rect 17267 8616 17279 8619
rect 17586 8616 17592 8628
rect 17267 8588 17592 8616
rect 17267 8585 17279 8588
rect 17221 8579 17279 8585
rect 15102 8548 15108 8560
rect 14660 8520 15108 8548
rect 15102 8508 15108 8520
rect 15160 8508 15166 8560
rect 15286 8508 15292 8560
rect 15344 8508 15350 8560
rect 16868 8548 16896 8579
rect 17586 8576 17592 8588
rect 17644 8576 17650 8628
rect 17773 8619 17831 8625
rect 17773 8585 17785 8619
rect 17819 8616 17831 8619
rect 17862 8616 17868 8628
rect 17819 8588 17868 8616
rect 17819 8585 17831 8588
rect 17773 8579 17831 8585
rect 17862 8576 17868 8588
rect 17920 8576 17926 8628
rect 18230 8576 18236 8628
rect 18288 8576 18294 8628
rect 18877 8619 18935 8625
rect 18877 8585 18889 8619
rect 18923 8616 18935 8619
rect 19058 8616 19064 8628
rect 18923 8588 19064 8616
rect 18923 8585 18935 8588
rect 18877 8579 18935 8585
rect 19058 8576 19064 8588
rect 19116 8576 19122 8628
rect 19168 8588 19472 8616
rect 17310 8548 17316 8560
rect 16868 8520 17316 8548
rect 17310 8508 17316 8520
rect 17368 8508 17374 8560
rect 14734 8440 14740 8492
rect 14792 8440 14798 8492
rect 15933 8483 15991 8489
rect 15933 8449 15945 8483
rect 15979 8480 15991 8483
rect 16298 8480 16304 8492
rect 15979 8452 16304 8480
rect 15979 8449 15991 8452
rect 15933 8443 15991 8449
rect 16298 8440 16304 8452
rect 16356 8440 16362 8492
rect 16393 8483 16451 8489
rect 16393 8449 16405 8483
rect 16439 8480 16451 8483
rect 16758 8480 16764 8492
rect 16439 8452 16764 8480
rect 16439 8449 16451 8452
rect 16393 8443 16451 8449
rect 16758 8440 16764 8452
rect 16816 8440 16822 8492
rect 17037 8483 17095 8489
rect 17037 8449 17049 8483
rect 17083 8449 17095 8483
rect 17037 8443 17095 8449
rect 16942 8412 16948 8424
rect 13464 8384 13584 8412
rect 13648 8384 16948 8412
rect 11701 8347 11759 8353
rect 9692 8316 11652 8344
rect 11624 8276 11652 8316
rect 11701 8313 11713 8347
rect 11747 8313 11759 8347
rect 13556 8344 13584 8384
rect 16942 8372 16948 8384
rect 17000 8372 17006 8424
rect 17052 8412 17080 8443
rect 17402 8440 17408 8492
rect 17460 8440 17466 8492
rect 17865 8483 17923 8489
rect 17865 8449 17877 8483
rect 17911 8480 17923 8483
rect 18046 8480 18052 8492
rect 17911 8452 18052 8480
rect 17911 8449 17923 8452
rect 17865 8443 17923 8449
rect 18046 8440 18052 8452
rect 18104 8440 18110 8492
rect 18141 8483 18199 8489
rect 18141 8449 18153 8483
rect 18187 8449 18199 8483
rect 18141 8443 18199 8449
rect 18969 8483 19027 8489
rect 18969 8449 18981 8483
rect 19015 8449 19027 8483
rect 18969 8443 19027 8449
rect 17310 8412 17316 8424
rect 17052 8384 17316 8412
rect 17310 8372 17316 8384
rect 17368 8372 17374 8424
rect 17770 8372 17776 8424
rect 17828 8412 17834 8424
rect 18156 8412 18184 8443
rect 17828 8384 18184 8412
rect 18984 8412 19012 8443
rect 19058 8440 19064 8492
rect 19116 8480 19122 8492
rect 19168 8480 19196 8588
rect 19334 8548 19340 8560
rect 19260 8520 19340 8548
rect 19260 8489 19288 8520
rect 19334 8508 19340 8520
rect 19392 8508 19398 8560
rect 19444 8548 19472 8588
rect 19610 8576 19616 8628
rect 19668 8616 19674 8628
rect 19889 8619 19947 8625
rect 19889 8616 19901 8619
rect 19668 8588 19901 8616
rect 19668 8576 19674 8588
rect 19889 8585 19901 8588
rect 19935 8585 19947 8619
rect 19889 8579 19947 8585
rect 19978 8576 19984 8628
rect 20036 8616 20042 8628
rect 22462 8616 22468 8628
rect 20036 8588 22468 8616
rect 20036 8576 20042 8588
rect 22462 8576 22468 8588
rect 22520 8576 22526 8628
rect 22738 8576 22744 8628
rect 22796 8616 22802 8628
rect 25958 8616 25964 8628
rect 22796 8588 25964 8616
rect 22796 8576 22802 8588
rect 25958 8576 25964 8588
rect 26016 8576 26022 8628
rect 27062 8616 27068 8628
rect 26344 8588 27068 8616
rect 26344 8548 26372 8588
rect 27062 8576 27068 8588
rect 27120 8576 27126 8628
rect 29549 8619 29607 8625
rect 29549 8616 29561 8619
rect 28920 8588 29561 8616
rect 19444 8520 26372 8548
rect 26970 8508 26976 8560
rect 27028 8548 27034 8560
rect 27028 8520 27292 8548
rect 27028 8508 27034 8520
rect 19116 8452 19196 8480
rect 19251 8483 19309 8489
rect 19116 8440 19122 8452
rect 19251 8449 19263 8483
rect 19297 8449 19309 8483
rect 19251 8443 19309 8449
rect 19794 8440 19800 8492
rect 19852 8440 19858 8492
rect 20438 8440 20444 8492
rect 20496 8440 20502 8492
rect 20717 8483 20775 8489
rect 20717 8449 20729 8483
rect 20763 8480 20775 8483
rect 20898 8480 20904 8492
rect 20763 8452 20904 8480
rect 20763 8449 20775 8452
rect 20717 8443 20775 8449
rect 20898 8440 20904 8452
rect 20956 8440 20962 8492
rect 20993 8483 21051 8489
rect 20993 8449 21005 8483
rect 21039 8480 21051 8483
rect 21174 8480 21180 8492
rect 21039 8452 21180 8480
rect 21039 8449 21051 8452
rect 20993 8443 21051 8449
rect 21174 8440 21180 8452
rect 21232 8440 21238 8492
rect 21269 8483 21327 8489
rect 21269 8449 21281 8483
rect 21315 8480 21327 8483
rect 21450 8480 21456 8492
rect 21315 8452 21456 8480
rect 21315 8449 21327 8452
rect 21269 8443 21327 8449
rect 21450 8440 21456 8452
rect 21508 8440 21514 8492
rect 21542 8440 21548 8492
rect 21600 8440 21606 8492
rect 21726 8440 21732 8492
rect 21784 8480 21790 8492
rect 22005 8483 22063 8489
rect 22005 8480 22017 8483
rect 21784 8452 22017 8480
rect 21784 8440 21790 8452
rect 22005 8449 22017 8452
rect 22051 8449 22063 8483
rect 22005 8443 22063 8449
rect 22094 8440 22100 8492
rect 22152 8480 22158 8492
rect 22281 8483 22339 8489
rect 22281 8480 22293 8483
rect 22152 8452 22293 8480
rect 22152 8440 22158 8452
rect 22281 8449 22293 8452
rect 22327 8449 22339 8483
rect 22281 8443 22339 8449
rect 22554 8440 22560 8492
rect 22612 8440 22618 8492
rect 22830 8440 22836 8492
rect 22888 8440 22894 8492
rect 22922 8440 22928 8492
rect 22980 8480 22986 8492
rect 23109 8483 23167 8489
rect 23109 8480 23121 8483
rect 22980 8452 23121 8480
rect 22980 8440 22986 8452
rect 23109 8449 23121 8452
rect 23155 8449 23167 8483
rect 23109 8443 23167 8449
rect 23382 8440 23388 8492
rect 23440 8440 23446 8492
rect 23474 8440 23480 8492
rect 23532 8480 23538 8492
rect 23661 8483 23719 8489
rect 23661 8480 23673 8483
rect 23532 8452 23673 8480
rect 23532 8440 23538 8452
rect 23661 8449 23673 8452
rect 23707 8449 23719 8483
rect 23661 8443 23719 8449
rect 23934 8440 23940 8492
rect 23992 8440 23998 8492
rect 24026 8440 24032 8492
rect 24084 8480 24090 8492
rect 24213 8483 24271 8489
rect 24213 8480 24225 8483
rect 24084 8452 24225 8480
rect 24084 8440 24090 8452
rect 24213 8449 24225 8452
rect 24259 8449 24271 8483
rect 24213 8443 24271 8449
rect 24394 8440 24400 8492
rect 24452 8440 24458 8492
rect 24670 8440 24676 8492
rect 24728 8440 24734 8492
rect 24762 8440 24768 8492
rect 24820 8480 24826 8492
rect 24949 8483 25007 8489
rect 24949 8480 24961 8483
rect 24820 8452 24961 8480
rect 24820 8440 24826 8452
rect 24949 8449 24961 8452
rect 24995 8449 25007 8483
rect 24949 8443 25007 8449
rect 25222 8440 25228 8492
rect 25280 8440 25286 8492
rect 25314 8440 25320 8492
rect 25372 8480 25378 8492
rect 25685 8483 25743 8489
rect 25685 8480 25697 8483
rect 25372 8452 25697 8480
rect 25372 8440 25378 8452
rect 25685 8449 25697 8452
rect 25731 8449 25743 8483
rect 25685 8443 25743 8449
rect 25774 8440 25780 8492
rect 25832 8440 25838 8492
rect 26050 8440 26056 8492
rect 26108 8440 26114 8492
rect 26142 8440 26148 8492
rect 26200 8480 26206 8492
rect 26329 8483 26387 8489
rect 26329 8480 26341 8483
rect 26200 8452 26341 8480
rect 26200 8440 26206 8452
rect 26329 8449 26341 8452
rect 26375 8449 26387 8483
rect 26329 8443 26387 8449
rect 26602 8440 26608 8492
rect 26660 8440 26666 8492
rect 26694 8440 26700 8492
rect 26752 8480 26758 8492
rect 27264 8489 27292 8520
rect 28074 8508 28080 8560
rect 28132 8548 28138 8560
rect 28920 8548 28948 8588
rect 29549 8585 29561 8588
rect 29595 8585 29607 8619
rect 29549 8579 29607 8585
rect 29730 8576 29736 8628
rect 29788 8616 29794 8628
rect 29788 8588 30328 8616
rect 29788 8576 29794 8588
rect 28132 8520 28580 8548
rect 28132 8508 28138 8520
rect 27157 8483 27215 8489
rect 27157 8480 27169 8483
rect 26752 8452 27169 8480
rect 26752 8440 26758 8452
rect 27157 8449 27169 8452
rect 27203 8449 27215 8483
rect 27157 8443 27215 8449
rect 27249 8483 27307 8489
rect 27249 8449 27261 8483
rect 27295 8449 27307 8483
rect 27249 8443 27307 8449
rect 27522 8440 27528 8492
rect 27580 8440 27586 8492
rect 27614 8440 27620 8492
rect 27672 8480 27678 8492
rect 27801 8483 27859 8489
rect 27801 8480 27813 8483
rect 27672 8452 27813 8480
rect 27672 8440 27678 8452
rect 27801 8449 27813 8452
rect 27847 8449 27859 8483
rect 27801 8443 27859 8449
rect 27982 8440 27988 8492
rect 28040 8480 28046 8492
rect 28552 8489 28580 8520
rect 28736 8520 28948 8548
rect 28261 8483 28319 8489
rect 28261 8480 28273 8483
rect 28040 8452 28273 8480
rect 28040 8440 28046 8452
rect 28261 8449 28273 8452
rect 28307 8449 28319 8483
rect 28261 8443 28319 8449
rect 28537 8483 28595 8489
rect 28537 8449 28549 8483
rect 28583 8449 28595 8483
rect 28537 8443 28595 8449
rect 19334 8412 19340 8424
rect 18984 8384 19340 8412
rect 17828 8372 17834 8384
rect 19334 8372 19340 8384
rect 19392 8372 19398 8424
rect 25406 8412 25412 8424
rect 21468 8384 25412 8412
rect 11701 8307 11759 8313
rect 11808 8316 13492 8344
rect 13556 8316 16344 8344
rect 11808 8276 11836 8316
rect 11624 8248 11836 8276
rect 13464 8276 13492 8316
rect 14182 8276 14188 8288
rect 13464 8248 14188 8276
rect 14182 8236 14188 8248
rect 14240 8236 14246 8288
rect 16316 8276 16344 8316
rect 16390 8304 16396 8356
rect 16448 8344 16454 8356
rect 16448 8316 18644 8344
rect 16448 8304 16454 8316
rect 16574 8276 16580 8288
rect 16316 8248 16580 8276
rect 16574 8236 16580 8248
rect 16632 8236 16638 8288
rect 16666 8236 16672 8288
rect 16724 8276 16730 8288
rect 18322 8276 18328 8288
rect 16724 8248 18328 8276
rect 16724 8236 16730 8248
rect 18322 8236 18328 8248
rect 18380 8236 18386 8288
rect 18616 8276 18644 8316
rect 18690 8304 18696 8356
rect 18748 8344 18754 8356
rect 19429 8347 19487 8353
rect 19429 8344 19441 8347
rect 18748 8316 19441 8344
rect 18748 8304 18754 8316
rect 19429 8313 19441 8316
rect 19475 8313 19487 8347
rect 21361 8347 21419 8353
rect 21361 8344 21373 8347
rect 19429 8307 19487 8313
rect 19536 8316 21373 8344
rect 19536 8276 19564 8316
rect 21361 8313 21373 8316
rect 21407 8313 21419 8347
rect 21361 8307 21419 8313
rect 21468 8288 21496 8384
rect 25406 8372 25412 8384
rect 25464 8372 25470 8424
rect 28736 8412 28764 8520
rect 28994 8508 29000 8560
rect 29052 8548 29058 8560
rect 29052 8520 29408 8548
rect 29052 8508 29058 8520
rect 28813 8483 28871 8489
rect 28813 8449 28825 8483
rect 28859 8449 28871 8483
rect 28813 8443 28871 8449
rect 27816 8384 28764 8412
rect 22186 8304 22192 8356
rect 22244 8344 22250 8356
rect 22244 8316 22692 8344
rect 22244 8304 22250 8316
rect 18616 8248 19564 8276
rect 20070 8236 20076 8288
rect 20128 8276 20134 8288
rect 20257 8279 20315 8285
rect 20257 8276 20269 8279
rect 20128 8248 20269 8276
rect 20128 8236 20134 8248
rect 20257 8245 20269 8248
rect 20303 8245 20315 8279
rect 20257 8239 20315 8245
rect 20346 8236 20352 8288
rect 20404 8276 20410 8288
rect 20533 8279 20591 8285
rect 20533 8276 20545 8279
rect 20404 8248 20545 8276
rect 20404 8236 20410 8248
rect 20533 8245 20545 8248
rect 20579 8245 20591 8279
rect 20533 8239 20591 8245
rect 20806 8236 20812 8288
rect 20864 8236 20870 8288
rect 21082 8236 21088 8288
rect 21140 8236 21146 8288
rect 21450 8236 21456 8288
rect 21508 8236 21514 8288
rect 21542 8236 21548 8288
rect 21600 8276 21606 8288
rect 21821 8279 21879 8285
rect 21821 8276 21833 8279
rect 21600 8248 21833 8276
rect 21600 8236 21606 8248
rect 21821 8245 21833 8248
rect 21867 8245 21879 8279
rect 21821 8239 21879 8245
rect 22094 8236 22100 8288
rect 22152 8236 22158 8288
rect 22370 8236 22376 8288
rect 22428 8236 22434 8288
rect 22664 8285 22692 8316
rect 24946 8304 24952 8356
rect 25004 8344 25010 8356
rect 26142 8344 26148 8356
rect 25004 8316 26148 8344
rect 25004 8304 25010 8316
rect 26142 8304 26148 8316
rect 26200 8304 26206 8356
rect 27246 8304 27252 8356
rect 27304 8344 27310 8356
rect 27816 8344 27844 8384
rect 27304 8316 27844 8344
rect 27304 8304 27310 8316
rect 27890 8304 27896 8356
rect 27948 8344 27954 8356
rect 28353 8347 28411 8353
rect 28353 8344 28365 8347
rect 27948 8316 28365 8344
rect 27948 8304 27954 8316
rect 28353 8313 28365 8316
rect 28399 8313 28411 8347
rect 28353 8307 28411 8313
rect 28534 8304 28540 8356
rect 28592 8344 28598 8356
rect 28828 8344 28856 8443
rect 28902 8440 28908 8492
rect 28960 8480 28966 8492
rect 29380 8489 29408 8520
rect 29638 8508 29644 8560
rect 29696 8548 29702 8560
rect 29696 8520 30052 8548
rect 29696 8508 29702 8520
rect 29089 8483 29147 8489
rect 29089 8480 29101 8483
rect 28960 8452 29101 8480
rect 28960 8440 28966 8452
rect 29089 8449 29101 8452
rect 29135 8449 29147 8483
rect 29089 8443 29147 8449
rect 29365 8483 29423 8489
rect 29365 8449 29377 8483
rect 29411 8449 29423 8483
rect 29365 8443 29423 8449
rect 29733 8483 29791 8489
rect 29733 8449 29745 8483
rect 29779 8449 29791 8483
rect 29733 8443 29791 8449
rect 29178 8372 29184 8424
rect 29236 8412 29242 8424
rect 29748 8412 29776 8443
rect 29822 8440 29828 8492
rect 29880 8440 29886 8492
rect 30024 8489 30052 8520
rect 30300 8489 30328 8588
rect 30374 8576 30380 8628
rect 30432 8616 30438 8628
rect 30653 8619 30711 8625
rect 30653 8616 30665 8619
rect 30432 8588 30665 8616
rect 30432 8576 30438 8588
rect 30653 8585 30665 8588
rect 30699 8585 30711 8619
rect 30653 8579 30711 8585
rect 30834 8576 30840 8628
rect 30892 8616 30898 8628
rect 30892 8588 31432 8616
rect 30892 8576 30898 8588
rect 30742 8508 30748 8560
rect 30800 8548 30806 8560
rect 30800 8520 31156 8548
rect 30800 8508 30806 8520
rect 30009 8483 30067 8489
rect 30009 8449 30021 8483
rect 30055 8449 30067 8483
rect 30009 8443 30067 8449
rect 30285 8483 30343 8489
rect 30285 8449 30297 8483
rect 30331 8449 30343 8483
rect 30285 8443 30343 8449
rect 30374 8440 30380 8492
rect 30432 8480 30438 8492
rect 30561 8483 30619 8489
rect 30561 8480 30573 8483
rect 30432 8452 30573 8480
rect 30432 8440 30438 8452
rect 30561 8449 30573 8452
rect 30607 8449 30619 8483
rect 30561 8443 30619 8449
rect 30837 8483 30895 8489
rect 30837 8449 30849 8483
rect 30883 8449 30895 8483
rect 30837 8443 30895 8449
rect 29236 8384 29776 8412
rect 29236 8372 29242 8384
rect 28592 8316 28856 8344
rect 28592 8304 28598 8316
rect 28902 8304 28908 8356
rect 28960 8304 28966 8356
rect 29840 8344 29868 8440
rect 29012 8316 29776 8344
rect 29840 8316 30236 8344
rect 22649 8279 22707 8285
rect 22649 8245 22661 8279
rect 22695 8245 22707 8279
rect 22649 8239 22707 8245
rect 22922 8236 22928 8288
rect 22980 8236 22986 8288
rect 23198 8236 23204 8288
rect 23256 8236 23262 8288
rect 23474 8236 23480 8288
rect 23532 8236 23538 8288
rect 23566 8236 23572 8288
rect 23624 8276 23630 8288
rect 23753 8279 23811 8285
rect 23753 8276 23765 8279
rect 23624 8248 23765 8276
rect 23624 8236 23630 8248
rect 23753 8245 23765 8248
rect 23799 8245 23811 8279
rect 23753 8239 23811 8245
rect 24026 8236 24032 8288
rect 24084 8236 24090 8288
rect 24578 8236 24584 8288
rect 24636 8236 24642 8288
rect 24854 8236 24860 8288
rect 24912 8236 24918 8288
rect 25130 8236 25136 8288
rect 25188 8236 25194 8288
rect 25406 8236 25412 8288
rect 25464 8236 25470 8288
rect 25498 8236 25504 8288
rect 25556 8236 25562 8288
rect 25958 8236 25964 8288
rect 26016 8236 26022 8288
rect 26234 8236 26240 8288
rect 26292 8236 26298 8288
rect 26510 8236 26516 8288
rect 26568 8236 26574 8288
rect 26786 8236 26792 8288
rect 26844 8236 26850 8288
rect 26970 8236 26976 8288
rect 27028 8236 27034 8288
rect 27338 8236 27344 8288
rect 27396 8276 27402 8288
rect 27433 8279 27491 8285
rect 27433 8276 27445 8279
rect 27396 8248 27445 8276
rect 27396 8236 27402 8248
rect 27433 8245 27445 8248
rect 27479 8245 27491 8279
rect 27433 8239 27491 8245
rect 27709 8279 27767 8285
rect 27709 8245 27721 8279
rect 27755 8276 27767 8279
rect 27798 8276 27804 8288
rect 27755 8248 27804 8276
rect 27755 8245 27767 8248
rect 27709 8239 27767 8245
rect 27798 8236 27804 8248
rect 27856 8236 27862 8288
rect 27982 8236 27988 8288
rect 28040 8236 28046 8288
rect 28074 8236 28080 8288
rect 28132 8236 28138 8288
rect 28626 8236 28632 8288
rect 28684 8236 28690 8288
rect 28718 8236 28724 8288
rect 28776 8276 28782 8288
rect 29012 8276 29040 8316
rect 28776 8248 29040 8276
rect 28776 8236 28782 8248
rect 29178 8236 29184 8288
rect 29236 8236 29242 8288
rect 29748 8276 29776 8316
rect 29825 8279 29883 8285
rect 29825 8276 29837 8279
rect 29748 8248 29837 8276
rect 29825 8245 29837 8248
rect 29871 8245 29883 8279
rect 29825 8239 29883 8245
rect 29914 8236 29920 8288
rect 29972 8276 29978 8288
rect 30101 8279 30159 8285
rect 30101 8276 30113 8279
rect 29972 8248 30113 8276
rect 29972 8236 29978 8248
rect 30101 8245 30113 8248
rect 30147 8245 30159 8279
rect 30208 8276 30236 8316
rect 30282 8304 30288 8356
rect 30340 8344 30346 8356
rect 30852 8344 30880 8443
rect 31018 8440 31024 8492
rect 31076 8440 31082 8492
rect 31128 8489 31156 8520
rect 31404 8489 31432 8588
rect 31478 8576 31484 8628
rect 31536 8576 31542 8628
rect 31846 8576 31852 8628
rect 31904 8616 31910 8628
rect 32125 8619 32183 8625
rect 32125 8616 32137 8619
rect 31904 8588 32137 8616
rect 31904 8576 31910 8588
rect 32125 8585 32137 8588
rect 32171 8585 32183 8619
rect 32125 8579 32183 8585
rect 32398 8576 32404 8628
rect 32456 8576 32462 8628
rect 32490 8576 32496 8628
rect 32548 8616 32554 8628
rect 32548 8588 33180 8616
rect 32548 8576 32554 8588
rect 31754 8508 31760 8560
rect 31812 8548 31818 8560
rect 31812 8520 32076 8548
rect 31812 8508 31818 8520
rect 31113 8483 31171 8489
rect 31113 8449 31125 8483
rect 31159 8449 31171 8483
rect 31113 8443 31171 8449
rect 31389 8483 31447 8489
rect 31389 8449 31401 8483
rect 31435 8449 31447 8483
rect 31665 8483 31723 8489
rect 31665 8480 31677 8483
rect 31389 8443 31447 8449
rect 31496 8452 31677 8480
rect 30340 8316 30880 8344
rect 30340 8304 30346 8316
rect 30926 8304 30932 8356
rect 30984 8304 30990 8356
rect 31036 8344 31064 8440
rect 31294 8372 31300 8424
rect 31352 8412 31358 8424
rect 31496 8412 31524 8452
rect 31665 8449 31677 8452
rect 31711 8449 31723 8483
rect 31665 8443 31723 8449
rect 31941 8483 31999 8489
rect 31941 8449 31953 8483
rect 31987 8449 31999 8483
rect 32048 8480 32076 8520
rect 32214 8508 32220 8560
rect 32272 8548 32278 8560
rect 32272 8520 32904 8548
rect 32272 8508 32278 8520
rect 32876 8489 32904 8520
rect 33152 8489 33180 8588
rect 33502 8576 33508 8628
rect 33560 8576 33566 8628
rect 33870 8576 33876 8628
rect 33928 8616 33934 8628
rect 34149 8619 34207 8625
rect 34149 8616 34161 8619
rect 33928 8588 34161 8616
rect 33928 8576 33934 8588
rect 34149 8585 34161 8588
rect 34195 8585 34207 8619
rect 34149 8579 34207 8585
rect 34238 8576 34244 8628
rect 34296 8616 34302 8628
rect 34885 8619 34943 8625
rect 34885 8616 34897 8619
rect 34296 8588 34897 8616
rect 34296 8576 34302 8588
rect 34885 8585 34897 8588
rect 34931 8585 34943 8619
rect 34885 8579 34943 8585
rect 35066 8576 35072 8628
rect 35124 8616 35130 8628
rect 36173 8619 36231 8625
rect 36173 8616 36185 8619
rect 35124 8588 36185 8616
rect 35124 8576 35130 8588
rect 36173 8585 36185 8588
rect 36219 8585 36231 8619
rect 36173 8579 36231 8585
rect 36541 8619 36599 8625
rect 36541 8585 36553 8619
rect 36587 8585 36599 8619
rect 36541 8579 36599 8585
rect 33226 8508 33232 8560
rect 33284 8548 33290 8560
rect 33284 8520 33732 8548
rect 33284 8508 33290 8520
rect 33704 8489 33732 8520
rect 33778 8508 33784 8560
rect 33836 8548 33842 8560
rect 33836 8520 34560 8548
rect 33836 8508 33842 8520
rect 32309 8483 32367 8489
rect 32309 8480 32321 8483
rect 32048 8452 32321 8480
rect 31941 8443 31999 8449
rect 32309 8449 32321 8452
rect 32355 8449 32367 8483
rect 32309 8443 32367 8449
rect 32585 8483 32643 8489
rect 32585 8449 32597 8483
rect 32631 8449 32643 8483
rect 32585 8443 32643 8449
rect 32861 8483 32919 8489
rect 32861 8449 32873 8483
rect 32907 8449 32919 8483
rect 32861 8443 32919 8449
rect 33137 8483 33195 8489
rect 33137 8449 33149 8483
rect 33183 8449 33195 8483
rect 33137 8443 33195 8449
rect 33413 8483 33471 8489
rect 33413 8449 33425 8483
rect 33459 8449 33471 8483
rect 33413 8443 33471 8449
rect 33689 8483 33747 8489
rect 33689 8449 33701 8483
rect 33735 8449 33747 8483
rect 33689 8443 33747 8449
rect 31352 8384 31524 8412
rect 31352 8372 31358 8384
rect 31570 8372 31576 8424
rect 31628 8412 31634 8424
rect 31956 8412 31984 8443
rect 31628 8384 31984 8412
rect 31628 8372 31634 8384
rect 32030 8372 32036 8424
rect 32088 8412 32094 8424
rect 32600 8412 32628 8443
rect 32088 8384 32628 8412
rect 32088 8372 32094 8384
rect 32766 8372 32772 8424
rect 32824 8412 32830 8424
rect 33428 8412 33456 8443
rect 33962 8440 33968 8492
rect 34020 8440 34026 8492
rect 34532 8489 34560 8520
rect 34974 8508 34980 8560
rect 35032 8548 35038 8560
rect 36556 8548 36584 8579
rect 37458 8576 37464 8628
rect 37516 8616 37522 8628
rect 37516 8588 39068 8616
rect 37516 8576 37522 8588
rect 35032 8520 36584 8548
rect 35032 8508 35038 8520
rect 37550 8508 37556 8560
rect 37608 8548 37614 8560
rect 37921 8551 37979 8557
rect 37921 8548 37933 8551
rect 37608 8520 37933 8548
rect 37608 8508 37614 8520
rect 37921 8517 37933 8520
rect 37967 8517 37979 8551
rect 37921 8511 37979 8517
rect 38010 8508 38016 8560
rect 38068 8548 38074 8560
rect 39040 8557 39068 8588
rect 39298 8576 39304 8628
rect 39356 8576 39362 8628
rect 39666 8576 39672 8628
rect 39724 8616 39730 8628
rect 41141 8619 41199 8625
rect 41141 8616 41153 8619
rect 39724 8588 41153 8616
rect 39724 8576 39730 8588
rect 41141 8585 41153 8588
rect 41187 8585 41199 8619
rect 41141 8579 41199 8585
rect 38473 8551 38531 8557
rect 38473 8548 38485 8551
rect 38068 8520 38485 8548
rect 38068 8508 38074 8520
rect 38473 8517 38485 8520
rect 38519 8517 38531 8551
rect 38473 8511 38531 8517
rect 39025 8551 39083 8557
rect 39025 8517 39037 8551
rect 39071 8517 39083 8551
rect 40865 8551 40923 8557
rect 40865 8548 40877 8551
rect 39025 8511 39083 8517
rect 39132 8520 40877 8548
rect 34517 8483 34575 8489
rect 34517 8449 34529 8483
rect 34563 8449 34575 8483
rect 34517 8443 34575 8449
rect 34790 8440 34796 8492
rect 34848 8440 34854 8492
rect 35342 8440 35348 8492
rect 35400 8440 35406 8492
rect 35894 8440 35900 8492
rect 35952 8440 35958 8492
rect 36449 8483 36507 8489
rect 36449 8449 36461 8483
rect 36495 8449 36507 8483
rect 36449 8443 36507 8449
rect 36464 8412 36492 8443
rect 36630 8440 36636 8492
rect 36688 8480 36694 8492
rect 37369 8483 37427 8489
rect 37369 8480 37381 8483
rect 36688 8452 37381 8480
rect 36688 8440 36694 8452
rect 37369 8449 37381 8452
rect 37415 8449 37427 8483
rect 37369 8443 37427 8449
rect 38378 8440 38384 8492
rect 38436 8480 38442 8492
rect 39132 8480 39160 8520
rect 40865 8517 40877 8520
rect 40911 8517 40923 8551
rect 40865 8511 40923 8517
rect 38436 8452 39160 8480
rect 38436 8440 38442 8452
rect 39298 8440 39304 8492
rect 39356 8480 39362 8492
rect 39945 8483 40003 8489
rect 39945 8480 39957 8483
rect 39356 8452 39957 8480
rect 39356 8440 39362 8452
rect 39945 8449 39957 8452
rect 39991 8449 40003 8483
rect 39945 8443 40003 8449
rect 40497 8483 40555 8489
rect 40497 8449 40509 8483
rect 40543 8449 40555 8483
rect 40497 8443 40555 8449
rect 32824 8384 33456 8412
rect 33520 8384 36492 8412
rect 32824 8372 32830 8384
rect 31205 8347 31263 8353
rect 31205 8344 31217 8347
rect 31036 8316 31217 8344
rect 31205 8313 31217 8316
rect 31251 8313 31263 8347
rect 33520 8344 33548 8384
rect 36538 8372 36544 8424
rect 36596 8412 36602 8424
rect 36596 8384 38148 8412
rect 36596 8372 36602 8384
rect 31205 8307 31263 8313
rect 31404 8316 33548 8344
rect 31404 8288 31432 8316
rect 33594 8304 33600 8356
rect 33652 8344 33658 8356
rect 34333 8347 34391 8353
rect 34333 8344 34345 8347
rect 33652 8316 34345 8344
rect 33652 8304 33658 8316
rect 34333 8313 34345 8316
rect 34379 8313 34391 8347
rect 34333 8307 34391 8313
rect 34422 8304 34428 8356
rect 34480 8344 34486 8356
rect 35529 8347 35587 8353
rect 35529 8344 35541 8347
rect 34480 8316 35541 8344
rect 34480 8304 34486 8316
rect 35529 8313 35541 8316
rect 35575 8313 35587 8347
rect 35529 8307 35587 8313
rect 35802 8304 35808 8356
rect 35860 8344 35866 8356
rect 38120 8353 38148 8384
rect 38286 8372 38292 8424
rect 38344 8412 38350 8424
rect 38344 8384 39068 8412
rect 38344 8372 38350 8384
rect 37553 8347 37611 8353
rect 37553 8344 37565 8347
rect 35860 8316 37565 8344
rect 35860 8304 35866 8316
rect 37553 8313 37565 8316
rect 37599 8313 37611 8347
rect 37553 8307 37611 8313
rect 38105 8347 38163 8353
rect 38105 8313 38117 8347
rect 38151 8313 38163 8347
rect 38105 8307 38163 8313
rect 38654 8304 38660 8356
rect 38712 8304 38718 8356
rect 39040 8344 39068 8384
rect 39574 8372 39580 8424
rect 39632 8412 39638 8424
rect 40512 8412 40540 8443
rect 41046 8440 41052 8492
rect 41104 8440 41110 8492
rect 39632 8384 40540 8412
rect 39632 8372 39638 8384
rect 40129 8347 40187 8353
rect 40129 8344 40141 8347
rect 39040 8316 40141 8344
rect 40129 8313 40141 8316
rect 40175 8313 40187 8347
rect 40129 8307 40187 8313
rect 30377 8279 30435 8285
rect 30377 8276 30389 8279
rect 30208 8248 30389 8276
rect 30101 8239 30159 8245
rect 30377 8245 30389 8248
rect 30423 8245 30435 8279
rect 30377 8239 30435 8245
rect 31386 8236 31392 8288
rect 31444 8236 31450 8288
rect 31662 8236 31668 8288
rect 31720 8276 31726 8288
rect 31757 8279 31815 8285
rect 31757 8276 31769 8279
rect 31720 8248 31769 8276
rect 31720 8236 31726 8248
rect 31757 8245 31769 8248
rect 31803 8245 31815 8279
rect 31757 8239 31815 8245
rect 32122 8236 32128 8288
rect 32180 8276 32186 8288
rect 32677 8279 32735 8285
rect 32677 8276 32689 8279
rect 32180 8248 32689 8276
rect 32180 8236 32186 8248
rect 32677 8245 32689 8248
rect 32723 8245 32735 8279
rect 32677 8239 32735 8245
rect 32950 8236 32956 8288
rect 33008 8236 33014 8288
rect 33229 8279 33287 8285
rect 33229 8245 33241 8279
rect 33275 8276 33287 8279
rect 33410 8276 33416 8288
rect 33275 8248 33416 8276
rect 33275 8245 33287 8248
rect 33229 8239 33287 8245
rect 33410 8236 33416 8248
rect 33468 8236 33474 8288
rect 1104 8186 43516 8208
rect 1104 8134 6251 8186
rect 6303 8134 6315 8186
rect 6367 8134 6379 8186
rect 6431 8134 6443 8186
rect 6495 8134 6507 8186
rect 6559 8134 16854 8186
rect 16906 8134 16918 8186
rect 16970 8134 16982 8186
rect 17034 8134 17046 8186
rect 17098 8134 17110 8186
rect 17162 8134 27457 8186
rect 27509 8134 27521 8186
rect 27573 8134 27585 8186
rect 27637 8134 27649 8186
rect 27701 8134 27713 8186
rect 27765 8134 38060 8186
rect 38112 8134 38124 8186
rect 38176 8134 38188 8186
rect 38240 8134 38252 8186
rect 38304 8134 38316 8186
rect 38368 8134 43516 8186
rect 1104 8112 43516 8134
rect 5994 8032 6000 8084
rect 6052 8032 6058 8084
rect 6546 8032 6552 8084
rect 6604 8032 6610 8084
rect 7098 8032 7104 8084
rect 7156 8032 7162 8084
rect 8018 8032 8024 8084
rect 8076 8032 8082 8084
rect 8570 8032 8576 8084
rect 8628 8032 8634 8084
rect 9306 8032 9312 8084
rect 9364 8032 9370 8084
rect 10410 8032 10416 8084
rect 10468 8032 10474 8084
rect 10686 8032 10692 8084
rect 10744 8032 10750 8084
rect 11238 8032 11244 8084
rect 11296 8032 11302 8084
rect 11790 8032 11796 8084
rect 11848 8032 11854 8084
rect 12618 8032 12624 8084
rect 12676 8032 12682 8084
rect 13446 8032 13452 8084
rect 13504 8032 13510 8084
rect 14274 8032 14280 8084
rect 14332 8032 14338 8084
rect 14826 8032 14832 8084
rect 14884 8032 14890 8084
rect 15565 8075 15623 8081
rect 15565 8041 15577 8075
rect 15611 8072 15623 8075
rect 15654 8072 15660 8084
rect 15611 8044 15660 8072
rect 15611 8041 15623 8044
rect 15565 8035 15623 8041
rect 15654 8032 15660 8044
rect 15712 8032 15718 8084
rect 15930 8032 15936 8084
rect 15988 8032 15994 8084
rect 16482 8032 16488 8084
rect 16540 8032 16546 8084
rect 17586 8072 17592 8084
rect 16592 8044 17592 8072
rect 10045 8007 10103 8013
rect 10045 7973 10057 8007
rect 10091 8004 10103 8007
rect 10704 8004 10732 8032
rect 10091 7976 10732 8004
rect 10091 7973 10103 7976
rect 10045 7967 10103 7973
rect 12802 7964 12808 8016
rect 12860 8004 12866 8016
rect 16592 8004 16620 8044
rect 17586 8032 17592 8044
rect 17644 8032 17650 8084
rect 17770 8032 17776 8084
rect 17828 8032 17834 8084
rect 17954 8032 17960 8084
rect 18012 8072 18018 8084
rect 18141 8075 18199 8081
rect 18141 8072 18153 8075
rect 18012 8044 18153 8072
rect 18012 8032 18018 8044
rect 18141 8041 18153 8044
rect 18187 8041 18199 8075
rect 18141 8035 18199 8041
rect 18414 8032 18420 8084
rect 18472 8072 18478 8084
rect 18509 8075 18567 8081
rect 18509 8072 18521 8075
rect 18472 8044 18521 8072
rect 18472 8032 18478 8044
rect 18509 8041 18521 8044
rect 18555 8041 18567 8075
rect 20625 8075 20683 8081
rect 20625 8072 20637 8075
rect 18509 8035 18567 8041
rect 18616 8044 20637 8072
rect 12860 7976 16620 8004
rect 12860 7964 12866 7976
rect 17126 7964 17132 8016
rect 17184 7964 17190 8016
rect 18616 8004 18644 8044
rect 20625 8041 20637 8044
rect 20671 8041 20683 8075
rect 20625 8035 20683 8041
rect 20732 8044 21864 8072
rect 17512 7976 18644 8004
rect 18877 8007 18935 8013
rect 17034 7936 17040 7948
rect 15764 7908 17040 7936
rect 10229 7871 10287 7877
rect 10229 7837 10241 7871
rect 10275 7837 10287 7871
rect 10229 7831 10287 7837
rect 6270 7760 6276 7812
rect 6328 7760 6334 7812
rect 6822 7760 6828 7812
rect 6880 7760 6886 7812
rect 7377 7803 7435 7809
rect 7377 7769 7389 7803
rect 7423 7769 7435 7803
rect 7377 7763 7435 7769
rect 7392 7732 7420 7763
rect 8110 7760 8116 7812
rect 8168 7760 8174 7812
rect 8665 7803 8723 7809
rect 8665 7769 8677 7803
rect 8711 7800 8723 7803
rect 9490 7800 9496 7812
rect 8711 7772 9496 7800
rect 8711 7769 8723 7772
rect 8665 7763 8723 7769
rect 9490 7760 9496 7772
rect 9548 7760 9554 7812
rect 9582 7760 9588 7812
rect 9640 7760 9646 7812
rect 10244 7800 10272 7831
rect 10686 7828 10692 7880
rect 10744 7828 10750 7880
rect 11517 7871 11575 7877
rect 11517 7837 11529 7871
rect 11563 7868 11575 7871
rect 13630 7868 13636 7880
rect 11563 7840 13636 7868
rect 11563 7837 11575 7840
rect 11517 7831 11575 7837
rect 13630 7828 13636 7840
rect 13688 7828 13694 7880
rect 13722 7828 13728 7880
rect 13780 7828 13786 7880
rect 15764 7877 15792 7908
rect 17034 7896 17040 7908
rect 17092 7896 17098 7948
rect 14553 7871 14611 7877
rect 14553 7837 14565 7871
rect 14599 7868 14611 7871
rect 15749 7871 15807 7877
rect 14599 7840 15700 7868
rect 14599 7837 14611 7840
rect 14553 7831 14611 7837
rect 11882 7800 11888 7812
rect 10244 7772 11888 7800
rect 11882 7760 11888 7772
rect 11940 7760 11946 7812
rect 12069 7803 12127 7809
rect 12069 7769 12081 7803
rect 12115 7800 12127 7803
rect 12802 7800 12808 7812
rect 12115 7772 12808 7800
rect 12115 7769 12127 7772
rect 12069 7763 12127 7769
rect 12802 7760 12808 7772
rect 12860 7760 12866 7812
rect 12894 7760 12900 7812
rect 12952 7760 12958 7812
rect 15102 7760 15108 7812
rect 15160 7760 15166 7812
rect 15672 7800 15700 7840
rect 15749 7837 15761 7871
rect 15795 7837 15807 7871
rect 15749 7831 15807 7837
rect 16209 7871 16267 7877
rect 16209 7837 16221 7871
rect 16255 7868 16267 7871
rect 16390 7868 16396 7880
rect 16255 7840 16396 7868
rect 16255 7837 16267 7840
rect 16209 7831 16267 7837
rect 16390 7828 16396 7840
rect 16448 7828 16454 7880
rect 16761 7871 16819 7877
rect 16761 7837 16773 7871
rect 16807 7868 16819 7871
rect 17512 7868 17540 7976
rect 18877 7973 18889 8007
rect 18923 7973 18935 8007
rect 18877 7967 18935 7973
rect 18506 7936 18512 7948
rect 17880 7908 18512 7936
rect 16807 7840 17540 7868
rect 17597 7867 17655 7873
rect 16807 7837 16819 7840
rect 16761 7831 16819 7837
rect 17597 7833 17609 7867
rect 17643 7844 17655 7867
rect 17880 7844 17908 7908
rect 18506 7896 18512 7908
rect 18564 7896 18570 7948
rect 17643 7833 17908 7844
rect 17597 7827 17908 7833
rect 18049 7871 18107 7877
rect 18049 7837 18061 7871
rect 18095 7868 18107 7871
rect 18230 7868 18236 7880
rect 18095 7840 18236 7868
rect 18095 7837 18107 7840
rect 18049 7831 18107 7837
rect 18230 7828 18236 7840
rect 18288 7828 18294 7880
rect 18322 7828 18328 7880
rect 18380 7828 18386 7880
rect 18690 7828 18696 7880
rect 18748 7828 18754 7880
rect 18782 7828 18788 7880
rect 18840 7868 18846 7880
rect 18892 7868 18920 7967
rect 19058 7964 19064 8016
rect 19116 8004 19122 8016
rect 19245 8007 19303 8013
rect 19245 8004 19257 8007
rect 19116 7976 19257 8004
rect 19116 7964 19122 7976
rect 19245 7973 19257 7976
rect 19291 7973 19303 8007
rect 19245 7967 19303 7973
rect 19521 8007 19579 8013
rect 19521 7973 19533 8007
rect 19567 8004 19579 8007
rect 20254 8004 20260 8016
rect 19567 7976 19656 8004
rect 19567 7973 19579 7976
rect 19521 7967 19579 7973
rect 18840 7840 18920 7868
rect 18840 7828 18846 7840
rect 19058 7828 19064 7880
rect 19116 7828 19122 7880
rect 19150 7828 19156 7880
rect 19208 7868 19214 7880
rect 19334 7868 19340 7880
rect 19208 7840 19340 7868
rect 19208 7828 19214 7840
rect 19334 7828 19340 7840
rect 19392 7828 19398 7880
rect 19429 7871 19487 7877
rect 19429 7837 19441 7871
rect 19475 7868 19487 7871
rect 19475 7864 19564 7868
rect 19628 7864 19656 7976
rect 19904 7976 20260 8004
rect 19475 7840 19656 7864
rect 19475 7837 19487 7840
rect 19429 7831 19487 7837
rect 19536 7836 19656 7840
rect 19705 7871 19763 7877
rect 19705 7837 19717 7871
rect 19751 7868 19763 7871
rect 19904 7868 19932 7976
rect 20254 7964 20260 7976
rect 20312 7964 20318 8016
rect 20438 7964 20444 8016
rect 20496 8004 20502 8016
rect 20732 8004 20760 8044
rect 20496 7976 20760 8004
rect 20496 7964 20502 7976
rect 20898 7964 20904 8016
rect 20956 7964 20962 8016
rect 21082 7964 21088 8016
rect 21140 7964 21146 8016
rect 21174 7964 21180 8016
rect 21232 7964 21238 8016
rect 21726 7964 21732 8016
rect 21784 7964 21790 8016
rect 21836 8004 21864 8044
rect 24946 8032 24952 8084
rect 25004 8072 25010 8084
rect 25501 8075 25559 8081
rect 25501 8072 25513 8075
rect 25004 8044 25513 8072
rect 25004 8032 25010 8044
rect 25501 8041 25513 8044
rect 25547 8041 25559 8075
rect 25777 8075 25835 8081
rect 25777 8072 25789 8075
rect 25501 8035 25559 8041
rect 25608 8044 25789 8072
rect 25608 8004 25636 8044
rect 25777 8041 25789 8044
rect 25823 8041 25835 8075
rect 25777 8035 25835 8041
rect 25866 8032 25872 8084
rect 25924 8072 25930 8084
rect 26053 8075 26111 8081
rect 26053 8072 26065 8075
rect 25924 8044 26065 8072
rect 25924 8032 25930 8044
rect 26053 8041 26065 8044
rect 26099 8041 26111 8075
rect 26053 8035 26111 8041
rect 27890 8032 27896 8084
rect 27948 8032 27954 8084
rect 28074 8032 28080 8084
rect 28132 8032 28138 8084
rect 29362 8032 29368 8084
rect 29420 8072 29426 8084
rect 32950 8072 32956 8084
rect 29420 8044 32956 8072
rect 29420 8032 29426 8044
rect 32950 8032 32956 8044
rect 33008 8032 33014 8084
rect 36078 8032 36084 8084
rect 36136 8072 36142 8084
rect 36357 8075 36415 8081
rect 36357 8072 36369 8075
rect 36136 8044 36369 8072
rect 36136 8032 36142 8044
rect 36357 8041 36369 8044
rect 36403 8041 36415 8075
rect 36357 8035 36415 8041
rect 36814 8032 36820 8084
rect 36872 8072 36878 8084
rect 37461 8075 37519 8081
rect 37461 8072 37473 8075
rect 36872 8044 37473 8072
rect 36872 8032 36878 8044
rect 37461 8041 37473 8044
rect 37507 8041 37519 8075
rect 37461 8035 37519 8041
rect 37734 8032 37740 8084
rect 37792 8072 37798 8084
rect 38013 8075 38071 8081
rect 38013 8072 38025 8075
rect 37792 8044 38025 8072
rect 37792 8032 37798 8044
rect 38013 8041 38025 8044
rect 38059 8041 38071 8075
rect 38013 8035 38071 8041
rect 38838 8032 38844 8084
rect 38896 8072 38902 8084
rect 40037 8075 40095 8081
rect 40037 8072 40049 8075
rect 38896 8044 40049 8072
rect 38896 8032 38902 8044
rect 40037 8041 40049 8044
rect 40083 8041 40095 8075
rect 40037 8035 40095 8041
rect 40589 8075 40647 8081
rect 40589 8041 40601 8075
rect 40635 8041 40647 8075
rect 40589 8035 40647 8041
rect 27908 8004 27936 8032
rect 21836 7976 25636 8004
rect 25700 7976 27936 8004
rect 21100 7936 21128 7964
rect 22370 7936 22376 7948
rect 20548 7908 21128 7936
rect 21836 7908 22376 7936
rect 19751 7840 19932 7868
rect 19981 7871 20039 7877
rect 19751 7837 19763 7840
rect 19705 7831 19763 7837
rect 19981 7837 19993 7871
rect 20027 7868 20039 7871
rect 20070 7868 20076 7880
rect 20027 7840 20076 7868
rect 20027 7837 20039 7840
rect 19981 7831 20039 7837
rect 20070 7828 20076 7840
rect 20128 7828 20134 7880
rect 20257 7871 20315 7877
rect 20257 7837 20269 7871
rect 20303 7868 20315 7871
rect 20346 7868 20352 7880
rect 20303 7840 20352 7868
rect 20303 7837 20315 7840
rect 20257 7831 20315 7837
rect 20346 7828 20352 7840
rect 20404 7828 20410 7880
rect 20548 7877 20576 7908
rect 20533 7871 20591 7877
rect 20533 7837 20545 7871
rect 20579 7837 20591 7871
rect 20533 7831 20591 7837
rect 20809 7871 20867 7877
rect 20809 7837 20821 7871
rect 20855 7868 20867 7871
rect 20990 7868 20996 7880
rect 20855 7840 20996 7868
rect 20855 7837 20867 7840
rect 20809 7831 20867 7837
rect 20990 7828 20996 7840
rect 21048 7828 21054 7880
rect 21085 7871 21143 7877
rect 21085 7837 21097 7871
rect 21131 7868 21143 7871
rect 21174 7868 21180 7880
rect 21131 7840 21180 7868
rect 21131 7837 21143 7840
rect 21085 7831 21143 7837
rect 21174 7828 21180 7840
rect 21232 7828 21238 7880
rect 21358 7828 21364 7880
rect 21416 7828 21422 7880
rect 21637 7871 21695 7877
rect 21637 7837 21649 7871
rect 21683 7864 21695 7871
rect 21836 7864 21864 7908
rect 22370 7896 22376 7908
rect 22428 7896 22434 7948
rect 22646 7936 22652 7948
rect 22480 7908 22652 7936
rect 22480 7877 22508 7908
rect 22646 7896 22652 7908
rect 22704 7896 22710 7948
rect 23382 7936 23388 7948
rect 22756 7908 23388 7936
rect 22756 7877 22784 7908
rect 23382 7896 23388 7908
rect 23440 7896 23446 7948
rect 24136 7908 24808 7936
rect 21683 7837 21864 7864
rect 21637 7836 21864 7837
rect 21913 7871 21971 7877
rect 21913 7837 21925 7871
rect 21959 7868 21971 7871
rect 22189 7871 22247 7877
rect 21959 7840 22140 7868
rect 21959 7837 21971 7840
rect 21637 7831 21695 7836
rect 21913 7831 21971 7837
rect 17604 7816 17908 7827
rect 16942 7800 16948 7812
rect 15672 7772 16948 7800
rect 16942 7760 16948 7772
rect 17000 7760 17006 7812
rect 17313 7803 17371 7809
rect 17313 7769 17325 7803
rect 17359 7800 17371 7803
rect 17494 7800 17500 7812
rect 17359 7772 17500 7800
rect 17359 7769 17371 7772
rect 17313 7763 17371 7769
rect 17494 7760 17500 7772
rect 17552 7760 17558 7812
rect 18414 7760 18420 7812
rect 18472 7800 18478 7812
rect 18472 7772 21496 7800
rect 18472 7760 18478 7772
rect 11974 7732 11980 7744
rect 7392 7704 11980 7732
rect 11974 7692 11980 7704
rect 12032 7692 12038 7744
rect 14366 7692 14372 7744
rect 14424 7732 14430 7744
rect 17865 7735 17923 7741
rect 17865 7732 17877 7735
rect 14424 7704 17877 7732
rect 14424 7692 14430 7704
rect 17865 7701 17877 7704
rect 17911 7701 17923 7735
rect 17865 7695 17923 7701
rect 17954 7692 17960 7744
rect 18012 7732 18018 7744
rect 19797 7735 19855 7741
rect 19797 7732 19809 7735
rect 18012 7704 19809 7732
rect 18012 7692 18018 7704
rect 19797 7701 19809 7704
rect 19843 7701 19855 7735
rect 19797 7695 19855 7701
rect 20073 7735 20131 7741
rect 20073 7701 20085 7735
rect 20119 7732 20131 7735
rect 20254 7732 20260 7744
rect 20119 7704 20260 7732
rect 20119 7701 20131 7704
rect 20073 7695 20131 7701
rect 20254 7692 20260 7704
rect 20312 7692 20318 7744
rect 20346 7692 20352 7744
rect 20404 7692 20410 7744
rect 21468 7741 21496 7772
rect 21453 7735 21511 7741
rect 21453 7701 21465 7735
rect 21499 7701 21511 7735
rect 21453 7695 21511 7701
rect 21818 7692 21824 7744
rect 21876 7732 21882 7744
rect 22005 7735 22063 7741
rect 22005 7732 22017 7735
rect 21876 7704 22017 7732
rect 21876 7692 21882 7704
rect 22005 7701 22017 7704
rect 22051 7701 22063 7735
rect 22112 7732 22140 7840
rect 22189 7837 22201 7871
rect 22235 7837 22247 7871
rect 22189 7831 22247 7837
rect 22465 7871 22523 7877
rect 22465 7837 22477 7871
rect 22511 7837 22523 7871
rect 22465 7831 22523 7837
rect 22741 7871 22799 7877
rect 22741 7837 22753 7871
rect 22787 7837 22799 7871
rect 22741 7831 22799 7837
rect 22204 7800 22232 7831
rect 22922 7828 22928 7880
rect 22980 7828 22986 7880
rect 23017 7871 23075 7877
rect 23017 7837 23029 7871
rect 23063 7837 23075 7871
rect 23017 7831 23075 7837
rect 22940 7800 22968 7828
rect 22204 7772 22968 7800
rect 23032 7800 23060 7831
rect 23290 7828 23296 7880
rect 23348 7828 23354 7880
rect 23474 7828 23480 7880
rect 23532 7828 23538 7880
rect 23569 7871 23627 7877
rect 23569 7837 23581 7871
rect 23615 7837 23627 7871
rect 23569 7831 23627 7837
rect 23492 7800 23520 7828
rect 23032 7772 23520 7800
rect 23584 7800 23612 7831
rect 23842 7828 23848 7880
rect 23900 7828 23906 7880
rect 24026 7828 24032 7880
rect 24084 7828 24090 7880
rect 24136 7877 24164 7908
rect 24780 7880 24808 7908
rect 24121 7871 24179 7877
rect 24121 7837 24133 7871
rect 24167 7837 24179 7871
rect 24121 7831 24179 7837
rect 24578 7828 24584 7880
rect 24636 7828 24642 7880
rect 24762 7828 24768 7880
rect 24820 7828 24826 7880
rect 24854 7828 24860 7880
rect 24912 7828 24918 7880
rect 25130 7828 25136 7880
rect 25188 7828 25194 7880
rect 25406 7828 25412 7880
rect 25464 7828 25470 7880
rect 25700 7877 25728 7976
rect 25774 7896 25780 7948
rect 25832 7936 25838 7948
rect 28092 7936 28120 8032
rect 35802 7964 35808 8016
rect 35860 8004 35866 8016
rect 35897 8007 35955 8013
rect 35897 8004 35909 8007
rect 35860 7976 35909 8004
rect 35860 7964 35866 7976
rect 35897 7973 35909 7976
rect 35943 7973 35955 8007
rect 35897 7967 35955 7973
rect 39206 7964 39212 8016
rect 39264 8004 39270 8016
rect 40604 8004 40632 8035
rect 39264 7976 40632 8004
rect 39264 7964 39270 7976
rect 25832 7908 26648 7936
rect 25832 7896 25838 7908
rect 25685 7871 25743 7877
rect 25685 7837 25697 7871
rect 25731 7837 25743 7871
rect 25685 7831 25743 7837
rect 25958 7828 25964 7880
rect 26016 7828 26022 7880
rect 26234 7828 26240 7880
rect 26292 7828 26298 7880
rect 26510 7828 26516 7880
rect 26568 7828 26574 7880
rect 24044 7800 24072 7828
rect 23584 7772 24072 7800
rect 24136 7772 24992 7800
rect 24136 7744 24164 7772
rect 22186 7732 22192 7744
rect 22112 7704 22192 7732
rect 22005 7695 22063 7701
rect 22186 7692 22192 7704
rect 22244 7692 22250 7744
rect 22278 7692 22284 7744
rect 22336 7692 22342 7744
rect 22554 7692 22560 7744
rect 22612 7692 22618 7744
rect 22830 7692 22836 7744
rect 22888 7692 22894 7744
rect 23014 7692 23020 7744
rect 23072 7732 23078 7744
rect 23109 7735 23167 7741
rect 23109 7732 23121 7735
rect 23072 7704 23121 7732
rect 23072 7692 23078 7704
rect 23109 7701 23121 7704
rect 23155 7701 23167 7735
rect 23109 7695 23167 7701
rect 23382 7692 23388 7744
rect 23440 7692 23446 7744
rect 23658 7692 23664 7744
rect 23716 7692 23722 7744
rect 23934 7692 23940 7744
rect 23992 7692 23998 7744
rect 24118 7692 24124 7744
rect 24176 7692 24182 7744
rect 24394 7692 24400 7744
rect 24452 7692 24458 7744
rect 24670 7692 24676 7744
rect 24728 7692 24734 7744
rect 24964 7741 24992 7772
rect 24949 7735 25007 7741
rect 24949 7701 24961 7735
rect 24995 7701 25007 7735
rect 24949 7695 25007 7701
rect 25222 7692 25228 7744
rect 25280 7692 25286 7744
rect 26142 7692 26148 7744
rect 26200 7732 26206 7744
rect 26620 7741 26648 7908
rect 27080 7908 28120 7936
rect 26786 7828 26792 7880
rect 26844 7828 26850 7880
rect 27080 7877 27108 7908
rect 32674 7896 32680 7948
rect 32732 7936 32738 7948
rect 32732 7908 37412 7936
rect 32732 7896 32738 7908
rect 27065 7871 27123 7877
rect 27065 7837 27077 7871
rect 27111 7837 27123 7871
rect 27065 7831 27123 7837
rect 27338 7828 27344 7880
rect 27396 7828 27402 7880
rect 27617 7871 27675 7877
rect 27617 7837 27629 7871
rect 27663 7868 27675 7871
rect 27798 7868 27804 7880
rect 27663 7840 27804 7868
rect 27663 7837 27675 7840
rect 27617 7831 27675 7837
rect 27798 7828 27804 7840
rect 27856 7828 27862 7880
rect 27893 7871 27951 7877
rect 27893 7837 27905 7871
rect 27939 7868 27951 7871
rect 27982 7868 27988 7880
rect 27939 7840 27988 7868
rect 27939 7837 27951 7840
rect 27893 7831 27951 7837
rect 27982 7828 27988 7840
rect 28040 7828 28046 7880
rect 33318 7828 33324 7880
rect 33376 7868 33382 7880
rect 37384 7877 37412 7908
rect 33597 7871 33655 7877
rect 33597 7868 33609 7871
rect 33376 7840 33609 7868
rect 33376 7828 33382 7840
rect 33597 7837 33609 7840
rect 33643 7837 33655 7871
rect 37369 7871 37427 7877
rect 33597 7831 33655 7837
rect 33704 7840 35894 7868
rect 28074 7760 28080 7812
rect 28132 7800 28138 7812
rect 33704 7800 33732 7840
rect 28132 7772 33732 7800
rect 28132 7760 28138 7772
rect 35710 7760 35716 7812
rect 35768 7760 35774 7812
rect 35866 7800 35894 7840
rect 36188 7840 37228 7868
rect 36188 7800 36216 7840
rect 35866 7772 36216 7800
rect 36262 7760 36268 7812
rect 36320 7760 36326 7812
rect 36814 7760 36820 7812
rect 36872 7760 36878 7812
rect 37200 7800 37228 7840
rect 37369 7837 37381 7871
rect 37415 7837 37427 7871
rect 38473 7871 38531 7877
rect 38473 7868 38485 7871
rect 37369 7831 37427 7837
rect 37476 7840 38485 7868
rect 37476 7800 37504 7840
rect 38473 7837 38485 7840
rect 38519 7837 38531 7871
rect 38473 7831 38531 7837
rect 39850 7828 39856 7880
rect 39908 7868 39914 7880
rect 39908 7840 40540 7868
rect 39908 7828 39914 7840
rect 37200 7772 37504 7800
rect 37918 7760 37924 7812
rect 37976 7760 37982 7812
rect 38378 7760 38384 7812
rect 38436 7800 38442 7812
rect 39025 7803 39083 7809
rect 39025 7800 39037 7803
rect 38436 7772 39037 7800
rect 38436 7760 38442 7772
rect 39025 7769 39037 7772
rect 39071 7769 39083 7803
rect 39025 7763 39083 7769
rect 39942 7760 39948 7812
rect 40000 7760 40006 7812
rect 40512 7809 40540 7840
rect 40497 7803 40555 7809
rect 40497 7769 40509 7803
rect 40543 7769 40555 7803
rect 40497 7763 40555 7769
rect 26329 7735 26387 7741
rect 26329 7732 26341 7735
rect 26200 7704 26341 7732
rect 26200 7692 26206 7704
rect 26329 7701 26341 7704
rect 26375 7701 26387 7735
rect 26329 7695 26387 7701
rect 26605 7735 26663 7741
rect 26605 7701 26617 7735
rect 26651 7701 26663 7735
rect 26605 7695 26663 7701
rect 26878 7692 26884 7744
rect 26936 7692 26942 7744
rect 27154 7692 27160 7744
rect 27212 7692 27218 7744
rect 27430 7692 27436 7744
rect 27488 7692 27494 7744
rect 27709 7735 27767 7741
rect 27709 7701 27721 7735
rect 27755 7732 27767 7735
rect 28166 7732 28172 7744
rect 27755 7704 28172 7732
rect 27755 7701 27767 7704
rect 27709 7695 27767 7701
rect 28166 7692 28172 7704
rect 28224 7692 28230 7744
rect 33410 7692 33416 7744
rect 33468 7692 33474 7744
rect 35250 7692 35256 7744
rect 35308 7732 35314 7744
rect 36909 7735 36967 7741
rect 36909 7732 36921 7735
rect 35308 7704 36921 7732
rect 35308 7692 35314 7704
rect 36909 7701 36921 7704
rect 36955 7701 36967 7735
rect 36909 7695 36967 7701
rect 38746 7692 38752 7744
rect 38804 7692 38810 7744
rect 39114 7692 39120 7744
rect 39172 7692 39178 7744
rect 1104 7642 43675 7664
rect 1104 7590 11552 7642
rect 11604 7590 11616 7642
rect 11668 7590 11680 7642
rect 11732 7590 11744 7642
rect 11796 7590 11808 7642
rect 11860 7590 22155 7642
rect 22207 7590 22219 7642
rect 22271 7590 22283 7642
rect 22335 7590 22347 7642
rect 22399 7590 22411 7642
rect 22463 7590 32758 7642
rect 32810 7590 32822 7642
rect 32874 7590 32886 7642
rect 32938 7590 32950 7642
rect 33002 7590 33014 7642
rect 33066 7590 43361 7642
rect 43413 7590 43425 7642
rect 43477 7590 43489 7642
rect 43541 7590 43553 7642
rect 43605 7590 43617 7642
rect 43669 7590 43675 7642
rect 1104 7568 43675 7590
rect 6270 7488 6276 7540
rect 6328 7528 6334 7540
rect 14366 7528 14372 7540
rect 6328 7500 14372 7528
rect 6328 7488 6334 7500
rect 14366 7488 14372 7500
rect 14424 7488 14430 7540
rect 14461 7531 14519 7537
rect 14461 7497 14473 7531
rect 14507 7528 14519 7531
rect 14550 7528 14556 7540
rect 14507 7500 14556 7528
rect 14507 7497 14519 7500
rect 14461 7491 14519 7497
rect 14550 7488 14556 7500
rect 14608 7488 14614 7540
rect 17218 7488 17224 7540
rect 17276 7528 17282 7540
rect 17681 7531 17739 7537
rect 17681 7528 17693 7531
rect 17276 7500 17693 7528
rect 17276 7488 17282 7500
rect 17681 7497 17693 7500
rect 17727 7497 17739 7531
rect 17681 7491 17739 7497
rect 18046 7488 18052 7540
rect 18104 7528 18110 7540
rect 18233 7531 18291 7537
rect 18233 7528 18245 7531
rect 18104 7500 18245 7528
rect 18104 7488 18110 7500
rect 18233 7497 18245 7500
rect 18279 7497 18291 7531
rect 18233 7491 18291 7497
rect 18690 7488 18696 7540
rect 18748 7528 18754 7540
rect 18785 7531 18843 7537
rect 18785 7528 18797 7531
rect 18748 7500 18797 7528
rect 18748 7488 18754 7500
rect 18785 7497 18797 7500
rect 18831 7497 18843 7531
rect 18785 7491 18843 7497
rect 19058 7488 19064 7540
rect 19116 7488 19122 7540
rect 19242 7488 19248 7540
rect 19300 7488 19306 7540
rect 19521 7531 19579 7537
rect 19521 7497 19533 7531
rect 19567 7528 19579 7531
rect 19794 7528 19800 7540
rect 19567 7500 19800 7528
rect 19567 7497 19579 7500
rect 19521 7491 19579 7497
rect 19794 7488 19800 7500
rect 19852 7488 19858 7540
rect 20257 7531 20315 7537
rect 20257 7528 20269 7531
rect 19904 7500 20269 7528
rect 9030 7460 9036 7472
rect 8680 7432 9036 7460
rect 7282 7352 7288 7404
rect 7340 7352 7346 7404
rect 7101 7259 7159 7265
rect 7101 7225 7113 7259
rect 7147 7256 7159 7259
rect 7374 7256 7380 7268
rect 7147 7228 7380 7256
rect 7147 7225 7159 7228
rect 7101 7219 7159 7225
rect 7374 7216 7380 7228
rect 7432 7216 7438 7268
rect 8573 7259 8631 7265
rect 8573 7225 8585 7259
rect 8619 7256 8631 7259
rect 8680 7256 8708 7432
rect 9030 7420 9036 7432
rect 9088 7420 9094 7472
rect 9490 7420 9496 7472
rect 9548 7460 9554 7472
rect 16666 7460 16672 7472
rect 9548 7432 16672 7460
rect 9548 7420 9554 7432
rect 16666 7420 16672 7432
rect 16724 7420 16730 7472
rect 17770 7460 17776 7472
rect 17696 7432 17776 7460
rect 17696 7416 17724 7432
rect 17770 7420 17776 7432
rect 17828 7420 17834 7472
rect 19076 7460 19104 7488
rect 19904 7460 19932 7500
rect 20257 7497 20269 7500
rect 20303 7497 20315 7531
rect 20257 7491 20315 7497
rect 20806 7488 20812 7540
rect 20864 7488 20870 7540
rect 21453 7531 21511 7537
rect 21453 7528 21465 7531
rect 20916 7500 21465 7528
rect 19076 7432 19932 7460
rect 20070 7420 20076 7472
rect 20128 7460 20134 7472
rect 20128 7432 20484 7460
rect 20128 7420 20134 7432
rect 8757 7395 8815 7401
rect 8757 7361 8769 7395
rect 8803 7361 8815 7395
rect 8757 7355 8815 7361
rect 8619 7228 8708 7256
rect 8619 7225 8631 7228
rect 8573 7219 8631 7225
rect 8772 7188 8800 7355
rect 9582 7352 9588 7404
rect 9640 7352 9646 7404
rect 14642 7352 14648 7404
rect 14700 7352 14706 7404
rect 15102 7352 15108 7404
rect 15160 7392 15166 7404
rect 17494 7392 17500 7404
rect 15160 7364 17500 7392
rect 15160 7352 15166 7364
rect 17494 7352 17500 7364
rect 17552 7352 17558 7404
rect 17604 7401 17724 7416
rect 17589 7395 17724 7401
rect 17589 7361 17601 7395
rect 17635 7388 17724 7395
rect 17635 7361 17647 7388
rect 17589 7355 17647 7361
rect 17862 7352 17868 7404
rect 17920 7352 17926 7404
rect 18138 7352 18144 7404
rect 18196 7352 18202 7404
rect 18417 7395 18475 7401
rect 18417 7361 18429 7395
rect 18463 7392 18475 7395
rect 18598 7392 18604 7404
rect 18463 7364 18604 7392
rect 18463 7361 18475 7364
rect 18417 7355 18475 7361
rect 18598 7352 18604 7364
rect 18656 7352 18662 7404
rect 18966 7352 18972 7404
rect 19024 7352 19030 7404
rect 19058 7352 19064 7404
rect 19116 7352 19122 7404
rect 19337 7395 19395 7401
rect 19337 7361 19349 7395
rect 19383 7392 19395 7395
rect 19702 7392 19708 7404
rect 19383 7364 19708 7392
rect 19383 7361 19395 7364
rect 19337 7355 19395 7361
rect 19702 7352 19708 7364
rect 19760 7352 19766 7404
rect 19794 7352 19800 7404
rect 19852 7352 19858 7404
rect 19978 7352 19984 7404
rect 20036 7392 20042 7404
rect 20456 7401 20484 7432
rect 20824 7401 20852 7488
rect 20165 7395 20223 7401
rect 20165 7392 20177 7395
rect 20036 7364 20177 7392
rect 20036 7352 20042 7364
rect 20165 7361 20177 7364
rect 20211 7361 20223 7395
rect 20165 7355 20223 7361
rect 20441 7395 20499 7401
rect 20441 7361 20453 7395
rect 20487 7361 20499 7395
rect 20441 7355 20499 7361
rect 20809 7395 20867 7401
rect 20809 7361 20821 7395
rect 20855 7361 20867 7395
rect 20809 7355 20867 7361
rect 9600 7324 9628 7352
rect 16758 7324 16764 7336
rect 9600 7296 16764 7324
rect 16758 7284 16764 7296
rect 16816 7284 16822 7336
rect 18046 7284 18052 7336
rect 18104 7324 18110 7336
rect 20916 7324 20944 7500
rect 21453 7497 21465 7500
rect 21499 7497 21511 7531
rect 21453 7491 21511 7497
rect 21542 7488 21548 7540
rect 21600 7488 21606 7540
rect 22002 7528 22008 7540
rect 21652 7500 22008 7528
rect 21174 7460 21180 7472
rect 18104 7296 20944 7324
rect 21008 7432 21180 7460
rect 21008 7324 21036 7432
rect 21174 7420 21180 7432
rect 21232 7420 21238 7472
rect 21085 7395 21143 7401
rect 21085 7361 21097 7395
rect 21131 7392 21143 7395
rect 21266 7392 21272 7404
rect 21131 7364 21272 7392
rect 21131 7361 21143 7364
rect 21085 7355 21143 7361
rect 21266 7352 21272 7364
rect 21324 7352 21330 7404
rect 21361 7395 21419 7401
rect 21361 7361 21373 7395
rect 21407 7392 21419 7395
rect 21560 7392 21588 7488
rect 21652 7401 21680 7500
rect 22002 7488 22008 7500
rect 22060 7488 22066 7540
rect 22557 7531 22615 7537
rect 22557 7497 22569 7531
rect 22603 7528 22615 7531
rect 22646 7528 22652 7540
rect 22603 7500 22652 7528
rect 22603 7497 22615 7500
rect 22557 7491 22615 7497
rect 22646 7488 22652 7500
rect 22704 7488 22710 7540
rect 23198 7488 23204 7540
rect 23256 7488 23262 7540
rect 23290 7488 23296 7540
rect 23348 7528 23354 7540
rect 29178 7528 29184 7540
rect 23348 7500 29184 7528
rect 23348 7488 23354 7500
rect 29178 7488 29184 7500
rect 29236 7488 29242 7540
rect 33410 7488 33416 7540
rect 33468 7488 33474 7540
rect 23106 7460 23112 7472
rect 22020 7432 23112 7460
rect 22020 7401 22048 7432
rect 23106 7420 23112 7432
rect 23164 7420 23170 7472
rect 21407 7364 21588 7392
rect 21637 7395 21695 7401
rect 21407 7361 21419 7364
rect 21361 7355 21419 7361
rect 21637 7361 21649 7395
rect 21683 7361 21695 7395
rect 21637 7355 21695 7361
rect 22005 7395 22063 7401
rect 22005 7361 22017 7395
rect 22051 7361 22063 7395
rect 22005 7355 22063 7361
rect 22741 7395 22799 7401
rect 22741 7361 22753 7395
rect 22787 7392 22799 7395
rect 23216 7392 23244 7488
rect 25498 7460 25504 7472
rect 24964 7432 25504 7460
rect 24964 7401 24992 7432
rect 25498 7420 25504 7432
rect 25556 7420 25562 7472
rect 26970 7460 26976 7472
rect 26344 7432 26976 7460
rect 26344 7401 26372 7432
rect 26970 7420 26976 7432
rect 27028 7420 27034 7472
rect 22787 7364 23244 7392
rect 24949 7395 25007 7401
rect 22787 7361 22799 7364
rect 22741 7355 22799 7361
rect 24949 7361 24961 7395
rect 24995 7361 25007 7395
rect 24949 7355 25007 7361
rect 26329 7395 26387 7401
rect 26329 7361 26341 7395
rect 26375 7361 26387 7395
rect 26329 7355 26387 7361
rect 21008 7296 31754 7324
rect 18104 7284 18110 7296
rect 17862 7216 17868 7268
rect 17920 7256 17926 7268
rect 17957 7259 18015 7265
rect 17957 7256 17969 7259
rect 17920 7228 17969 7256
rect 17920 7216 17926 7228
rect 17957 7225 17969 7228
rect 18003 7225 18015 7259
rect 17957 7219 18015 7225
rect 19334 7216 19340 7268
rect 19392 7216 19398 7268
rect 19426 7216 19432 7268
rect 19484 7256 19490 7268
rect 19484 7228 19748 7256
rect 19484 7216 19490 7228
rect 14458 7188 14464 7200
rect 8772 7160 14464 7188
rect 14458 7148 14464 7160
rect 14516 7148 14522 7200
rect 17402 7148 17408 7200
rect 17460 7148 17466 7200
rect 19352 7188 19380 7216
rect 19613 7191 19671 7197
rect 19613 7188 19625 7191
rect 19352 7160 19625 7188
rect 19613 7157 19625 7160
rect 19659 7157 19671 7191
rect 19720 7188 19748 7228
rect 21174 7216 21180 7268
rect 21232 7216 21238 7268
rect 23842 7216 23848 7268
rect 23900 7256 23906 7268
rect 28626 7256 28632 7268
rect 23900 7228 28632 7256
rect 23900 7216 23906 7228
rect 28626 7216 28632 7228
rect 28684 7216 28690 7268
rect 19981 7191 20039 7197
rect 19981 7188 19993 7191
rect 19720 7160 19993 7188
rect 19613 7151 19671 7157
rect 19981 7157 19993 7160
rect 20027 7157 20039 7191
rect 19981 7151 20039 7157
rect 20622 7148 20628 7200
rect 20680 7148 20686 7200
rect 20714 7148 20720 7200
rect 20772 7188 20778 7200
rect 20901 7191 20959 7197
rect 20901 7188 20913 7191
rect 20772 7160 20913 7188
rect 20772 7148 20778 7160
rect 20901 7157 20913 7160
rect 20947 7157 20959 7191
rect 20901 7151 20959 7157
rect 21450 7148 21456 7200
rect 21508 7188 21514 7200
rect 21821 7191 21879 7197
rect 21821 7188 21833 7191
rect 21508 7160 21833 7188
rect 21508 7148 21514 7160
rect 21821 7157 21833 7160
rect 21867 7157 21879 7191
rect 21821 7151 21879 7157
rect 24762 7148 24768 7200
rect 24820 7148 24826 7200
rect 26050 7148 26056 7200
rect 26108 7188 26114 7200
rect 26145 7191 26203 7197
rect 26145 7188 26157 7191
rect 26108 7160 26157 7188
rect 26108 7148 26114 7160
rect 26145 7157 26157 7160
rect 26191 7157 26203 7191
rect 31726 7188 31754 7296
rect 33428 7188 33456 7488
rect 31726 7160 33456 7188
rect 26145 7151 26203 7157
rect 1104 7098 43516 7120
rect 1104 7046 6251 7098
rect 6303 7046 6315 7098
rect 6367 7046 6379 7098
rect 6431 7046 6443 7098
rect 6495 7046 6507 7098
rect 6559 7046 16854 7098
rect 16906 7046 16918 7098
rect 16970 7046 16982 7098
rect 17034 7046 17046 7098
rect 17098 7046 17110 7098
rect 17162 7046 27457 7098
rect 27509 7046 27521 7098
rect 27573 7046 27585 7098
rect 27637 7046 27649 7098
rect 27701 7046 27713 7098
rect 27765 7046 38060 7098
rect 38112 7046 38124 7098
rect 38176 7046 38188 7098
rect 38240 7046 38252 7098
rect 38304 7046 38316 7098
rect 38368 7046 43516 7098
rect 1104 7024 43516 7046
rect 7282 6944 7288 6996
rect 7340 6984 7346 6996
rect 12342 6984 12348 6996
rect 7340 6956 12348 6984
rect 7340 6944 7346 6956
rect 12342 6944 12348 6956
rect 12400 6944 12406 6996
rect 14642 6944 14648 6996
rect 14700 6984 14706 6996
rect 24762 6984 24768 6996
rect 14700 6956 24768 6984
rect 14700 6944 14706 6956
rect 24762 6944 24768 6956
rect 24820 6944 24826 6996
rect 25222 6944 25228 6996
rect 25280 6944 25286 6996
rect 8110 6876 8116 6928
rect 8168 6916 8174 6928
rect 8168 6888 16528 6916
rect 8168 6876 8174 6888
rect 9214 6808 9220 6860
rect 9272 6848 9278 6860
rect 10134 6848 10140 6860
rect 9272 6820 10140 6848
rect 9272 6808 9278 6820
rect 10134 6808 10140 6820
rect 10192 6808 10198 6860
rect 10686 6808 10692 6860
rect 10744 6808 10750 6860
rect 16500 6848 16528 6888
rect 17494 6876 17500 6928
rect 17552 6916 17558 6928
rect 25240 6916 25268 6944
rect 17552 6888 25268 6916
rect 17552 6876 17558 6888
rect 21818 6848 21824 6860
rect 16500 6820 21824 6848
rect 21818 6808 21824 6820
rect 21876 6808 21882 6860
rect 38562 6808 38568 6860
rect 38620 6848 38626 6860
rect 39114 6848 39120 6860
rect 38620 6820 39120 6848
rect 38620 6808 38626 6820
rect 39114 6808 39120 6820
rect 39172 6808 39178 6860
rect 10704 6780 10732 6808
rect 17954 6780 17960 6792
rect 10704 6752 17960 6780
rect 17954 6740 17960 6752
rect 18012 6740 18018 6792
rect 18046 6740 18052 6792
rect 18104 6740 18110 6792
rect 18230 6740 18236 6792
rect 18288 6740 18294 6792
rect 18322 6740 18328 6792
rect 18380 6740 18386 6792
rect 19610 6740 19616 6792
rect 19668 6780 19674 6792
rect 19797 6783 19855 6789
rect 19797 6780 19809 6783
rect 19668 6752 19809 6780
rect 19668 6740 19674 6752
rect 19797 6749 19809 6752
rect 19843 6749 19855 6783
rect 19797 6743 19855 6749
rect 19886 6740 19892 6792
rect 19944 6780 19950 6792
rect 19944 6752 20024 6780
rect 19944 6740 19950 6752
rect 14458 6672 14464 6724
rect 14516 6712 14522 6724
rect 18064 6712 18092 6740
rect 14516 6684 18092 6712
rect 14516 6672 14522 6684
rect 18248 6644 18276 6740
rect 18340 6712 18368 6740
rect 19996 6712 20024 6752
rect 20070 6740 20076 6792
rect 20128 6740 20134 6792
rect 36906 6740 36912 6792
rect 36964 6780 36970 6792
rect 38654 6780 38660 6792
rect 36964 6752 38660 6780
rect 36964 6740 36970 6752
rect 38654 6740 38660 6752
rect 38712 6740 38718 6792
rect 28718 6712 28724 6724
rect 18340 6684 19932 6712
rect 19996 6684 28724 6712
rect 19904 6653 19932 6684
rect 28718 6672 28724 6684
rect 28776 6672 28782 6724
rect 37182 6672 37188 6724
rect 37240 6712 37246 6724
rect 38746 6712 38752 6724
rect 37240 6684 38752 6712
rect 37240 6672 37246 6684
rect 38746 6672 38752 6684
rect 38804 6672 38810 6724
rect 19613 6647 19671 6653
rect 19613 6644 19625 6647
rect 18248 6616 19625 6644
rect 19613 6613 19625 6616
rect 19659 6613 19671 6647
rect 19613 6607 19671 6613
rect 19889 6647 19947 6653
rect 19889 6613 19901 6647
rect 19935 6613 19947 6647
rect 19889 6607 19947 6613
rect 1104 6554 43675 6576
rect 1104 6502 11552 6554
rect 11604 6502 11616 6554
rect 11668 6502 11680 6554
rect 11732 6502 11744 6554
rect 11796 6502 11808 6554
rect 11860 6502 22155 6554
rect 22207 6502 22219 6554
rect 22271 6502 22283 6554
rect 22335 6502 22347 6554
rect 22399 6502 22411 6554
rect 22463 6502 32758 6554
rect 32810 6502 32822 6554
rect 32874 6502 32886 6554
rect 32938 6502 32950 6554
rect 33002 6502 33014 6554
rect 33066 6502 43361 6554
rect 43413 6502 43425 6554
rect 43477 6502 43489 6554
rect 43541 6502 43553 6554
rect 43605 6502 43617 6554
rect 43669 6502 43675 6554
rect 1104 6480 43675 6502
rect 15194 6400 15200 6452
rect 15252 6440 15258 6452
rect 20254 6440 20260 6452
rect 15252 6412 20260 6440
rect 15252 6400 15258 6412
rect 20254 6400 20260 6412
rect 20312 6400 20318 6452
rect 16114 6332 16120 6384
rect 16172 6372 16178 6384
rect 20346 6372 20352 6384
rect 16172 6344 20352 6372
rect 16172 6332 16178 6344
rect 20346 6332 20352 6344
rect 20404 6332 20410 6384
rect 16574 6264 16580 6316
rect 16632 6304 16638 6316
rect 20622 6304 20628 6316
rect 16632 6276 20628 6304
rect 16632 6264 16638 6276
rect 20622 6264 20628 6276
rect 20680 6264 20686 6316
rect 1104 6010 43516 6032
rect 1104 5958 6251 6010
rect 6303 5958 6315 6010
rect 6367 5958 6379 6010
rect 6431 5958 6443 6010
rect 6495 5958 6507 6010
rect 6559 5958 16854 6010
rect 16906 5958 16918 6010
rect 16970 5958 16982 6010
rect 17034 5958 17046 6010
rect 17098 5958 17110 6010
rect 17162 5958 27457 6010
rect 27509 5958 27521 6010
rect 27573 5958 27585 6010
rect 27637 5958 27649 6010
rect 27701 5958 27713 6010
rect 27765 5958 38060 6010
rect 38112 5958 38124 6010
rect 38176 5958 38188 6010
rect 38240 5958 38252 6010
rect 38304 5958 38316 6010
rect 38368 5958 43516 6010
rect 1104 5936 43516 5958
rect 25958 5652 25964 5704
rect 26016 5692 26022 5704
rect 30466 5692 30472 5704
rect 26016 5664 30472 5692
rect 26016 5652 26022 5664
rect 30466 5652 30472 5664
rect 30524 5652 30530 5704
rect 23014 5584 23020 5636
rect 23072 5624 23078 5636
rect 35342 5624 35348 5636
rect 23072 5596 35348 5624
rect 23072 5584 23078 5596
rect 35342 5584 35348 5596
rect 35400 5584 35406 5636
rect 1104 5466 43675 5488
rect 1104 5414 11552 5466
rect 11604 5414 11616 5466
rect 11668 5414 11680 5466
rect 11732 5414 11744 5466
rect 11796 5414 11808 5466
rect 11860 5414 22155 5466
rect 22207 5414 22219 5466
rect 22271 5414 22283 5466
rect 22335 5414 22347 5466
rect 22399 5414 22411 5466
rect 22463 5414 32758 5466
rect 32810 5414 32822 5466
rect 32874 5414 32886 5466
rect 32938 5414 32950 5466
rect 33002 5414 33014 5466
rect 33066 5414 43361 5466
rect 43413 5414 43425 5466
rect 43477 5414 43489 5466
rect 43541 5414 43553 5466
rect 43605 5414 43617 5466
rect 43669 5414 43675 5466
rect 1104 5392 43675 5414
rect 37553 5355 37611 5361
rect 37553 5321 37565 5355
rect 37599 5352 37611 5355
rect 39298 5352 39304 5364
rect 37599 5324 39304 5352
rect 37599 5321 37611 5324
rect 37553 5315 37611 5321
rect 39298 5312 39304 5324
rect 39356 5312 39362 5364
rect 37366 5176 37372 5228
rect 37424 5176 37430 5228
rect 23842 5108 23848 5160
rect 23900 5148 23906 5160
rect 32674 5148 32680 5160
rect 23900 5120 32680 5148
rect 23900 5108 23906 5120
rect 32674 5108 32680 5120
rect 32732 5108 32738 5160
rect 1104 4922 43516 4944
rect 1104 4870 6251 4922
rect 6303 4870 6315 4922
rect 6367 4870 6379 4922
rect 6431 4870 6443 4922
rect 6495 4870 6507 4922
rect 6559 4870 16854 4922
rect 16906 4870 16918 4922
rect 16970 4870 16982 4922
rect 17034 4870 17046 4922
rect 17098 4870 17110 4922
rect 17162 4870 27457 4922
rect 27509 4870 27521 4922
rect 27573 4870 27585 4922
rect 27637 4870 27649 4922
rect 27701 4870 27713 4922
rect 27765 4870 38060 4922
rect 38112 4870 38124 4922
rect 38176 4870 38188 4922
rect 38240 4870 38252 4922
rect 38304 4870 38316 4922
rect 38368 4870 43516 4922
rect 1104 4848 43516 4870
rect 23014 4768 23020 4820
rect 23072 4768 23078 4820
rect 23842 4768 23848 4820
rect 23900 4768 23906 4820
rect 25958 4768 25964 4820
rect 26016 4768 26022 4820
rect 28074 4768 28080 4820
rect 28132 4768 28138 4820
rect 36814 4808 36820 4820
rect 31726 4780 36820 4808
rect 22741 4743 22799 4749
rect 22741 4709 22753 4743
rect 22787 4709 22799 4743
rect 22741 4703 22799 4709
rect 23293 4743 23351 4749
rect 23293 4709 23305 4743
rect 23339 4740 23351 4743
rect 31726 4740 31754 4780
rect 36814 4768 36820 4780
rect 36872 4768 36878 4820
rect 36909 4811 36967 4817
rect 36909 4777 36921 4811
rect 36955 4808 36967 4811
rect 37366 4808 37372 4820
rect 36955 4780 37372 4808
rect 36955 4777 36967 4780
rect 36909 4771 36967 4777
rect 37366 4768 37372 4780
rect 37424 4768 37430 4820
rect 38197 4811 38255 4817
rect 38197 4777 38209 4811
rect 38243 4808 38255 4811
rect 38378 4808 38384 4820
rect 38243 4780 38384 4808
rect 38243 4777 38255 4780
rect 38197 4771 38255 4777
rect 38378 4768 38384 4780
rect 38436 4768 38442 4820
rect 23339 4712 31754 4740
rect 32309 4743 32367 4749
rect 23339 4709 23351 4712
rect 23293 4703 23351 4709
rect 32309 4709 32321 4743
rect 32355 4740 32367 4743
rect 37918 4740 37924 4752
rect 32355 4712 37924 4740
rect 32355 4709 32367 4712
rect 32309 4703 32367 4709
rect 22756 4672 22784 4703
rect 37918 4700 37924 4712
rect 37976 4700 37982 4752
rect 31110 4672 31116 4684
rect 22756 4644 31116 4672
rect 31110 4632 31116 4644
rect 31168 4632 31174 4684
rect 21542 4564 21548 4616
rect 21600 4564 21606 4616
rect 22554 4564 22560 4616
rect 22612 4564 22618 4616
rect 22830 4564 22836 4616
rect 22888 4564 22894 4616
rect 23109 4607 23167 4613
rect 23109 4573 23121 4607
rect 23155 4573 23167 4607
rect 23109 4567 23167 4573
rect 22646 4496 22652 4548
rect 22704 4536 22710 4548
rect 23124 4536 23152 4567
rect 23658 4564 23664 4616
rect 23716 4564 23722 4616
rect 25774 4564 25780 4616
rect 25832 4564 25838 4616
rect 27890 4564 27896 4616
rect 27948 4564 27954 4616
rect 32122 4564 32128 4616
rect 32180 4564 32186 4616
rect 34514 4564 34520 4616
rect 34572 4604 34578 4616
rect 36725 4607 36783 4613
rect 36725 4604 36737 4607
rect 34572 4576 36737 4604
rect 34572 4564 34578 4576
rect 36725 4573 36737 4576
rect 36771 4573 36783 4607
rect 36725 4567 36783 4573
rect 38010 4564 38016 4616
rect 38068 4564 38074 4616
rect 22704 4508 23152 4536
rect 22704 4496 22710 4508
rect 21729 4471 21787 4477
rect 21729 4437 21741 4471
rect 21775 4468 21787 4471
rect 29270 4468 29276 4480
rect 21775 4440 29276 4468
rect 21775 4437 21787 4440
rect 21729 4431 21787 4437
rect 29270 4428 29276 4440
rect 29328 4428 29334 4480
rect 1104 4378 43675 4400
rect 1104 4326 11552 4378
rect 11604 4326 11616 4378
rect 11668 4326 11680 4378
rect 11732 4326 11744 4378
rect 11796 4326 11808 4378
rect 11860 4326 22155 4378
rect 22207 4326 22219 4378
rect 22271 4326 22283 4378
rect 22335 4326 22347 4378
rect 22399 4326 22411 4378
rect 22463 4326 32758 4378
rect 32810 4326 32822 4378
rect 32874 4326 32886 4378
rect 32938 4326 32950 4378
rect 33002 4326 33014 4378
rect 33066 4326 43361 4378
rect 43413 4326 43425 4378
rect 43477 4326 43489 4378
rect 43541 4326 43553 4378
rect 43605 4326 43617 4378
rect 43669 4326 43675 4378
rect 1104 4304 43675 4326
rect 20901 4267 20959 4273
rect 20901 4233 20913 4267
rect 20947 4264 20959 4267
rect 21542 4264 21548 4276
rect 20947 4236 21548 4264
rect 20947 4233 20959 4236
rect 20901 4227 20959 4233
rect 21542 4224 21548 4236
rect 21600 4224 21606 4276
rect 22005 4267 22063 4273
rect 22005 4233 22017 4267
rect 22051 4264 22063 4267
rect 22554 4264 22560 4276
rect 22051 4236 22560 4264
rect 22051 4233 22063 4236
rect 22005 4227 22063 4233
rect 22554 4224 22560 4236
rect 22612 4224 22618 4276
rect 25133 4267 25191 4273
rect 25133 4233 25145 4267
rect 25179 4264 25191 4267
rect 25774 4264 25780 4276
rect 25179 4236 25780 4264
rect 25179 4233 25191 4236
rect 25133 4227 25191 4233
rect 25774 4224 25780 4236
rect 25832 4224 25838 4276
rect 37645 4267 37703 4273
rect 37645 4233 37657 4267
rect 37691 4264 37703 4267
rect 38010 4264 38016 4276
rect 37691 4236 38016 4264
rect 37691 4233 37703 4236
rect 37645 4227 37703 4233
rect 38010 4224 38016 4236
rect 38068 4224 38074 4276
rect 20438 4088 20444 4140
rect 20496 4128 20502 4140
rect 20717 4131 20775 4137
rect 20717 4128 20729 4131
rect 20496 4100 20729 4128
rect 20496 4088 20502 4100
rect 20717 4097 20729 4100
rect 20763 4097 20775 4131
rect 20717 4091 20775 4097
rect 21821 4131 21879 4137
rect 21821 4097 21833 4131
rect 21867 4097 21879 4131
rect 21821 4091 21879 4097
rect 22097 4131 22155 4137
rect 22097 4097 22109 4131
rect 22143 4097 22155 4131
rect 22097 4091 22155 4097
rect 22373 4131 22431 4137
rect 22373 4097 22385 4131
rect 22419 4097 22431 4131
rect 22373 4091 22431 4097
rect 7742 4020 7748 4072
rect 7800 4060 7806 4072
rect 21836 4060 21864 4091
rect 7800 4032 21864 4060
rect 7800 4020 7806 4032
rect 5626 3952 5632 4004
rect 5684 3992 5690 4004
rect 22112 3992 22140 4091
rect 22388 3992 22416 4091
rect 22462 4088 22468 4140
rect 22520 4128 22526 4140
rect 22649 4131 22707 4137
rect 22649 4128 22661 4131
rect 22520 4100 22661 4128
rect 22520 4088 22526 4100
rect 22649 4097 22661 4100
rect 22695 4097 22707 4131
rect 22649 4091 22707 4097
rect 24762 4088 24768 4140
rect 24820 4128 24826 4140
rect 24949 4131 25007 4137
rect 24949 4128 24961 4131
rect 24820 4100 24961 4128
rect 24820 4088 24826 4100
rect 24949 4097 24961 4100
rect 24995 4097 25007 4131
rect 24949 4091 25007 4097
rect 27062 4088 27068 4140
rect 27120 4088 27126 4140
rect 31294 4088 31300 4140
rect 31352 4088 31358 4140
rect 37458 4088 37464 4140
rect 37516 4088 37522 4140
rect 39758 4088 39764 4140
rect 39816 4088 39822 4140
rect 22830 4020 22836 4072
rect 22888 4020 22894 4072
rect 27890 4060 27896 4072
rect 27264 4032 27896 4060
rect 22848 3992 22876 4020
rect 27264 4001 27292 4032
rect 27890 4020 27896 4032
rect 27948 4020 27954 4072
rect 32122 4020 32128 4072
rect 32180 4020 32186 4072
rect 5684 3964 22140 3992
rect 22204 3964 22416 3992
rect 22480 3964 22876 3992
rect 27249 3995 27307 4001
rect 5684 3952 5690 3964
rect 19518 3884 19524 3936
rect 19576 3924 19582 3936
rect 22204 3924 22232 3964
rect 19576 3896 22232 3924
rect 22281 3927 22339 3933
rect 19576 3884 19582 3896
rect 22281 3893 22293 3927
rect 22327 3924 22339 3927
rect 22480 3924 22508 3964
rect 27249 3961 27261 3995
rect 27295 3961 27307 3995
rect 27249 3955 27307 3961
rect 31481 3995 31539 4001
rect 31481 3961 31493 3995
rect 31527 3992 31539 3995
rect 32140 3992 32168 4020
rect 31527 3964 32168 3992
rect 31527 3961 31539 3964
rect 31481 3955 31539 3961
rect 22327 3896 22508 3924
rect 22557 3927 22615 3933
rect 22327 3893 22339 3896
rect 22281 3887 22339 3893
rect 22557 3893 22569 3927
rect 22603 3924 22615 3927
rect 22646 3924 22652 3936
rect 22603 3896 22652 3924
rect 22603 3893 22615 3896
rect 22557 3887 22615 3893
rect 22646 3884 22652 3896
rect 22704 3884 22710 3936
rect 22833 3927 22891 3933
rect 22833 3893 22845 3927
rect 22879 3924 22891 3927
rect 31386 3924 31392 3936
rect 22879 3896 31392 3924
rect 22879 3893 22891 3896
rect 22833 3887 22891 3893
rect 31386 3884 31392 3896
rect 31444 3884 31450 3936
rect 39850 3884 39856 3936
rect 39908 3924 39914 3936
rect 39945 3927 40003 3933
rect 39945 3924 39957 3927
rect 39908 3896 39957 3924
rect 39908 3884 39914 3896
rect 39945 3893 39957 3896
rect 39991 3893 40003 3927
rect 39945 3887 40003 3893
rect 1104 3834 43516 3856
rect 1104 3782 6251 3834
rect 6303 3782 6315 3834
rect 6367 3782 6379 3834
rect 6431 3782 6443 3834
rect 6495 3782 6507 3834
rect 6559 3782 16854 3834
rect 16906 3782 16918 3834
rect 16970 3782 16982 3834
rect 17034 3782 17046 3834
rect 17098 3782 17110 3834
rect 17162 3782 27457 3834
rect 27509 3782 27521 3834
rect 27573 3782 27585 3834
rect 27637 3782 27649 3834
rect 27701 3782 27713 3834
rect 27765 3782 38060 3834
rect 38112 3782 38124 3834
rect 38176 3782 38188 3834
rect 38240 3782 38252 3834
rect 38304 3782 38316 3834
rect 38368 3782 43516 3834
rect 1104 3760 43516 3782
rect 22097 3723 22155 3729
rect 22097 3689 22109 3723
rect 22143 3720 22155 3723
rect 22462 3720 22468 3732
rect 22143 3692 22468 3720
rect 22143 3689 22155 3692
rect 22097 3683 22155 3689
rect 22462 3680 22468 3692
rect 22520 3680 22526 3732
rect 23017 3723 23075 3729
rect 23017 3689 23029 3723
rect 23063 3720 23075 3723
rect 23658 3720 23664 3732
rect 23063 3692 23664 3720
rect 23063 3689 23075 3692
rect 23017 3683 23075 3689
rect 23658 3680 23664 3692
rect 23716 3680 23722 3732
rect 30193 3723 30251 3729
rect 30193 3689 30205 3723
rect 30239 3720 30251 3723
rect 34606 3720 34612 3732
rect 30239 3692 34612 3720
rect 30239 3689 30251 3692
rect 30193 3683 30251 3689
rect 34606 3680 34612 3692
rect 34664 3680 34670 3732
rect 37277 3723 37335 3729
rect 37277 3689 37289 3723
rect 37323 3720 37335 3723
rect 39574 3720 39580 3732
rect 37323 3692 39580 3720
rect 37323 3689 37335 3692
rect 37277 3683 37335 3689
rect 39574 3680 39580 3692
rect 39632 3680 39638 3732
rect 39758 3680 39764 3732
rect 39816 3720 39822 3732
rect 40497 3723 40555 3729
rect 40497 3720 40509 3723
rect 39816 3692 40509 3720
rect 39816 3680 39822 3692
rect 40497 3689 40509 3692
rect 40543 3689 40555 3723
rect 40497 3683 40555 3689
rect 19613 3655 19671 3661
rect 19613 3621 19625 3655
rect 19659 3652 19671 3655
rect 36262 3652 36268 3664
rect 19659 3624 36268 3652
rect 19659 3621 19671 3624
rect 19613 3615 19671 3621
rect 36262 3612 36268 3624
rect 36320 3612 36326 3664
rect 19426 3476 19432 3528
rect 19484 3476 19490 3528
rect 21913 3519 21971 3525
rect 21913 3516 21925 3519
rect 19536 3488 21925 3516
rect 19242 3408 19248 3460
rect 19300 3448 19306 3460
rect 19536 3448 19564 3488
rect 21913 3485 21925 3488
rect 21959 3485 21971 3519
rect 21913 3479 21971 3485
rect 22002 3476 22008 3528
rect 22060 3516 22066 3528
rect 22189 3519 22247 3525
rect 22189 3516 22201 3519
rect 22060 3488 22201 3516
rect 22060 3476 22066 3488
rect 22189 3485 22201 3488
rect 22235 3485 22247 3519
rect 22189 3479 22247 3485
rect 22465 3519 22523 3525
rect 22465 3485 22477 3519
rect 22511 3485 22523 3519
rect 22465 3479 22523 3485
rect 19300 3420 19564 3448
rect 19300 3408 19306 3420
rect 21266 3408 21272 3460
rect 21324 3448 21330 3460
rect 22480 3448 22508 3479
rect 22830 3476 22836 3528
rect 22888 3476 22894 3528
rect 30006 3476 30012 3528
rect 30064 3476 30070 3528
rect 35710 3476 35716 3528
rect 35768 3476 35774 3528
rect 37090 3476 37096 3528
rect 37148 3476 37154 3528
rect 40678 3476 40684 3528
rect 40736 3476 40742 3528
rect 35728 3448 35756 3476
rect 21324 3420 22508 3448
rect 22572 3420 35756 3448
rect 21324 3408 21330 3420
rect 22373 3383 22431 3389
rect 22373 3349 22385 3383
rect 22419 3380 22431 3383
rect 22572 3380 22600 3420
rect 22419 3352 22600 3380
rect 22649 3383 22707 3389
rect 22419 3349 22431 3352
rect 22373 3343 22431 3349
rect 22649 3349 22661 3383
rect 22695 3380 22707 3383
rect 36630 3380 36636 3392
rect 22695 3352 36636 3380
rect 22695 3349 22707 3352
rect 22649 3343 22707 3349
rect 36630 3340 36636 3352
rect 36688 3340 36694 3392
rect 1104 3290 43675 3312
rect 1104 3238 11552 3290
rect 11604 3238 11616 3290
rect 11668 3238 11680 3290
rect 11732 3238 11744 3290
rect 11796 3238 11808 3290
rect 11860 3238 22155 3290
rect 22207 3238 22219 3290
rect 22271 3238 22283 3290
rect 22335 3238 22347 3290
rect 22399 3238 22411 3290
rect 22463 3238 32758 3290
rect 32810 3238 32822 3290
rect 32874 3238 32886 3290
rect 32938 3238 32950 3290
rect 33002 3238 33014 3290
rect 33066 3238 43361 3290
rect 43413 3238 43425 3290
rect 43477 3238 43489 3290
rect 43541 3238 43553 3290
rect 43605 3238 43617 3290
rect 43669 3238 43675 3290
rect 1104 3216 43675 3238
rect 18785 3179 18843 3185
rect 18785 3145 18797 3179
rect 18831 3176 18843 3179
rect 19426 3176 19432 3188
rect 18831 3148 19432 3176
rect 18831 3145 18843 3148
rect 18785 3139 18843 3145
rect 19426 3136 19432 3148
rect 19484 3136 19490 3188
rect 21266 3136 21272 3188
rect 21324 3136 21330 3188
rect 21545 3179 21603 3185
rect 21545 3145 21557 3179
rect 21591 3176 21603 3179
rect 22002 3176 22008 3188
rect 21591 3148 22008 3176
rect 21591 3145 21603 3148
rect 21545 3139 21603 3145
rect 22002 3136 22008 3148
rect 22060 3136 22066 3188
rect 29365 3179 29423 3185
rect 29365 3145 29377 3179
rect 29411 3176 29423 3179
rect 30006 3176 30012 3188
rect 29411 3148 30012 3176
rect 29411 3145 29423 3148
rect 29365 3139 29423 3145
rect 30006 3136 30012 3148
rect 30064 3136 30070 3188
rect 36173 3179 36231 3185
rect 36173 3145 36185 3179
rect 36219 3176 36231 3179
rect 37090 3176 37096 3188
rect 36219 3148 37096 3176
rect 36219 3145 36231 3148
rect 36173 3139 36231 3145
rect 37090 3136 37096 3148
rect 37148 3136 37154 3188
rect 39945 3179 40003 3185
rect 39945 3145 39957 3179
rect 39991 3176 40003 3179
rect 41046 3176 41052 3188
rect 39991 3148 41052 3176
rect 39991 3145 40003 3148
rect 39945 3139 40003 3145
rect 41046 3136 41052 3148
rect 41104 3136 41110 3188
rect 18598 3000 18604 3052
rect 18656 3000 18662 3052
rect 21085 3043 21143 3049
rect 21085 3009 21097 3043
rect 21131 3009 21143 3043
rect 21085 3003 21143 3009
rect 16206 2932 16212 2984
rect 16264 2972 16270 2984
rect 21100 2972 21128 3003
rect 21358 3000 21364 3052
rect 21416 3000 21422 3052
rect 22646 3000 22652 3052
rect 22704 3000 22710 3052
rect 28902 3000 28908 3052
rect 28960 3040 28966 3052
rect 29181 3043 29239 3049
rect 29181 3040 29193 3043
rect 28960 3012 29193 3040
rect 28960 3000 28966 3012
rect 29181 3009 29193 3012
rect 29227 3009 29239 3043
rect 29181 3003 29239 3009
rect 35250 3000 35256 3052
rect 35308 3040 35314 3052
rect 35989 3043 36047 3049
rect 35989 3040 36001 3043
rect 35308 3012 36001 3040
rect 35308 3000 35314 3012
rect 35989 3009 36001 3012
rect 36035 3009 36047 3043
rect 35989 3003 36047 3009
rect 39761 3043 39819 3049
rect 39761 3009 39773 3043
rect 39807 3040 39819 3043
rect 40218 3040 40224 3052
rect 39807 3012 40224 3040
rect 39807 3009 39819 3012
rect 39761 3003 39819 3009
rect 40218 3000 40224 3012
rect 40276 3000 40282 3052
rect 16264 2944 21128 2972
rect 16264 2932 16270 2944
rect 22833 2907 22891 2913
rect 22833 2873 22845 2907
rect 22879 2904 22891 2907
rect 23382 2904 23388 2916
rect 22879 2876 23388 2904
rect 22879 2873 22891 2876
rect 22833 2867 22891 2873
rect 23382 2864 23388 2876
rect 23440 2864 23446 2916
rect 1104 2746 43516 2768
rect 1104 2694 6251 2746
rect 6303 2694 6315 2746
rect 6367 2694 6379 2746
rect 6431 2694 6443 2746
rect 6495 2694 6507 2746
rect 6559 2694 16854 2746
rect 16906 2694 16918 2746
rect 16970 2694 16982 2746
rect 17034 2694 17046 2746
rect 17098 2694 17110 2746
rect 17162 2694 27457 2746
rect 27509 2694 27521 2746
rect 27573 2694 27585 2746
rect 27637 2694 27649 2746
rect 27701 2694 27713 2746
rect 27765 2694 38060 2746
rect 38112 2694 38124 2746
rect 38176 2694 38188 2746
rect 38240 2694 38252 2746
rect 38304 2694 38316 2746
rect 38368 2694 43516 2746
rect 1104 2672 43516 2694
rect 22097 2635 22155 2641
rect 22097 2601 22109 2635
rect 22143 2632 22155 2635
rect 22646 2632 22652 2644
rect 22143 2604 22652 2632
rect 22143 2601 22155 2604
rect 22097 2595 22155 2601
rect 22646 2592 22652 2604
rect 22704 2592 22710 2644
rect 39209 2635 39267 2641
rect 39209 2601 39221 2635
rect 39255 2632 39267 2635
rect 39942 2632 39948 2644
rect 39255 2604 39948 2632
rect 39255 2601 39267 2604
rect 39209 2595 39267 2601
rect 39942 2592 39948 2604
rect 40000 2592 40006 2644
rect 40218 2592 40224 2644
rect 40276 2592 40282 2644
rect 3510 2388 3516 2440
rect 3568 2428 3574 2440
rect 21913 2431 21971 2437
rect 21913 2428 21925 2431
rect 3568 2400 21925 2428
rect 3568 2388 3574 2400
rect 21913 2397 21925 2400
rect 21959 2397 21971 2431
rect 21913 2391 21971 2397
rect 39022 2388 39028 2440
rect 39080 2388 39086 2440
rect 40405 2431 40463 2437
rect 40405 2397 40417 2431
rect 40451 2428 40463 2431
rect 42978 2428 42984 2440
rect 40451 2400 42984 2428
rect 40451 2397 40463 2400
rect 40405 2391 40463 2397
rect 42978 2388 42984 2400
rect 43036 2388 43042 2440
rect 1104 2202 43675 2224
rect 1104 2150 11552 2202
rect 11604 2150 11616 2202
rect 11668 2150 11680 2202
rect 11732 2150 11744 2202
rect 11796 2150 11808 2202
rect 11860 2150 22155 2202
rect 22207 2150 22219 2202
rect 22271 2150 22283 2202
rect 22335 2150 22347 2202
rect 22399 2150 22411 2202
rect 22463 2150 32758 2202
rect 32810 2150 32822 2202
rect 32874 2150 32886 2202
rect 32938 2150 32950 2202
rect 33002 2150 33014 2202
rect 33066 2150 43361 2202
rect 43413 2150 43425 2202
rect 43477 2150 43489 2202
rect 43541 2150 43553 2202
rect 43605 2150 43617 2202
rect 43669 2150 43675 2202
rect 1104 2128 43675 2150
rect 39022 2048 39028 2100
rect 39080 2048 39086 2100
rect 1578 1912 1584 1964
rect 1636 1952 1642 1964
rect 21361 1955 21419 1961
rect 21361 1952 21373 1955
rect 1636 1924 21373 1952
rect 1636 1912 1642 1924
rect 21361 1921 21373 1924
rect 21407 1921 21419 1955
rect 21361 1915 21419 1921
rect 38838 1912 38844 1964
rect 38896 1912 38902 1964
rect 21545 1751 21603 1757
rect 21545 1717 21557 1751
rect 21591 1748 21603 1751
rect 33962 1748 33968 1760
rect 21591 1720 33968 1748
rect 21591 1717 21603 1720
rect 21545 1711 21603 1717
rect 33962 1708 33968 1720
rect 34020 1708 34026 1760
rect 1104 1658 43516 1680
rect 1104 1606 6251 1658
rect 6303 1606 6315 1658
rect 6367 1606 6379 1658
rect 6431 1606 6443 1658
rect 6495 1606 6507 1658
rect 6559 1606 16854 1658
rect 16906 1606 16918 1658
rect 16970 1606 16982 1658
rect 17034 1606 17046 1658
rect 17098 1606 17110 1658
rect 17162 1606 27457 1658
rect 27509 1606 27521 1658
rect 27573 1606 27585 1658
rect 27637 1606 27649 1658
rect 27701 1606 27713 1658
rect 27765 1606 38060 1658
rect 38112 1606 38124 1658
rect 38176 1606 38188 1658
rect 38240 1606 38252 1658
rect 38304 1606 38316 1658
rect 38368 1606 43516 1658
rect 1104 1584 43516 1606
rect 1578 1504 1584 1556
rect 1636 1504 1642 1556
rect 3510 1504 3516 1556
rect 3568 1504 3574 1556
rect 38838 1504 38844 1556
rect 38896 1544 38902 1556
rect 39301 1547 39359 1553
rect 39301 1544 39313 1547
rect 38896 1516 39313 1544
rect 38896 1504 38902 1516
rect 39301 1513 39313 1516
rect 39347 1513 39359 1547
rect 39301 1507 39359 1513
rect 42978 1504 42984 1556
rect 43036 1504 43042 1556
rect 14277 1479 14335 1485
rect 14277 1445 14289 1479
rect 14323 1445 14335 1479
rect 14277 1439 14335 1445
rect 1118 1300 1124 1352
rect 1176 1340 1182 1352
rect 1397 1343 1455 1349
rect 1397 1340 1409 1343
rect 1176 1312 1409 1340
rect 1176 1300 1182 1312
rect 1397 1309 1409 1312
rect 1443 1309 1455 1343
rect 1397 1303 1455 1309
rect 3326 1300 3332 1352
rect 3384 1300 3390 1352
rect 5442 1300 5448 1352
rect 5500 1300 5506 1352
rect 5626 1300 5632 1352
rect 5684 1300 5690 1352
rect 7558 1300 7564 1352
rect 7616 1300 7622 1352
rect 9674 1300 9680 1352
rect 9732 1300 9738 1352
rect 11790 1300 11796 1352
rect 11848 1300 11854 1352
rect 14090 1300 14096 1352
rect 14148 1300 14154 1352
rect 14292 1340 14320 1439
rect 15948 1380 16160 1408
rect 15948 1340 15976 1380
rect 14292 1312 15976 1340
rect 16022 1300 16028 1352
rect 16080 1300 16086 1352
rect 16132 1340 16160 1380
rect 18064 1380 18276 1408
rect 18064 1340 18092 1380
rect 16132 1312 18092 1340
rect 18138 1300 18144 1352
rect 18196 1300 18202 1352
rect 18248 1316 18276 1380
rect 5644 1213 5672 1300
rect 18248 1288 18368 1316
rect 18414 1300 18420 1352
rect 18472 1340 18478 1352
rect 19518 1340 19524 1352
rect 18472 1312 19524 1340
rect 18472 1300 18478 1312
rect 19518 1300 19524 1312
rect 19576 1300 19582 1352
rect 20254 1300 20260 1352
rect 20312 1300 20318 1352
rect 21358 1300 21364 1352
rect 21416 1300 21422 1352
rect 22370 1300 22376 1352
rect 22428 1300 22434 1352
rect 22738 1300 22744 1352
rect 22796 1300 22802 1352
rect 24486 1300 24492 1352
rect 24544 1300 24550 1352
rect 26602 1300 26608 1352
rect 26660 1300 26666 1352
rect 27062 1300 27068 1352
rect 27120 1300 27126 1352
rect 28718 1300 28724 1352
rect 28776 1300 28782 1352
rect 28902 1300 28908 1352
rect 28960 1300 28966 1352
rect 30834 1300 30840 1352
rect 30892 1300 30898 1352
rect 31294 1300 31300 1352
rect 31352 1300 31358 1352
rect 32674 1300 32680 1352
rect 32732 1340 32738 1352
rect 32953 1343 33011 1349
rect 32953 1340 32965 1343
rect 32732 1312 32965 1340
rect 32732 1300 32738 1312
rect 32953 1309 32965 1312
rect 32999 1309 33011 1343
rect 32953 1303 33011 1309
rect 34514 1300 34520 1352
rect 34572 1300 34578 1352
rect 35066 1300 35072 1352
rect 35124 1300 35130 1352
rect 35250 1300 35256 1352
rect 35308 1300 35314 1352
rect 37274 1300 37280 1352
rect 37332 1300 37338 1352
rect 37458 1300 37464 1352
rect 37516 1300 37522 1352
rect 39482 1300 39488 1352
rect 39540 1300 39546 1352
rect 40678 1300 40684 1352
rect 40736 1300 40742 1352
rect 41322 1300 41328 1352
rect 41380 1340 41386 1352
rect 41601 1343 41659 1349
rect 41601 1340 41613 1343
rect 41380 1312 41613 1340
rect 41380 1300 41386 1312
rect 41601 1309 41613 1312
rect 41647 1309 41659 1343
rect 41601 1303 41659 1309
rect 43162 1300 43168 1352
rect 43220 1300 43226 1352
rect 18340 1272 18368 1288
rect 21376 1272 21404 1300
rect 16132 1244 16574 1272
rect 18340 1244 21404 1272
rect 5629 1207 5687 1213
rect 5629 1173 5641 1207
rect 5675 1173 5687 1207
rect 5629 1167 5687 1173
rect 7742 1164 7748 1216
rect 7800 1164 7806 1216
rect 9858 1164 9864 1216
rect 9916 1164 9922 1216
rect 11977 1207 12035 1213
rect 11977 1173 11989 1207
rect 12023 1204 12035 1207
rect 16132 1204 16160 1244
rect 12023 1176 16160 1204
rect 12023 1173 12035 1176
rect 11977 1167 12035 1173
rect 16206 1164 16212 1216
rect 16264 1164 16270 1216
rect 16546 1204 16574 1244
rect 18230 1204 18236 1216
rect 16546 1176 18236 1204
rect 18230 1164 18236 1176
rect 18288 1164 18294 1216
rect 18325 1207 18383 1213
rect 18325 1173 18337 1207
rect 18371 1204 18383 1207
rect 18598 1204 18604 1216
rect 18371 1176 18604 1204
rect 18371 1173 18383 1176
rect 18325 1167 18383 1173
rect 18598 1164 18604 1176
rect 18656 1164 18662 1216
rect 20438 1164 20444 1216
rect 20496 1164 20502 1216
rect 22557 1207 22615 1213
rect 22557 1173 22569 1207
rect 22603 1204 22615 1207
rect 22756 1204 22784 1300
rect 24762 1232 24768 1284
rect 24820 1232 24826 1284
rect 22603 1176 22784 1204
rect 24673 1207 24731 1213
rect 22603 1173 22615 1176
rect 22557 1167 22615 1173
rect 24673 1173 24685 1207
rect 24719 1204 24731 1207
rect 24780 1204 24808 1232
rect 24719 1176 24808 1204
rect 26789 1207 26847 1213
rect 24719 1173 24731 1176
rect 24673 1167 24731 1173
rect 26789 1173 26801 1207
rect 26835 1204 26847 1207
rect 27080 1204 27108 1300
rect 28920 1213 28948 1300
rect 26835 1176 27108 1204
rect 28905 1207 28963 1213
rect 26835 1173 26847 1176
rect 26789 1167 26847 1173
rect 28905 1173 28917 1207
rect 28951 1173 28963 1207
rect 28905 1167 28963 1173
rect 31021 1207 31079 1213
rect 31021 1173 31033 1207
rect 31067 1204 31079 1207
rect 31312 1204 31340 1300
rect 31067 1176 31340 1204
rect 33137 1207 33195 1213
rect 31067 1173 31079 1176
rect 31021 1167 31079 1173
rect 33137 1173 33149 1207
rect 33183 1204 33195 1207
rect 34532 1204 34560 1300
rect 35268 1213 35296 1300
rect 37476 1213 37504 1300
rect 33183 1176 34560 1204
rect 35253 1207 35311 1213
rect 33183 1173 33195 1176
rect 33137 1167 33195 1173
rect 35253 1173 35265 1207
rect 35299 1173 35311 1207
rect 35253 1167 35311 1173
rect 37461 1207 37519 1213
rect 37461 1173 37473 1207
rect 37507 1173 37519 1207
rect 40696 1204 40724 1300
rect 41417 1207 41475 1213
rect 41417 1204 41429 1207
rect 40696 1176 41429 1204
rect 37461 1167 37519 1173
rect 41417 1173 41429 1176
rect 41463 1173 41475 1207
rect 41417 1167 41475 1173
rect 1104 1114 43675 1136
rect 1104 1062 11552 1114
rect 11604 1062 11616 1114
rect 11668 1062 11680 1114
rect 11732 1062 11744 1114
rect 11796 1062 11808 1114
rect 11860 1062 22155 1114
rect 22207 1062 22219 1114
rect 22271 1062 22283 1114
rect 22335 1062 22347 1114
rect 22399 1062 22411 1114
rect 22463 1062 32758 1114
rect 32810 1062 32822 1114
rect 32874 1062 32886 1114
rect 32938 1062 32950 1114
rect 33002 1062 33014 1114
rect 33066 1062 43361 1114
rect 43413 1062 43425 1114
rect 43477 1062 43489 1114
rect 43541 1062 43553 1114
rect 43605 1062 43617 1114
rect 43669 1062 43675 1114
rect 1104 1040 43675 1062
rect 9858 960 9864 1012
rect 9916 1000 9922 1012
rect 19242 1000 19248 1012
rect 9916 972 19248 1000
rect 9916 960 9922 972
rect 19242 960 19248 972
rect 19300 960 19306 1012
<< via1 >>
rect 11152 9936 11204 9988
rect 23020 9936 23072 9988
rect 23204 9936 23256 9988
rect 27160 9936 27212 9988
rect 19984 9868 20036 9920
rect 20168 9868 20220 9920
rect 23572 9868 23624 9920
rect 29276 9868 29328 9920
rect 17224 9800 17276 9852
rect 22100 9800 22152 9852
rect 22192 9800 22244 9852
rect 28172 9800 28224 9852
rect 8576 9596 8628 9648
rect 10784 9596 10836 9648
rect 16856 9596 16908 9648
rect 17776 9664 17828 9716
rect 18328 9664 18380 9716
rect 20168 9596 20220 9648
rect 17500 9528 17552 9580
rect 20720 9528 20772 9580
rect 21088 9732 21140 9784
rect 26792 9732 26844 9784
rect 33416 9800 33468 9852
rect 21548 9664 21600 9716
rect 30472 9664 30524 9716
rect 21916 9596 21968 9648
rect 22928 9596 22980 9648
rect 26884 9596 26936 9648
rect 20996 9528 21048 9580
rect 21824 9528 21876 9580
rect 31484 9528 31536 9580
rect 5540 9460 5592 9512
rect 14648 9460 14700 9512
rect 14740 9460 14792 9512
rect 21364 9460 21416 9512
rect 7288 9392 7340 9444
rect 17960 9392 18012 9444
rect 18604 9392 18656 9444
rect 31024 9460 31076 9512
rect 22192 9392 22244 9444
rect 31852 9392 31904 9444
rect 4712 9188 4764 9240
rect 22928 9324 22980 9376
rect 26792 9324 26844 9376
rect 37556 9392 37608 9444
rect 17224 9256 17276 9308
rect 18880 9256 18932 9308
rect 20996 9256 21048 9308
rect 23296 9256 23348 9308
rect 29920 9256 29972 9308
rect 38016 9324 38068 9376
rect 32128 9256 32180 9308
rect 12532 9188 12584 9240
rect 13820 9188 13872 9240
rect 13912 9188 13964 9240
rect 21640 9188 21692 9240
rect 24584 9188 24636 9240
rect 30748 9188 30800 9240
rect 34704 9188 34756 9240
rect 35072 9188 35124 9240
rect 11336 9120 11388 9172
rect 12256 9120 12308 9172
rect 12992 9120 13044 9172
rect 21824 9120 21876 9172
rect 21916 9120 21968 9172
rect 6184 8780 6236 8832
rect 8392 8984 8444 9036
rect 13636 8984 13688 9036
rect 13820 9052 13872 9104
rect 22100 9052 22152 9104
rect 22192 9052 22244 9104
rect 24952 9052 25004 9104
rect 25412 9120 25464 9172
rect 29368 9120 29420 9172
rect 24124 8984 24176 9036
rect 8668 8848 8720 8900
rect 16120 8916 16172 8968
rect 16304 8916 16356 8968
rect 17500 8916 17552 8968
rect 18512 8916 18564 8968
rect 30932 8984 30984 9036
rect 31576 8984 31628 9036
rect 34612 8984 34664 9036
rect 37464 8984 37516 9036
rect 9680 8780 9732 8832
rect 15200 8848 15252 8900
rect 15292 8848 15344 8900
rect 20812 8848 20864 8900
rect 20996 8848 21048 8900
rect 13360 8780 13412 8832
rect 21640 8780 21692 8832
rect 23112 8848 23164 8900
rect 24584 8848 24636 8900
rect 29828 8916 29880 8968
rect 31116 8916 31168 8968
rect 35900 8916 35952 8968
rect 27068 8848 27120 8900
rect 30380 8848 30432 8900
rect 37648 8780 37700 8832
rect 39304 8780 39356 8832
rect 11552 8678 11604 8730
rect 11616 8678 11668 8730
rect 11680 8678 11732 8730
rect 11744 8678 11796 8730
rect 11808 8678 11860 8730
rect 22155 8678 22207 8730
rect 22219 8678 22271 8730
rect 22283 8678 22335 8730
rect 22347 8678 22399 8730
rect 22411 8678 22463 8730
rect 32758 8678 32810 8730
rect 32822 8678 32874 8730
rect 32886 8678 32938 8730
rect 32950 8678 33002 8730
rect 33014 8678 33066 8730
rect 43361 8678 43413 8730
rect 43425 8678 43477 8730
rect 43489 8678 43541 8730
rect 43553 8678 43605 8730
rect 43617 8678 43669 8730
rect 5448 8576 5500 8628
rect 5540 8576 5592 8628
rect 5724 8576 5776 8628
rect 6276 8576 6328 8628
rect 6828 8576 6880 8628
rect 7288 8576 7340 8628
rect 7932 8576 7984 8628
rect 8484 8576 8536 8628
rect 4712 8483 4764 8492
rect 4712 8449 4721 8483
rect 4721 8449 4755 8483
rect 4755 8449 4764 8483
rect 4712 8440 4764 8449
rect 8392 8508 8444 8560
rect 9864 8576 9916 8628
rect 9588 8508 9640 8560
rect 10968 8576 11020 8628
rect 12072 8576 12124 8628
rect 12348 8576 12400 8628
rect 13084 8576 13136 8628
rect 13544 8576 13596 8628
rect 13636 8576 13688 8628
rect 14004 8576 14056 8628
rect 11428 8508 11480 8560
rect 6184 8483 6236 8492
rect 6184 8449 6193 8483
rect 6193 8449 6227 8483
rect 6227 8449 6236 8483
rect 6184 8440 6236 8449
rect 7196 8440 7248 8492
rect 8576 8440 8628 8492
rect 8668 8483 8720 8492
rect 8668 8449 8677 8483
rect 8677 8449 8711 8483
rect 8711 8449 8720 8483
rect 8668 8440 8720 8449
rect 9680 8440 9732 8492
rect 10784 8440 10836 8492
rect 11152 8440 11204 8492
rect 11336 8483 11388 8492
rect 11336 8449 11345 8483
rect 11345 8449 11379 8483
rect 11379 8449 11388 8483
rect 11336 8440 11388 8449
rect 12256 8440 12308 8492
rect 12532 8440 12584 8492
rect 12992 8483 13044 8492
rect 12992 8449 13001 8483
rect 13001 8449 13035 8483
rect 13035 8449 13044 8483
rect 12992 8440 13044 8449
rect 13360 8483 13412 8492
rect 13360 8449 13369 8483
rect 13369 8449 13403 8483
rect 13403 8449 13412 8483
rect 13360 8440 13412 8449
rect 5172 8304 5224 8356
rect 7656 8304 7708 8356
rect 9128 8347 9180 8356
rect 9128 8313 9137 8347
rect 9137 8313 9171 8347
rect 9171 8313 9180 8347
rect 9128 8304 9180 8313
rect 12716 8372 12768 8424
rect 13820 8551 13872 8560
rect 13820 8517 13829 8551
rect 13829 8517 13863 8551
rect 13863 8517 13872 8551
rect 13820 8508 13872 8517
rect 15384 8576 15436 8628
rect 16212 8576 16264 8628
rect 16764 8576 16816 8628
rect 15108 8508 15160 8560
rect 15292 8551 15344 8560
rect 15292 8517 15301 8551
rect 15301 8517 15335 8551
rect 15335 8517 15344 8551
rect 15292 8508 15344 8517
rect 17592 8576 17644 8628
rect 17868 8576 17920 8628
rect 18236 8619 18288 8628
rect 18236 8585 18245 8619
rect 18245 8585 18279 8619
rect 18279 8585 18288 8619
rect 18236 8576 18288 8585
rect 19064 8576 19116 8628
rect 17316 8508 17368 8560
rect 14740 8483 14792 8492
rect 14740 8449 14749 8483
rect 14749 8449 14783 8483
rect 14783 8449 14792 8483
rect 14740 8440 14792 8449
rect 16304 8440 16356 8492
rect 16764 8440 16816 8492
rect 16948 8372 17000 8424
rect 17408 8483 17460 8492
rect 17408 8449 17417 8483
rect 17417 8449 17451 8483
rect 17451 8449 17460 8483
rect 17408 8440 17460 8449
rect 18052 8440 18104 8492
rect 17316 8372 17368 8424
rect 17776 8372 17828 8424
rect 19064 8440 19116 8492
rect 19340 8508 19392 8560
rect 19616 8576 19668 8628
rect 19984 8576 20036 8628
rect 22468 8576 22520 8628
rect 22744 8576 22796 8628
rect 25964 8576 26016 8628
rect 27068 8576 27120 8628
rect 26976 8508 27028 8560
rect 19800 8483 19852 8492
rect 19800 8449 19809 8483
rect 19809 8449 19843 8483
rect 19843 8449 19852 8483
rect 19800 8440 19852 8449
rect 20444 8483 20496 8492
rect 20444 8449 20453 8483
rect 20453 8449 20487 8483
rect 20487 8449 20496 8483
rect 20444 8440 20496 8449
rect 20904 8440 20956 8492
rect 21180 8440 21232 8492
rect 21456 8440 21508 8492
rect 21548 8483 21600 8492
rect 21548 8449 21557 8483
rect 21557 8449 21591 8483
rect 21591 8449 21600 8483
rect 21548 8440 21600 8449
rect 21732 8440 21784 8492
rect 22100 8440 22152 8492
rect 22560 8483 22612 8492
rect 22560 8449 22569 8483
rect 22569 8449 22603 8483
rect 22603 8449 22612 8483
rect 22560 8440 22612 8449
rect 22836 8483 22888 8492
rect 22836 8449 22845 8483
rect 22845 8449 22879 8483
rect 22879 8449 22888 8483
rect 22836 8440 22888 8449
rect 22928 8440 22980 8492
rect 23388 8483 23440 8492
rect 23388 8449 23397 8483
rect 23397 8449 23431 8483
rect 23431 8449 23440 8483
rect 23388 8440 23440 8449
rect 23480 8440 23532 8492
rect 23940 8483 23992 8492
rect 23940 8449 23949 8483
rect 23949 8449 23983 8483
rect 23983 8449 23992 8483
rect 23940 8440 23992 8449
rect 24032 8440 24084 8492
rect 24400 8483 24452 8492
rect 24400 8449 24409 8483
rect 24409 8449 24443 8483
rect 24443 8449 24452 8483
rect 24400 8440 24452 8449
rect 24676 8483 24728 8492
rect 24676 8449 24685 8483
rect 24685 8449 24719 8483
rect 24719 8449 24728 8483
rect 24676 8440 24728 8449
rect 24768 8440 24820 8492
rect 25228 8483 25280 8492
rect 25228 8449 25237 8483
rect 25237 8449 25271 8483
rect 25271 8449 25280 8483
rect 25228 8440 25280 8449
rect 25320 8440 25372 8492
rect 25780 8483 25832 8492
rect 25780 8449 25789 8483
rect 25789 8449 25823 8483
rect 25823 8449 25832 8483
rect 25780 8440 25832 8449
rect 26056 8483 26108 8492
rect 26056 8449 26065 8483
rect 26065 8449 26099 8483
rect 26099 8449 26108 8483
rect 26056 8440 26108 8449
rect 26148 8440 26200 8492
rect 26608 8483 26660 8492
rect 26608 8449 26617 8483
rect 26617 8449 26651 8483
rect 26651 8449 26660 8483
rect 26608 8440 26660 8449
rect 26700 8440 26752 8492
rect 28080 8508 28132 8560
rect 29736 8576 29788 8628
rect 27528 8483 27580 8492
rect 27528 8449 27537 8483
rect 27537 8449 27571 8483
rect 27571 8449 27580 8483
rect 27528 8440 27580 8449
rect 27620 8440 27672 8492
rect 27988 8440 28040 8492
rect 19340 8372 19392 8424
rect 14188 8236 14240 8288
rect 16396 8304 16448 8356
rect 16580 8236 16632 8288
rect 16672 8236 16724 8288
rect 18328 8236 18380 8288
rect 18696 8304 18748 8356
rect 25412 8372 25464 8424
rect 29000 8508 29052 8560
rect 22192 8304 22244 8356
rect 20076 8236 20128 8288
rect 20352 8236 20404 8288
rect 20812 8279 20864 8288
rect 20812 8245 20821 8279
rect 20821 8245 20855 8279
rect 20855 8245 20864 8279
rect 20812 8236 20864 8245
rect 21088 8279 21140 8288
rect 21088 8245 21097 8279
rect 21097 8245 21131 8279
rect 21131 8245 21140 8279
rect 21088 8236 21140 8245
rect 21456 8236 21508 8288
rect 21548 8236 21600 8288
rect 22100 8279 22152 8288
rect 22100 8245 22109 8279
rect 22109 8245 22143 8279
rect 22143 8245 22152 8279
rect 22100 8236 22152 8245
rect 22376 8279 22428 8288
rect 22376 8245 22385 8279
rect 22385 8245 22419 8279
rect 22419 8245 22428 8279
rect 22376 8236 22428 8245
rect 24952 8304 25004 8356
rect 26148 8304 26200 8356
rect 27252 8304 27304 8356
rect 27896 8304 27948 8356
rect 28540 8304 28592 8356
rect 28908 8440 28960 8492
rect 29644 8508 29696 8560
rect 29184 8372 29236 8424
rect 29828 8440 29880 8492
rect 30380 8576 30432 8628
rect 30840 8576 30892 8628
rect 30748 8508 30800 8560
rect 30380 8440 30432 8492
rect 28908 8347 28960 8356
rect 28908 8313 28917 8347
rect 28917 8313 28951 8347
rect 28951 8313 28960 8347
rect 28908 8304 28960 8313
rect 22928 8279 22980 8288
rect 22928 8245 22937 8279
rect 22937 8245 22971 8279
rect 22971 8245 22980 8279
rect 22928 8236 22980 8245
rect 23204 8279 23256 8288
rect 23204 8245 23213 8279
rect 23213 8245 23247 8279
rect 23247 8245 23256 8279
rect 23204 8236 23256 8245
rect 23480 8279 23532 8288
rect 23480 8245 23489 8279
rect 23489 8245 23523 8279
rect 23523 8245 23532 8279
rect 23480 8236 23532 8245
rect 23572 8236 23624 8288
rect 24032 8279 24084 8288
rect 24032 8245 24041 8279
rect 24041 8245 24075 8279
rect 24075 8245 24084 8279
rect 24032 8236 24084 8245
rect 24584 8279 24636 8288
rect 24584 8245 24593 8279
rect 24593 8245 24627 8279
rect 24627 8245 24636 8279
rect 24584 8236 24636 8245
rect 24860 8279 24912 8288
rect 24860 8245 24869 8279
rect 24869 8245 24903 8279
rect 24903 8245 24912 8279
rect 24860 8236 24912 8245
rect 25136 8279 25188 8288
rect 25136 8245 25145 8279
rect 25145 8245 25179 8279
rect 25179 8245 25188 8279
rect 25136 8236 25188 8245
rect 25412 8279 25464 8288
rect 25412 8245 25421 8279
rect 25421 8245 25455 8279
rect 25455 8245 25464 8279
rect 25412 8236 25464 8245
rect 25504 8279 25556 8288
rect 25504 8245 25513 8279
rect 25513 8245 25547 8279
rect 25547 8245 25556 8279
rect 25504 8236 25556 8245
rect 25964 8279 26016 8288
rect 25964 8245 25973 8279
rect 25973 8245 26007 8279
rect 26007 8245 26016 8279
rect 25964 8236 26016 8245
rect 26240 8279 26292 8288
rect 26240 8245 26249 8279
rect 26249 8245 26283 8279
rect 26283 8245 26292 8279
rect 26240 8236 26292 8245
rect 26516 8279 26568 8288
rect 26516 8245 26525 8279
rect 26525 8245 26559 8279
rect 26559 8245 26568 8279
rect 26516 8236 26568 8245
rect 26792 8279 26844 8288
rect 26792 8245 26801 8279
rect 26801 8245 26835 8279
rect 26835 8245 26844 8279
rect 26792 8236 26844 8245
rect 26976 8279 27028 8288
rect 26976 8245 26985 8279
rect 26985 8245 27019 8279
rect 27019 8245 27028 8279
rect 26976 8236 27028 8245
rect 27344 8236 27396 8288
rect 27804 8236 27856 8288
rect 27988 8279 28040 8288
rect 27988 8245 27997 8279
rect 27997 8245 28031 8279
rect 28031 8245 28040 8279
rect 27988 8236 28040 8245
rect 28080 8279 28132 8288
rect 28080 8245 28089 8279
rect 28089 8245 28123 8279
rect 28123 8245 28132 8279
rect 28080 8236 28132 8245
rect 28632 8279 28684 8288
rect 28632 8245 28641 8279
rect 28641 8245 28675 8279
rect 28675 8245 28684 8279
rect 28632 8236 28684 8245
rect 28724 8236 28776 8288
rect 29184 8279 29236 8288
rect 29184 8245 29193 8279
rect 29193 8245 29227 8279
rect 29227 8245 29236 8279
rect 29184 8236 29236 8245
rect 29920 8236 29972 8288
rect 30288 8304 30340 8356
rect 31024 8440 31076 8492
rect 31484 8619 31536 8628
rect 31484 8585 31493 8619
rect 31493 8585 31527 8619
rect 31527 8585 31536 8619
rect 31484 8576 31536 8585
rect 31852 8576 31904 8628
rect 32404 8619 32456 8628
rect 32404 8585 32413 8619
rect 32413 8585 32447 8619
rect 32447 8585 32456 8619
rect 32404 8576 32456 8585
rect 32496 8576 32548 8628
rect 31760 8508 31812 8560
rect 30932 8347 30984 8356
rect 30932 8313 30941 8347
rect 30941 8313 30975 8347
rect 30975 8313 30984 8347
rect 30932 8304 30984 8313
rect 31300 8372 31352 8424
rect 32220 8508 32272 8560
rect 33508 8619 33560 8628
rect 33508 8585 33517 8619
rect 33517 8585 33551 8619
rect 33551 8585 33560 8619
rect 33508 8576 33560 8585
rect 33876 8576 33928 8628
rect 34244 8576 34296 8628
rect 35072 8576 35124 8628
rect 33232 8508 33284 8560
rect 33784 8508 33836 8560
rect 31576 8372 31628 8424
rect 32036 8372 32088 8424
rect 32772 8372 32824 8424
rect 33968 8483 34020 8492
rect 33968 8449 33977 8483
rect 33977 8449 34011 8483
rect 34011 8449 34020 8483
rect 33968 8440 34020 8449
rect 34980 8508 35032 8560
rect 37464 8576 37516 8628
rect 37556 8508 37608 8560
rect 38016 8508 38068 8560
rect 39304 8619 39356 8628
rect 39304 8585 39313 8619
rect 39313 8585 39347 8619
rect 39347 8585 39356 8619
rect 39304 8576 39356 8585
rect 39672 8576 39724 8628
rect 34796 8483 34848 8492
rect 34796 8449 34805 8483
rect 34805 8449 34839 8483
rect 34839 8449 34848 8483
rect 34796 8440 34848 8449
rect 35348 8483 35400 8492
rect 35348 8449 35357 8483
rect 35357 8449 35391 8483
rect 35391 8449 35400 8483
rect 35348 8440 35400 8449
rect 35900 8483 35952 8492
rect 35900 8449 35909 8483
rect 35909 8449 35943 8483
rect 35943 8449 35952 8483
rect 35900 8440 35952 8449
rect 36636 8440 36688 8492
rect 38384 8440 38436 8492
rect 39304 8440 39356 8492
rect 36544 8372 36596 8424
rect 33600 8304 33652 8356
rect 34428 8304 34480 8356
rect 35808 8304 35860 8356
rect 38292 8372 38344 8424
rect 38660 8347 38712 8356
rect 38660 8313 38669 8347
rect 38669 8313 38703 8347
rect 38703 8313 38712 8347
rect 38660 8304 38712 8313
rect 39580 8372 39632 8424
rect 41052 8483 41104 8492
rect 41052 8449 41061 8483
rect 41061 8449 41095 8483
rect 41095 8449 41104 8483
rect 41052 8440 41104 8449
rect 31392 8236 31444 8288
rect 31668 8236 31720 8288
rect 32128 8236 32180 8288
rect 32956 8279 33008 8288
rect 32956 8245 32965 8279
rect 32965 8245 32999 8279
rect 32999 8245 33008 8279
rect 32956 8236 33008 8245
rect 33416 8236 33468 8288
rect 6251 8134 6303 8186
rect 6315 8134 6367 8186
rect 6379 8134 6431 8186
rect 6443 8134 6495 8186
rect 6507 8134 6559 8186
rect 16854 8134 16906 8186
rect 16918 8134 16970 8186
rect 16982 8134 17034 8186
rect 17046 8134 17098 8186
rect 17110 8134 17162 8186
rect 27457 8134 27509 8186
rect 27521 8134 27573 8186
rect 27585 8134 27637 8186
rect 27649 8134 27701 8186
rect 27713 8134 27765 8186
rect 38060 8134 38112 8186
rect 38124 8134 38176 8186
rect 38188 8134 38240 8186
rect 38252 8134 38304 8186
rect 38316 8134 38368 8186
rect 6000 8075 6052 8084
rect 6000 8041 6009 8075
rect 6009 8041 6043 8075
rect 6043 8041 6052 8075
rect 6000 8032 6052 8041
rect 6552 8075 6604 8084
rect 6552 8041 6561 8075
rect 6561 8041 6595 8075
rect 6595 8041 6604 8075
rect 6552 8032 6604 8041
rect 7104 8075 7156 8084
rect 7104 8041 7113 8075
rect 7113 8041 7147 8075
rect 7147 8041 7156 8075
rect 7104 8032 7156 8041
rect 8024 8075 8076 8084
rect 8024 8041 8033 8075
rect 8033 8041 8067 8075
rect 8067 8041 8076 8075
rect 8024 8032 8076 8041
rect 8576 8075 8628 8084
rect 8576 8041 8585 8075
rect 8585 8041 8619 8075
rect 8619 8041 8628 8075
rect 8576 8032 8628 8041
rect 9312 8075 9364 8084
rect 9312 8041 9321 8075
rect 9321 8041 9355 8075
rect 9355 8041 9364 8075
rect 9312 8032 9364 8041
rect 10416 8075 10468 8084
rect 10416 8041 10425 8075
rect 10425 8041 10459 8075
rect 10459 8041 10468 8075
rect 10416 8032 10468 8041
rect 10692 8032 10744 8084
rect 11244 8075 11296 8084
rect 11244 8041 11253 8075
rect 11253 8041 11287 8075
rect 11287 8041 11296 8075
rect 11244 8032 11296 8041
rect 11796 8075 11848 8084
rect 11796 8041 11805 8075
rect 11805 8041 11839 8075
rect 11839 8041 11848 8075
rect 11796 8032 11848 8041
rect 12624 8075 12676 8084
rect 12624 8041 12633 8075
rect 12633 8041 12667 8075
rect 12667 8041 12676 8075
rect 12624 8032 12676 8041
rect 13452 8075 13504 8084
rect 13452 8041 13461 8075
rect 13461 8041 13495 8075
rect 13495 8041 13504 8075
rect 13452 8032 13504 8041
rect 14280 8075 14332 8084
rect 14280 8041 14289 8075
rect 14289 8041 14323 8075
rect 14323 8041 14332 8075
rect 14280 8032 14332 8041
rect 14832 8075 14884 8084
rect 14832 8041 14841 8075
rect 14841 8041 14875 8075
rect 14875 8041 14884 8075
rect 14832 8032 14884 8041
rect 15660 8032 15712 8084
rect 15936 8075 15988 8084
rect 15936 8041 15945 8075
rect 15945 8041 15979 8075
rect 15979 8041 15988 8075
rect 15936 8032 15988 8041
rect 16488 8075 16540 8084
rect 16488 8041 16497 8075
rect 16497 8041 16531 8075
rect 16531 8041 16540 8075
rect 16488 8032 16540 8041
rect 12808 7964 12860 8016
rect 17592 8032 17644 8084
rect 17776 8075 17828 8084
rect 17776 8041 17785 8075
rect 17785 8041 17819 8075
rect 17819 8041 17828 8075
rect 17776 8032 17828 8041
rect 17960 8032 18012 8084
rect 18420 8032 18472 8084
rect 17132 8007 17184 8016
rect 17132 7973 17141 8007
rect 17141 7973 17175 8007
rect 17175 7973 17184 8007
rect 17132 7964 17184 7973
rect 6276 7803 6328 7812
rect 6276 7769 6285 7803
rect 6285 7769 6319 7803
rect 6319 7769 6328 7803
rect 6276 7760 6328 7769
rect 6828 7803 6880 7812
rect 6828 7769 6837 7803
rect 6837 7769 6871 7803
rect 6871 7769 6880 7803
rect 6828 7760 6880 7769
rect 8116 7803 8168 7812
rect 8116 7769 8125 7803
rect 8125 7769 8159 7803
rect 8159 7769 8168 7803
rect 8116 7760 8168 7769
rect 9496 7760 9548 7812
rect 9588 7803 9640 7812
rect 9588 7769 9597 7803
rect 9597 7769 9631 7803
rect 9631 7769 9640 7803
rect 9588 7760 9640 7769
rect 10692 7871 10744 7880
rect 10692 7837 10701 7871
rect 10701 7837 10735 7871
rect 10735 7837 10744 7871
rect 10692 7828 10744 7837
rect 13636 7828 13688 7880
rect 13728 7871 13780 7880
rect 13728 7837 13737 7871
rect 13737 7837 13771 7871
rect 13771 7837 13780 7871
rect 13728 7828 13780 7837
rect 17040 7896 17092 7948
rect 11888 7760 11940 7812
rect 12808 7760 12860 7812
rect 12900 7803 12952 7812
rect 12900 7769 12909 7803
rect 12909 7769 12943 7803
rect 12943 7769 12952 7803
rect 12900 7760 12952 7769
rect 15108 7803 15160 7812
rect 15108 7769 15117 7803
rect 15117 7769 15151 7803
rect 15151 7769 15160 7803
rect 15108 7760 15160 7769
rect 16396 7828 16448 7880
rect 18512 7896 18564 7948
rect 18236 7828 18288 7880
rect 18328 7871 18380 7880
rect 18328 7837 18337 7871
rect 18337 7837 18371 7871
rect 18371 7837 18380 7871
rect 18328 7828 18380 7837
rect 18696 7871 18748 7880
rect 18696 7837 18705 7871
rect 18705 7837 18739 7871
rect 18739 7837 18748 7871
rect 18696 7828 18748 7837
rect 18788 7828 18840 7880
rect 19064 7964 19116 8016
rect 19064 7871 19116 7880
rect 19064 7837 19073 7871
rect 19073 7837 19107 7871
rect 19107 7837 19116 7871
rect 19064 7828 19116 7837
rect 19156 7828 19208 7880
rect 19340 7828 19392 7880
rect 20260 7964 20312 8016
rect 20444 7964 20496 8016
rect 20904 8007 20956 8016
rect 20904 7973 20913 8007
rect 20913 7973 20947 8007
rect 20947 7973 20956 8007
rect 20904 7964 20956 7973
rect 21088 7964 21140 8016
rect 21180 8007 21232 8016
rect 21180 7973 21189 8007
rect 21189 7973 21223 8007
rect 21223 7973 21232 8007
rect 21180 7964 21232 7973
rect 21732 8007 21784 8016
rect 21732 7973 21741 8007
rect 21741 7973 21775 8007
rect 21775 7973 21784 8007
rect 21732 7964 21784 7973
rect 24952 8032 25004 8084
rect 25872 8032 25924 8084
rect 27896 8032 27948 8084
rect 28080 8032 28132 8084
rect 29368 8032 29420 8084
rect 32956 8032 33008 8084
rect 36084 8032 36136 8084
rect 36820 8032 36872 8084
rect 37740 8032 37792 8084
rect 38844 8032 38896 8084
rect 20076 7828 20128 7880
rect 20352 7828 20404 7880
rect 20996 7828 21048 7880
rect 21180 7828 21232 7880
rect 21364 7871 21416 7880
rect 21364 7837 21373 7871
rect 21373 7837 21407 7871
rect 21407 7837 21416 7871
rect 21364 7828 21416 7837
rect 22376 7896 22428 7948
rect 22652 7896 22704 7948
rect 23388 7896 23440 7948
rect 16948 7760 17000 7812
rect 17500 7760 17552 7812
rect 18420 7760 18472 7812
rect 11980 7692 12032 7744
rect 14372 7692 14424 7744
rect 17960 7692 18012 7744
rect 20260 7692 20312 7744
rect 20352 7735 20404 7744
rect 20352 7701 20361 7735
rect 20361 7701 20395 7735
rect 20395 7701 20404 7735
rect 20352 7692 20404 7701
rect 21824 7692 21876 7744
rect 22928 7828 22980 7880
rect 23296 7871 23348 7880
rect 23296 7837 23305 7871
rect 23305 7837 23339 7871
rect 23339 7837 23348 7871
rect 23296 7828 23348 7837
rect 23480 7828 23532 7880
rect 23848 7871 23900 7880
rect 23848 7837 23857 7871
rect 23857 7837 23891 7871
rect 23891 7837 23900 7871
rect 23848 7828 23900 7837
rect 24032 7828 24084 7880
rect 24584 7871 24636 7880
rect 24584 7837 24593 7871
rect 24593 7837 24627 7871
rect 24627 7837 24636 7871
rect 24584 7828 24636 7837
rect 24768 7828 24820 7880
rect 24860 7871 24912 7880
rect 24860 7837 24869 7871
rect 24869 7837 24903 7871
rect 24903 7837 24912 7871
rect 24860 7828 24912 7837
rect 25136 7871 25188 7880
rect 25136 7837 25145 7871
rect 25145 7837 25179 7871
rect 25179 7837 25188 7871
rect 25136 7828 25188 7837
rect 25412 7871 25464 7880
rect 25412 7837 25421 7871
rect 25421 7837 25455 7871
rect 25455 7837 25464 7871
rect 25412 7828 25464 7837
rect 25780 7896 25832 7948
rect 35808 7964 35860 8016
rect 39212 7964 39264 8016
rect 25964 7871 26016 7880
rect 25964 7837 25973 7871
rect 25973 7837 26007 7871
rect 26007 7837 26016 7871
rect 25964 7828 26016 7837
rect 26240 7871 26292 7880
rect 26240 7837 26249 7871
rect 26249 7837 26283 7871
rect 26283 7837 26292 7871
rect 26240 7828 26292 7837
rect 26516 7871 26568 7880
rect 26516 7837 26525 7871
rect 26525 7837 26559 7871
rect 26559 7837 26568 7871
rect 26516 7828 26568 7837
rect 22192 7692 22244 7744
rect 22284 7735 22336 7744
rect 22284 7701 22293 7735
rect 22293 7701 22327 7735
rect 22327 7701 22336 7735
rect 22284 7692 22336 7701
rect 22560 7735 22612 7744
rect 22560 7701 22569 7735
rect 22569 7701 22603 7735
rect 22603 7701 22612 7735
rect 22560 7692 22612 7701
rect 22836 7735 22888 7744
rect 22836 7701 22845 7735
rect 22845 7701 22879 7735
rect 22879 7701 22888 7735
rect 22836 7692 22888 7701
rect 23020 7692 23072 7744
rect 23388 7735 23440 7744
rect 23388 7701 23397 7735
rect 23397 7701 23431 7735
rect 23431 7701 23440 7735
rect 23388 7692 23440 7701
rect 23664 7735 23716 7744
rect 23664 7701 23673 7735
rect 23673 7701 23707 7735
rect 23707 7701 23716 7735
rect 23664 7692 23716 7701
rect 23940 7735 23992 7744
rect 23940 7701 23949 7735
rect 23949 7701 23983 7735
rect 23983 7701 23992 7735
rect 23940 7692 23992 7701
rect 24124 7692 24176 7744
rect 24400 7735 24452 7744
rect 24400 7701 24409 7735
rect 24409 7701 24443 7735
rect 24443 7701 24452 7735
rect 24400 7692 24452 7701
rect 24676 7735 24728 7744
rect 24676 7701 24685 7735
rect 24685 7701 24719 7735
rect 24719 7701 24728 7735
rect 24676 7692 24728 7701
rect 25228 7735 25280 7744
rect 25228 7701 25237 7735
rect 25237 7701 25271 7735
rect 25271 7701 25280 7735
rect 25228 7692 25280 7701
rect 26148 7692 26200 7744
rect 26792 7871 26844 7880
rect 26792 7837 26801 7871
rect 26801 7837 26835 7871
rect 26835 7837 26844 7871
rect 26792 7828 26844 7837
rect 32680 7896 32732 7948
rect 27344 7871 27396 7880
rect 27344 7837 27353 7871
rect 27353 7837 27387 7871
rect 27387 7837 27396 7871
rect 27344 7828 27396 7837
rect 27804 7828 27856 7880
rect 27988 7828 28040 7880
rect 33324 7828 33376 7880
rect 28080 7760 28132 7812
rect 35716 7803 35768 7812
rect 35716 7769 35725 7803
rect 35725 7769 35759 7803
rect 35759 7769 35768 7803
rect 35716 7760 35768 7769
rect 36268 7803 36320 7812
rect 36268 7769 36277 7803
rect 36277 7769 36311 7803
rect 36311 7769 36320 7803
rect 36268 7760 36320 7769
rect 36820 7803 36872 7812
rect 36820 7769 36829 7803
rect 36829 7769 36863 7803
rect 36863 7769 36872 7803
rect 36820 7760 36872 7769
rect 39856 7828 39908 7880
rect 37924 7803 37976 7812
rect 37924 7769 37933 7803
rect 37933 7769 37967 7803
rect 37967 7769 37976 7803
rect 37924 7760 37976 7769
rect 38384 7760 38436 7812
rect 39948 7803 40000 7812
rect 39948 7769 39957 7803
rect 39957 7769 39991 7803
rect 39991 7769 40000 7803
rect 39948 7760 40000 7769
rect 26884 7735 26936 7744
rect 26884 7701 26893 7735
rect 26893 7701 26927 7735
rect 26927 7701 26936 7735
rect 26884 7692 26936 7701
rect 27160 7735 27212 7744
rect 27160 7701 27169 7735
rect 27169 7701 27203 7735
rect 27203 7701 27212 7735
rect 27160 7692 27212 7701
rect 27436 7735 27488 7744
rect 27436 7701 27445 7735
rect 27445 7701 27479 7735
rect 27479 7701 27488 7735
rect 27436 7692 27488 7701
rect 28172 7692 28224 7744
rect 33416 7735 33468 7744
rect 33416 7701 33425 7735
rect 33425 7701 33459 7735
rect 33459 7701 33468 7735
rect 33416 7692 33468 7701
rect 35256 7692 35308 7744
rect 38752 7735 38804 7744
rect 38752 7701 38761 7735
rect 38761 7701 38795 7735
rect 38795 7701 38804 7735
rect 38752 7692 38804 7701
rect 39120 7735 39172 7744
rect 39120 7701 39129 7735
rect 39129 7701 39163 7735
rect 39163 7701 39172 7735
rect 39120 7692 39172 7701
rect 11552 7590 11604 7642
rect 11616 7590 11668 7642
rect 11680 7590 11732 7642
rect 11744 7590 11796 7642
rect 11808 7590 11860 7642
rect 22155 7590 22207 7642
rect 22219 7590 22271 7642
rect 22283 7590 22335 7642
rect 22347 7590 22399 7642
rect 22411 7590 22463 7642
rect 32758 7590 32810 7642
rect 32822 7590 32874 7642
rect 32886 7590 32938 7642
rect 32950 7590 33002 7642
rect 33014 7590 33066 7642
rect 43361 7590 43413 7642
rect 43425 7590 43477 7642
rect 43489 7590 43541 7642
rect 43553 7590 43605 7642
rect 43617 7590 43669 7642
rect 6276 7488 6328 7540
rect 14372 7488 14424 7540
rect 14556 7488 14608 7540
rect 17224 7488 17276 7540
rect 18052 7488 18104 7540
rect 18696 7488 18748 7540
rect 19064 7488 19116 7540
rect 19248 7531 19300 7540
rect 19248 7497 19257 7531
rect 19257 7497 19291 7531
rect 19291 7497 19300 7531
rect 19248 7488 19300 7497
rect 19800 7488 19852 7540
rect 7288 7395 7340 7404
rect 7288 7361 7297 7395
rect 7297 7361 7331 7395
rect 7331 7361 7340 7395
rect 7288 7352 7340 7361
rect 7380 7216 7432 7268
rect 9036 7420 9088 7472
rect 9496 7420 9548 7472
rect 16672 7420 16724 7472
rect 17776 7420 17828 7472
rect 20812 7488 20864 7540
rect 20076 7420 20128 7472
rect 9588 7352 9640 7404
rect 14648 7395 14700 7404
rect 14648 7361 14657 7395
rect 14657 7361 14691 7395
rect 14691 7361 14700 7395
rect 14648 7352 14700 7361
rect 15108 7352 15160 7404
rect 17500 7352 17552 7404
rect 17868 7395 17920 7404
rect 17868 7361 17877 7395
rect 17877 7361 17911 7395
rect 17911 7361 17920 7395
rect 17868 7352 17920 7361
rect 18144 7395 18196 7404
rect 18144 7361 18153 7395
rect 18153 7361 18187 7395
rect 18187 7361 18196 7395
rect 18144 7352 18196 7361
rect 18604 7352 18656 7404
rect 18972 7395 19024 7404
rect 18972 7361 18981 7395
rect 18981 7361 19015 7395
rect 19015 7361 19024 7395
rect 18972 7352 19024 7361
rect 19064 7395 19116 7404
rect 19064 7361 19073 7395
rect 19073 7361 19107 7395
rect 19107 7361 19116 7395
rect 19064 7352 19116 7361
rect 19708 7352 19760 7404
rect 19800 7395 19852 7404
rect 19800 7361 19809 7395
rect 19809 7361 19843 7395
rect 19843 7361 19852 7395
rect 19800 7352 19852 7361
rect 19984 7352 20036 7404
rect 16764 7284 16816 7336
rect 18052 7284 18104 7336
rect 21548 7488 21600 7540
rect 21180 7420 21232 7472
rect 21272 7352 21324 7404
rect 22008 7488 22060 7540
rect 22652 7488 22704 7540
rect 23204 7488 23256 7540
rect 23296 7488 23348 7540
rect 29184 7488 29236 7540
rect 33416 7488 33468 7540
rect 23112 7420 23164 7472
rect 25504 7420 25556 7472
rect 26976 7420 27028 7472
rect 17868 7216 17920 7268
rect 19340 7216 19392 7268
rect 19432 7216 19484 7268
rect 14464 7148 14516 7200
rect 17408 7191 17460 7200
rect 17408 7157 17417 7191
rect 17417 7157 17451 7191
rect 17451 7157 17460 7191
rect 17408 7148 17460 7157
rect 21180 7259 21232 7268
rect 21180 7225 21189 7259
rect 21189 7225 21223 7259
rect 21223 7225 21232 7259
rect 21180 7216 21232 7225
rect 23848 7216 23900 7268
rect 28632 7216 28684 7268
rect 20628 7191 20680 7200
rect 20628 7157 20637 7191
rect 20637 7157 20671 7191
rect 20671 7157 20680 7191
rect 20628 7148 20680 7157
rect 20720 7148 20772 7200
rect 21456 7148 21508 7200
rect 24768 7191 24820 7200
rect 24768 7157 24777 7191
rect 24777 7157 24811 7191
rect 24811 7157 24820 7191
rect 24768 7148 24820 7157
rect 26056 7148 26108 7200
rect 6251 7046 6303 7098
rect 6315 7046 6367 7098
rect 6379 7046 6431 7098
rect 6443 7046 6495 7098
rect 6507 7046 6559 7098
rect 16854 7046 16906 7098
rect 16918 7046 16970 7098
rect 16982 7046 17034 7098
rect 17046 7046 17098 7098
rect 17110 7046 17162 7098
rect 27457 7046 27509 7098
rect 27521 7046 27573 7098
rect 27585 7046 27637 7098
rect 27649 7046 27701 7098
rect 27713 7046 27765 7098
rect 38060 7046 38112 7098
rect 38124 7046 38176 7098
rect 38188 7046 38240 7098
rect 38252 7046 38304 7098
rect 38316 7046 38368 7098
rect 7288 6944 7340 6996
rect 12348 6944 12400 6996
rect 14648 6944 14700 6996
rect 24768 6944 24820 6996
rect 25228 6944 25280 6996
rect 8116 6876 8168 6928
rect 9220 6808 9272 6860
rect 10140 6808 10192 6860
rect 10692 6808 10744 6860
rect 17500 6876 17552 6928
rect 21824 6808 21876 6860
rect 38568 6808 38620 6860
rect 39120 6808 39172 6860
rect 17960 6740 18012 6792
rect 18052 6740 18104 6792
rect 18236 6740 18288 6792
rect 18328 6740 18380 6792
rect 19616 6740 19668 6792
rect 19892 6740 19944 6792
rect 14464 6672 14516 6724
rect 20076 6783 20128 6792
rect 20076 6749 20085 6783
rect 20085 6749 20119 6783
rect 20119 6749 20128 6783
rect 20076 6740 20128 6749
rect 36912 6740 36964 6792
rect 38660 6740 38712 6792
rect 28724 6672 28776 6724
rect 37188 6672 37240 6724
rect 38752 6672 38804 6724
rect 11552 6502 11604 6554
rect 11616 6502 11668 6554
rect 11680 6502 11732 6554
rect 11744 6502 11796 6554
rect 11808 6502 11860 6554
rect 22155 6502 22207 6554
rect 22219 6502 22271 6554
rect 22283 6502 22335 6554
rect 22347 6502 22399 6554
rect 22411 6502 22463 6554
rect 32758 6502 32810 6554
rect 32822 6502 32874 6554
rect 32886 6502 32938 6554
rect 32950 6502 33002 6554
rect 33014 6502 33066 6554
rect 43361 6502 43413 6554
rect 43425 6502 43477 6554
rect 43489 6502 43541 6554
rect 43553 6502 43605 6554
rect 43617 6502 43669 6554
rect 15200 6400 15252 6452
rect 20260 6400 20312 6452
rect 16120 6332 16172 6384
rect 20352 6332 20404 6384
rect 16580 6264 16632 6316
rect 20628 6264 20680 6316
rect 6251 5958 6303 6010
rect 6315 5958 6367 6010
rect 6379 5958 6431 6010
rect 6443 5958 6495 6010
rect 6507 5958 6559 6010
rect 16854 5958 16906 6010
rect 16918 5958 16970 6010
rect 16982 5958 17034 6010
rect 17046 5958 17098 6010
rect 17110 5958 17162 6010
rect 27457 5958 27509 6010
rect 27521 5958 27573 6010
rect 27585 5958 27637 6010
rect 27649 5958 27701 6010
rect 27713 5958 27765 6010
rect 38060 5958 38112 6010
rect 38124 5958 38176 6010
rect 38188 5958 38240 6010
rect 38252 5958 38304 6010
rect 38316 5958 38368 6010
rect 25964 5652 26016 5704
rect 30472 5652 30524 5704
rect 23020 5584 23072 5636
rect 35348 5584 35400 5636
rect 11552 5414 11604 5466
rect 11616 5414 11668 5466
rect 11680 5414 11732 5466
rect 11744 5414 11796 5466
rect 11808 5414 11860 5466
rect 22155 5414 22207 5466
rect 22219 5414 22271 5466
rect 22283 5414 22335 5466
rect 22347 5414 22399 5466
rect 22411 5414 22463 5466
rect 32758 5414 32810 5466
rect 32822 5414 32874 5466
rect 32886 5414 32938 5466
rect 32950 5414 33002 5466
rect 33014 5414 33066 5466
rect 43361 5414 43413 5466
rect 43425 5414 43477 5466
rect 43489 5414 43541 5466
rect 43553 5414 43605 5466
rect 43617 5414 43669 5466
rect 39304 5312 39356 5364
rect 37372 5219 37424 5228
rect 37372 5185 37381 5219
rect 37381 5185 37415 5219
rect 37415 5185 37424 5219
rect 37372 5176 37424 5185
rect 23848 5108 23900 5160
rect 32680 5108 32732 5160
rect 6251 4870 6303 4922
rect 6315 4870 6367 4922
rect 6379 4870 6431 4922
rect 6443 4870 6495 4922
rect 6507 4870 6559 4922
rect 16854 4870 16906 4922
rect 16918 4870 16970 4922
rect 16982 4870 17034 4922
rect 17046 4870 17098 4922
rect 17110 4870 17162 4922
rect 27457 4870 27509 4922
rect 27521 4870 27573 4922
rect 27585 4870 27637 4922
rect 27649 4870 27701 4922
rect 27713 4870 27765 4922
rect 38060 4870 38112 4922
rect 38124 4870 38176 4922
rect 38188 4870 38240 4922
rect 38252 4870 38304 4922
rect 38316 4870 38368 4922
rect 23020 4811 23072 4820
rect 23020 4777 23029 4811
rect 23029 4777 23063 4811
rect 23063 4777 23072 4811
rect 23020 4768 23072 4777
rect 23848 4811 23900 4820
rect 23848 4777 23857 4811
rect 23857 4777 23891 4811
rect 23891 4777 23900 4811
rect 23848 4768 23900 4777
rect 25964 4811 26016 4820
rect 25964 4777 25973 4811
rect 25973 4777 26007 4811
rect 26007 4777 26016 4811
rect 25964 4768 26016 4777
rect 28080 4811 28132 4820
rect 28080 4777 28089 4811
rect 28089 4777 28123 4811
rect 28123 4777 28132 4811
rect 28080 4768 28132 4777
rect 36820 4768 36872 4820
rect 37372 4768 37424 4820
rect 38384 4768 38436 4820
rect 37924 4700 37976 4752
rect 31116 4632 31168 4684
rect 21548 4607 21600 4616
rect 21548 4573 21557 4607
rect 21557 4573 21591 4607
rect 21591 4573 21600 4607
rect 21548 4564 21600 4573
rect 22560 4607 22612 4616
rect 22560 4573 22569 4607
rect 22569 4573 22603 4607
rect 22603 4573 22612 4607
rect 22560 4564 22612 4573
rect 22836 4607 22888 4616
rect 22836 4573 22845 4607
rect 22845 4573 22879 4607
rect 22879 4573 22888 4607
rect 22836 4564 22888 4573
rect 22652 4496 22704 4548
rect 23664 4607 23716 4616
rect 23664 4573 23673 4607
rect 23673 4573 23707 4607
rect 23707 4573 23716 4607
rect 23664 4564 23716 4573
rect 25780 4607 25832 4616
rect 25780 4573 25789 4607
rect 25789 4573 25823 4607
rect 25823 4573 25832 4607
rect 25780 4564 25832 4573
rect 27896 4607 27948 4616
rect 27896 4573 27905 4607
rect 27905 4573 27939 4607
rect 27939 4573 27948 4607
rect 27896 4564 27948 4573
rect 32128 4607 32180 4616
rect 32128 4573 32137 4607
rect 32137 4573 32171 4607
rect 32171 4573 32180 4607
rect 32128 4564 32180 4573
rect 34520 4564 34572 4616
rect 38016 4607 38068 4616
rect 38016 4573 38025 4607
rect 38025 4573 38059 4607
rect 38059 4573 38068 4607
rect 38016 4564 38068 4573
rect 29276 4428 29328 4480
rect 11552 4326 11604 4378
rect 11616 4326 11668 4378
rect 11680 4326 11732 4378
rect 11744 4326 11796 4378
rect 11808 4326 11860 4378
rect 22155 4326 22207 4378
rect 22219 4326 22271 4378
rect 22283 4326 22335 4378
rect 22347 4326 22399 4378
rect 22411 4326 22463 4378
rect 32758 4326 32810 4378
rect 32822 4326 32874 4378
rect 32886 4326 32938 4378
rect 32950 4326 33002 4378
rect 33014 4326 33066 4378
rect 43361 4326 43413 4378
rect 43425 4326 43477 4378
rect 43489 4326 43541 4378
rect 43553 4326 43605 4378
rect 43617 4326 43669 4378
rect 21548 4224 21600 4276
rect 22560 4224 22612 4276
rect 25780 4224 25832 4276
rect 38016 4224 38068 4276
rect 20444 4088 20496 4140
rect 7748 4020 7800 4072
rect 5632 3952 5684 4004
rect 22468 4088 22520 4140
rect 24768 4088 24820 4140
rect 27068 4131 27120 4140
rect 27068 4097 27077 4131
rect 27077 4097 27111 4131
rect 27111 4097 27120 4131
rect 27068 4088 27120 4097
rect 31300 4131 31352 4140
rect 31300 4097 31309 4131
rect 31309 4097 31343 4131
rect 31343 4097 31352 4131
rect 31300 4088 31352 4097
rect 37464 4131 37516 4140
rect 37464 4097 37473 4131
rect 37473 4097 37507 4131
rect 37507 4097 37516 4131
rect 37464 4088 37516 4097
rect 39764 4131 39816 4140
rect 39764 4097 39773 4131
rect 39773 4097 39807 4131
rect 39807 4097 39816 4131
rect 39764 4088 39816 4097
rect 22836 4020 22888 4072
rect 27896 4020 27948 4072
rect 32128 4020 32180 4072
rect 19524 3884 19576 3936
rect 22652 3884 22704 3936
rect 31392 3884 31444 3936
rect 39856 3884 39908 3936
rect 6251 3782 6303 3834
rect 6315 3782 6367 3834
rect 6379 3782 6431 3834
rect 6443 3782 6495 3834
rect 6507 3782 6559 3834
rect 16854 3782 16906 3834
rect 16918 3782 16970 3834
rect 16982 3782 17034 3834
rect 17046 3782 17098 3834
rect 17110 3782 17162 3834
rect 27457 3782 27509 3834
rect 27521 3782 27573 3834
rect 27585 3782 27637 3834
rect 27649 3782 27701 3834
rect 27713 3782 27765 3834
rect 38060 3782 38112 3834
rect 38124 3782 38176 3834
rect 38188 3782 38240 3834
rect 38252 3782 38304 3834
rect 38316 3782 38368 3834
rect 22468 3680 22520 3732
rect 23664 3680 23716 3732
rect 34612 3680 34664 3732
rect 39580 3680 39632 3732
rect 39764 3680 39816 3732
rect 36268 3612 36320 3664
rect 19432 3519 19484 3528
rect 19432 3485 19441 3519
rect 19441 3485 19475 3519
rect 19475 3485 19484 3519
rect 19432 3476 19484 3485
rect 19248 3408 19300 3460
rect 22008 3476 22060 3528
rect 21272 3408 21324 3460
rect 22836 3519 22888 3528
rect 22836 3485 22845 3519
rect 22845 3485 22879 3519
rect 22879 3485 22888 3519
rect 22836 3476 22888 3485
rect 30012 3519 30064 3528
rect 30012 3485 30021 3519
rect 30021 3485 30055 3519
rect 30055 3485 30064 3519
rect 30012 3476 30064 3485
rect 35716 3476 35768 3528
rect 37096 3519 37148 3528
rect 37096 3485 37105 3519
rect 37105 3485 37139 3519
rect 37139 3485 37148 3519
rect 37096 3476 37148 3485
rect 40684 3519 40736 3528
rect 40684 3485 40693 3519
rect 40693 3485 40727 3519
rect 40727 3485 40736 3519
rect 40684 3476 40736 3485
rect 36636 3340 36688 3392
rect 11552 3238 11604 3290
rect 11616 3238 11668 3290
rect 11680 3238 11732 3290
rect 11744 3238 11796 3290
rect 11808 3238 11860 3290
rect 22155 3238 22207 3290
rect 22219 3238 22271 3290
rect 22283 3238 22335 3290
rect 22347 3238 22399 3290
rect 22411 3238 22463 3290
rect 32758 3238 32810 3290
rect 32822 3238 32874 3290
rect 32886 3238 32938 3290
rect 32950 3238 33002 3290
rect 33014 3238 33066 3290
rect 43361 3238 43413 3290
rect 43425 3238 43477 3290
rect 43489 3238 43541 3290
rect 43553 3238 43605 3290
rect 43617 3238 43669 3290
rect 19432 3136 19484 3188
rect 21272 3179 21324 3188
rect 21272 3145 21281 3179
rect 21281 3145 21315 3179
rect 21315 3145 21324 3179
rect 21272 3136 21324 3145
rect 22008 3136 22060 3188
rect 30012 3136 30064 3188
rect 37096 3136 37148 3188
rect 41052 3136 41104 3188
rect 18604 3043 18656 3052
rect 18604 3009 18613 3043
rect 18613 3009 18647 3043
rect 18647 3009 18656 3043
rect 18604 3000 18656 3009
rect 16212 2932 16264 2984
rect 21364 3043 21416 3052
rect 21364 3009 21373 3043
rect 21373 3009 21407 3043
rect 21407 3009 21416 3043
rect 21364 3000 21416 3009
rect 22652 3043 22704 3052
rect 22652 3009 22661 3043
rect 22661 3009 22695 3043
rect 22695 3009 22704 3043
rect 22652 3000 22704 3009
rect 28908 3000 28960 3052
rect 35256 3000 35308 3052
rect 40224 3000 40276 3052
rect 23388 2864 23440 2916
rect 6251 2694 6303 2746
rect 6315 2694 6367 2746
rect 6379 2694 6431 2746
rect 6443 2694 6495 2746
rect 6507 2694 6559 2746
rect 16854 2694 16906 2746
rect 16918 2694 16970 2746
rect 16982 2694 17034 2746
rect 17046 2694 17098 2746
rect 17110 2694 17162 2746
rect 27457 2694 27509 2746
rect 27521 2694 27573 2746
rect 27585 2694 27637 2746
rect 27649 2694 27701 2746
rect 27713 2694 27765 2746
rect 38060 2694 38112 2746
rect 38124 2694 38176 2746
rect 38188 2694 38240 2746
rect 38252 2694 38304 2746
rect 38316 2694 38368 2746
rect 22652 2592 22704 2644
rect 39948 2592 40000 2644
rect 40224 2635 40276 2644
rect 40224 2601 40233 2635
rect 40233 2601 40267 2635
rect 40267 2601 40276 2635
rect 40224 2592 40276 2601
rect 3516 2388 3568 2440
rect 39028 2431 39080 2440
rect 39028 2397 39037 2431
rect 39037 2397 39071 2431
rect 39071 2397 39080 2431
rect 39028 2388 39080 2397
rect 42984 2388 43036 2440
rect 11552 2150 11604 2202
rect 11616 2150 11668 2202
rect 11680 2150 11732 2202
rect 11744 2150 11796 2202
rect 11808 2150 11860 2202
rect 22155 2150 22207 2202
rect 22219 2150 22271 2202
rect 22283 2150 22335 2202
rect 22347 2150 22399 2202
rect 22411 2150 22463 2202
rect 32758 2150 32810 2202
rect 32822 2150 32874 2202
rect 32886 2150 32938 2202
rect 32950 2150 33002 2202
rect 33014 2150 33066 2202
rect 43361 2150 43413 2202
rect 43425 2150 43477 2202
rect 43489 2150 43541 2202
rect 43553 2150 43605 2202
rect 43617 2150 43669 2202
rect 39028 2091 39080 2100
rect 39028 2057 39037 2091
rect 39037 2057 39071 2091
rect 39071 2057 39080 2091
rect 39028 2048 39080 2057
rect 1584 1912 1636 1964
rect 38844 1955 38896 1964
rect 38844 1921 38853 1955
rect 38853 1921 38887 1955
rect 38887 1921 38896 1955
rect 38844 1912 38896 1921
rect 33968 1708 34020 1760
rect 6251 1606 6303 1658
rect 6315 1606 6367 1658
rect 6379 1606 6431 1658
rect 6443 1606 6495 1658
rect 6507 1606 6559 1658
rect 16854 1606 16906 1658
rect 16918 1606 16970 1658
rect 16982 1606 17034 1658
rect 17046 1606 17098 1658
rect 17110 1606 17162 1658
rect 27457 1606 27509 1658
rect 27521 1606 27573 1658
rect 27585 1606 27637 1658
rect 27649 1606 27701 1658
rect 27713 1606 27765 1658
rect 38060 1606 38112 1658
rect 38124 1606 38176 1658
rect 38188 1606 38240 1658
rect 38252 1606 38304 1658
rect 38316 1606 38368 1658
rect 1584 1547 1636 1556
rect 1584 1513 1593 1547
rect 1593 1513 1627 1547
rect 1627 1513 1636 1547
rect 1584 1504 1636 1513
rect 3516 1547 3568 1556
rect 3516 1513 3525 1547
rect 3525 1513 3559 1547
rect 3559 1513 3568 1547
rect 3516 1504 3568 1513
rect 38844 1504 38896 1556
rect 42984 1547 43036 1556
rect 42984 1513 42993 1547
rect 42993 1513 43027 1547
rect 43027 1513 43036 1547
rect 42984 1504 43036 1513
rect 1124 1300 1176 1352
rect 3332 1343 3384 1352
rect 3332 1309 3341 1343
rect 3341 1309 3375 1343
rect 3375 1309 3384 1343
rect 3332 1300 3384 1309
rect 5448 1343 5500 1352
rect 5448 1309 5457 1343
rect 5457 1309 5491 1343
rect 5491 1309 5500 1343
rect 5448 1300 5500 1309
rect 5632 1300 5684 1352
rect 7564 1343 7616 1352
rect 7564 1309 7573 1343
rect 7573 1309 7607 1343
rect 7607 1309 7616 1343
rect 7564 1300 7616 1309
rect 9680 1343 9732 1352
rect 9680 1309 9689 1343
rect 9689 1309 9723 1343
rect 9723 1309 9732 1343
rect 9680 1300 9732 1309
rect 11796 1343 11848 1352
rect 11796 1309 11805 1343
rect 11805 1309 11839 1343
rect 11839 1309 11848 1343
rect 11796 1300 11848 1309
rect 14096 1343 14148 1352
rect 14096 1309 14105 1343
rect 14105 1309 14139 1343
rect 14139 1309 14148 1343
rect 14096 1300 14148 1309
rect 16028 1343 16080 1352
rect 16028 1309 16037 1343
rect 16037 1309 16071 1343
rect 16071 1309 16080 1343
rect 16028 1300 16080 1309
rect 18144 1343 18196 1352
rect 18144 1309 18153 1343
rect 18153 1309 18187 1343
rect 18187 1309 18196 1343
rect 18144 1300 18196 1309
rect 18420 1300 18472 1352
rect 19524 1300 19576 1352
rect 20260 1343 20312 1352
rect 20260 1309 20269 1343
rect 20269 1309 20303 1343
rect 20303 1309 20312 1343
rect 20260 1300 20312 1309
rect 21364 1300 21416 1352
rect 22376 1343 22428 1352
rect 22376 1309 22385 1343
rect 22385 1309 22419 1343
rect 22419 1309 22428 1343
rect 22376 1300 22428 1309
rect 22744 1300 22796 1352
rect 24492 1343 24544 1352
rect 24492 1309 24501 1343
rect 24501 1309 24535 1343
rect 24535 1309 24544 1343
rect 24492 1300 24544 1309
rect 26608 1343 26660 1352
rect 26608 1309 26617 1343
rect 26617 1309 26651 1343
rect 26651 1309 26660 1343
rect 26608 1300 26660 1309
rect 27068 1300 27120 1352
rect 28724 1343 28776 1352
rect 28724 1309 28733 1343
rect 28733 1309 28767 1343
rect 28767 1309 28776 1343
rect 28724 1300 28776 1309
rect 28908 1300 28960 1352
rect 30840 1343 30892 1352
rect 30840 1309 30849 1343
rect 30849 1309 30883 1343
rect 30883 1309 30892 1343
rect 30840 1300 30892 1309
rect 31300 1300 31352 1352
rect 32680 1300 32732 1352
rect 34520 1300 34572 1352
rect 35072 1343 35124 1352
rect 35072 1309 35081 1343
rect 35081 1309 35115 1343
rect 35115 1309 35124 1343
rect 35072 1300 35124 1309
rect 35256 1300 35308 1352
rect 37280 1343 37332 1352
rect 37280 1309 37289 1343
rect 37289 1309 37323 1343
rect 37323 1309 37332 1343
rect 37280 1300 37332 1309
rect 37464 1300 37516 1352
rect 39488 1343 39540 1352
rect 39488 1309 39497 1343
rect 39497 1309 39531 1343
rect 39531 1309 39540 1343
rect 39488 1300 39540 1309
rect 40684 1300 40736 1352
rect 41328 1300 41380 1352
rect 43168 1343 43220 1352
rect 43168 1309 43177 1343
rect 43177 1309 43211 1343
rect 43211 1309 43220 1343
rect 43168 1300 43220 1309
rect 7748 1207 7800 1216
rect 7748 1173 7757 1207
rect 7757 1173 7791 1207
rect 7791 1173 7800 1207
rect 7748 1164 7800 1173
rect 9864 1207 9916 1216
rect 9864 1173 9873 1207
rect 9873 1173 9907 1207
rect 9907 1173 9916 1207
rect 9864 1164 9916 1173
rect 16212 1207 16264 1216
rect 16212 1173 16221 1207
rect 16221 1173 16255 1207
rect 16255 1173 16264 1207
rect 16212 1164 16264 1173
rect 18236 1164 18288 1216
rect 18604 1164 18656 1216
rect 20444 1207 20496 1216
rect 20444 1173 20453 1207
rect 20453 1173 20487 1207
rect 20487 1173 20496 1207
rect 20444 1164 20496 1173
rect 24768 1232 24820 1284
rect 11552 1062 11604 1114
rect 11616 1062 11668 1114
rect 11680 1062 11732 1114
rect 11744 1062 11796 1114
rect 11808 1062 11860 1114
rect 22155 1062 22207 1114
rect 22219 1062 22271 1114
rect 22283 1062 22335 1114
rect 22347 1062 22399 1114
rect 22411 1062 22463 1114
rect 32758 1062 32810 1114
rect 32822 1062 32874 1114
rect 32886 1062 32938 1114
rect 32950 1062 33002 1114
rect 33014 1062 33066 1114
rect 43361 1062 43413 1114
rect 43425 1062 43477 1114
rect 43489 1062 43541 1114
rect 43553 1062 43605 1114
rect 43617 1062 43669 1114
rect 9864 960 9916 1012
rect 19248 960 19300 1012
<< metal2 >>
rect 5170 9840 5226 10300
rect 5446 9840 5502 10300
rect 5722 9840 5778 10300
rect 5998 9840 6054 10300
rect 6274 9840 6330 10300
rect 6550 9840 6606 10300
rect 6826 9840 6882 10300
rect 7102 9840 7158 10300
rect 7378 9840 7434 10300
rect 7654 9840 7710 10300
rect 7930 9840 7986 10300
rect 8206 9840 8262 10300
rect 8482 9840 8538 10300
rect 8758 9840 8814 10300
rect 9034 9840 9090 10300
rect 9310 9840 9366 10300
rect 9586 9840 9642 10300
rect 9862 9840 9918 10300
rect 10138 9840 10194 10300
rect 10414 9840 10470 10300
rect 10690 9840 10746 10300
rect 10966 9840 11022 10300
rect 11152 9988 11204 9994
rect 11152 9930 11204 9936
rect 4712 9240 4764 9246
rect 4712 9182 4764 9188
rect 4724 8498 4752 9182
rect 4712 8492 4764 8498
rect 4712 8434 4764 8440
rect 5184 8362 5212 9840
rect 5460 8634 5488 9840
rect 5540 9512 5592 9518
rect 5540 9454 5592 9460
rect 5552 8634 5580 9454
rect 5736 8634 5764 9840
rect 5448 8628 5500 8634
rect 5448 8570 5500 8576
rect 5540 8628 5592 8634
rect 5540 8570 5592 8576
rect 5724 8628 5776 8634
rect 5724 8570 5776 8576
rect 5172 8356 5224 8362
rect 5172 8298 5224 8304
rect 6012 8090 6040 9840
rect 6184 8832 6236 8838
rect 6184 8774 6236 8780
rect 6196 8498 6224 8774
rect 6288 8634 6316 9840
rect 6564 8820 6592 9840
rect 6564 8792 6684 8820
rect 6276 8628 6328 8634
rect 6276 8570 6328 8576
rect 6184 8492 6236 8498
rect 6184 8434 6236 8440
rect 6251 8188 6559 8197
rect 6251 8186 6257 8188
rect 6313 8186 6337 8188
rect 6393 8186 6417 8188
rect 6473 8186 6497 8188
rect 6553 8186 6559 8188
rect 6313 8134 6315 8186
rect 6495 8134 6497 8186
rect 6251 8132 6257 8134
rect 6313 8132 6337 8134
rect 6393 8132 6417 8134
rect 6473 8132 6497 8134
rect 6553 8132 6559 8134
rect 6251 8123 6559 8132
rect 6000 8084 6052 8090
rect 6000 8026 6052 8032
rect 6552 8084 6604 8090
rect 6656 8072 6684 8792
rect 6840 8634 6868 9840
rect 6828 8628 6880 8634
rect 6828 8570 6880 8576
rect 7116 8090 7144 9840
rect 7288 9444 7340 9450
rect 7288 9386 7340 9392
rect 7300 8634 7328 9386
rect 7288 8628 7340 8634
rect 7288 8570 7340 8576
rect 7196 8492 7248 8498
rect 7196 8434 7248 8440
rect 6604 8044 6684 8072
rect 7104 8084 7156 8090
rect 6552 8026 6604 8032
rect 7104 8026 7156 8032
rect 6276 7812 6328 7818
rect 6276 7754 6328 7760
rect 6828 7812 6880 7818
rect 6828 7754 6880 7760
rect 6288 7546 6316 7754
rect 6276 7540 6328 7546
rect 6276 7482 6328 7488
rect 6251 7100 6559 7109
rect 6251 7098 6257 7100
rect 6313 7098 6337 7100
rect 6393 7098 6417 7100
rect 6473 7098 6497 7100
rect 6553 7098 6559 7100
rect 6313 7046 6315 7098
rect 6495 7046 6497 7098
rect 6251 7044 6257 7046
rect 6313 7044 6337 7046
rect 6393 7044 6417 7046
rect 6473 7044 6497 7046
rect 6553 7044 6559 7046
rect 6251 7035 6559 7044
rect 6840 6361 6868 7754
rect 6826 6352 6882 6361
rect 6826 6287 6882 6296
rect 7208 6225 7236 8434
rect 7288 7404 7340 7410
rect 7288 7346 7340 7352
rect 7300 7002 7328 7346
rect 7392 7274 7420 9840
rect 7668 8362 7696 9840
rect 7944 8634 7972 9840
rect 7932 8628 7984 8634
rect 7932 8570 7984 8576
rect 7656 8356 7708 8362
rect 7656 8298 7708 8304
rect 8024 8084 8076 8090
rect 8220 8072 8248 9840
rect 8392 9036 8444 9042
rect 8392 8978 8444 8984
rect 8404 8566 8432 8978
rect 8496 8634 8524 9840
rect 8576 9648 8628 9654
rect 8576 9590 8628 9596
rect 8484 8628 8536 8634
rect 8484 8570 8536 8576
rect 8392 8560 8444 8566
rect 8392 8502 8444 8508
rect 8588 8498 8616 9590
rect 8668 8900 8720 8906
rect 8668 8842 8720 8848
rect 8680 8498 8708 8842
rect 8576 8492 8628 8498
rect 8576 8434 8628 8440
rect 8668 8492 8720 8498
rect 8668 8434 8720 8440
rect 8076 8044 8248 8072
rect 8576 8084 8628 8090
rect 8024 8026 8076 8032
rect 8772 8072 8800 9840
rect 8628 8044 8800 8072
rect 8576 8026 8628 8032
rect 8116 7812 8168 7818
rect 8116 7754 8168 7760
rect 7380 7268 7432 7274
rect 7380 7210 7432 7216
rect 7288 6996 7340 7002
rect 7288 6938 7340 6944
rect 8128 6934 8156 7754
rect 9048 7478 9076 9840
rect 9128 8356 9180 8362
rect 9180 8316 9260 8344
rect 9128 8298 9180 8304
rect 9036 7472 9088 7478
rect 9036 7414 9088 7420
rect 8116 6928 8168 6934
rect 8116 6870 8168 6876
rect 9232 6866 9260 8316
rect 9324 8090 9352 9840
rect 9600 8566 9628 9840
rect 9680 8832 9732 8838
rect 9680 8774 9732 8780
rect 9588 8560 9640 8566
rect 9588 8502 9640 8508
rect 9692 8498 9720 8774
rect 9876 8634 9904 9840
rect 9864 8628 9916 8634
rect 9864 8570 9916 8576
rect 9680 8492 9732 8498
rect 9680 8434 9732 8440
rect 9312 8084 9364 8090
rect 9312 8026 9364 8032
rect 9496 7812 9548 7818
rect 9496 7754 9548 7760
rect 9588 7812 9640 7818
rect 9588 7754 9640 7760
rect 9508 7478 9536 7754
rect 9496 7472 9548 7478
rect 9496 7414 9548 7420
rect 9600 7410 9628 7754
rect 9588 7404 9640 7410
rect 9588 7346 9640 7352
rect 10152 6866 10180 9840
rect 10428 8090 10456 9840
rect 10704 8090 10732 9840
rect 10784 9648 10836 9654
rect 10784 9590 10836 9596
rect 10796 8498 10824 9590
rect 10980 8634 11008 9840
rect 10968 8628 11020 8634
rect 10968 8570 11020 8576
rect 11164 8498 11192 9930
rect 11242 9840 11298 10300
rect 11518 9840 11574 10300
rect 11794 9840 11850 10300
rect 12070 9840 12126 10300
rect 12346 9840 12402 10300
rect 12622 9840 12678 10300
rect 12898 9840 12954 10300
rect 13174 9840 13230 10300
rect 13450 9840 13506 10300
rect 13726 9840 13782 10300
rect 14002 9840 14058 10300
rect 14278 9840 14334 10300
rect 14554 9840 14610 10300
rect 14830 9840 14886 10300
rect 15106 9840 15162 10300
rect 15382 9840 15438 10300
rect 15658 9840 15714 10300
rect 15934 9840 15990 10300
rect 16210 9840 16266 10300
rect 16486 9840 16542 10300
rect 16762 9840 16818 10300
rect 17038 9840 17094 10300
rect 17224 9852 17276 9858
rect 10784 8492 10836 8498
rect 10784 8434 10836 8440
rect 11152 8492 11204 8498
rect 11152 8434 11204 8440
rect 11256 8090 11284 9840
rect 11336 9172 11388 9178
rect 11336 9114 11388 9120
rect 11348 8498 11376 9114
rect 11532 8820 11560 9840
rect 11440 8792 11560 8820
rect 11808 8820 11836 9840
rect 11808 8792 11928 8820
rect 11440 8566 11468 8792
rect 11552 8732 11860 8741
rect 11552 8730 11558 8732
rect 11614 8730 11638 8732
rect 11694 8730 11718 8732
rect 11774 8730 11798 8732
rect 11854 8730 11860 8732
rect 11614 8678 11616 8730
rect 11796 8678 11798 8730
rect 11552 8676 11558 8678
rect 11614 8676 11638 8678
rect 11694 8676 11718 8678
rect 11774 8676 11798 8678
rect 11854 8676 11860 8678
rect 11552 8667 11860 8676
rect 11428 8560 11480 8566
rect 11428 8502 11480 8508
rect 11336 8492 11388 8498
rect 11336 8434 11388 8440
rect 10416 8084 10468 8090
rect 10416 8026 10468 8032
rect 10692 8084 10744 8090
rect 10692 8026 10744 8032
rect 11244 8084 11296 8090
rect 11244 8026 11296 8032
rect 11796 8084 11848 8090
rect 11900 8072 11928 8792
rect 12084 8634 12112 9840
rect 12256 9172 12308 9178
rect 12256 9114 12308 9120
rect 12072 8628 12124 8634
rect 12072 8570 12124 8576
rect 12268 8498 12296 9114
rect 12360 8634 12388 9840
rect 12532 9240 12584 9246
rect 12532 9182 12584 9188
rect 12348 8628 12400 8634
rect 12348 8570 12400 8576
rect 12544 8498 12572 9182
rect 12256 8492 12308 8498
rect 12256 8434 12308 8440
rect 12532 8492 12584 8498
rect 12532 8434 12584 8440
rect 12636 8090 12664 9840
rect 12912 9160 12940 9840
rect 12728 9132 12940 9160
rect 12992 9172 13044 9178
rect 12728 8430 12756 9132
rect 12992 9114 13044 9120
rect 13004 8498 13032 9114
rect 13084 8628 13136 8634
rect 13188 8616 13216 9840
rect 13360 8832 13412 8838
rect 13360 8774 13412 8780
rect 13136 8588 13216 8616
rect 13084 8570 13136 8576
rect 13372 8498 13400 8774
rect 12992 8492 13044 8498
rect 12992 8434 13044 8440
rect 13360 8492 13412 8498
rect 13360 8434 13412 8440
rect 12716 8424 12768 8430
rect 12716 8366 12768 8372
rect 13464 8090 13492 9840
rect 13740 9160 13768 9840
rect 13820 9240 13872 9246
rect 13820 9182 13872 9188
rect 13912 9240 13964 9246
rect 13912 9182 13964 9188
rect 13556 9132 13768 9160
rect 13556 8634 13584 9132
rect 13832 9110 13860 9182
rect 13820 9104 13872 9110
rect 13820 9046 13872 9052
rect 13636 9036 13688 9042
rect 13636 8978 13688 8984
rect 13648 8634 13676 8978
rect 13924 8956 13952 9182
rect 13832 8928 13952 8956
rect 13544 8628 13596 8634
rect 13544 8570 13596 8576
rect 13636 8628 13688 8634
rect 13636 8570 13688 8576
rect 13832 8566 13860 8928
rect 14016 8634 14044 9840
rect 14004 8628 14056 8634
rect 14004 8570 14056 8576
rect 13820 8560 13872 8566
rect 13820 8502 13872 8508
rect 14188 8288 14240 8294
rect 14188 8230 14240 8236
rect 11848 8044 11928 8072
rect 12624 8084 12676 8090
rect 11796 8026 11848 8032
rect 12624 8026 12676 8032
rect 13452 8084 13504 8090
rect 13452 8026 13504 8032
rect 12808 8016 12860 8022
rect 12808 7958 12860 7964
rect 13726 7984 13782 7993
rect 10692 7880 10744 7886
rect 10692 7822 10744 7828
rect 11886 7848 11942 7857
rect 10704 6866 10732 7822
rect 12820 7818 12848 7958
rect 13726 7919 13782 7928
rect 13740 7886 13768 7919
rect 13636 7880 13688 7886
rect 13636 7822 13688 7828
rect 13728 7880 13780 7886
rect 13728 7822 13780 7828
rect 11886 7783 11888 7792
rect 11940 7783 11942 7792
rect 12808 7812 12860 7818
rect 11888 7754 11940 7760
rect 12808 7754 12860 7760
rect 12900 7812 12952 7818
rect 12900 7754 12952 7760
rect 11980 7744 12032 7750
rect 11980 7686 12032 7692
rect 11552 7644 11860 7653
rect 11552 7642 11558 7644
rect 11614 7642 11638 7644
rect 11694 7642 11718 7644
rect 11774 7642 11798 7644
rect 11854 7642 11860 7644
rect 11614 7590 11616 7642
rect 11796 7590 11798 7642
rect 11552 7588 11558 7590
rect 11614 7588 11638 7590
rect 11694 7588 11718 7590
rect 11774 7588 11798 7590
rect 11854 7588 11860 7590
rect 11552 7579 11860 7588
rect 11992 6905 12020 7686
rect 12912 7585 12940 7754
rect 13648 7732 13676 7822
rect 13648 7704 13860 7732
rect 12898 7576 12954 7585
rect 12898 7511 12954 7520
rect 13832 7041 13860 7704
rect 13818 7032 13874 7041
rect 12348 6996 12400 7002
rect 13818 6967 13874 6976
rect 12348 6938 12400 6944
rect 11978 6896 12034 6905
rect 9220 6860 9272 6866
rect 9220 6802 9272 6808
rect 10140 6860 10192 6866
rect 10140 6802 10192 6808
rect 10692 6860 10744 6866
rect 11978 6831 12034 6840
rect 10692 6802 10744 6808
rect 11552 6556 11860 6565
rect 11552 6554 11558 6556
rect 11614 6554 11638 6556
rect 11694 6554 11718 6556
rect 11774 6554 11798 6556
rect 11854 6554 11860 6556
rect 11614 6502 11616 6554
rect 11796 6502 11798 6554
rect 11552 6500 11558 6502
rect 11614 6500 11638 6502
rect 11694 6500 11718 6502
rect 11774 6500 11798 6502
rect 11854 6500 11860 6502
rect 11552 6491 11860 6500
rect 7194 6216 7250 6225
rect 7194 6151 7250 6160
rect 6251 6012 6559 6021
rect 6251 6010 6257 6012
rect 6313 6010 6337 6012
rect 6393 6010 6417 6012
rect 6473 6010 6497 6012
rect 6553 6010 6559 6012
rect 6313 5958 6315 6010
rect 6495 5958 6497 6010
rect 6251 5956 6257 5958
rect 6313 5956 6337 5958
rect 6393 5956 6417 5958
rect 6473 5956 6497 5958
rect 6553 5956 6559 5958
rect 6251 5947 6559 5956
rect 12360 5817 12388 6938
rect 14200 6746 14228 8230
rect 14292 8090 14320 9840
rect 14280 8084 14332 8090
rect 14280 8026 14332 8032
rect 14372 7744 14424 7750
rect 14372 7686 14424 7692
rect 14384 7546 14412 7686
rect 14568 7546 14596 9840
rect 14648 9512 14700 9518
rect 14648 9454 14700 9460
rect 14740 9512 14792 9518
rect 14740 9454 14792 9460
rect 14660 8673 14688 9454
rect 14646 8664 14702 8673
rect 14646 8599 14702 8608
rect 14752 8498 14780 9454
rect 14740 8492 14792 8498
rect 14740 8434 14792 8440
rect 14844 8090 14872 9840
rect 15120 8566 15148 9840
rect 15200 8900 15252 8906
rect 15200 8842 15252 8848
rect 15292 8900 15344 8906
rect 15292 8842 15344 8848
rect 15108 8560 15160 8566
rect 15108 8502 15160 8508
rect 14832 8084 14884 8090
rect 14832 8026 14884 8032
rect 15108 7812 15160 7818
rect 15108 7754 15160 7760
rect 14372 7540 14424 7546
rect 14372 7482 14424 7488
rect 14556 7540 14608 7546
rect 14556 7482 14608 7488
rect 15120 7410 15148 7754
rect 14648 7404 14700 7410
rect 14648 7346 14700 7352
rect 15108 7404 15160 7410
rect 15108 7346 15160 7352
rect 14464 7200 14516 7206
rect 14464 7142 14516 7148
rect 14278 6760 14334 6769
rect 14200 6718 14278 6746
rect 14476 6730 14504 7142
rect 14660 7002 14688 7346
rect 14648 6996 14700 7002
rect 14648 6938 14700 6944
rect 14278 6695 14334 6704
rect 14464 6724 14516 6730
rect 14464 6666 14516 6672
rect 15212 6458 15240 8842
rect 15304 8566 15332 8842
rect 15396 8634 15424 9840
rect 15384 8628 15436 8634
rect 15384 8570 15436 8576
rect 15292 8560 15344 8566
rect 15292 8502 15344 8508
rect 15672 8090 15700 9840
rect 15948 8090 15976 9840
rect 16120 8968 16172 8974
rect 16120 8910 16172 8916
rect 15660 8084 15712 8090
rect 15660 8026 15712 8032
rect 15936 8084 15988 8090
rect 15936 8026 15988 8032
rect 15200 6452 15252 6458
rect 15200 6394 15252 6400
rect 16132 6390 16160 8910
rect 16224 8634 16252 9840
rect 16304 8968 16356 8974
rect 16304 8910 16356 8916
rect 16212 8628 16264 8634
rect 16212 8570 16264 8576
rect 16316 8498 16344 8910
rect 16304 8492 16356 8498
rect 16304 8434 16356 8440
rect 16396 8356 16448 8362
rect 16396 8298 16448 8304
rect 16408 7886 16436 8298
rect 16500 8090 16528 9840
rect 16776 8634 16804 9840
rect 16856 9648 16908 9654
rect 16856 9590 16908 9596
rect 16764 8628 16816 8634
rect 16764 8570 16816 8576
rect 16764 8492 16816 8498
rect 16764 8434 16816 8440
rect 16580 8288 16632 8294
rect 16580 8230 16632 8236
rect 16672 8288 16724 8294
rect 16672 8230 16724 8236
rect 16488 8084 16540 8090
rect 16488 8026 16540 8032
rect 16396 7880 16448 7886
rect 16396 7822 16448 7828
rect 16120 6384 16172 6390
rect 16120 6326 16172 6332
rect 16592 6322 16620 8230
rect 16684 7478 16712 8230
rect 16672 7472 16724 7478
rect 16776 7449 16804 8434
rect 16868 8401 16896 9590
rect 17052 8786 17080 9840
rect 17314 9840 17370 10300
rect 17590 9840 17646 10300
rect 17866 9840 17922 10300
rect 18142 9840 18198 10300
rect 18418 9840 18474 10300
rect 18694 9840 18750 10300
rect 18970 9840 19026 10300
rect 19076 9846 19196 9874
rect 17224 9794 17276 9800
rect 17236 9314 17264 9794
rect 17224 9308 17276 9314
rect 17224 9250 17276 9256
rect 17052 8758 17264 8786
rect 16946 8528 17002 8537
rect 16946 8463 17002 8472
rect 16960 8430 16988 8463
rect 16948 8424 17000 8430
rect 16854 8392 16910 8401
rect 16948 8366 17000 8372
rect 16854 8327 16910 8336
rect 16854 8188 17162 8197
rect 16854 8186 16860 8188
rect 16916 8186 16940 8188
rect 16996 8186 17020 8188
rect 17076 8186 17100 8188
rect 17156 8186 17162 8188
rect 16916 8134 16918 8186
rect 17098 8134 17100 8186
rect 16854 8132 16860 8134
rect 16916 8132 16940 8134
rect 16996 8132 17020 8134
rect 17076 8132 17100 8134
rect 17156 8132 17162 8134
rect 16854 8123 17162 8132
rect 17132 8016 17184 8022
rect 17236 8004 17264 8758
rect 17328 8566 17356 9840
rect 17500 9580 17552 9586
rect 17500 9522 17552 9528
rect 17512 8974 17540 9522
rect 17500 8968 17552 8974
rect 17500 8910 17552 8916
rect 17604 8634 17632 9840
rect 17776 9716 17828 9722
rect 17776 9658 17828 9664
rect 17682 9344 17738 9353
rect 17682 9279 17738 9288
rect 17592 8628 17644 8634
rect 17592 8570 17644 8576
rect 17316 8560 17368 8566
rect 17316 8502 17368 8508
rect 17408 8492 17460 8498
rect 17408 8434 17460 8440
rect 17316 8424 17368 8430
rect 17316 8366 17368 8372
rect 17184 7976 17264 8004
rect 17132 7958 17184 7964
rect 17040 7948 17092 7954
rect 17328 7936 17356 8366
rect 17040 7890 17092 7896
rect 17236 7908 17356 7936
rect 16948 7812 17000 7818
rect 16948 7754 17000 7760
rect 16960 7721 16988 7754
rect 16946 7712 17002 7721
rect 16946 7647 17002 7656
rect 16672 7414 16724 7420
rect 16762 7440 16818 7449
rect 16762 7375 16818 7384
rect 16764 7336 16816 7342
rect 16762 7304 16764 7313
rect 16816 7304 16818 7313
rect 16762 7239 16818 7248
rect 17052 7188 17080 7890
rect 17236 7546 17264 7908
rect 17224 7540 17276 7546
rect 17224 7482 17276 7488
rect 17420 7206 17448 8434
rect 17590 8120 17646 8129
rect 17590 8055 17592 8064
rect 17644 8055 17646 8064
rect 17592 8026 17644 8032
rect 17696 7970 17724 9279
rect 17788 8514 17816 9658
rect 17880 8634 17908 9840
rect 17960 9444 18012 9450
rect 17960 9386 18012 9392
rect 17868 8628 17920 8634
rect 17868 8570 17920 8576
rect 17788 8486 17908 8514
rect 17776 8424 17828 8430
rect 17776 8366 17828 8372
rect 17788 8090 17816 8366
rect 17776 8084 17828 8090
rect 17776 8026 17828 8032
rect 17696 7942 17816 7970
rect 17500 7812 17552 7818
rect 17500 7754 17552 7760
rect 17512 7528 17540 7754
rect 17512 7500 17632 7528
rect 17500 7404 17552 7410
rect 17500 7346 17552 7352
rect 17408 7200 17460 7206
rect 17052 7160 17264 7188
rect 17236 7154 17264 7160
rect 17314 7168 17370 7177
rect 17236 7126 17314 7154
rect 17408 7142 17460 7148
rect 16854 7100 17162 7109
rect 17314 7103 17370 7112
rect 16854 7098 16860 7100
rect 16916 7098 16940 7100
rect 16996 7098 17020 7100
rect 17076 7098 17100 7100
rect 17156 7098 17162 7100
rect 16916 7046 16918 7098
rect 17098 7046 17100 7098
rect 16854 7044 16860 7046
rect 16916 7044 16940 7046
rect 16996 7044 17020 7046
rect 17076 7044 17100 7046
rect 17156 7044 17162 7046
rect 16670 7032 16726 7041
rect 16854 7035 17162 7044
rect 17314 7032 17370 7041
rect 16726 6976 17314 6984
rect 16670 6967 17370 6976
rect 16684 6956 17356 6967
rect 17512 6934 17540 7346
rect 17604 7256 17632 7500
rect 17788 7478 17816 7942
rect 17776 7472 17828 7478
rect 17776 7414 17828 7420
rect 17880 7410 17908 8486
rect 17972 8090 18000 9386
rect 18156 8616 18184 9840
rect 18328 9716 18380 9722
rect 18328 9658 18380 9664
rect 18236 8628 18288 8634
rect 18156 8588 18236 8616
rect 18236 8570 18288 8576
rect 18340 8514 18368 9658
rect 18052 8492 18104 8498
rect 18052 8434 18104 8440
rect 18156 8486 18368 8514
rect 17960 8084 18012 8090
rect 17960 8026 18012 8032
rect 17960 7744 18012 7750
rect 17960 7686 18012 7692
rect 17868 7404 17920 7410
rect 17868 7346 17920 7352
rect 17868 7268 17920 7274
rect 17604 7228 17868 7256
rect 17868 7210 17920 7216
rect 17500 6928 17552 6934
rect 17500 6870 17552 6876
rect 17972 6798 18000 7686
rect 18064 7546 18092 8434
rect 18052 7540 18104 7546
rect 18052 7482 18104 7488
rect 18156 7410 18184 8486
rect 18328 8288 18380 8294
rect 18328 8230 18380 8236
rect 18340 7970 18368 8230
rect 18432 8090 18460 9840
rect 18604 9444 18656 9450
rect 18604 9386 18656 9392
rect 18512 8968 18564 8974
rect 18512 8910 18564 8916
rect 18420 8084 18472 8090
rect 18420 8026 18472 8032
rect 18340 7942 18460 7970
rect 18524 7954 18552 8910
rect 18236 7880 18288 7886
rect 18236 7822 18288 7828
rect 18328 7880 18380 7886
rect 18328 7822 18380 7828
rect 18144 7404 18196 7410
rect 18144 7346 18196 7352
rect 18052 7336 18104 7342
rect 18052 7278 18104 7284
rect 18064 6798 18092 7278
rect 18248 6798 18276 7822
rect 18340 6798 18368 7822
rect 18432 7818 18460 7942
rect 18512 7948 18564 7954
rect 18512 7890 18564 7896
rect 18420 7812 18472 7818
rect 18420 7754 18472 7760
rect 18616 7410 18644 9386
rect 18708 8362 18736 9840
rect 18880 9308 18932 9314
rect 18880 9250 18932 9256
rect 18786 8664 18842 8673
rect 18786 8599 18842 8608
rect 18696 8356 18748 8362
rect 18696 8298 18748 8304
rect 18800 7886 18828 8599
rect 18696 7880 18748 7886
rect 18696 7822 18748 7828
rect 18788 7880 18840 7886
rect 18788 7822 18840 7828
rect 18708 7546 18736 7822
rect 18696 7540 18748 7546
rect 18696 7482 18748 7488
rect 18604 7404 18656 7410
rect 18604 7346 18656 7352
rect 18892 7290 18920 9250
rect 18984 9081 19012 9840
rect 18970 9072 19026 9081
rect 18970 9007 19026 9016
rect 19076 8634 19104 9846
rect 19168 9840 19196 9846
rect 19246 9840 19302 10300
rect 19522 9840 19578 10300
rect 19614 9888 19670 9897
rect 19168 9812 19288 9840
rect 19536 9832 19614 9840
rect 19798 9840 19854 10300
rect 19984 9920 20036 9926
rect 19984 9862 20036 9868
rect 19536 9823 19670 9832
rect 19536 9812 19656 9823
rect 19246 9072 19302 9081
rect 19246 9007 19302 9016
rect 19260 8956 19288 9007
rect 19260 8928 19380 8956
rect 19352 8809 19380 8928
rect 19338 8800 19394 8809
rect 19338 8735 19394 8744
rect 19614 8800 19670 8809
rect 19614 8735 19670 8744
rect 19628 8634 19656 8735
rect 19706 8664 19762 8673
rect 19064 8628 19116 8634
rect 19064 8570 19116 8576
rect 19616 8628 19668 8634
rect 19706 8599 19762 8608
rect 19812 8616 19840 9840
rect 19996 8634 20024 9862
rect 20074 9840 20130 10300
rect 20168 9920 20220 9926
rect 20168 9862 20220 9868
rect 20088 8650 20116 9840
rect 20180 9654 20208 9862
rect 20350 9840 20406 10300
rect 20626 9840 20682 10300
rect 20902 9840 20958 10300
rect 21178 9840 21234 10300
rect 21454 9840 21510 10300
rect 21730 9840 21786 10300
rect 22006 9840 22062 10300
rect 22098 9888 22154 9897
rect 20168 9648 20220 9654
rect 20168 9590 20220 9596
rect 20364 8888 20392 9840
rect 20272 8860 20392 8888
rect 19984 8628 20036 8634
rect 19616 8570 19668 8576
rect 19340 8560 19392 8566
rect 19260 8508 19340 8514
rect 19260 8502 19392 8508
rect 19064 8492 19116 8498
rect 18984 8452 19064 8480
rect 18984 7410 19012 8452
rect 19064 8434 19116 8440
rect 19260 8486 19380 8502
rect 19062 8392 19118 8401
rect 19062 8327 19118 8336
rect 19076 8022 19104 8327
rect 19064 8016 19116 8022
rect 19064 7958 19116 7964
rect 19064 7880 19116 7886
rect 19064 7822 19116 7828
rect 19156 7880 19208 7886
rect 19156 7822 19208 7828
rect 19076 7546 19104 7822
rect 19168 7721 19196 7822
rect 19154 7712 19210 7721
rect 19154 7647 19210 7656
rect 19260 7546 19288 8486
rect 19340 8424 19392 8430
rect 19338 8392 19340 8401
rect 19392 8392 19394 8401
rect 19338 8327 19394 8336
rect 19430 7984 19486 7993
rect 19430 7919 19486 7928
rect 19340 7880 19392 7886
rect 19444 7868 19472 7919
rect 19392 7840 19472 7868
rect 19340 7822 19392 7828
rect 19338 7712 19394 7721
rect 19338 7647 19394 7656
rect 19064 7540 19116 7546
rect 19064 7482 19116 7488
rect 19248 7540 19300 7546
rect 19248 7482 19300 7488
rect 18972 7404 19024 7410
rect 18972 7346 19024 7352
rect 19064 7404 19116 7410
rect 19064 7346 19116 7352
rect 19076 7290 19104 7346
rect 18892 7262 19104 7290
rect 19352 7274 19380 7647
rect 19430 7440 19486 7449
rect 19430 7375 19486 7384
rect 19614 7440 19670 7449
rect 19720 7410 19748 8599
rect 19812 8588 19932 8616
rect 19800 8492 19852 8498
rect 19800 8434 19852 8440
rect 19812 7546 19840 8434
rect 19800 7540 19852 7546
rect 19800 7482 19852 7488
rect 19614 7375 19670 7384
rect 19708 7404 19760 7410
rect 19444 7274 19472 7375
rect 19340 7268 19392 7274
rect 19340 7210 19392 7216
rect 19432 7268 19484 7274
rect 19432 7210 19484 7216
rect 19628 6798 19656 7375
rect 19708 7346 19760 7352
rect 19800 7404 19852 7410
rect 19800 7346 19852 7352
rect 17960 6792 18012 6798
rect 17960 6734 18012 6740
rect 18052 6792 18104 6798
rect 18052 6734 18104 6740
rect 18236 6792 18288 6798
rect 18236 6734 18288 6740
rect 18328 6792 18380 6798
rect 18328 6734 18380 6740
rect 19616 6792 19668 6798
rect 19812 6780 19840 7346
rect 19904 7290 19932 8588
rect 20088 8622 20208 8650
rect 19984 8570 20036 8576
rect 20076 8288 20128 8294
rect 20076 8230 20128 8236
rect 20088 7886 20116 8230
rect 20076 7880 20128 7886
rect 20076 7822 20128 7828
rect 20180 7732 20208 8622
rect 20272 8022 20300 8860
rect 20444 8492 20496 8498
rect 20640 8480 20668 9840
rect 20720 9580 20772 9586
rect 20720 9522 20772 9528
rect 20496 8452 20668 8480
rect 20444 8434 20496 8440
rect 20352 8288 20404 8294
rect 20352 8230 20404 8236
rect 20260 8016 20312 8022
rect 20260 7958 20312 7964
rect 20364 7886 20392 8230
rect 20444 8016 20496 8022
rect 20442 7984 20444 7993
rect 20496 7984 20498 7993
rect 20442 7919 20498 7928
rect 20352 7880 20404 7886
rect 20352 7822 20404 7828
rect 19982 7712 20038 7721
rect 19982 7647 20038 7656
rect 20088 7704 20208 7732
rect 20260 7744 20312 7750
rect 19996 7410 20024 7647
rect 20088 7478 20116 7704
rect 20260 7686 20312 7692
rect 20352 7744 20404 7750
rect 20352 7686 20404 7692
rect 20076 7472 20128 7478
rect 20076 7414 20128 7420
rect 19984 7404 20036 7410
rect 19984 7346 20036 7352
rect 19904 7262 20116 7290
rect 20088 6798 20116 7262
rect 19892 6792 19944 6798
rect 19812 6752 19892 6780
rect 19616 6734 19668 6740
rect 19892 6734 19944 6740
rect 20076 6792 20128 6798
rect 20076 6734 20128 6740
rect 20272 6458 20300 7686
rect 20260 6452 20312 6458
rect 20260 6394 20312 6400
rect 20364 6390 20392 7686
rect 20732 7206 20760 9522
rect 20812 8900 20864 8906
rect 20812 8842 20864 8848
rect 20824 8378 20852 8842
rect 20916 8498 20944 9840
rect 21088 9784 21140 9790
rect 21088 9726 21140 9732
rect 20994 9616 21050 9625
rect 20994 9551 20996 9560
rect 21048 9551 21050 9560
rect 20996 9522 21048 9528
rect 20996 9308 21048 9314
rect 20996 9250 21048 9256
rect 21008 8906 21036 9250
rect 20996 8900 21048 8906
rect 20996 8842 21048 8848
rect 20904 8492 20956 8498
rect 20904 8434 20956 8440
rect 21100 8378 21128 9726
rect 21192 8498 21220 9840
rect 21364 9512 21416 9518
rect 21364 9454 21416 9460
rect 21180 8492 21232 8498
rect 21180 8434 21232 8440
rect 20824 8350 20944 8378
rect 20812 8288 20864 8294
rect 20812 8230 20864 8236
rect 20824 7546 20852 8230
rect 20916 8022 20944 8350
rect 21008 8350 21128 8378
rect 20904 8016 20956 8022
rect 20904 7958 20956 7964
rect 21008 7886 21036 8350
rect 21088 8288 21140 8294
rect 21088 8230 21140 8236
rect 21100 8022 21128 8230
rect 21376 8106 21404 9454
rect 21468 8498 21496 9840
rect 21548 9716 21600 9722
rect 21548 9658 21600 9664
rect 21560 8498 21588 9658
rect 21638 9480 21694 9489
rect 21638 9415 21694 9424
rect 21652 9246 21680 9415
rect 21640 9240 21692 9246
rect 21640 9182 21692 9188
rect 21638 8936 21694 8945
rect 21638 8871 21694 8880
rect 21652 8838 21680 8871
rect 21640 8832 21692 8838
rect 21640 8774 21692 8780
rect 21638 8528 21694 8537
rect 21456 8492 21508 8498
rect 21456 8434 21508 8440
rect 21548 8492 21600 8498
rect 21744 8498 21772 9840
rect 21916 9648 21968 9654
rect 21916 9590 21968 9596
rect 21824 9580 21876 9586
rect 21824 9522 21876 9528
rect 21836 9353 21864 9522
rect 21822 9344 21878 9353
rect 21822 9279 21878 9288
rect 21822 9208 21878 9217
rect 21928 9178 21956 9590
rect 21822 9143 21824 9152
rect 21876 9143 21878 9152
rect 21916 9172 21968 9178
rect 21824 9114 21876 9120
rect 21916 9114 21968 9120
rect 21638 8463 21694 8472
rect 21732 8492 21784 8498
rect 21548 8434 21600 8440
rect 21456 8288 21508 8294
rect 21456 8230 21508 8236
rect 21548 8288 21600 8294
rect 21548 8230 21600 8236
rect 21192 8078 21404 8106
rect 21192 8022 21220 8078
rect 21088 8016 21140 8022
rect 21088 7958 21140 7964
rect 21180 8016 21232 8022
rect 21180 7958 21232 7964
rect 21362 7984 21418 7993
rect 21362 7919 21418 7928
rect 21376 7886 21404 7919
rect 20996 7880 21048 7886
rect 20996 7822 21048 7828
rect 21180 7880 21232 7886
rect 21180 7822 21232 7828
rect 21364 7880 21416 7886
rect 21364 7822 21416 7828
rect 20812 7540 20864 7546
rect 20812 7482 20864 7488
rect 21192 7478 21220 7822
rect 21180 7472 21232 7478
rect 21180 7414 21232 7420
rect 21272 7404 21324 7410
rect 21468 7392 21496 8230
rect 21560 7546 21588 8230
rect 21652 8004 21680 8463
rect 22020 8480 22048 9840
rect 22098 9823 22100 9832
rect 22152 9823 22154 9832
rect 22192 9852 22244 9858
rect 22100 9794 22152 9800
rect 22282 9840 22338 10300
rect 22558 9840 22614 10300
rect 22834 9840 22890 10300
rect 23020 9988 23072 9994
rect 23020 9930 23072 9936
rect 22192 9794 22244 9800
rect 22204 9738 22232 9794
rect 22112 9710 22232 9738
rect 22112 9110 22140 9710
rect 22190 9616 22246 9625
rect 22190 9551 22246 9560
rect 22204 9450 22232 9551
rect 22192 9444 22244 9450
rect 22192 9386 22244 9392
rect 22296 9194 22324 9840
rect 22572 9296 22600 9840
rect 22572 9268 22692 9296
rect 22296 9166 22600 9194
rect 22100 9104 22152 9110
rect 22192 9104 22244 9110
rect 22100 9046 22152 9052
rect 22190 9072 22192 9081
rect 22244 9072 22246 9081
rect 22190 9007 22246 9016
rect 22155 8732 22463 8741
rect 22155 8730 22161 8732
rect 22217 8730 22241 8732
rect 22297 8730 22321 8732
rect 22377 8730 22401 8732
rect 22457 8730 22463 8732
rect 22217 8678 22219 8730
rect 22399 8678 22401 8730
rect 22155 8676 22161 8678
rect 22217 8676 22241 8678
rect 22297 8676 22321 8678
rect 22377 8676 22401 8678
rect 22457 8676 22463 8678
rect 22155 8667 22463 8676
rect 22468 8628 22520 8634
rect 22468 8570 22520 8576
rect 22100 8492 22152 8498
rect 22020 8452 22100 8480
rect 21732 8434 21784 8440
rect 22100 8434 22152 8440
rect 22192 8356 22244 8362
rect 22192 8298 22244 8304
rect 22100 8288 22152 8294
rect 22100 8230 22152 8236
rect 21732 8016 21784 8022
rect 21652 7976 21732 8004
rect 21732 7958 21784 7964
rect 22112 7834 22140 8230
rect 22020 7806 22140 7834
rect 21824 7744 21876 7750
rect 21824 7686 21876 7692
rect 21548 7540 21600 7546
rect 21548 7482 21600 7488
rect 21324 7364 21496 7392
rect 21272 7346 21324 7352
rect 21178 7304 21234 7313
rect 21178 7239 21180 7248
rect 21232 7239 21234 7248
rect 21180 7210 21232 7216
rect 20628 7200 20680 7206
rect 20628 7142 20680 7148
rect 20720 7200 20772 7206
rect 21456 7200 21508 7206
rect 20720 7142 20772 7148
rect 21362 7168 21418 7177
rect 20352 6384 20404 6390
rect 20352 6326 20404 6332
rect 20640 6322 20668 7142
rect 21418 7148 21456 7154
rect 21418 7142 21508 7148
rect 21418 7126 21496 7142
rect 21362 7103 21418 7112
rect 21836 6866 21864 7686
rect 22020 7546 22048 7806
rect 22204 7750 22232 8298
rect 22376 8288 22428 8294
rect 22376 8230 22428 8236
rect 22388 7954 22416 8230
rect 22376 7948 22428 7954
rect 22376 7890 22428 7896
rect 22282 7848 22338 7857
rect 22480 7834 22508 8570
rect 22572 8498 22600 9166
rect 22560 8492 22612 8498
rect 22664 8480 22692 9268
rect 22742 9208 22798 9217
rect 22848 9194 22876 9840
rect 22928 9648 22980 9654
rect 22928 9590 22980 9596
rect 22940 9382 22968 9590
rect 22928 9376 22980 9382
rect 22928 9318 22980 9324
rect 22848 9166 22968 9194
rect 22742 9143 22798 9152
rect 22756 8634 22784 9143
rect 22744 8628 22796 8634
rect 22744 8570 22796 8576
rect 22940 8498 22968 9166
rect 22836 8492 22888 8498
rect 22664 8452 22836 8480
rect 22560 8434 22612 8440
rect 22836 8434 22888 8440
rect 22928 8492 22980 8498
rect 22928 8434 22980 8440
rect 22650 8392 22706 8401
rect 22650 8327 22706 8336
rect 22664 7954 22692 8327
rect 22928 8288 22980 8294
rect 22928 8230 22980 8236
rect 22652 7948 22704 7954
rect 22652 7890 22704 7896
rect 22940 7886 22968 8230
rect 22928 7880 22980 7886
rect 22480 7806 22692 7834
rect 22928 7822 22980 7828
rect 22282 7783 22338 7792
rect 22296 7750 22324 7783
rect 22192 7744 22244 7750
rect 22192 7686 22244 7692
rect 22284 7744 22336 7750
rect 22284 7686 22336 7692
rect 22560 7744 22612 7750
rect 22560 7686 22612 7692
rect 22155 7644 22463 7653
rect 22155 7642 22161 7644
rect 22217 7642 22241 7644
rect 22297 7642 22321 7644
rect 22377 7642 22401 7644
rect 22457 7642 22463 7644
rect 22217 7590 22219 7642
rect 22399 7590 22401 7642
rect 22155 7588 22161 7590
rect 22217 7588 22241 7590
rect 22297 7588 22321 7590
rect 22377 7588 22401 7590
rect 22457 7588 22463 7590
rect 22155 7579 22463 7588
rect 22008 7540 22060 7546
rect 22008 7482 22060 7488
rect 21824 6860 21876 6866
rect 21824 6802 21876 6808
rect 22572 6769 22600 7686
rect 22664 7546 22692 7806
rect 23032 7750 23060 9930
rect 23110 9840 23166 10300
rect 23204 9988 23256 9994
rect 23204 9930 23256 9936
rect 23124 9194 23152 9840
rect 23216 9761 23244 9930
rect 23386 9840 23442 10300
rect 23572 9920 23624 9926
rect 23572 9862 23624 9868
rect 23202 9752 23258 9761
rect 23202 9687 23258 9696
rect 23296 9308 23348 9314
rect 23296 9250 23348 9256
rect 23124 9166 23244 9194
rect 23112 8900 23164 8906
rect 23112 8842 23164 8848
rect 22836 7744 22888 7750
rect 22836 7686 22888 7692
rect 23020 7744 23072 7750
rect 23020 7686 23072 7692
rect 22652 7540 22704 7546
rect 22652 7482 22704 7488
rect 22558 6760 22614 6769
rect 22558 6695 22614 6704
rect 22155 6556 22463 6565
rect 22155 6554 22161 6556
rect 22217 6554 22241 6556
rect 22297 6554 22321 6556
rect 22377 6554 22401 6556
rect 22457 6554 22463 6556
rect 22217 6502 22219 6554
rect 22399 6502 22401 6554
rect 22155 6500 22161 6502
rect 22217 6500 22241 6502
rect 22297 6500 22321 6502
rect 22377 6500 22401 6502
rect 22457 6500 22463 6502
rect 22155 6491 22463 6500
rect 16580 6316 16632 6322
rect 16580 6258 16632 6264
rect 20628 6316 20680 6322
rect 20628 6258 20680 6264
rect 16854 6012 17162 6021
rect 16854 6010 16860 6012
rect 16916 6010 16940 6012
rect 16996 6010 17020 6012
rect 17076 6010 17100 6012
rect 17156 6010 17162 6012
rect 16916 5958 16918 6010
rect 17098 5958 17100 6010
rect 16854 5956 16860 5958
rect 16916 5956 16940 5958
rect 16996 5956 17020 5958
rect 17076 5956 17100 5958
rect 17156 5956 17162 5958
rect 16854 5947 17162 5956
rect 22848 5817 22876 7686
rect 23124 7478 23152 8842
rect 23216 8480 23244 9166
rect 23308 8945 23336 9250
rect 23400 9194 23428 9840
rect 23400 9166 23520 9194
rect 23294 8936 23350 8945
rect 23294 8871 23350 8880
rect 23492 8498 23520 9166
rect 23388 8492 23440 8498
rect 23216 8452 23388 8480
rect 23388 8434 23440 8440
rect 23480 8492 23532 8498
rect 23480 8434 23532 8440
rect 23584 8378 23612 9862
rect 23662 9840 23718 10300
rect 23938 9840 23994 10300
rect 24214 9840 24270 10300
rect 24490 9840 24546 10300
rect 24766 9840 24822 10300
rect 25042 9840 25098 10300
rect 25318 9840 25374 10300
rect 25594 9840 25650 10300
rect 25870 9840 25926 10300
rect 26146 9840 26202 10300
rect 26422 9840 26478 10300
rect 26698 9840 26754 10300
rect 26974 9840 27030 10300
rect 27160 9988 27212 9994
rect 27160 9930 27212 9936
rect 23676 9194 23704 9840
rect 23952 9194 23980 9840
rect 23676 9166 23796 9194
rect 23952 9166 24072 9194
rect 23768 8480 23796 9166
rect 24044 8498 24072 9166
rect 24124 9036 24176 9042
rect 24124 8978 24176 8984
rect 23940 8492 23992 8498
rect 23768 8452 23940 8480
rect 23940 8434 23992 8440
rect 24032 8492 24084 8498
rect 24032 8434 24084 8440
rect 23584 8350 23704 8378
rect 23204 8288 23256 8294
rect 23204 8230 23256 8236
rect 23480 8288 23532 8294
rect 23480 8230 23532 8236
rect 23572 8288 23624 8294
rect 23572 8230 23624 8236
rect 23216 7546 23244 8230
rect 23492 8106 23520 8230
rect 23400 8078 23520 8106
rect 23400 7954 23428 8078
rect 23584 7970 23612 8230
rect 23388 7948 23440 7954
rect 23388 7890 23440 7896
rect 23492 7942 23612 7970
rect 23492 7886 23520 7942
rect 23296 7880 23348 7886
rect 23296 7822 23348 7828
rect 23480 7880 23532 7886
rect 23480 7822 23532 7828
rect 23308 7546 23336 7822
rect 23676 7750 23704 8350
rect 24032 8288 24084 8294
rect 24032 8230 24084 8236
rect 24044 7886 24072 8230
rect 23848 7880 23900 7886
rect 23848 7822 23900 7828
rect 24032 7880 24084 7886
rect 24032 7822 24084 7828
rect 23388 7744 23440 7750
rect 23388 7686 23440 7692
rect 23664 7744 23716 7750
rect 23664 7686 23716 7692
rect 23204 7540 23256 7546
rect 23204 7482 23256 7488
rect 23296 7540 23348 7546
rect 23296 7482 23348 7488
rect 23112 7472 23164 7478
rect 23112 7414 23164 7420
rect 23400 6905 23428 7686
rect 23860 7274 23888 7822
rect 24136 7750 24164 8978
rect 24228 8480 24256 9840
rect 24400 8492 24452 8498
rect 24228 8452 24400 8480
rect 24504 8480 24532 9840
rect 24584 9240 24636 9246
rect 24584 9182 24636 9188
rect 24596 8906 24624 9182
rect 24584 8900 24636 8906
rect 24584 8842 24636 8848
rect 24780 8498 24808 9840
rect 24952 9104 25004 9110
rect 24952 9046 25004 9052
rect 24676 8492 24728 8498
rect 24504 8452 24676 8480
rect 24400 8434 24452 8440
rect 24676 8434 24728 8440
rect 24768 8492 24820 8498
rect 24768 8434 24820 8440
rect 24964 8362 24992 9046
rect 25056 8480 25084 9840
rect 25332 8498 25360 9840
rect 25412 9172 25464 9178
rect 25412 9114 25464 9120
rect 25228 8492 25280 8498
rect 25056 8452 25228 8480
rect 25228 8434 25280 8440
rect 25320 8492 25372 8498
rect 25320 8434 25372 8440
rect 25424 8430 25452 9114
rect 25608 8480 25636 9840
rect 25686 9480 25742 9489
rect 25686 9415 25742 9424
rect 25700 8616 25728 9415
rect 25884 9194 25912 9840
rect 25884 9166 26096 9194
rect 25964 8628 26016 8634
rect 25700 8588 25912 8616
rect 25780 8492 25832 8498
rect 25608 8452 25780 8480
rect 25780 8434 25832 8440
rect 25412 8424 25464 8430
rect 25412 8366 25464 8372
rect 24952 8356 25004 8362
rect 24952 8298 25004 8304
rect 24584 8288 24636 8294
rect 24584 8230 24636 8236
rect 24860 8288 24912 8294
rect 24860 8230 24912 8236
rect 25136 8288 25188 8294
rect 25136 8230 25188 8236
rect 25412 8288 25464 8294
rect 25412 8230 25464 8236
rect 25504 8288 25556 8294
rect 25504 8230 25556 8236
rect 25594 8256 25650 8265
rect 24596 7886 24624 8230
rect 24872 7886 24900 8230
rect 24950 8120 25006 8129
rect 24950 8055 24952 8064
rect 25004 8055 25006 8064
rect 24952 8026 25004 8032
rect 25148 7886 25176 8230
rect 25424 7886 25452 8230
rect 24584 7880 24636 7886
rect 24768 7880 24820 7886
rect 24584 7822 24636 7828
rect 24766 7848 24768 7857
rect 24860 7880 24912 7886
rect 24820 7848 24822 7857
rect 24860 7822 24912 7828
rect 25136 7880 25188 7886
rect 25136 7822 25188 7828
rect 25412 7880 25464 7886
rect 25412 7822 25464 7828
rect 24766 7783 24822 7792
rect 23940 7744 23992 7750
rect 23940 7686 23992 7692
rect 24124 7744 24176 7750
rect 24124 7686 24176 7692
rect 24400 7744 24452 7750
rect 24400 7686 24452 7692
rect 24676 7744 24728 7750
rect 24676 7686 24728 7692
rect 25228 7744 25280 7750
rect 25228 7686 25280 7692
rect 23848 7268 23900 7274
rect 23848 7210 23900 7216
rect 23952 7041 23980 7686
rect 23938 7032 23994 7041
rect 23938 6967 23994 6976
rect 23386 6896 23442 6905
rect 23386 6831 23442 6840
rect 24412 6225 24440 7686
rect 24688 6361 24716 7686
rect 24768 7200 24820 7206
rect 24768 7142 24820 7148
rect 24780 7002 24808 7142
rect 25240 7002 25268 7686
rect 25516 7478 25544 8230
rect 25594 8191 25650 8200
rect 25608 7970 25636 8191
rect 25884 8090 25912 8588
rect 25964 8570 26016 8576
rect 25976 8378 26004 8570
rect 26068 8498 26096 9166
rect 26160 8498 26188 9840
rect 26056 8492 26108 8498
rect 26056 8434 26108 8440
rect 26148 8492 26200 8498
rect 26436 8480 26464 9840
rect 26712 8498 26740 9840
rect 26792 9784 26844 9790
rect 26792 9726 26844 9732
rect 26804 9382 26832 9726
rect 26884 9648 26936 9654
rect 26884 9590 26936 9596
rect 26792 9376 26844 9382
rect 26792 9318 26844 9324
rect 26608 8492 26660 8498
rect 26436 8452 26608 8480
rect 26148 8434 26200 8440
rect 26608 8434 26660 8440
rect 26700 8492 26752 8498
rect 26700 8434 26752 8440
rect 25976 8350 26096 8378
rect 25964 8288 26016 8294
rect 25964 8230 26016 8236
rect 25872 8084 25924 8090
rect 25872 8026 25924 8032
rect 25608 7954 25820 7970
rect 25608 7948 25832 7954
rect 25608 7942 25780 7948
rect 25780 7890 25832 7896
rect 25976 7886 26004 8230
rect 25964 7880 26016 7886
rect 25964 7822 26016 7828
rect 25504 7472 25556 7478
rect 25504 7414 25556 7420
rect 26068 7206 26096 8350
rect 26148 8356 26200 8362
rect 26148 8298 26200 8304
rect 26160 7750 26188 8298
rect 26240 8288 26292 8294
rect 26240 8230 26292 8236
rect 26516 8288 26568 8294
rect 26516 8230 26568 8236
rect 26792 8288 26844 8294
rect 26792 8230 26844 8236
rect 26252 7886 26280 8230
rect 26528 7886 26556 8230
rect 26804 7886 26832 8230
rect 26240 7880 26292 7886
rect 26240 7822 26292 7828
rect 26516 7880 26568 7886
rect 26516 7822 26568 7828
rect 26792 7880 26844 7886
rect 26792 7822 26844 7828
rect 26896 7750 26924 9590
rect 26988 8566 27016 9840
rect 27068 8900 27120 8906
rect 27068 8842 27120 8848
rect 27080 8634 27108 8842
rect 27068 8628 27120 8634
rect 27068 8570 27120 8576
rect 26976 8560 27028 8566
rect 26976 8502 27028 8508
rect 26976 8288 27028 8294
rect 26976 8230 27028 8236
rect 26148 7744 26200 7750
rect 26148 7686 26200 7692
rect 26884 7744 26936 7750
rect 26884 7686 26936 7692
rect 26988 7478 27016 8230
rect 27172 7750 27200 9930
rect 27250 9840 27306 10300
rect 27526 9840 27582 10300
rect 27802 9840 27858 10300
rect 28078 9840 28134 10300
rect 28172 9852 28224 9858
rect 27264 8480 27292 9840
rect 27540 8616 27568 9840
rect 27540 8588 27660 8616
rect 27632 8498 27660 8588
rect 27528 8492 27580 8498
rect 27264 8452 27528 8480
rect 27528 8434 27580 8440
rect 27620 8492 27672 8498
rect 27816 8480 27844 9840
rect 28092 8566 28120 9840
rect 28354 9840 28410 10300
rect 28460 9846 28580 9874
rect 28460 9840 28488 9846
rect 28368 9812 28488 9840
rect 28172 9794 28224 9800
rect 28080 8560 28132 8566
rect 28080 8502 28132 8508
rect 27988 8492 28040 8498
rect 27816 8452 27988 8480
rect 27620 8434 27672 8440
rect 27988 8434 28040 8440
rect 27250 8392 27306 8401
rect 27250 8327 27252 8336
rect 27304 8327 27306 8336
rect 27896 8356 27948 8362
rect 27252 8298 27304 8304
rect 27896 8298 27948 8304
rect 27344 8288 27396 8294
rect 27344 8230 27396 8236
rect 27804 8288 27856 8294
rect 27804 8230 27856 8236
rect 27356 7886 27384 8230
rect 27457 8188 27765 8197
rect 27457 8186 27463 8188
rect 27519 8186 27543 8188
rect 27599 8186 27623 8188
rect 27679 8186 27703 8188
rect 27759 8186 27765 8188
rect 27519 8134 27521 8186
rect 27701 8134 27703 8186
rect 27457 8132 27463 8134
rect 27519 8132 27543 8134
rect 27599 8132 27623 8134
rect 27679 8132 27703 8134
rect 27759 8132 27765 8134
rect 27457 8123 27765 8132
rect 27816 7886 27844 8230
rect 27908 8090 27936 8298
rect 27988 8288 28040 8294
rect 27988 8230 28040 8236
rect 28080 8288 28132 8294
rect 28080 8230 28132 8236
rect 27896 8084 27948 8090
rect 27896 8026 27948 8032
rect 28000 7886 28028 8230
rect 28092 8090 28120 8230
rect 28080 8084 28132 8090
rect 28080 8026 28132 8032
rect 27344 7880 27396 7886
rect 27344 7822 27396 7828
rect 27804 7880 27856 7886
rect 27804 7822 27856 7828
rect 27988 7880 28040 7886
rect 27988 7822 28040 7828
rect 28080 7812 28132 7818
rect 28080 7754 28132 7760
rect 27160 7744 27212 7750
rect 27160 7686 27212 7692
rect 27436 7744 27488 7750
rect 27436 7686 27488 7692
rect 26976 7472 27028 7478
rect 26976 7414 27028 7420
rect 27448 7313 27476 7686
rect 27434 7304 27490 7313
rect 27434 7239 27490 7248
rect 26056 7200 26108 7206
rect 26056 7142 26108 7148
rect 27457 7100 27765 7109
rect 27457 7098 27463 7100
rect 27519 7098 27543 7100
rect 27599 7098 27623 7100
rect 27679 7098 27703 7100
rect 27759 7098 27765 7100
rect 27519 7046 27521 7098
rect 27701 7046 27703 7098
rect 27457 7044 27463 7046
rect 27519 7044 27543 7046
rect 27599 7044 27623 7046
rect 27679 7044 27703 7046
rect 27759 7044 27765 7046
rect 27457 7035 27765 7044
rect 24768 6996 24820 7002
rect 24768 6938 24820 6944
rect 25228 6996 25280 7002
rect 25228 6938 25280 6944
rect 24674 6352 24730 6361
rect 24674 6287 24730 6296
rect 24398 6216 24454 6225
rect 24398 6151 24454 6160
rect 27457 6012 27765 6021
rect 27457 6010 27463 6012
rect 27519 6010 27543 6012
rect 27599 6010 27623 6012
rect 27679 6010 27703 6012
rect 27759 6010 27765 6012
rect 27519 5958 27521 6010
rect 27701 5958 27703 6010
rect 27457 5956 27463 5958
rect 27519 5956 27543 5958
rect 27599 5956 27623 5958
rect 27679 5956 27703 5958
rect 27759 5956 27765 5958
rect 27457 5947 27765 5956
rect 12346 5808 12402 5817
rect 12346 5743 12402 5752
rect 22834 5808 22890 5817
rect 22834 5743 22890 5752
rect 25964 5704 26016 5710
rect 25964 5646 26016 5652
rect 23020 5636 23072 5642
rect 23020 5578 23072 5584
rect 11552 5468 11860 5477
rect 11552 5466 11558 5468
rect 11614 5466 11638 5468
rect 11694 5466 11718 5468
rect 11774 5466 11798 5468
rect 11854 5466 11860 5468
rect 11614 5414 11616 5466
rect 11796 5414 11798 5466
rect 11552 5412 11558 5414
rect 11614 5412 11638 5414
rect 11694 5412 11718 5414
rect 11774 5412 11798 5414
rect 11854 5412 11860 5414
rect 11552 5403 11860 5412
rect 22155 5468 22463 5477
rect 22155 5466 22161 5468
rect 22217 5466 22241 5468
rect 22297 5466 22321 5468
rect 22377 5466 22401 5468
rect 22457 5466 22463 5468
rect 22217 5414 22219 5466
rect 22399 5414 22401 5466
rect 22155 5412 22161 5414
rect 22217 5412 22241 5414
rect 22297 5412 22321 5414
rect 22377 5412 22401 5414
rect 22457 5412 22463 5414
rect 22155 5403 22463 5412
rect 6251 4924 6559 4933
rect 6251 4922 6257 4924
rect 6313 4922 6337 4924
rect 6393 4922 6417 4924
rect 6473 4922 6497 4924
rect 6553 4922 6559 4924
rect 6313 4870 6315 4922
rect 6495 4870 6497 4922
rect 6251 4868 6257 4870
rect 6313 4868 6337 4870
rect 6393 4868 6417 4870
rect 6473 4868 6497 4870
rect 6553 4868 6559 4870
rect 6251 4859 6559 4868
rect 16854 4924 17162 4933
rect 16854 4922 16860 4924
rect 16916 4922 16940 4924
rect 16996 4922 17020 4924
rect 17076 4922 17100 4924
rect 17156 4922 17162 4924
rect 16916 4870 16918 4922
rect 17098 4870 17100 4922
rect 16854 4868 16860 4870
rect 16916 4868 16940 4870
rect 16996 4868 17020 4870
rect 17076 4868 17100 4870
rect 17156 4868 17162 4870
rect 16854 4859 17162 4868
rect 23032 4826 23060 5578
rect 23848 5160 23900 5166
rect 23848 5102 23900 5108
rect 23860 4826 23888 5102
rect 25976 4826 26004 5646
rect 27457 4924 27765 4933
rect 27457 4922 27463 4924
rect 27519 4922 27543 4924
rect 27599 4922 27623 4924
rect 27679 4922 27703 4924
rect 27759 4922 27765 4924
rect 27519 4870 27521 4922
rect 27701 4870 27703 4922
rect 27457 4868 27463 4870
rect 27519 4868 27543 4870
rect 27599 4868 27623 4870
rect 27679 4868 27703 4870
rect 27759 4868 27765 4870
rect 27457 4859 27765 4868
rect 28092 4826 28120 7754
rect 28184 7750 28212 9794
rect 28552 8362 28580 9846
rect 28630 9840 28686 10300
rect 28906 9840 28962 10300
rect 29182 9840 29238 10300
rect 29276 9920 29328 9926
rect 29276 9862 29328 9868
rect 28644 8480 28672 9840
rect 28920 9194 28948 9840
rect 28920 9166 29040 9194
rect 29012 8566 29040 9166
rect 29000 8560 29052 8566
rect 29000 8502 29052 8508
rect 28908 8492 28960 8498
rect 28644 8452 28908 8480
rect 28908 8434 28960 8440
rect 29196 8430 29224 9840
rect 29184 8424 29236 8430
rect 29184 8366 29236 8372
rect 28540 8356 28592 8362
rect 28540 8298 28592 8304
rect 28908 8356 28960 8362
rect 28908 8298 28960 8304
rect 28632 8288 28684 8294
rect 28632 8230 28684 8236
rect 28724 8288 28776 8294
rect 28724 8230 28776 8236
rect 28172 7744 28224 7750
rect 28172 7686 28224 7692
rect 28644 7274 28672 8230
rect 28632 7268 28684 7274
rect 28632 7210 28684 7216
rect 28736 6730 28764 8230
rect 28920 7857 28948 8298
rect 29184 8288 29236 8294
rect 29184 8230 29236 8236
rect 28906 7848 28962 7857
rect 28906 7783 28962 7792
rect 29196 7546 29224 8230
rect 29184 7540 29236 7546
rect 29184 7482 29236 7488
rect 28724 6724 28776 6730
rect 28724 6666 28776 6672
rect 23020 4820 23072 4826
rect 23020 4762 23072 4768
rect 23848 4820 23900 4826
rect 23848 4762 23900 4768
rect 25964 4820 26016 4826
rect 25964 4762 26016 4768
rect 28080 4820 28132 4826
rect 28080 4762 28132 4768
rect 21548 4616 21600 4622
rect 21548 4558 21600 4564
rect 22560 4616 22612 4622
rect 22560 4558 22612 4564
rect 22836 4616 22888 4622
rect 22836 4558 22888 4564
rect 23664 4616 23716 4622
rect 23664 4558 23716 4564
rect 25780 4616 25832 4622
rect 25780 4558 25832 4564
rect 27896 4616 27948 4622
rect 27896 4558 27948 4564
rect 11552 4380 11860 4389
rect 11552 4378 11558 4380
rect 11614 4378 11638 4380
rect 11694 4378 11718 4380
rect 11774 4378 11798 4380
rect 11854 4378 11860 4380
rect 11614 4326 11616 4378
rect 11796 4326 11798 4378
rect 11552 4324 11558 4326
rect 11614 4324 11638 4326
rect 11694 4324 11718 4326
rect 11774 4324 11798 4326
rect 11854 4324 11860 4326
rect 11552 4315 11860 4324
rect 21560 4282 21588 4558
rect 22155 4380 22463 4389
rect 22155 4378 22161 4380
rect 22217 4378 22241 4380
rect 22297 4378 22321 4380
rect 22377 4378 22401 4380
rect 22457 4378 22463 4380
rect 22217 4326 22219 4378
rect 22399 4326 22401 4378
rect 22155 4324 22161 4326
rect 22217 4324 22241 4326
rect 22297 4324 22321 4326
rect 22377 4324 22401 4326
rect 22457 4324 22463 4326
rect 22155 4315 22463 4324
rect 22572 4282 22600 4558
rect 22652 4548 22704 4554
rect 22652 4490 22704 4496
rect 21548 4276 21600 4282
rect 21548 4218 21600 4224
rect 22560 4276 22612 4282
rect 22560 4218 22612 4224
rect 20444 4140 20496 4146
rect 20444 4082 20496 4088
rect 22468 4140 22520 4146
rect 22468 4082 22520 4088
rect 7748 4072 7800 4078
rect 7748 4014 7800 4020
rect 5632 4004 5684 4010
rect 5632 3946 5684 3952
rect 3516 2440 3568 2446
rect 3516 2382 3568 2388
rect 1584 1964 1636 1970
rect 1584 1906 1636 1912
rect 1596 1562 1624 1906
rect 3528 1562 3556 2382
rect 1584 1556 1636 1562
rect 1584 1498 1636 1504
rect 3516 1556 3568 1562
rect 3516 1498 3568 1504
rect 5644 1358 5672 3946
rect 6251 3836 6559 3845
rect 6251 3834 6257 3836
rect 6313 3834 6337 3836
rect 6393 3834 6417 3836
rect 6473 3834 6497 3836
rect 6553 3834 6559 3836
rect 6313 3782 6315 3834
rect 6495 3782 6497 3834
rect 6251 3780 6257 3782
rect 6313 3780 6337 3782
rect 6393 3780 6417 3782
rect 6473 3780 6497 3782
rect 6553 3780 6559 3782
rect 6251 3771 6559 3780
rect 6251 2748 6559 2757
rect 6251 2746 6257 2748
rect 6313 2746 6337 2748
rect 6393 2746 6417 2748
rect 6473 2746 6497 2748
rect 6553 2746 6559 2748
rect 6313 2694 6315 2746
rect 6495 2694 6497 2746
rect 6251 2692 6257 2694
rect 6313 2692 6337 2694
rect 6393 2692 6417 2694
rect 6473 2692 6497 2694
rect 6553 2692 6559 2694
rect 6251 2683 6559 2692
rect 6251 1660 6559 1669
rect 6251 1658 6257 1660
rect 6313 1658 6337 1660
rect 6393 1658 6417 1660
rect 6473 1658 6497 1660
rect 6553 1658 6559 1660
rect 6313 1606 6315 1658
rect 6495 1606 6497 1658
rect 6251 1604 6257 1606
rect 6313 1604 6337 1606
rect 6393 1604 6417 1606
rect 6473 1604 6497 1606
rect 6553 1604 6559 1606
rect 6251 1595 6559 1604
rect 1124 1352 1176 1358
rect 1124 1294 1176 1300
rect 3332 1352 3384 1358
rect 3332 1294 3384 1300
rect 5448 1352 5500 1358
rect 5448 1294 5500 1300
rect 5632 1352 5684 1358
rect 5632 1294 5684 1300
rect 7564 1352 7616 1358
rect 7564 1294 7616 1300
rect 1136 160 1164 1294
rect 1122 -300 1178 160
rect 3238 82 3294 160
rect 3344 82 3372 1294
rect 3238 54 3372 82
rect 5354 82 5410 160
rect 5460 82 5488 1294
rect 5354 54 5488 82
rect 7470 82 7526 160
rect 7576 82 7604 1294
rect 7760 1222 7788 4014
rect 19524 3936 19576 3942
rect 19524 3878 19576 3884
rect 16854 3836 17162 3845
rect 16854 3834 16860 3836
rect 16916 3834 16940 3836
rect 16996 3834 17020 3836
rect 17076 3834 17100 3836
rect 17156 3834 17162 3836
rect 16916 3782 16918 3834
rect 17098 3782 17100 3834
rect 16854 3780 16860 3782
rect 16916 3780 16940 3782
rect 16996 3780 17020 3782
rect 17076 3780 17100 3782
rect 17156 3780 17162 3782
rect 16854 3771 17162 3780
rect 19432 3528 19484 3534
rect 19432 3470 19484 3476
rect 19248 3460 19300 3466
rect 19248 3402 19300 3408
rect 11552 3292 11860 3301
rect 11552 3290 11558 3292
rect 11614 3290 11638 3292
rect 11694 3290 11718 3292
rect 11774 3290 11798 3292
rect 11854 3290 11860 3292
rect 11614 3238 11616 3290
rect 11796 3238 11798 3290
rect 11552 3236 11558 3238
rect 11614 3236 11638 3238
rect 11694 3236 11718 3238
rect 11774 3236 11798 3238
rect 11854 3236 11860 3238
rect 11552 3227 11860 3236
rect 18604 3052 18656 3058
rect 18604 2994 18656 3000
rect 16212 2984 16264 2990
rect 16212 2926 16264 2932
rect 11552 2204 11860 2213
rect 11552 2202 11558 2204
rect 11614 2202 11638 2204
rect 11694 2202 11718 2204
rect 11774 2202 11798 2204
rect 11854 2202 11860 2204
rect 11614 2150 11616 2202
rect 11796 2150 11798 2202
rect 11552 2148 11558 2150
rect 11614 2148 11638 2150
rect 11694 2148 11718 2150
rect 11774 2148 11798 2150
rect 11854 2148 11860 2150
rect 11552 2139 11860 2148
rect 9680 1352 9732 1358
rect 9680 1294 9732 1300
rect 11796 1352 11848 1358
rect 14096 1352 14148 1358
rect 11848 1300 11928 1306
rect 11796 1294 11928 1300
rect 14096 1294 14148 1300
rect 16028 1352 16080 1358
rect 16028 1294 16080 1300
rect 7748 1216 7800 1222
rect 7748 1158 7800 1164
rect 7470 54 7604 82
rect 9586 82 9642 160
rect 9692 82 9720 1294
rect 11808 1278 11928 1294
rect 9864 1216 9916 1222
rect 9864 1158 9916 1164
rect 9876 1018 9904 1158
rect 11552 1116 11860 1125
rect 11552 1114 11558 1116
rect 11614 1114 11638 1116
rect 11694 1114 11718 1116
rect 11774 1114 11798 1116
rect 11854 1114 11860 1116
rect 11614 1062 11616 1114
rect 11796 1062 11798 1114
rect 11552 1060 11558 1062
rect 11614 1060 11638 1062
rect 11694 1060 11718 1062
rect 11774 1060 11798 1062
rect 11854 1060 11860 1062
rect 11552 1051 11860 1060
rect 9864 1012 9916 1018
rect 9864 954 9916 960
rect 9586 54 9720 82
rect 11702 82 11758 160
rect 11900 82 11928 1278
rect 11702 54 11928 82
rect 13818 82 13874 160
rect 14108 82 14136 1294
rect 13818 54 14136 82
rect 15934 82 15990 160
rect 16040 82 16068 1294
rect 16224 1222 16252 2926
rect 16854 2748 17162 2757
rect 16854 2746 16860 2748
rect 16916 2746 16940 2748
rect 16996 2746 17020 2748
rect 17076 2746 17100 2748
rect 17156 2746 17162 2748
rect 16916 2694 16918 2746
rect 17098 2694 17100 2746
rect 16854 2692 16860 2694
rect 16916 2692 16940 2694
rect 16996 2692 17020 2694
rect 17076 2692 17100 2694
rect 17156 2692 17162 2694
rect 16854 2683 17162 2692
rect 16854 1660 17162 1669
rect 16854 1658 16860 1660
rect 16916 1658 16940 1660
rect 16996 1658 17020 1660
rect 17076 1658 17100 1660
rect 17156 1658 17162 1660
rect 16916 1606 16918 1658
rect 17098 1606 17100 1658
rect 16854 1604 16860 1606
rect 16916 1604 16940 1606
rect 16996 1604 17020 1606
rect 17076 1604 17100 1606
rect 17156 1604 17162 1606
rect 16854 1595 17162 1604
rect 18144 1352 18196 1358
rect 18420 1352 18472 1358
rect 18144 1294 18196 1300
rect 18248 1312 18420 1340
rect 16212 1216 16264 1222
rect 16212 1158 16264 1164
rect 15934 54 16068 82
rect 18050 82 18106 160
rect 18156 82 18184 1294
rect 18248 1222 18276 1312
rect 18420 1294 18472 1300
rect 18616 1222 18644 2994
rect 18236 1216 18288 1222
rect 18236 1158 18288 1164
rect 18604 1216 18656 1222
rect 18604 1158 18656 1164
rect 19260 1018 19288 3402
rect 19444 3194 19472 3470
rect 19432 3188 19484 3194
rect 19432 3130 19484 3136
rect 19536 1358 19564 3878
rect 19524 1352 19576 1358
rect 19524 1294 19576 1300
rect 20260 1352 20312 1358
rect 20260 1294 20312 1300
rect 19248 1012 19300 1018
rect 19248 954 19300 960
rect 18050 54 18184 82
rect 20166 82 20222 160
rect 20272 82 20300 1294
rect 20456 1222 20484 4082
rect 22480 3738 22508 4082
rect 22664 3942 22692 4490
rect 22848 4078 22876 4558
rect 22836 4072 22888 4078
rect 22836 4014 22888 4020
rect 22652 3936 22704 3942
rect 22652 3878 22704 3884
rect 23676 3738 23704 4558
rect 25792 4282 25820 4558
rect 25780 4276 25832 4282
rect 25780 4218 25832 4224
rect 24768 4140 24820 4146
rect 24768 4082 24820 4088
rect 27068 4140 27120 4146
rect 27068 4082 27120 4088
rect 22468 3732 22520 3738
rect 22468 3674 22520 3680
rect 23664 3732 23716 3738
rect 23664 3674 23716 3680
rect 22008 3528 22060 3534
rect 22008 3470 22060 3476
rect 22836 3528 22888 3534
rect 22836 3470 22888 3476
rect 21272 3460 21324 3466
rect 21272 3402 21324 3408
rect 21284 3194 21312 3402
rect 22020 3194 22048 3470
rect 22155 3292 22463 3301
rect 22155 3290 22161 3292
rect 22217 3290 22241 3292
rect 22297 3290 22321 3292
rect 22377 3290 22401 3292
rect 22457 3290 22463 3292
rect 22217 3238 22219 3290
rect 22399 3238 22401 3290
rect 22155 3236 22161 3238
rect 22217 3236 22241 3238
rect 22297 3236 22321 3238
rect 22377 3236 22401 3238
rect 22457 3236 22463 3238
rect 22155 3227 22463 3236
rect 21272 3188 21324 3194
rect 21272 3130 21324 3136
rect 22008 3188 22060 3194
rect 22008 3130 22060 3136
rect 21364 3052 21416 3058
rect 21364 2994 21416 3000
rect 22652 3052 22704 3058
rect 22652 2994 22704 3000
rect 21376 1358 21404 2994
rect 22664 2650 22692 2994
rect 22848 2774 22876 3470
rect 23386 2952 23442 2961
rect 23386 2887 23388 2896
rect 23440 2887 23442 2896
rect 23388 2858 23440 2864
rect 22756 2746 22876 2774
rect 22652 2644 22704 2650
rect 22652 2586 22704 2592
rect 22155 2204 22463 2213
rect 22155 2202 22161 2204
rect 22217 2202 22241 2204
rect 22297 2202 22321 2204
rect 22377 2202 22401 2204
rect 22457 2202 22463 2204
rect 22217 2150 22219 2202
rect 22399 2150 22401 2202
rect 22155 2148 22161 2150
rect 22217 2148 22241 2150
rect 22297 2148 22321 2150
rect 22377 2148 22401 2150
rect 22457 2148 22463 2150
rect 22155 2139 22463 2148
rect 22756 1358 22784 2746
rect 21364 1352 21416 1358
rect 21364 1294 21416 1300
rect 22376 1352 22428 1358
rect 22744 1352 22796 1358
rect 22428 1312 22600 1340
rect 22376 1294 22428 1300
rect 20444 1216 20496 1222
rect 20444 1158 20496 1164
rect 22155 1116 22463 1125
rect 22155 1114 22161 1116
rect 22217 1114 22241 1116
rect 22297 1114 22321 1116
rect 22377 1114 22401 1116
rect 22457 1114 22463 1116
rect 22217 1062 22219 1114
rect 22399 1062 22401 1114
rect 22155 1060 22161 1062
rect 22217 1060 22241 1062
rect 22297 1060 22321 1062
rect 22377 1060 22401 1062
rect 22457 1060 22463 1062
rect 22155 1051 22463 1060
rect 20166 54 20300 82
rect 22282 82 22338 160
rect 22572 82 22600 1312
rect 22744 1294 22796 1300
rect 24492 1352 24544 1358
rect 24492 1294 24544 1300
rect 22282 54 22600 82
rect 24398 82 24454 160
rect 24504 82 24532 1294
rect 24780 1290 24808 4082
rect 27080 1358 27108 4082
rect 27908 4078 27936 4558
rect 29288 4486 29316 9862
rect 29458 9840 29514 10300
rect 29734 9840 29790 10300
rect 30010 9840 30066 10300
rect 30286 9840 30342 10300
rect 30562 9840 30618 10300
rect 30838 9840 30894 10300
rect 31114 9840 31170 10300
rect 31390 9840 31446 10300
rect 31666 9840 31722 10300
rect 31942 9840 31998 10300
rect 32218 9840 32274 10300
rect 32494 9840 32550 10300
rect 32770 9840 32826 10300
rect 33046 9840 33102 10300
rect 33322 9840 33378 10300
rect 33416 9852 33468 9858
rect 29472 9194 29500 9840
rect 29368 9172 29420 9178
rect 29472 9166 29592 9194
rect 29368 9114 29420 9120
rect 29380 8090 29408 9114
rect 29564 8548 29592 9166
rect 29748 8634 29776 9840
rect 29920 9308 29972 9314
rect 29920 9250 29972 9256
rect 29828 8968 29880 8974
rect 29828 8910 29880 8916
rect 29736 8628 29788 8634
rect 29736 8570 29788 8576
rect 29644 8560 29696 8566
rect 29564 8520 29644 8548
rect 29644 8502 29696 8508
rect 29840 8498 29868 8910
rect 29828 8492 29880 8498
rect 29828 8434 29880 8440
rect 29932 8294 29960 9250
rect 30024 8537 30052 9840
rect 30010 8528 30066 8537
rect 30010 8463 30066 8472
rect 30300 8362 30328 9840
rect 30472 9716 30524 9722
rect 30472 9658 30524 9664
rect 30380 8900 30432 8906
rect 30380 8842 30432 8848
rect 30392 8634 30420 8842
rect 30380 8628 30432 8634
rect 30380 8570 30432 8576
rect 30378 8528 30434 8537
rect 30378 8463 30380 8472
rect 30432 8463 30434 8472
rect 30380 8434 30432 8440
rect 30288 8356 30340 8362
rect 30288 8298 30340 8304
rect 29920 8288 29972 8294
rect 29920 8230 29972 8236
rect 29368 8084 29420 8090
rect 29368 8026 29420 8032
rect 30484 5710 30512 9658
rect 30576 8548 30604 9840
rect 30748 9240 30800 9246
rect 30748 9182 30800 9188
rect 30760 8945 30788 9182
rect 30746 8936 30802 8945
rect 30746 8871 30802 8880
rect 30852 8634 30880 9840
rect 31024 9512 31076 9518
rect 31024 9454 31076 9460
rect 30932 9036 30984 9042
rect 30932 8978 30984 8984
rect 30840 8628 30892 8634
rect 30840 8570 30892 8576
rect 30748 8560 30800 8566
rect 30576 8520 30748 8548
rect 30748 8502 30800 8508
rect 30944 8362 30972 8978
rect 31036 8498 31064 9454
rect 31128 9194 31156 9840
rect 31128 9166 31340 9194
rect 31116 8968 31168 8974
rect 31116 8910 31168 8916
rect 31024 8492 31076 8498
rect 31024 8434 31076 8440
rect 30932 8356 30984 8362
rect 30932 8298 30984 8304
rect 30472 5704 30524 5710
rect 30472 5646 30524 5652
rect 31128 4690 31156 8910
rect 31312 8430 31340 9166
rect 31300 8424 31352 8430
rect 31404 8412 31432 9840
rect 31484 9580 31536 9586
rect 31484 9522 31536 9528
rect 31496 8634 31524 9522
rect 31576 9036 31628 9042
rect 31576 8978 31628 8984
rect 31484 8628 31536 8634
rect 31484 8570 31536 8576
rect 31588 8514 31616 8978
rect 31680 8650 31708 9840
rect 31852 9444 31904 9450
rect 31852 9386 31904 9392
rect 31680 8622 31800 8650
rect 31864 8634 31892 9386
rect 31956 9194 31984 9840
rect 32128 9308 32180 9314
rect 32128 9250 32180 9256
rect 31956 9166 32076 9194
rect 31772 8566 31800 8622
rect 31852 8628 31904 8634
rect 31852 8570 31904 8576
rect 31760 8560 31812 8566
rect 31588 8486 31708 8514
rect 31760 8502 31812 8508
rect 31576 8424 31628 8430
rect 31404 8384 31576 8412
rect 31300 8366 31352 8372
rect 31576 8366 31628 8372
rect 31680 8294 31708 8486
rect 32048 8430 32076 9166
rect 32036 8424 32088 8430
rect 32036 8366 32088 8372
rect 32140 8294 32168 9250
rect 32232 8566 32260 9840
rect 32508 8634 32536 9840
rect 32784 9194 32812 9840
rect 32692 9166 32812 9194
rect 32404 8628 32456 8634
rect 32404 8570 32456 8576
rect 32496 8628 32548 8634
rect 32496 8570 32548 8576
rect 32220 8560 32272 8566
rect 32220 8502 32272 8508
rect 31392 8288 31444 8294
rect 31392 8230 31444 8236
rect 31668 8288 31720 8294
rect 31668 8230 31720 8236
rect 32128 8288 32180 8294
rect 32128 8230 32180 8236
rect 31116 4684 31168 4690
rect 31116 4626 31168 4632
rect 29276 4480 29328 4486
rect 29276 4422 29328 4428
rect 31300 4140 31352 4146
rect 31300 4082 31352 4088
rect 27896 4072 27948 4078
rect 27896 4014 27948 4020
rect 27457 3836 27765 3845
rect 27457 3834 27463 3836
rect 27519 3834 27543 3836
rect 27599 3834 27623 3836
rect 27679 3834 27703 3836
rect 27759 3834 27765 3836
rect 27519 3782 27521 3834
rect 27701 3782 27703 3834
rect 27457 3780 27463 3782
rect 27519 3780 27543 3782
rect 27599 3780 27623 3782
rect 27679 3780 27703 3782
rect 27759 3780 27765 3782
rect 27457 3771 27765 3780
rect 30012 3528 30064 3534
rect 30012 3470 30064 3476
rect 30024 3194 30052 3470
rect 30012 3188 30064 3194
rect 30012 3130 30064 3136
rect 28908 3052 28960 3058
rect 28908 2994 28960 3000
rect 27457 2748 27765 2757
rect 27457 2746 27463 2748
rect 27519 2746 27543 2748
rect 27599 2746 27623 2748
rect 27679 2746 27703 2748
rect 27759 2746 27765 2748
rect 27519 2694 27521 2746
rect 27701 2694 27703 2746
rect 27457 2692 27463 2694
rect 27519 2692 27543 2694
rect 27599 2692 27623 2694
rect 27679 2692 27703 2694
rect 27759 2692 27765 2694
rect 27457 2683 27765 2692
rect 27457 1660 27765 1669
rect 27457 1658 27463 1660
rect 27519 1658 27543 1660
rect 27599 1658 27623 1660
rect 27679 1658 27703 1660
rect 27759 1658 27765 1660
rect 27519 1606 27521 1658
rect 27701 1606 27703 1658
rect 27457 1604 27463 1606
rect 27519 1604 27543 1606
rect 27599 1604 27623 1606
rect 27679 1604 27703 1606
rect 27759 1604 27765 1606
rect 27457 1595 27765 1604
rect 28920 1358 28948 2994
rect 31312 1358 31340 4082
rect 31404 3942 31432 8230
rect 32416 7449 32444 8570
rect 32692 8514 32720 9166
rect 33060 8922 33088 9840
rect 33060 8894 33272 8922
rect 32758 8732 33066 8741
rect 32758 8730 32764 8732
rect 32820 8730 32844 8732
rect 32900 8730 32924 8732
rect 32980 8730 33004 8732
rect 33060 8730 33066 8732
rect 32820 8678 32822 8730
rect 33002 8678 33004 8730
rect 32758 8676 32764 8678
rect 32820 8676 32844 8678
rect 32900 8676 32924 8678
rect 32980 8676 33004 8678
rect 33060 8676 33066 8678
rect 32758 8667 33066 8676
rect 33244 8566 33272 8894
rect 33232 8560 33284 8566
rect 32692 8486 32812 8514
rect 33232 8502 33284 8508
rect 32784 8430 32812 8486
rect 32772 8424 32824 8430
rect 32772 8366 32824 8372
rect 32956 8288 33008 8294
rect 32956 8230 33008 8236
rect 32968 8090 32996 8230
rect 32956 8084 33008 8090
rect 32956 8026 33008 8032
rect 32680 7948 32732 7954
rect 32680 7890 32732 7896
rect 32402 7440 32458 7449
rect 32402 7375 32458 7384
rect 32692 5166 32720 7890
rect 33336 7886 33364 9840
rect 33598 9840 33654 10300
rect 33874 9840 33930 10300
rect 34150 9840 34206 10300
rect 34426 9840 34482 10300
rect 34702 9840 34758 10300
rect 34978 9840 35034 10300
rect 35254 9840 35310 10300
rect 35530 9840 35586 10300
rect 35806 9840 35862 10300
rect 36082 9840 36138 10300
rect 36358 9840 36414 10300
rect 36634 9840 36690 10300
rect 36910 9840 36966 10300
rect 37186 9840 37242 10300
rect 37462 9840 37518 10300
rect 37738 9840 37794 10300
rect 38014 9840 38070 10300
rect 38290 9840 38346 10300
rect 38566 9840 38622 10300
rect 38842 9840 38898 10300
rect 39118 9840 39174 10300
rect 39394 9840 39450 10300
rect 39500 9846 39712 9874
rect 33416 9794 33468 9800
rect 33428 8294 33456 9794
rect 33612 9194 33640 9840
rect 33612 9166 33824 9194
rect 33506 8936 33562 8945
rect 33506 8871 33562 8880
rect 33520 8634 33548 8871
rect 33508 8628 33560 8634
rect 33508 8570 33560 8576
rect 33796 8566 33824 9166
rect 33888 8634 33916 9840
rect 34164 9058 34192 9840
rect 34164 9030 34284 9058
rect 34256 8634 34284 9030
rect 33876 8628 33928 8634
rect 33876 8570 33928 8576
rect 34244 8628 34296 8634
rect 34244 8570 34296 8576
rect 33784 8560 33836 8566
rect 33784 8502 33836 8508
rect 33968 8492 34020 8498
rect 33968 8434 34020 8440
rect 33600 8356 33652 8362
rect 33600 8298 33652 8304
rect 33416 8288 33468 8294
rect 33416 8230 33468 8236
rect 33612 7993 33640 8298
rect 33598 7984 33654 7993
rect 33598 7919 33654 7928
rect 33324 7880 33376 7886
rect 33324 7822 33376 7828
rect 33416 7744 33468 7750
rect 33416 7686 33468 7692
rect 32758 7644 33066 7653
rect 32758 7642 32764 7644
rect 32820 7642 32844 7644
rect 32900 7642 32924 7644
rect 32980 7642 33004 7644
rect 33060 7642 33066 7644
rect 32820 7590 32822 7642
rect 33002 7590 33004 7642
rect 32758 7588 32764 7590
rect 32820 7588 32844 7590
rect 32900 7588 32924 7590
rect 32980 7588 33004 7590
rect 33060 7588 33066 7590
rect 32758 7579 33066 7588
rect 33428 7546 33456 7686
rect 33416 7540 33468 7546
rect 33416 7482 33468 7488
rect 32758 6556 33066 6565
rect 32758 6554 32764 6556
rect 32820 6554 32844 6556
rect 32900 6554 32924 6556
rect 32980 6554 33004 6556
rect 33060 6554 33066 6556
rect 32820 6502 32822 6554
rect 33002 6502 33004 6554
rect 32758 6500 32764 6502
rect 32820 6500 32844 6502
rect 32900 6500 32924 6502
rect 32980 6500 33004 6502
rect 33060 6500 33066 6502
rect 32758 6491 33066 6500
rect 32758 5468 33066 5477
rect 32758 5466 32764 5468
rect 32820 5466 32844 5468
rect 32900 5466 32924 5468
rect 32980 5466 33004 5468
rect 33060 5466 33066 5468
rect 32820 5414 32822 5466
rect 33002 5414 33004 5466
rect 32758 5412 32764 5414
rect 32820 5412 32844 5414
rect 32900 5412 32924 5414
rect 32980 5412 33004 5414
rect 33060 5412 33066 5414
rect 32758 5403 33066 5412
rect 32680 5160 32732 5166
rect 32680 5102 32732 5108
rect 32128 4616 32180 4622
rect 32128 4558 32180 4564
rect 32140 4078 32168 4558
rect 32758 4380 33066 4389
rect 32758 4378 32764 4380
rect 32820 4378 32844 4380
rect 32900 4378 32924 4380
rect 32980 4378 33004 4380
rect 33060 4378 33066 4380
rect 32820 4326 32822 4378
rect 33002 4326 33004 4378
rect 32758 4324 32764 4326
rect 32820 4324 32844 4326
rect 32900 4324 32924 4326
rect 32980 4324 33004 4326
rect 33060 4324 33066 4326
rect 32758 4315 33066 4324
rect 32128 4072 32180 4078
rect 32128 4014 32180 4020
rect 31392 3936 31444 3942
rect 31392 3878 31444 3884
rect 32758 3292 33066 3301
rect 32758 3290 32764 3292
rect 32820 3290 32844 3292
rect 32900 3290 32924 3292
rect 32980 3290 33004 3292
rect 33060 3290 33066 3292
rect 32820 3238 32822 3290
rect 33002 3238 33004 3290
rect 32758 3236 32764 3238
rect 32820 3236 32844 3238
rect 32900 3236 32924 3238
rect 32980 3236 33004 3238
rect 33060 3236 33066 3238
rect 32758 3227 33066 3236
rect 32758 2204 33066 2213
rect 32758 2202 32764 2204
rect 32820 2202 32844 2204
rect 32900 2202 32924 2204
rect 32980 2202 33004 2204
rect 33060 2202 33066 2204
rect 32820 2150 32822 2202
rect 33002 2150 33004 2202
rect 32758 2148 32764 2150
rect 32820 2148 32844 2150
rect 32900 2148 32924 2150
rect 32980 2148 33004 2150
rect 33060 2148 33066 2150
rect 32758 2139 33066 2148
rect 33980 1766 34008 8434
rect 34440 8362 34468 9840
rect 34716 9246 34744 9840
rect 34704 9240 34756 9246
rect 34704 9182 34756 9188
rect 34612 9036 34664 9042
rect 34612 8978 34664 8984
rect 34428 8356 34480 8362
rect 34428 8298 34480 8304
rect 34520 4616 34572 4622
rect 34520 4558 34572 4564
rect 33968 1760 34020 1766
rect 33968 1702 34020 1708
rect 34532 1358 34560 4558
rect 34624 3738 34652 8978
rect 34992 8566 35020 9840
rect 35072 9240 35124 9246
rect 35072 9182 35124 9188
rect 35084 8634 35112 9182
rect 35072 8628 35124 8634
rect 35072 8570 35124 8576
rect 34980 8560 35032 8566
rect 34980 8502 35032 8508
rect 34796 8492 34848 8498
rect 34796 8434 34848 8440
rect 34808 8401 34836 8434
rect 34794 8392 34850 8401
rect 34794 8327 34850 8336
rect 35268 7750 35296 9840
rect 35348 8492 35400 8498
rect 35348 8434 35400 8440
rect 35256 7744 35308 7750
rect 35256 7686 35308 7692
rect 35360 5642 35388 8434
rect 35544 8242 35572 9840
rect 35820 8362 35848 9840
rect 35900 8968 35952 8974
rect 35900 8910 35952 8916
rect 35912 8498 35940 8910
rect 35900 8492 35952 8498
rect 35900 8434 35952 8440
rect 35808 8356 35860 8362
rect 35808 8298 35860 8304
rect 35544 8214 35848 8242
rect 35820 8022 35848 8214
rect 36096 8090 36124 9840
rect 36372 9058 36400 9840
rect 36648 9194 36676 9840
rect 36648 9166 36860 9194
rect 36372 9030 36584 9058
rect 36556 8430 36584 9030
rect 36636 8492 36688 8498
rect 36636 8434 36688 8440
rect 36544 8424 36596 8430
rect 36544 8366 36596 8372
rect 36084 8084 36136 8090
rect 36084 8026 36136 8032
rect 35808 8016 35860 8022
rect 35808 7958 35860 7964
rect 35716 7812 35768 7818
rect 35716 7754 35768 7760
rect 36268 7812 36320 7818
rect 36268 7754 36320 7760
rect 35348 5636 35400 5642
rect 35348 5578 35400 5584
rect 34612 3732 34664 3738
rect 34612 3674 34664 3680
rect 35728 3534 35756 7754
rect 36280 3670 36308 7754
rect 36268 3664 36320 3670
rect 36268 3606 36320 3612
rect 35716 3528 35768 3534
rect 35716 3470 35768 3476
rect 36648 3398 36676 8434
rect 36832 8090 36860 9166
rect 36820 8084 36872 8090
rect 36820 8026 36872 8032
rect 36820 7812 36872 7818
rect 36820 7754 36872 7760
rect 36832 4826 36860 7754
rect 36924 6798 36952 9840
rect 36912 6792 36964 6798
rect 36912 6734 36964 6740
rect 37200 6730 37228 9840
rect 37476 9602 37504 9840
rect 37476 9574 37688 9602
rect 37556 9444 37608 9450
rect 37556 9386 37608 9392
rect 37464 9036 37516 9042
rect 37464 8978 37516 8984
rect 37476 8634 37504 8978
rect 37464 8628 37516 8634
rect 37464 8570 37516 8576
rect 37568 8566 37596 9386
rect 37660 8838 37688 9574
rect 37648 8832 37700 8838
rect 37648 8774 37700 8780
rect 37556 8560 37608 8566
rect 37556 8502 37608 8508
rect 37752 8090 37780 9840
rect 38028 9466 38056 9840
rect 38304 9738 38332 9840
rect 38304 9710 38424 9738
rect 38028 9438 38332 9466
rect 38016 9376 38068 9382
rect 38016 9318 38068 9324
rect 38028 8566 38056 9318
rect 38016 8560 38068 8566
rect 38016 8502 38068 8508
rect 38304 8430 38332 9438
rect 38396 8498 38424 9710
rect 38384 8492 38436 8498
rect 38384 8434 38436 8440
rect 38292 8424 38344 8430
rect 38292 8366 38344 8372
rect 38060 8188 38368 8197
rect 38060 8186 38066 8188
rect 38122 8186 38146 8188
rect 38202 8186 38226 8188
rect 38282 8186 38306 8188
rect 38362 8186 38368 8188
rect 38122 8134 38124 8186
rect 38304 8134 38306 8186
rect 38060 8132 38066 8134
rect 38122 8132 38146 8134
rect 38202 8132 38226 8134
rect 38282 8132 38306 8134
rect 38362 8132 38368 8134
rect 38060 8123 38368 8132
rect 37740 8084 37792 8090
rect 37740 8026 37792 8032
rect 37924 7812 37976 7818
rect 37924 7754 37976 7760
rect 38384 7812 38436 7818
rect 38384 7754 38436 7760
rect 37188 6724 37240 6730
rect 37188 6666 37240 6672
rect 37372 5228 37424 5234
rect 37372 5170 37424 5176
rect 37384 4826 37412 5170
rect 36820 4820 36872 4826
rect 36820 4762 36872 4768
rect 37372 4820 37424 4826
rect 37372 4762 37424 4768
rect 37936 4758 37964 7754
rect 38060 7100 38368 7109
rect 38060 7098 38066 7100
rect 38122 7098 38146 7100
rect 38202 7098 38226 7100
rect 38282 7098 38306 7100
rect 38362 7098 38368 7100
rect 38122 7046 38124 7098
rect 38304 7046 38306 7098
rect 38060 7044 38066 7046
rect 38122 7044 38146 7046
rect 38202 7044 38226 7046
rect 38282 7044 38306 7046
rect 38362 7044 38368 7046
rect 38060 7035 38368 7044
rect 38060 6012 38368 6021
rect 38060 6010 38066 6012
rect 38122 6010 38146 6012
rect 38202 6010 38226 6012
rect 38282 6010 38306 6012
rect 38362 6010 38368 6012
rect 38122 5958 38124 6010
rect 38304 5958 38306 6010
rect 38060 5956 38066 5958
rect 38122 5956 38146 5958
rect 38202 5956 38226 5958
rect 38282 5956 38306 5958
rect 38362 5956 38368 5958
rect 38060 5947 38368 5956
rect 38060 4924 38368 4933
rect 38060 4922 38066 4924
rect 38122 4922 38146 4924
rect 38202 4922 38226 4924
rect 38282 4922 38306 4924
rect 38362 4922 38368 4924
rect 38122 4870 38124 4922
rect 38304 4870 38306 4922
rect 38060 4868 38066 4870
rect 38122 4868 38146 4870
rect 38202 4868 38226 4870
rect 38282 4868 38306 4870
rect 38362 4868 38368 4870
rect 38060 4859 38368 4868
rect 38396 4826 38424 7754
rect 38580 6866 38608 9840
rect 38660 8356 38712 8362
rect 38660 8298 38712 8304
rect 38568 6860 38620 6866
rect 38568 6802 38620 6808
rect 38672 6798 38700 8298
rect 38856 8090 38884 9840
rect 38844 8084 38896 8090
rect 38844 8026 38896 8032
rect 39132 8004 39160 9840
rect 39408 9738 39436 9840
rect 39500 9738 39528 9846
rect 39408 9710 39528 9738
rect 39304 8832 39356 8838
rect 39304 8774 39356 8780
rect 39316 8634 39344 8774
rect 39684 8634 39712 9846
rect 43361 8732 43669 8741
rect 43361 8730 43367 8732
rect 43423 8730 43447 8732
rect 43503 8730 43527 8732
rect 43583 8730 43607 8732
rect 43663 8730 43669 8732
rect 43423 8678 43425 8730
rect 43605 8678 43607 8730
rect 43361 8676 43367 8678
rect 43423 8676 43447 8678
rect 43503 8676 43527 8678
rect 43583 8676 43607 8678
rect 43663 8676 43669 8678
rect 43361 8667 43669 8676
rect 39304 8628 39356 8634
rect 39304 8570 39356 8576
rect 39672 8628 39724 8634
rect 39672 8570 39724 8576
rect 39304 8492 39356 8498
rect 39304 8434 39356 8440
rect 41052 8492 41104 8498
rect 41052 8434 41104 8440
rect 39212 8016 39264 8022
rect 39132 7976 39212 8004
rect 39212 7958 39264 7964
rect 38752 7744 38804 7750
rect 38752 7686 38804 7692
rect 39120 7744 39172 7750
rect 39120 7686 39172 7692
rect 38660 6792 38712 6798
rect 38660 6734 38712 6740
rect 38764 6730 38792 7686
rect 39132 6866 39160 7686
rect 39120 6860 39172 6866
rect 39120 6802 39172 6808
rect 38752 6724 38804 6730
rect 38752 6666 38804 6672
rect 39316 5370 39344 8434
rect 39580 8424 39632 8430
rect 39580 8366 39632 8372
rect 39304 5364 39356 5370
rect 39304 5306 39356 5312
rect 38384 4820 38436 4826
rect 38384 4762 38436 4768
rect 37924 4752 37976 4758
rect 37924 4694 37976 4700
rect 38016 4616 38068 4622
rect 38016 4558 38068 4564
rect 38028 4282 38056 4558
rect 38016 4276 38068 4282
rect 38016 4218 38068 4224
rect 37464 4140 37516 4146
rect 37464 4082 37516 4088
rect 37096 3528 37148 3534
rect 37096 3470 37148 3476
rect 36636 3392 36688 3398
rect 36636 3334 36688 3340
rect 37108 3194 37136 3470
rect 37096 3188 37148 3194
rect 37096 3130 37148 3136
rect 35256 3052 35308 3058
rect 35256 2994 35308 3000
rect 35268 1358 35296 2994
rect 37476 1358 37504 4082
rect 38060 3836 38368 3845
rect 38060 3834 38066 3836
rect 38122 3834 38146 3836
rect 38202 3834 38226 3836
rect 38282 3834 38306 3836
rect 38362 3834 38368 3836
rect 38122 3782 38124 3834
rect 38304 3782 38306 3834
rect 38060 3780 38066 3782
rect 38122 3780 38146 3782
rect 38202 3780 38226 3782
rect 38282 3780 38306 3782
rect 38362 3780 38368 3782
rect 38060 3771 38368 3780
rect 39592 3738 39620 8366
rect 39856 7880 39908 7886
rect 39856 7822 39908 7828
rect 39764 4140 39816 4146
rect 39764 4082 39816 4088
rect 39776 3738 39804 4082
rect 39868 3942 39896 7822
rect 39948 7812 40000 7818
rect 39948 7754 40000 7760
rect 39856 3936 39908 3942
rect 39856 3878 39908 3884
rect 39580 3732 39632 3738
rect 39580 3674 39632 3680
rect 39764 3732 39816 3738
rect 39764 3674 39816 3680
rect 38060 2748 38368 2757
rect 38060 2746 38066 2748
rect 38122 2746 38146 2748
rect 38202 2746 38226 2748
rect 38282 2746 38306 2748
rect 38362 2746 38368 2748
rect 38122 2694 38124 2746
rect 38304 2694 38306 2746
rect 38060 2692 38066 2694
rect 38122 2692 38146 2694
rect 38202 2692 38226 2694
rect 38282 2692 38306 2694
rect 38362 2692 38368 2694
rect 38060 2683 38368 2692
rect 39960 2650 39988 7754
rect 40684 3528 40736 3534
rect 40684 3470 40736 3476
rect 40224 3052 40276 3058
rect 40224 2994 40276 3000
rect 40236 2650 40264 2994
rect 39948 2644 40000 2650
rect 39948 2586 40000 2592
rect 40224 2644 40276 2650
rect 40224 2586 40276 2592
rect 39028 2440 39080 2446
rect 39028 2382 39080 2388
rect 39040 2106 39068 2382
rect 39028 2100 39080 2106
rect 39028 2042 39080 2048
rect 38844 1964 38896 1970
rect 38844 1906 38896 1912
rect 38060 1660 38368 1669
rect 38060 1658 38066 1660
rect 38122 1658 38146 1660
rect 38202 1658 38226 1660
rect 38282 1658 38306 1660
rect 38362 1658 38368 1660
rect 38122 1606 38124 1658
rect 38304 1606 38306 1658
rect 38060 1604 38066 1606
rect 38122 1604 38146 1606
rect 38202 1604 38226 1606
rect 38282 1604 38306 1606
rect 38362 1604 38368 1606
rect 38060 1595 38368 1604
rect 38856 1562 38884 1906
rect 38844 1556 38896 1562
rect 38844 1498 38896 1504
rect 40696 1358 40724 3470
rect 41064 3194 41092 8434
rect 43361 7644 43669 7653
rect 43361 7642 43367 7644
rect 43423 7642 43447 7644
rect 43503 7642 43527 7644
rect 43583 7642 43607 7644
rect 43663 7642 43669 7644
rect 43423 7590 43425 7642
rect 43605 7590 43607 7642
rect 43361 7588 43367 7590
rect 43423 7588 43447 7590
rect 43503 7588 43527 7590
rect 43583 7588 43607 7590
rect 43663 7588 43669 7590
rect 43361 7579 43669 7588
rect 43361 6556 43669 6565
rect 43361 6554 43367 6556
rect 43423 6554 43447 6556
rect 43503 6554 43527 6556
rect 43583 6554 43607 6556
rect 43663 6554 43669 6556
rect 43423 6502 43425 6554
rect 43605 6502 43607 6554
rect 43361 6500 43367 6502
rect 43423 6500 43447 6502
rect 43503 6500 43527 6502
rect 43583 6500 43607 6502
rect 43663 6500 43669 6502
rect 43361 6491 43669 6500
rect 43361 5468 43669 5477
rect 43361 5466 43367 5468
rect 43423 5466 43447 5468
rect 43503 5466 43527 5468
rect 43583 5466 43607 5468
rect 43663 5466 43669 5468
rect 43423 5414 43425 5466
rect 43605 5414 43607 5466
rect 43361 5412 43367 5414
rect 43423 5412 43447 5414
rect 43503 5412 43527 5414
rect 43583 5412 43607 5414
rect 43663 5412 43669 5414
rect 43361 5403 43669 5412
rect 43361 4380 43669 4389
rect 43361 4378 43367 4380
rect 43423 4378 43447 4380
rect 43503 4378 43527 4380
rect 43583 4378 43607 4380
rect 43663 4378 43669 4380
rect 43423 4326 43425 4378
rect 43605 4326 43607 4378
rect 43361 4324 43367 4326
rect 43423 4324 43447 4326
rect 43503 4324 43527 4326
rect 43583 4324 43607 4326
rect 43663 4324 43669 4326
rect 43361 4315 43669 4324
rect 43361 3292 43669 3301
rect 43361 3290 43367 3292
rect 43423 3290 43447 3292
rect 43503 3290 43527 3292
rect 43583 3290 43607 3292
rect 43663 3290 43669 3292
rect 43423 3238 43425 3290
rect 43605 3238 43607 3290
rect 43361 3236 43367 3238
rect 43423 3236 43447 3238
rect 43503 3236 43527 3238
rect 43583 3236 43607 3238
rect 43663 3236 43669 3238
rect 43361 3227 43669 3236
rect 41052 3188 41104 3194
rect 41052 3130 41104 3136
rect 42984 2440 43036 2446
rect 42984 2382 43036 2388
rect 42996 1562 43024 2382
rect 43361 2204 43669 2213
rect 43361 2202 43367 2204
rect 43423 2202 43447 2204
rect 43503 2202 43527 2204
rect 43583 2202 43607 2204
rect 43663 2202 43669 2204
rect 43423 2150 43425 2202
rect 43605 2150 43607 2202
rect 43361 2148 43367 2150
rect 43423 2148 43447 2150
rect 43503 2148 43527 2150
rect 43583 2148 43607 2150
rect 43663 2148 43669 2150
rect 43361 2139 43669 2148
rect 42984 1556 43036 1562
rect 42984 1498 43036 1504
rect 26608 1352 26660 1358
rect 26608 1294 26660 1300
rect 27068 1352 27120 1358
rect 27068 1294 27120 1300
rect 28724 1352 28776 1358
rect 28724 1294 28776 1300
rect 28908 1352 28960 1358
rect 28908 1294 28960 1300
rect 30840 1352 30892 1358
rect 30840 1294 30892 1300
rect 31300 1352 31352 1358
rect 31300 1294 31352 1300
rect 32680 1352 32732 1358
rect 32680 1294 32732 1300
rect 34520 1352 34572 1358
rect 34520 1294 34572 1300
rect 35072 1352 35124 1358
rect 35072 1294 35124 1300
rect 35256 1352 35308 1358
rect 35256 1294 35308 1300
rect 37280 1352 37332 1358
rect 37280 1294 37332 1300
rect 37464 1352 37516 1358
rect 37464 1294 37516 1300
rect 39488 1352 39540 1358
rect 39488 1294 39540 1300
rect 40684 1352 40736 1358
rect 40684 1294 40736 1300
rect 41328 1352 41380 1358
rect 41328 1294 41380 1300
rect 43168 1352 43220 1358
rect 43168 1294 43220 1300
rect 24768 1284 24820 1290
rect 24768 1226 24820 1232
rect 24398 54 24532 82
rect 26514 82 26570 160
rect 26620 82 26648 1294
rect 26514 54 26648 82
rect 28630 82 28686 160
rect 28736 82 28764 1294
rect 28630 54 28764 82
rect 30746 82 30802 160
rect 30852 82 30880 1294
rect 30746 54 30880 82
rect 32692 82 32720 1294
rect 32758 1116 33066 1125
rect 32758 1114 32764 1116
rect 32820 1114 32844 1116
rect 32900 1114 32924 1116
rect 32980 1114 33004 1116
rect 33060 1114 33066 1116
rect 32820 1062 32822 1114
rect 33002 1062 33004 1114
rect 32758 1060 32764 1062
rect 32820 1060 32844 1062
rect 32900 1060 32924 1062
rect 32980 1060 33004 1062
rect 33060 1060 33066 1062
rect 32758 1051 33066 1060
rect 32862 82 32918 160
rect 32692 54 32918 82
rect 3238 -300 3294 54
rect 5354 -300 5410 54
rect 7470 -300 7526 54
rect 9586 -300 9642 54
rect 11702 -300 11758 54
rect 13818 -300 13874 54
rect 15934 -300 15990 54
rect 18050 -300 18106 54
rect 20166 -300 20222 54
rect 22282 -300 22338 54
rect 24398 -300 24454 54
rect 26514 -300 26570 54
rect 28630 -300 28686 54
rect 30746 -300 30802 54
rect 32862 -300 32918 54
rect 34978 82 35034 160
rect 35084 82 35112 1294
rect 37292 762 37320 1294
rect 37108 734 37320 762
rect 37108 160 37136 734
rect 34978 54 35112 82
rect 34978 -300 35034 54
rect 37094 -300 37150 160
rect 39210 82 39266 160
rect 39500 82 39528 1294
rect 41340 160 41368 1294
rect 39210 54 39528 82
rect 39210 -300 39266 54
rect 41326 -300 41382 160
rect 43180 82 43208 1294
rect 43361 1116 43669 1125
rect 43361 1114 43367 1116
rect 43423 1114 43447 1116
rect 43503 1114 43527 1116
rect 43583 1114 43607 1116
rect 43663 1114 43669 1116
rect 43423 1062 43425 1114
rect 43605 1062 43607 1114
rect 43361 1060 43367 1062
rect 43423 1060 43447 1062
rect 43503 1060 43527 1062
rect 43583 1060 43607 1062
rect 43663 1060 43669 1062
rect 43361 1051 43669 1060
rect 43442 82 43498 160
rect 43180 54 43498 82
rect 43442 -300 43498 54
<< via2 >>
rect 6257 8186 6313 8188
rect 6337 8186 6393 8188
rect 6417 8186 6473 8188
rect 6497 8186 6553 8188
rect 6257 8134 6303 8186
rect 6303 8134 6313 8186
rect 6337 8134 6367 8186
rect 6367 8134 6379 8186
rect 6379 8134 6393 8186
rect 6417 8134 6431 8186
rect 6431 8134 6443 8186
rect 6443 8134 6473 8186
rect 6497 8134 6507 8186
rect 6507 8134 6553 8186
rect 6257 8132 6313 8134
rect 6337 8132 6393 8134
rect 6417 8132 6473 8134
rect 6497 8132 6553 8134
rect 6257 7098 6313 7100
rect 6337 7098 6393 7100
rect 6417 7098 6473 7100
rect 6497 7098 6553 7100
rect 6257 7046 6303 7098
rect 6303 7046 6313 7098
rect 6337 7046 6367 7098
rect 6367 7046 6379 7098
rect 6379 7046 6393 7098
rect 6417 7046 6431 7098
rect 6431 7046 6443 7098
rect 6443 7046 6473 7098
rect 6497 7046 6507 7098
rect 6507 7046 6553 7098
rect 6257 7044 6313 7046
rect 6337 7044 6393 7046
rect 6417 7044 6473 7046
rect 6497 7044 6553 7046
rect 6826 6296 6882 6352
rect 11558 8730 11614 8732
rect 11638 8730 11694 8732
rect 11718 8730 11774 8732
rect 11798 8730 11854 8732
rect 11558 8678 11604 8730
rect 11604 8678 11614 8730
rect 11638 8678 11668 8730
rect 11668 8678 11680 8730
rect 11680 8678 11694 8730
rect 11718 8678 11732 8730
rect 11732 8678 11744 8730
rect 11744 8678 11774 8730
rect 11798 8678 11808 8730
rect 11808 8678 11854 8730
rect 11558 8676 11614 8678
rect 11638 8676 11694 8678
rect 11718 8676 11774 8678
rect 11798 8676 11854 8678
rect 11886 7812 11942 7848
rect 13726 7928 13782 7984
rect 11886 7792 11888 7812
rect 11888 7792 11940 7812
rect 11940 7792 11942 7812
rect 11558 7642 11614 7644
rect 11638 7642 11694 7644
rect 11718 7642 11774 7644
rect 11798 7642 11854 7644
rect 11558 7590 11604 7642
rect 11604 7590 11614 7642
rect 11638 7590 11668 7642
rect 11668 7590 11680 7642
rect 11680 7590 11694 7642
rect 11718 7590 11732 7642
rect 11732 7590 11744 7642
rect 11744 7590 11774 7642
rect 11798 7590 11808 7642
rect 11808 7590 11854 7642
rect 11558 7588 11614 7590
rect 11638 7588 11694 7590
rect 11718 7588 11774 7590
rect 11798 7588 11854 7590
rect 12898 7520 12954 7576
rect 13818 6976 13874 7032
rect 11978 6840 12034 6896
rect 11558 6554 11614 6556
rect 11638 6554 11694 6556
rect 11718 6554 11774 6556
rect 11798 6554 11854 6556
rect 11558 6502 11604 6554
rect 11604 6502 11614 6554
rect 11638 6502 11668 6554
rect 11668 6502 11680 6554
rect 11680 6502 11694 6554
rect 11718 6502 11732 6554
rect 11732 6502 11744 6554
rect 11744 6502 11774 6554
rect 11798 6502 11808 6554
rect 11808 6502 11854 6554
rect 11558 6500 11614 6502
rect 11638 6500 11694 6502
rect 11718 6500 11774 6502
rect 11798 6500 11854 6502
rect 7194 6160 7250 6216
rect 6257 6010 6313 6012
rect 6337 6010 6393 6012
rect 6417 6010 6473 6012
rect 6497 6010 6553 6012
rect 6257 5958 6303 6010
rect 6303 5958 6313 6010
rect 6337 5958 6367 6010
rect 6367 5958 6379 6010
rect 6379 5958 6393 6010
rect 6417 5958 6431 6010
rect 6431 5958 6443 6010
rect 6443 5958 6473 6010
rect 6497 5958 6507 6010
rect 6507 5958 6553 6010
rect 6257 5956 6313 5958
rect 6337 5956 6393 5958
rect 6417 5956 6473 5958
rect 6497 5956 6553 5958
rect 14646 8608 14702 8664
rect 14278 6704 14334 6760
rect 16946 8472 17002 8528
rect 16854 8336 16910 8392
rect 16860 8186 16916 8188
rect 16940 8186 16996 8188
rect 17020 8186 17076 8188
rect 17100 8186 17156 8188
rect 16860 8134 16906 8186
rect 16906 8134 16916 8186
rect 16940 8134 16970 8186
rect 16970 8134 16982 8186
rect 16982 8134 16996 8186
rect 17020 8134 17034 8186
rect 17034 8134 17046 8186
rect 17046 8134 17076 8186
rect 17100 8134 17110 8186
rect 17110 8134 17156 8186
rect 16860 8132 16916 8134
rect 16940 8132 16996 8134
rect 17020 8132 17076 8134
rect 17100 8132 17156 8134
rect 17682 9288 17738 9344
rect 16946 7656 17002 7712
rect 16762 7384 16818 7440
rect 16762 7284 16764 7304
rect 16764 7284 16816 7304
rect 16816 7284 16818 7304
rect 16762 7248 16818 7284
rect 17590 8084 17646 8120
rect 17590 8064 17592 8084
rect 17592 8064 17644 8084
rect 17644 8064 17646 8084
rect 17314 7112 17370 7168
rect 16860 7098 16916 7100
rect 16940 7098 16996 7100
rect 17020 7098 17076 7100
rect 17100 7098 17156 7100
rect 16860 7046 16906 7098
rect 16906 7046 16916 7098
rect 16940 7046 16970 7098
rect 16970 7046 16982 7098
rect 16982 7046 16996 7098
rect 17020 7046 17034 7098
rect 17034 7046 17046 7098
rect 17046 7046 17076 7098
rect 17100 7046 17110 7098
rect 17110 7046 17156 7098
rect 16860 7044 16916 7046
rect 16940 7044 16996 7046
rect 17020 7044 17076 7046
rect 17100 7044 17156 7046
rect 16670 6976 16726 7032
rect 17314 6976 17370 7032
rect 18786 8608 18842 8664
rect 18970 9016 19026 9072
rect 19614 9832 19670 9888
rect 19246 9016 19302 9072
rect 19338 8744 19394 8800
rect 19614 8744 19670 8800
rect 19706 8608 19762 8664
rect 22098 9852 22154 9888
rect 19062 8336 19118 8392
rect 19154 7656 19210 7712
rect 19338 8372 19340 8392
rect 19340 8372 19392 8392
rect 19392 8372 19394 8392
rect 19338 8336 19394 8372
rect 19430 7928 19486 7984
rect 19338 7656 19394 7712
rect 19430 7384 19486 7440
rect 19614 7384 19670 7440
rect 20442 7964 20444 7984
rect 20444 7964 20496 7984
rect 20496 7964 20498 7984
rect 20442 7928 20498 7964
rect 19982 7656 20038 7712
rect 20994 9580 21050 9616
rect 20994 9560 20996 9580
rect 20996 9560 21048 9580
rect 21048 9560 21050 9580
rect 21638 9424 21694 9480
rect 21638 8880 21694 8936
rect 21638 8472 21694 8528
rect 21822 9288 21878 9344
rect 21822 9172 21878 9208
rect 21822 9152 21824 9172
rect 21824 9152 21876 9172
rect 21876 9152 21878 9172
rect 21362 7928 21418 7984
rect 22098 9832 22100 9852
rect 22100 9832 22152 9852
rect 22152 9832 22154 9852
rect 22190 9560 22246 9616
rect 22190 9052 22192 9072
rect 22192 9052 22244 9072
rect 22244 9052 22246 9072
rect 22190 9016 22246 9052
rect 22161 8730 22217 8732
rect 22241 8730 22297 8732
rect 22321 8730 22377 8732
rect 22401 8730 22457 8732
rect 22161 8678 22207 8730
rect 22207 8678 22217 8730
rect 22241 8678 22271 8730
rect 22271 8678 22283 8730
rect 22283 8678 22297 8730
rect 22321 8678 22335 8730
rect 22335 8678 22347 8730
rect 22347 8678 22377 8730
rect 22401 8678 22411 8730
rect 22411 8678 22457 8730
rect 22161 8676 22217 8678
rect 22241 8676 22297 8678
rect 22321 8676 22377 8678
rect 22401 8676 22457 8678
rect 21178 7268 21234 7304
rect 21178 7248 21180 7268
rect 21180 7248 21232 7268
rect 21232 7248 21234 7268
rect 21362 7112 21418 7168
rect 22282 7792 22338 7848
rect 22742 9152 22798 9208
rect 22650 8336 22706 8392
rect 22161 7642 22217 7644
rect 22241 7642 22297 7644
rect 22321 7642 22377 7644
rect 22401 7642 22457 7644
rect 22161 7590 22207 7642
rect 22207 7590 22217 7642
rect 22241 7590 22271 7642
rect 22271 7590 22283 7642
rect 22283 7590 22297 7642
rect 22321 7590 22335 7642
rect 22335 7590 22347 7642
rect 22347 7590 22377 7642
rect 22401 7590 22411 7642
rect 22411 7590 22457 7642
rect 22161 7588 22217 7590
rect 22241 7588 22297 7590
rect 22321 7588 22377 7590
rect 22401 7588 22457 7590
rect 23202 9696 23258 9752
rect 22558 6704 22614 6760
rect 22161 6554 22217 6556
rect 22241 6554 22297 6556
rect 22321 6554 22377 6556
rect 22401 6554 22457 6556
rect 22161 6502 22207 6554
rect 22207 6502 22217 6554
rect 22241 6502 22271 6554
rect 22271 6502 22283 6554
rect 22283 6502 22297 6554
rect 22321 6502 22335 6554
rect 22335 6502 22347 6554
rect 22347 6502 22377 6554
rect 22401 6502 22411 6554
rect 22411 6502 22457 6554
rect 22161 6500 22217 6502
rect 22241 6500 22297 6502
rect 22321 6500 22377 6502
rect 22401 6500 22457 6502
rect 16860 6010 16916 6012
rect 16940 6010 16996 6012
rect 17020 6010 17076 6012
rect 17100 6010 17156 6012
rect 16860 5958 16906 6010
rect 16906 5958 16916 6010
rect 16940 5958 16970 6010
rect 16970 5958 16982 6010
rect 16982 5958 16996 6010
rect 17020 5958 17034 6010
rect 17034 5958 17046 6010
rect 17046 5958 17076 6010
rect 17100 5958 17110 6010
rect 17110 5958 17156 6010
rect 16860 5956 16916 5958
rect 16940 5956 16996 5958
rect 17020 5956 17076 5958
rect 17100 5956 17156 5958
rect 23294 8880 23350 8936
rect 25686 9424 25742 9480
rect 24950 8084 25006 8120
rect 24950 8064 24952 8084
rect 24952 8064 25004 8084
rect 25004 8064 25006 8084
rect 24766 7828 24768 7848
rect 24768 7828 24820 7848
rect 24820 7828 24822 7848
rect 24766 7792 24822 7828
rect 23938 6976 23994 7032
rect 23386 6840 23442 6896
rect 25594 8200 25650 8256
rect 27250 8356 27306 8392
rect 27250 8336 27252 8356
rect 27252 8336 27304 8356
rect 27304 8336 27306 8356
rect 27463 8186 27519 8188
rect 27543 8186 27599 8188
rect 27623 8186 27679 8188
rect 27703 8186 27759 8188
rect 27463 8134 27509 8186
rect 27509 8134 27519 8186
rect 27543 8134 27573 8186
rect 27573 8134 27585 8186
rect 27585 8134 27599 8186
rect 27623 8134 27637 8186
rect 27637 8134 27649 8186
rect 27649 8134 27679 8186
rect 27703 8134 27713 8186
rect 27713 8134 27759 8186
rect 27463 8132 27519 8134
rect 27543 8132 27599 8134
rect 27623 8132 27679 8134
rect 27703 8132 27759 8134
rect 27434 7248 27490 7304
rect 27463 7098 27519 7100
rect 27543 7098 27599 7100
rect 27623 7098 27679 7100
rect 27703 7098 27759 7100
rect 27463 7046 27509 7098
rect 27509 7046 27519 7098
rect 27543 7046 27573 7098
rect 27573 7046 27585 7098
rect 27585 7046 27599 7098
rect 27623 7046 27637 7098
rect 27637 7046 27649 7098
rect 27649 7046 27679 7098
rect 27703 7046 27713 7098
rect 27713 7046 27759 7098
rect 27463 7044 27519 7046
rect 27543 7044 27599 7046
rect 27623 7044 27679 7046
rect 27703 7044 27759 7046
rect 24674 6296 24730 6352
rect 24398 6160 24454 6216
rect 27463 6010 27519 6012
rect 27543 6010 27599 6012
rect 27623 6010 27679 6012
rect 27703 6010 27759 6012
rect 27463 5958 27509 6010
rect 27509 5958 27519 6010
rect 27543 5958 27573 6010
rect 27573 5958 27585 6010
rect 27585 5958 27599 6010
rect 27623 5958 27637 6010
rect 27637 5958 27649 6010
rect 27649 5958 27679 6010
rect 27703 5958 27713 6010
rect 27713 5958 27759 6010
rect 27463 5956 27519 5958
rect 27543 5956 27599 5958
rect 27623 5956 27679 5958
rect 27703 5956 27759 5958
rect 12346 5752 12402 5808
rect 22834 5752 22890 5808
rect 11558 5466 11614 5468
rect 11638 5466 11694 5468
rect 11718 5466 11774 5468
rect 11798 5466 11854 5468
rect 11558 5414 11604 5466
rect 11604 5414 11614 5466
rect 11638 5414 11668 5466
rect 11668 5414 11680 5466
rect 11680 5414 11694 5466
rect 11718 5414 11732 5466
rect 11732 5414 11744 5466
rect 11744 5414 11774 5466
rect 11798 5414 11808 5466
rect 11808 5414 11854 5466
rect 11558 5412 11614 5414
rect 11638 5412 11694 5414
rect 11718 5412 11774 5414
rect 11798 5412 11854 5414
rect 22161 5466 22217 5468
rect 22241 5466 22297 5468
rect 22321 5466 22377 5468
rect 22401 5466 22457 5468
rect 22161 5414 22207 5466
rect 22207 5414 22217 5466
rect 22241 5414 22271 5466
rect 22271 5414 22283 5466
rect 22283 5414 22297 5466
rect 22321 5414 22335 5466
rect 22335 5414 22347 5466
rect 22347 5414 22377 5466
rect 22401 5414 22411 5466
rect 22411 5414 22457 5466
rect 22161 5412 22217 5414
rect 22241 5412 22297 5414
rect 22321 5412 22377 5414
rect 22401 5412 22457 5414
rect 6257 4922 6313 4924
rect 6337 4922 6393 4924
rect 6417 4922 6473 4924
rect 6497 4922 6553 4924
rect 6257 4870 6303 4922
rect 6303 4870 6313 4922
rect 6337 4870 6367 4922
rect 6367 4870 6379 4922
rect 6379 4870 6393 4922
rect 6417 4870 6431 4922
rect 6431 4870 6443 4922
rect 6443 4870 6473 4922
rect 6497 4870 6507 4922
rect 6507 4870 6553 4922
rect 6257 4868 6313 4870
rect 6337 4868 6393 4870
rect 6417 4868 6473 4870
rect 6497 4868 6553 4870
rect 16860 4922 16916 4924
rect 16940 4922 16996 4924
rect 17020 4922 17076 4924
rect 17100 4922 17156 4924
rect 16860 4870 16906 4922
rect 16906 4870 16916 4922
rect 16940 4870 16970 4922
rect 16970 4870 16982 4922
rect 16982 4870 16996 4922
rect 17020 4870 17034 4922
rect 17034 4870 17046 4922
rect 17046 4870 17076 4922
rect 17100 4870 17110 4922
rect 17110 4870 17156 4922
rect 16860 4868 16916 4870
rect 16940 4868 16996 4870
rect 17020 4868 17076 4870
rect 17100 4868 17156 4870
rect 27463 4922 27519 4924
rect 27543 4922 27599 4924
rect 27623 4922 27679 4924
rect 27703 4922 27759 4924
rect 27463 4870 27509 4922
rect 27509 4870 27519 4922
rect 27543 4870 27573 4922
rect 27573 4870 27585 4922
rect 27585 4870 27599 4922
rect 27623 4870 27637 4922
rect 27637 4870 27649 4922
rect 27649 4870 27679 4922
rect 27703 4870 27713 4922
rect 27713 4870 27759 4922
rect 27463 4868 27519 4870
rect 27543 4868 27599 4870
rect 27623 4868 27679 4870
rect 27703 4868 27759 4870
rect 28906 7792 28962 7848
rect 11558 4378 11614 4380
rect 11638 4378 11694 4380
rect 11718 4378 11774 4380
rect 11798 4378 11854 4380
rect 11558 4326 11604 4378
rect 11604 4326 11614 4378
rect 11638 4326 11668 4378
rect 11668 4326 11680 4378
rect 11680 4326 11694 4378
rect 11718 4326 11732 4378
rect 11732 4326 11744 4378
rect 11744 4326 11774 4378
rect 11798 4326 11808 4378
rect 11808 4326 11854 4378
rect 11558 4324 11614 4326
rect 11638 4324 11694 4326
rect 11718 4324 11774 4326
rect 11798 4324 11854 4326
rect 22161 4378 22217 4380
rect 22241 4378 22297 4380
rect 22321 4378 22377 4380
rect 22401 4378 22457 4380
rect 22161 4326 22207 4378
rect 22207 4326 22217 4378
rect 22241 4326 22271 4378
rect 22271 4326 22283 4378
rect 22283 4326 22297 4378
rect 22321 4326 22335 4378
rect 22335 4326 22347 4378
rect 22347 4326 22377 4378
rect 22401 4326 22411 4378
rect 22411 4326 22457 4378
rect 22161 4324 22217 4326
rect 22241 4324 22297 4326
rect 22321 4324 22377 4326
rect 22401 4324 22457 4326
rect 6257 3834 6313 3836
rect 6337 3834 6393 3836
rect 6417 3834 6473 3836
rect 6497 3834 6553 3836
rect 6257 3782 6303 3834
rect 6303 3782 6313 3834
rect 6337 3782 6367 3834
rect 6367 3782 6379 3834
rect 6379 3782 6393 3834
rect 6417 3782 6431 3834
rect 6431 3782 6443 3834
rect 6443 3782 6473 3834
rect 6497 3782 6507 3834
rect 6507 3782 6553 3834
rect 6257 3780 6313 3782
rect 6337 3780 6393 3782
rect 6417 3780 6473 3782
rect 6497 3780 6553 3782
rect 6257 2746 6313 2748
rect 6337 2746 6393 2748
rect 6417 2746 6473 2748
rect 6497 2746 6553 2748
rect 6257 2694 6303 2746
rect 6303 2694 6313 2746
rect 6337 2694 6367 2746
rect 6367 2694 6379 2746
rect 6379 2694 6393 2746
rect 6417 2694 6431 2746
rect 6431 2694 6443 2746
rect 6443 2694 6473 2746
rect 6497 2694 6507 2746
rect 6507 2694 6553 2746
rect 6257 2692 6313 2694
rect 6337 2692 6393 2694
rect 6417 2692 6473 2694
rect 6497 2692 6553 2694
rect 6257 1658 6313 1660
rect 6337 1658 6393 1660
rect 6417 1658 6473 1660
rect 6497 1658 6553 1660
rect 6257 1606 6303 1658
rect 6303 1606 6313 1658
rect 6337 1606 6367 1658
rect 6367 1606 6379 1658
rect 6379 1606 6393 1658
rect 6417 1606 6431 1658
rect 6431 1606 6443 1658
rect 6443 1606 6473 1658
rect 6497 1606 6507 1658
rect 6507 1606 6553 1658
rect 6257 1604 6313 1606
rect 6337 1604 6393 1606
rect 6417 1604 6473 1606
rect 6497 1604 6553 1606
rect 16860 3834 16916 3836
rect 16940 3834 16996 3836
rect 17020 3834 17076 3836
rect 17100 3834 17156 3836
rect 16860 3782 16906 3834
rect 16906 3782 16916 3834
rect 16940 3782 16970 3834
rect 16970 3782 16982 3834
rect 16982 3782 16996 3834
rect 17020 3782 17034 3834
rect 17034 3782 17046 3834
rect 17046 3782 17076 3834
rect 17100 3782 17110 3834
rect 17110 3782 17156 3834
rect 16860 3780 16916 3782
rect 16940 3780 16996 3782
rect 17020 3780 17076 3782
rect 17100 3780 17156 3782
rect 11558 3290 11614 3292
rect 11638 3290 11694 3292
rect 11718 3290 11774 3292
rect 11798 3290 11854 3292
rect 11558 3238 11604 3290
rect 11604 3238 11614 3290
rect 11638 3238 11668 3290
rect 11668 3238 11680 3290
rect 11680 3238 11694 3290
rect 11718 3238 11732 3290
rect 11732 3238 11744 3290
rect 11744 3238 11774 3290
rect 11798 3238 11808 3290
rect 11808 3238 11854 3290
rect 11558 3236 11614 3238
rect 11638 3236 11694 3238
rect 11718 3236 11774 3238
rect 11798 3236 11854 3238
rect 11558 2202 11614 2204
rect 11638 2202 11694 2204
rect 11718 2202 11774 2204
rect 11798 2202 11854 2204
rect 11558 2150 11604 2202
rect 11604 2150 11614 2202
rect 11638 2150 11668 2202
rect 11668 2150 11680 2202
rect 11680 2150 11694 2202
rect 11718 2150 11732 2202
rect 11732 2150 11744 2202
rect 11744 2150 11774 2202
rect 11798 2150 11808 2202
rect 11808 2150 11854 2202
rect 11558 2148 11614 2150
rect 11638 2148 11694 2150
rect 11718 2148 11774 2150
rect 11798 2148 11854 2150
rect 11558 1114 11614 1116
rect 11638 1114 11694 1116
rect 11718 1114 11774 1116
rect 11798 1114 11854 1116
rect 11558 1062 11604 1114
rect 11604 1062 11614 1114
rect 11638 1062 11668 1114
rect 11668 1062 11680 1114
rect 11680 1062 11694 1114
rect 11718 1062 11732 1114
rect 11732 1062 11744 1114
rect 11744 1062 11774 1114
rect 11798 1062 11808 1114
rect 11808 1062 11854 1114
rect 11558 1060 11614 1062
rect 11638 1060 11694 1062
rect 11718 1060 11774 1062
rect 11798 1060 11854 1062
rect 16860 2746 16916 2748
rect 16940 2746 16996 2748
rect 17020 2746 17076 2748
rect 17100 2746 17156 2748
rect 16860 2694 16906 2746
rect 16906 2694 16916 2746
rect 16940 2694 16970 2746
rect 16970 2694 16982 2746
rect 16982 2694 16996 2746
rect 17020 2694 17034 2746
rect 17034 2694 17046 2746
rect 17046 2694 17076 2746
rect 17100 2694 17110 2746
rect 17110 2694 17156 2746
rect 16860 2692 16916 2694
rect 16940 2692 16996 2694
rect 17020 2692 17076 2694
rect 17100 2692 17156 2694
rect 16860 1658 16916 1660
rect 16940 1658 16996 1660
rect 17020 1658 17076 1660
rect 17100 1658 17156 1660
rect 16860 1606 16906 1658
rect 16906 1606 16916 1658
rect 16940 1606 16970 1658
rect 16970 1606 16982 1658
rect 16982 1606 16996 1658
rect 17020 1606 17034 1658
rect 17034 1606 17046 1658
rect 17046 1606 17076 1658
rect 17100 1606 17110 1658
rect 17110 1606 17156 1658
rect 16860 1604 16916 1606
rect 16940 1604 16996 1606
rect 17020 1604 17076 1606
rect 17100 1604 17156 1606
rect 22161 3290 22217 3292
rect 22241 3290 22297 3292
rect 22321 3290 22377 3292
rect 22401 3290 22457 3292
rect 22161 3238 22207 3290
rect 22207 3238 22217 3290
rect 22241 3238 22271 3290
rect 22271 3238 22283 3290
rect 22283 3238 22297 3290
rect 22321 3238 22335 3290
rect 22335 3238 22347 3290
rect 22347 3238 22377 3290
rect 22401 3238 22411 3290
rect 22411 3238 22457 3290
rect 22161 3236 22217 3238
rect 22241 3236 22297 3238
rect 22321 3236 22377 3238
rect 22401 3236 22457 3238
rect 23386 2916 23442 2952
rect 23386 2896 23388 2916
rect 23388 2896 23440 2916
rect 23440 2896 23442 2916
rect 22161 2202 22217 2204
rect 22241 2202 22297 2204
rect 22321 2202 22377 2204
rect 22401 2202 22457 2204
rect 22161 2150 22207 2202
rect 22207 2150 22217 2202
rect 22241 2150 22271 2202
rect 22271 2150 22283 2202
rect 22283 2150 22297 2202
rect 22321 2150 22335 2202
rect 22335 2150 22347 2202
rect 22347 2150 22377 2202
rect 22401 2150 22411 2202
rect 22411 2150 22457 2202
rect 22161 2148 22217 2150
rect 22241 2148 22297 2150
rect 22321 2148 22377 2150
rect 22401 2148 22457 2150
rect 22161 1114 22217 1116
rect 22241 1114 22297 1116
rect 22321 1114 22377 1116
rect 22401 1114 22457 1116
rect 22161 1062 22207 1114
rect 22207 1062 22217 1114
rect 22241 1062 22271 1114
rect 22271 1062 22283 1114
rect 22283 1062 22297 1114
rect 22321 1062 22335 1114
rect 22335 1062 22347 1114
rect 22347 1062 22377 1114
rect 22401 1062 22411 1114
rect 22411 1062 22457 1114
rect 22161 1060 22217 1062
rect 22241 1060 22297 1062
rect 22321 1060 22377 1062
rect 22401 1060 22457 1062
rect 30010 8472 30066 8528
rect 30378 8492 30434 8528
rect 30378 8472 30380 8492
rect 30380 8472 30432 8492
rect 30432 8472 30434 8492
rect 30746 8880 30802 8936
rect 27463 3834 27519 3836
rect 27543 3834 27599 3836
rect 27623 3834 27679 3836
rect 27703 3834 27759 3836
rect 27463 3782 27509 3834
rect 27509 3782 27519 3834
rect 27543 3782 27573 3834
rect 27573 3782 27585 3834
rect 27585 3782 27599 3834
rect 27623 3782 27637 3834
rect 27637 3782 27649 3834
rect 27649 3782 27679 3834
rect 27703 3782 27713 3834
rect 27713 3782 27759 3834
rect 27463 3780 27519 3782
rect 27543 3780 27599 3782
rect 27623 3780 27679 3782
rect 27703 3780 27759 3782
rect 27463 2746 27519 2748
rect 27543 2746 27599 2748
rect 27623 2746 27679 2748
rect 27703 2746 27759 2748
rect 27463 2694 27509 2746
rect 27509 2694 27519 2746
rect 27543 2694 27573 2746
rect 27573 2694 27585 2746
rect 27585 2694 27599 2746
rect 27623 2694 27637 2746
rect 27637 2694 27649 2746
rect 27649 2694 27679 2746
rect 27703 2694 27713 2746
rect 27713 2694 27759 2746
rect 27463 2692 27519 2694
rect 27543 2692 27599 2694
rect 27623 2692 27679 2694
rect 27703 2692 27759 2694
rect 27463 1658 27519 1660
rect 27543 1658 27599 1660
rect 27623 1658 27679 1660
rect 27703 1658 27759 1660
rect 27463 1606 27509 1658
rect 27509 1606 27519 1658
rect 27543 1606 27573 1658
rect 27573 1606 27585 1658
rect 27585 1606 27599 1658
rect 27623 1606 27637 1658
rect 27637 1606 27649 1658
rect 27649 1606 27679 1658
rect 27703 1606 27713 1658
rect 27713 1606 27759 1658
rect 27463 1604 27519 1606
rect 27543 1604 27599 1606
rect 27623 1604 27679 1606
rect 27703 1604 27759 1606
rect 32764 8730 32820 8732
rect 32844 8730 32900 8732
rect 32924 8730 32980 8732
rect 33004 8730 33060 8732
rect 32764 8678 32810 8730
rect 32810 8678 32820 8730
rect 32844 8678 32874 8730
rect 32874 8678 32886 8730
rect 32886 8678 32900 8730
rect 32924 8678 32938 8730
rect 32938 8678 32950 8730
rect 32950 8678 32980 8730
rect 33004 8678 33014 8730
rect 33014 8678 33060 8730
rect 32764 8676 32820 8678
rect 32844 8676 32900 8678
rect 32924 8676 32980 8678
rect 33004 8676 33060 8678
rect 32402 7384 32458 7440
rect 33506 8880 33562 8936
rect 33598 7928 33654 7984
rect 32764 7642 32820 7644
rect 32844 7642 32900 7644
rect 32924 7642 32980 7644
rect 33004 7642 33060 7644
rect 32764 7590 32810 7642
rect 32810 7590 32820 7642
rect 32844 7590 32874 7642
rect 32874 7590 32886 7642
rect 32886 7590 32900 7642
rect 32924 7590 32938 7642
rect 32938 7590 32950 7642
rect 32950 7590 32980 7642
rect 33004 7590 33014 7642
rect 33014 7590 33060 7642
rect 32764 7588 32820 7590
rect 32844 7588 32900 7590
rect 32924 7588 32980 7590
rect 33004 7588 33060 7590
rect 32764 6554 32820 6556
rect 32844 6554 32900 6556
rect 32924 6554 32980 6556
rect 33004 6554 33060 6556
rect 32764 6502 32810 6554
rect 32810 6502 32820 6554
rect 32844 6502 32874 6554
rect 32874 6502 32886 6554
rect 32886 6502 32900 6554
rect 32924 6502 32938 6554
rect 32938 6502 32950 6554
rect 32950 6502 32980 6554
rect 33004 6502 33014 6554
rect 33014 6502 33060 6554
rect 32764 6500 32820 6502
rect 32844 6500 32900 6502
rect 32924 6500 32980 6502
rect 33004 6500 33060 6502
rect 32764 5466 32820 5468
rect 32844 5466 32900 5468
rect 32924 5466 32980 5468
rect 33004 5466 33060 5468
rect 32764 5414 32810 5466
rect 32810 5414 32820 5466
rect 32844 5414 32874 5466
rect 32874 5414 32886 5466
rect 32886 5414 32900 5466
rect 32924 5414 32938 5466
rect 32938 5414 32950 5466
rect 32950 5414 32980 5466
rect 33004 5414 33014 5466
rect 33014 5414 33060 5466
rect 32764 5412 32820 5414
rect 32844 5412 32900 5414
rect 32924 5412 32980 5414
rect 33004 5412 33060 5414
rect 32764 4378 32820 4380
rect 32844 4378 32900 4380
rect 32924 4378 32980 4380
rect 33004 4378 33060 4380
rect 32764 4326 32810 4378
rect 32810 4326 32820 4378
rect 32844 4326 32874 4378
rect 32874 4326 32886 4378
rect 32886 4326 32900 4378
rect 32924 4326 32938 4378
rect 32938 4326 32950 4378
rect 32950 4326 32980 4378
rect 33004 4326 33014 4378
rect 33014 4326 33060 4378
rect 32764 4324 32820 4326
rect 32844 4324 32900 4326
rect 32924 4324 32980 4326
rect 33004 4324 33060 4326
rect 32764 3290 32820 3292
rect 32844 3290 32900 3292
rect 32924 3290 32980 3292
rect 33004 3290 33060 3292
rect 32764 3238 32810 3290
rect 32810 3238 32820 3290
rect 32844 3238 32874 3290
rect 32874 3238 32886 3290
rect 32886 3238 32900 3290
rect 32924 3238 32938 3290
rect 32938 3238 32950 3290
rect 32950 3238 32980 3290
rect 33004 3238 33014 3290
rect 33014 3238 33060 3290
rect 32764 3236 32820 3238
rect 32844 3236 32900 3238
rect 32924 3236 32980 3238
rect 33004 3236 33060 3238
rect 32764 2202 32820 2204
rect 32844 2202 32900 2204
rect 32924 2202 32980 2204
rect 33004 2202 33060 2204
rect 32764 2150 32810 2202
rect 32810 2150 32820 2202
rect 32844 2150 32874 2202
rect 32874 2150 32886 2202
rect 32886 2150 32900 2202
rect 32924 2150 32938 2202
rect 32938 2150 32950 2202
rect 32950 2150 32980 2202
rect 33004 2150 33014 2202
rect 33014 2150 33060 2202
rect 32764 2148 32820 2150
rect 32844 2148 32900 2150
rect 32924 2148 32980 2150
rect 33004 2148 33060 2150
rect 34794 8336 34850 8392
rect 38066 8186 38122 8188
rect 38146 8186 38202 8188
rect 38226 8186 38282 8188
rect 38306 8186 38362 8188
rect 38066 8134 38112 8186
rect 38112 8134 38122 8186
rect 38146 8134 38176 8186
rect 38176 8134 38188 8186
rect 38188 8134 38202 8186
rect 38226 8134 38240 8186
rect 38240 8134 38252 8186
rect 38252 8134 38282 8186
rect 38306 8134 38316 8186
rect 38316 8134 38362 8186
rect 38066 8132 38122 8134
rect 38146 8132 38202 8134
rect 38226 8132 38282 8134
rect 38306 8132 38362 8134
rect 38066 7098 38122 7100
rect 38146 7098 38202 7100
rect 38226 7098 38282 7100
rect 38306 7098 38362 7100
rect 38066 7046 38112 7098
rect 38112 7046 38122 7098
rect 38146 7046 38176 7098
rect 38176 7046 38188 7098
rect 38188 7046 38202 7098
rect 38226 7046 38240 7098
rect 38240 7046 38252 7098
rect 38252 7046 38282 7098
rect 38306 7046 38316 7098
rect 38316 7046 38362 7098
rect 38066 7044 38122 7046
rect 38146 7044 38202 7046
rect 38226 7044 38282 7046
rect 38306 7044 38362 7046
rect 38066 6010 38122 6012
rect 38146 6010 38202 6012
rect 38226 6010 38282 6012
rect 38306 6010 38362 6012
rect 38066 5958 38112 6010
rect 38112 5958 38122 6010
rect 38146 5958 38176 6010
rect 38176 5958 38188 6010
rect 38188 5958 38202 6010
rect 38226 5958 38240 6010
rect 38240 5958 38252 6010
rect 38252 5958 38282 6010
rect 38306 5958 38316 6010
rect 38316 5958 38362 6010
rect 38066 5956 38122 5958
rect 38146 5956 38202 5958
rect 38226 5956 38282 5958
rect 38306 5956 38362 5958
rect 38066 4922 38122 4924
rect 38146 4922 38202 4924
rect 38226 4922 38282 4924
rect 38306 4922 38362 4924
rect 38066 4870 38112 4922
rect 38112 4870 38122 4922
rect 38146 4870 38176 4922
rect 38176 4870 38188 4922
rect 38188 4870 38202 4922
rect 38226 4870 38240 4922
rect 38240 4870 38252 4922
rect 38252 4870 38282 4922
rect 38306 4870 38316 4922
rect 38316 4870 38362 4922
rect 38066 4868 38122 4870
rect 38146 4868 38202 4870
rect 38226 4868 38282 4870
rect 38306 4868 38362 4870
rect 43367 8730 43423 8732
rect 43447 8730 43503 8732
rect 43527 8730 43583 8732
rect 43607 8730 43663 8732
rect 43367 8678 43413 8730
rect 43413 8678 43423 8730
rect 43447 8678 43477 8730
rect 43477 8678 43489 8730
rect 43489 8678 43503 8730
rect 43527 8678 43541 8730
rect 43541 8678 43553 8730
rect 43553 8678 43583 8730
rect 43607 8678 43617 8730
rect 43617 8678 43663 8730
rect 43367 8676 43423 8678
rect 43447 8676 43503 8678
rect 43527 8676 43583 8678
rect 43607 8676 43663 8678
rect 38066 3834 38122 3836
rect 38146 3834 38202 3836
rect 38226 3834 38282 3836
rect 38306 3834 38362 3836
rect 38066 3782 38112 3834
rect 38112 3782 38122 3834
rect 38146 3782 38176 3834
rect 38176 3782 38188 3834
rect 38188 3782 38202 3834
rect 38226 3782 38240 3834
rect 38240 3782 38252 3834
rect 38252 3782 38282 3834
rect 38306 3782 38316 3834
rect 38316 3782 38362 3834
rect 38066 3780 38122 3782
rect 38146 3780 38202 3782
rect 38226 3780 38282 3782
rect 38306 3780 38362 3782
rect 38066 2746 38122 2748
rect 38146 2746 38202 2748
rect 38226 2746 38282 2748
rect 38306 2746 38362 2748
rect 38066 2694 38112 2746
rect 38112 2694 38122 2746
rect 38146 2694 38176 2746
rect 38176 2694 38188 2746
rect 38188 2694 38202 2746
rect 38226 2694 38240 2746
rect 38240 2694 38252 2746
rect 38252 2694 38282 2746
rect 38306 2694 38316 2746
rect 38316 2694 38362 2746
rect 38066 2692 38122 2694
rect 38146 2692 38202 2694
rect 38226 2692 38282 2694
rect 38306 2692 38362 2694
rect 38066 1658 38122 1660
rect 38146 1658 38202 1660
rect 38226 1658 38282 1660
rect 38306 1658 38362 1660
rect 38066 1606 38112 1658
rect 38112 1606 38122 1658
rect 38146 1606 38176 1658
rect 38176 1606 38188 1658
rect 38188 1606 38202 1658
rect 38226 1606 38240 1658
rect 38240 1606 38252 1658
rect 38252 1606 38282 1658
rect 38306 1606 38316 1658
rect 38316 1606 38362 1658
rect 38066 1604 38122 1606
rect 38146 1604 38202 1606
rect 38226 1604 38282 1606
rect 38306 1604 38362 1606
rect 43367 7642 43423 7644
rect 43447 7642 43503 7644
rect 43527 7642 43583 7644
rect 43607 7642 43663 7644
rect 43367 7590 43413 7642
rect 43413 7590 43423 7642
rect 43447 7590 43477 7642
rect 43477 7590 43489 7642
rect 43489 7590 43503 7642
rect 43527 7590 43541 7642
rect 43541 7590 43553 7642
rect 43553 7590 43583 7642
rect 43607 7590 43617 7642
rect 43617 7590 43663 7642
rect 43367 7588 43423 7590
rect 43447 7588 43503 7590
rect 43527 7588 43583 7590
rect 43607 7588 43663 7590
rect 43367 6554 43423 6556
rect 43447 6554 43503 6556
rect 43527 6554 43583 6556
rect 43607 6554 43663 6556
rect 43367 6502 43413 6554
rect 43413 6502 43423 6554
rect 43447 6502 43477 6554
rect 43477 6502 43489 6554
rect 43489 6502 43503 6554
rect 43527 6502 43541 6554
rect 43541 6502 43553 6554
rect 43553 6502 43583 6554
rect 43607 6502 43617 6554
rect 43617 6502 43663 6554
rect 43367 6500 43423 6502
rect 43447 6500 43503 6502
rect 43527 6500 43583 6502
rect 43607 6500 43663 6502
rect 43367 5466 43423 5468
rect 43447 5466 43503 5468
rect 43527 5466 43583 5468
rect 43607 5466 43663 5468
rect 43367 5414 43413 5466
rect 43413 5414 43423 5466
rect 43447 5414 43477 5466
rect 43477 5414 43489 5466
rect 43489 5414 43503 5466
rect 43527 5414 43541 5466
rect 43541 5414 43553 5466
rect 43553 5414 43583 5466
rect 43607 5414 43617 5466
rect 43617 5414 43663 5466
rect 43367 5412 43423 5414
rect 43447 5412 43503 5414
rect 43527 5412 43583 5414
rect 43607 5412 43663 5414
rect 43367 4378 43423 4380
rect 43447 4378 43503 4380
rect 43527 4378 43583 4380
rect 43607 4378 43663 4380
rect 43367 4326 43413 4378
rect 43413 4326 43423 4378
rect 43447 4326 43477 4378
rect 43477 4326 43489 4378
rect 43489 4326 43503 4378
rect 43527 4326 43541 4378
rect 43541 4326 43553 4378
rect 43553 4326 43583 4378
rect 43607 4326 43617 4378
rect 43617 4326 43663 4378
rect 43367 4324 43423 4326
rect 43447 4324 43503 4326
rect 43527 4324 43583 4326
rect 43607 4324 43663 4326
rect 43367 3290 43423 3292
rect 43447 3290 43503 3292
rect 43527 3290 43583 3292
rect 43607 3290 43663 3292
rect 43367 3238 43413 3290
rect 43413 3238 43423 3290
rect 43447 3238 43477 3290
rect 43477 3238 43489 3290
rect 43489 3238 43503 3290
rect 43527 3238 43541 3290
rect 43541 3238 43553 3290
rect 43553 3238 43583 3290
rect 43607 3238 43617 3290
rect 43617 3238 43663 3290
rect 43367 3236 43423 3238
rect 43447 3236 43503 3238
rect 43527 3236 43583 3238
rect 43607 3236 43663 3238
rect 43367 2202 43423 2204
rect 43447 2202 43503 2204
rect 43527 2202 43583 2204
rect 43607 2202 43663 2204
rect 43367 2150 43413 2202
rect 43413 2150 43423 2202
rect 43447 2150 43477 2202
rect 43477 2150 43489 2202
rect 43489 2150 43503 2202
rect 43527 2150 43541 2202
rect 43541 2150 43553 2202
rect 43553 2150 43583 2202
rect 43607 2150 43617 2202
rect 43617 2150 43663 2202
rect 43367 2148 43423 2150
rect 43447 2148 43503 2150
rect 43527 2148 43583 2150
rect 43607 2148 43663 2150
rect 32764 1114 32820 1116
rect 32844 1114 32900 1116
rect 32924 1114 32980 1116
rect 33004 1114 33060 1116
rect 32764 1062 32810 1114
rect 32810 1062 32820 1114
rect 32844 1062 32874 1114
rect 32874 1062 32886 1114
rect 32886 1062 32900 1114
rect 32924 1062 32938 1114
rect 32938 1062 32950 1114
rect 32950 1062 32980 1114
rect 33004 1062 33014 1114
rect 33014 1062 33060 1114
rect 32764 1060 32820 1062
rect 32844 1060 32900 1062
rect 32924 1060 32980 1062
rect 33004 1060 33060 1062
rect 43367 1114 43423 1116
rect 43447 1114 43503 1116
rect 43527 1114 43583 1116
rect 43607 1114 43663 1116
rect 43367 1062 43413 1114
rect 43413 1062 43423 1114
rect 43447 1062 43477 1114
rect 43477 1062 43489 1114
rect 43489 1062 43503 1114
rect 43527 1062 43541 1114
rect 43541 1062 43553 1114
rect 43553 1062 43583 1114
rect 43607 1062 43617 1114
rect 43617 1062 43663 1114
rect 43367 1060 43423 1062
rect 43447 1060 43503 1062
rect 43527 1060 43583 1062
rect 43607 1060 43663 1062
<< metal3 >>
rect 19609 9892 19675 9893
rect 19558 9828 19564 9892
rect 19628 9890 19675 9892
rect 22093 9890 22159 9893
rect 19628 9888 19720 9890
rect 19670 9832 19720 9888
rect 19628 9830 19720 9832
rect 22093 9888 22754 9890
rect 22093 9832 22098 9888
rect 22154 9832 22754 9888
rect 22093 9830 22754 9832
rect 19628 9828 19675 9830
rect 19609 9827 19675 9828
rect 22093 9827 22159 9830
rect 22694 9754 22754 9830
rect 23197 9754 23263 9757
rect 22694 9752 23263 9754
rect 22694 9696 23202 9752
rect 23258 9696 23263 9752
rect 22694 9694 23263 9696
rect 23197 9691 23263 9694
rect 20989 9618 21055 9621
rect 22185 9618 22251 9621
rect 20989 9616 22251 9618
rect 20989 9560 20994 9616
rect 21050 9560 22190 9616
rect 22246 9560 22251 9616
rect 20989 9558 22251 9560
rect 20989 9555 21055 9558
rect 22185 9555 22251 9558
rect 21633 9482 21699 9485
rect 25681 9482 25747 9485
rect 21633 9480 25747 9482
rect 21633 9424 21638 9480
rect 21694 9424 25686 9480
rect 25742 9424 25747 9480
rect 21633 9422 25747 9424
rect 21633 9419 21699 9422
rect 25681 9419 25747 9422
rect 17677 9346 17743 9349
rect 21817 9346 21883 9349
rect 17677 9344 21883 9346
rect 17677 9288 17682 9344
rect 17738 9288 21822 9344
rect 21878 9288 21883 9344
rect 17677 9286 21883 9288
rect 17677 9283 17743 9286
rect 21817 9283 21883 9286
rect 21817 9210 21883 9213
rect 22737 9210 22803 9213
rect 21817 9208 22803 9210
rect 21817 9152 21822 9208
rect 21878 9152 22742 9208
rect 22798 9152 22803 9208
rect 21817 9150 22803 9152
rect 21817 9147 21883 9150
rect 22737 9147 22803 9150
rect 18965 9074 19031 9077
rect 19241 9074 19307 9077
rect 22185 9074 22251 9077
rect 18965 9072 19307 9074
rect 18965 9016 18970 9072
rect 19026 9016 19246 9072
rect 19302 9016 19307 9072
rect 18965 9014 19307 9016
rect 18965 9011 19031 9014
rect 19241 9011 19307 9014
rect 21774 9072 22251 9074
rect 21774 9016 22190 9072
rect 22246 9016 22251 9072
rect 21774 9014 22251 9016
rect 21633 8938 21699 8941
rect 21774 8938 21834 9014
rect 22185 9011 22251 9014
rect 23289 8938 23355 8941
rect 21633 8936 21834 8938
rect 21633 8880 21638 8936
rect 21694 8880 21834 8936
rect 21633 8878 21834 8880
rect 21958 8936 23355 8938
rect 21958 8880 23294 8936
rect 23350 8880 23355 8936
rect 21958 8878 23355 8880
rect 21633 8875 21699 8878
rect 19333 8802 19399 8805
rect 19609 8802 19675 8805
rect 21958 8802 22018 8878
rect 23289 8875 23355 8878
rect 30741 8938 30807 8941
rect 33501 8938 33567 8941
rect 30741 8936 33567 8938
rect 30741 8880 30746 8936
rect 30802 8880 33506 8936
rect 33562 8880 33567 8936
rect 30741 8878 33567 8880
rect 30741 8875 30807 8878
rect 33501 8875 33567 8878
rect 19333 8800 19675 8802
rect 19333 8744 19338 8800
rect 19394 8744 19614 8800
rect 19670 8744 19675 8800
rect 19333 8742 19675 8744
rect 19333 8739 19399 8742
rect 19609 8739 19675 8742
rect 21222 8742 22018 8802
rect 11548 8736 11864 8737
rect 11548 8672 11554 8736
rect 11618 8672 11634 8736
rect 11698 8672 11714 8736
rect 11778 8672 11794 8736
rect 11858 8672 11864 8736
rect 11548 8671 11864 8672
rect 14641 8666 14707 8669
rect 18781 8666 18847 8669
rect 14641 8664 18847 8666
rect 14641 8608 14646 8664
rect 14702 8608 18786 8664
rect 18842 8608 18847 8664
rect 14641 8606 18847 8608
rect 14641 8603 14707 8606
rect 18781 8603 18847 8606
rect 19701 8666 19767 8669
rect 21222 8666 21282 8742
rect 22151 8736 22467 8737
rect 22151 8672 22157 8736
rect 22221 8672 22237 8736
rect 22301 8672 22317 8736
rect 22381 8672 22397 8736
rect 22461 8672 22467 8736
rect 22151 8671 22467 8672
rect 32754 8736 33070 8737
rect 32754 8672 32760 8736
rect 32824 8672 32840 8736
rect 32904 8672 32920 8736
rect 32984 8672 33000 8736
rect 33064 8672 33070 8736
rect 32754 8671 33070 8672
rect 43357 8736 43673 8737
rect 43357 8672 43363 8736
rect 43427 8672 43443 8736
rect 43507 8672 43523 8736
rect 43587 8672 43603 8736
rect 43667 8672 43673 8736
rect 43357 8671 43673 8672
rect 19701 8664 21282 8666
rect 19701 8608 19706 8664
rect 19762 8608 21282 8664
rect 19701 8606 21282 8608
rect 19701 8603 19767 8606
rect 16941 8530 17007 8533
rect 21633 8530 21699 8533
rect 16941 8528 21699 8530
rect 16941 8472 16946 8528
rect 17002 8472 21638 8528
rect 21694 8472 21699 8528
rect 16941 8470 21699 8472
rect 16941 8467 17007 8470
rect 21633 8467 21699 8470
rect 30005 8530 30071 8533
rect 30373 8530 30439 8533
rect 30005 8528 30439 8530
rect 30005 8472 30010 8528
rect 30066 8472 30378 8528
rect 30434 8472 30439 8528
rect 30005 8470 30439 8472
rect 30005 8467 30071 8470
rect 30373 8467 30439 8470
rect 16849 8394 16915 8397
rect 19057 8394 19123 8397
rect 16849 8392 19123 8394
rect 16849 8336 16854 8392
rect 16910 8336 19062 8392
rect 19118 8336 19123 8392
rect 16849 8334 19123 8336
rect 16849 8331 16915 8334
rect 19057 8331 19123 8334
rect 19333 8396 19399 8397
rect 19333 8392 19380 8396
rect 19444 8394 19450 8396
rect 22645 8394 22711 8397
rect 27245 8394 27311 8397
rect 19333 8336 19338 8392
rect 19333 8332 19380 8336
rect 19444 8334 19490 8394
rect 22645 8392 27311 8394
rect 22645 8336 22650 8392
rect 22706 8336 27250 8392
rect 27306 8336 27311 8392
rect 22645 8334 27311 8336
rect 19444 8332 19450 8334
rect 19333 8331 19399 8332
rect 22645 8331 22711 8334
rect 27245 8331 27311 8334
rect 34462 8332 34468 8396
rect 34532 8394 34538 8396
rect 34789 8394 34855 8397
rect 34532 8392 34855 8394
rect 34532 8336 34794 8392
rect 34850 8336 34855 8392
rect 34532 8334 34855 8336
rect 34532 8332 34538 8334
rect 34789 8331 34855 8334
rect 25589 8258 25655 8261
rect 17358 8256 25655 8258
rect 17358 8200 25594 8256
rect 25650 8200 25655 8256
rect 17358 8198 25655 8200
rect 6247 8192 6563 8193
rect 6247 8128 6253 8192
rect 6317 8128 6333 8192
rect 6397 8128 6413 8192
rect 6477 8128 6493 8192
rect 6557 8128 6563 8192
rect 6247 8127 6563 8128
rect 16850 8192 17166 8193
rect 16850 8128 16856 8192
rect 16920 8128 16936 8192
rect 17000 8128 17016 8192
rect 17080 8128 17096 8192
rect 17160 8128 17166 8192
rect 16850 8127 17166 8128
rect 13721 7986 13787 7989
rect 17358 7986 17418 8198
rect 25589 8195 25655 8198
rect 27453 8192 27769 8193
rect 27453 8128 27459 8192
rect 27523 8128 27539 8192
rect 27603 8128 27619 8192
rect 27683 8128 27699 8192
rect 27763 8128 27769 8192
rect 27453 8127 27769 8128
rect 38056 8192 38372 8193
rect 38056 8128 38062 8192
rect 38126 8128 38142 8192
rect 38206 8128 38222 8192
rect 38286 8128 38302 8192
rect 38366 8128 38372 8192
rect 38056 8127 38372 8128
rect 17585 8122 17651 8125
rect 24945 8122 25011 8125
rect 17585 8120 25011 8122
rect 17585 8064 17590 8120
rect 17646 8064 24950 8120
rect 25006 8064 25011 8120
rect 17585 8062 25011 8064
rect 17585 8059 17651 8062
rect 24945 8059 25011 8062
rect 13721 7984 17418 7986
rect 13721 7928 13726 7984
rect 13782 7928 17418 7984
rect 13721 7926 17418 7928
rect 19425 7986 19491 7989
rect 20437 7986 20503 7989
rect 19425 7984 20503 7986
rect 19425 7928 19430 7984
rect 19486 7928 20442 7984
rect 20498 7928 20503 7984
rect 19425 7926 20503 7928
rect 13721 7923 13787 7926
rect 19425 7923 19491 7926
rect 20437 7923 20503 7926
rect 21357 7986 21423 7989
rect 33593 7986 33659 7989
rect 21357 7984 33659 7986
rect 21357 7928 21362 7984
rect 21418 7928 33598 7984
rect 33654 7928 33659 7984
rect 21357 7926 33659 7928
rect 21357 7923 21423 7926
rect 33593 7923 33659 7926
rect 11881 7850 11947 7853
rect 22277 7850 22343 7853
rect 11881 7848 22343 7850
rect 11881 7792 11886 7848
rect 11942 7792 22282 7848
rect 22338 7792 22343 7848
rect 11881 7790 22343 7792
rect 11881 7787 11947 7790
rect 22277 7787 22343 7790
rect 24761 7850 24827 7853
rect 28901 7850 28967 7853
rect 24761 7848 28967 7850
rect 24761 7792 24766 7848
rect 24822 7792 28906 7848
rect 28962 7792 28967 7848
rect 24761 7790 28967 7792
rect 24761 7787 24827 7790
rect 28901 7787 28967 7790
rect 16941 7714 17007 7717
rect 19149 7714 19215 7717
rect 16941 7712 19215 7714
rect 16941 7656 16946 7712
rect 17002 7656 19154 7712
rect 19210 7656 19215 7712
rect 16941 7654 19215 7656
rect 16941 7651 17007 7654
rect 19149 7651 19215 7654
rect 19333 7716 19399 7717
rect 19333 7712 19380 7716
rect 19444 7714 19450 7716
rect 19977 7714 20043 7717
rect 19333 7656 19338 7712
rect 19333 7652 19380 7656
rect 19444 7654 19490 7714
rect 19977 7712 21650 7714
rect 19977 7656 19982 7712
rect 20038 7656 21650 7712
rect 19977 7654 21650 7656
rect 19444 7652 19450 7654
rect 19333 7651 19399 7652
rect 19977 7651 20043 7654
rect 11548 7648 11864 7649
rect 11548 7584 11554 7648
rect 11618 7584 11634 7648
rect 11698 7584 11714 7648
rect 11778 7584 11794 7648
rect 11858 7584 11864 7648
rect 11548 7583 11864 7584
rect 12893 7578 12959 7581
rect 12893 7576 21466 7578
rect 12893 7520 12898 7576
rect 12954 7520 21466 7576
rect 12893 7518 21466 7520
rect 12893 7515 12959 7518
rect 16757 7442 16823 7445
rect 19425 7442 19491 7445
rect 19609 7444 19675 7445
rect 16757 7440 19491 7442
rect 16757 7384 16762 7440
rect 16818 7384 19430 7440
rect 19486 7384 19491 7440
rect 16757 7382 19491 7384
rect 16757 7379 16823 7382
rect 19425 7379 19491 7382
rect 19558 7380 19564 7444
rect 19628 7442 19675 7444
rect 19628 7440 19720 7442
rect 19670 7384 19720 7440
rect 19628 7382 19720 7384
rect 19628 7380 19675 7382
rect 19609 7379 19675 7380
rect 16757 7306 16823 7309
rect 21173 7306 21239 7309
rect 16757 7304 21239 7306
rect 16757 7248 16762 7304
rect 16818 7248 21178 7304
rect 21234 7248 21239 7304
rect 16757 7246 21239 7248
rect 21406 7306 21466 7518
rect 21590 7442 21650 7654
rect 22151 7648 22467 7649
rect 22151 7584 22157 7648
rect 22221 7584 22237 7648
rect 22301 7584 22317 7648
rect 22381 7584 22397 7648
rect 22461 7584 22467 7648
rect 22151 7583 22467 7584
rect 32754 7648 33070 7649
rect 32754 7584 32760 7648
rect 32824 7584 32840 7648
rect 32904 7584 32920 7648
rect 32984 7584 33000 7648
rect 33064 7584 33070 7648
rect 32754 7583 33070 7584
rect 43357 7648 43673 7649
rect 43357 7584 43363 7648
rect 43427 7584 43443 7648
rect 43507 7584 43523 7648
rect 43587 7584 43603 7648
rect 43667 7584 43673 7648
rect 43357 7583 43673 7584
rect 32397 7442 32463 7445
rect 21590 7440 32463 7442
rect 21590 7384 32402 7440
rect 32458 7384 32463 7440
rect 21590 7382 32463 7384
rect 32397 7379 32463 7382
rect 27429 7306 27495 7309
rect 21406 7304 27495 7306
rect 21406 7248 27434 7304
rect 27490 7248 27495 7304
rect 21406 7246 27495 7248
rect 16757 7243 16823 7246
rect 21173 7243 21239 7246
rect 27429 7243 27495 7246
rect 17309 7170 17375 7173
rect 21357 7170 21423 7173
rect 17309 7168 21423 7170
rect 17309 7112 17314 7168
rect 17370 7112 21362 7168
rect 21418 7112 21423 7168
rect 17309 7110 21423 7112
rect 17309 7107 17375 7110
rect 21357 7107 21423 7110
rect 6247 7104 6563 7105
rect 6247 7040 6253 7104
rect 6317 7040 6333 7104
rect 6397 7040 6413 7104
rect 6477 7040 6493 7104
rect 6557 7040 6563 7104
rect 6247 7039 6563 7040
rect 16850 7104 17166 7105
rect 16850 7040 16856 7104
rect 16920 7040 16936 7104
rect 17000 7040 17016 7104
rect 17080 7040 17096 7104
rect 17160 7040 17166 7104
rect 16850 7039 17166 7040
rect 27453 7104 27769 7105
rect 27453 7040 27459 7104
rect 27523 7040 27539 7104
rect 27603 7040 27619 7104
rect 27683 7040 27699 7104
rect 27763 7040 27769 7104
rect 27453 7039 27769 7040
rect 38056 7104 38372 7105
rect 38056 7040 38062 7104
rect 38126 7040 38142 7104
rect 38206 7040 38222 7104
rect 38286 7040 38302 7104
rect 38366 7040 38372 7104
rect 38056 7039 38372 7040
rect 13813 7034 13879 7037
rect 16665 7034 16731 7037
rect 13813 7032 16731 7034
rect 13813 6976 13818 7032
rect 13874 6976 16670 7032
rect 16726 6976 16731 7032
rect 13813 6974 16731 6976
rect 13813 6971 13879 6974
rect 16665 6971 16731 6974
rect 17309 7034 17375 7037
rect 23933 7034 23999 7037
rect 17309 7032 23999 7034
rect 17309 6976 17314 7032
rect 17370 6976 23938 7032
rect 23994 6976 23999 7032
rect 17309 6974 23999 6976
rect 17309 6971 17375 6974
rect 23933 6971 23999 6974
rect 11973 6898 12039 6901
rect 23381 6898 23447 6901
rect 11973 6896 23447 6898
rect 11973 6840 11978 6896
rect 12034 6840 23386 6896
rect 23442 6840 23447 6896
rect 11973 6838 23447 6840
rect 11973 6835 12039 6838
rect 23381 6835 23447 6838
rect 14273 6762 14339 6765
rect 22553 6762 22619 6765
rect 14273 6760 22619 6762
rect 14273 6704 14278 6760
rect 14334 6704 22558 6760
rect 22614 6704 22619 6760
rect 14273 6702 22619 6704
rect 14273 6699 14339 6702
rect 22553 6699 22619 6702
rect 11548 6560 11864 6561
rect 11548 6496 11554 6560
rect 11618 6496 11634 6560
rect 11698 6496 11714 6560
rect 11778 6496 11794 6560
rect 11858 6496 11864 6560
rect 11548 6495 11864 6496
rect 22151 6560 22467 6561
rect 22151 6496 22157 6560
rect 22221 6496 22237 6560
rect 22301 6496 22317 6560
rect 22381 6496 22397 6560
rect 22461 6496 22467 6560
rect 22151 6495 22467 6496
rect 32754 6560 33070 6561
rect 32754 6496 32760 6560
rect 32824 6496 32840 6560
rect 32904 6496 32920 6560
rect 32984 6496 33000 6560
rect 33064 6496 33070 6560
rect 32754 6495 33070 6496
rect 43357 6560 43673 6561
rect 43357 6496 43363 6560
rect 43427 6496 43443 6560
rect 43507 6496 43523 6560
rect 43587 6496 43603 6560
rect 43667 6496 43673 6560
rect 43357 6495 43673 6496
rect 6821 6354 6887 6357
rect 24669 6354 24735 6357
rect 6821 6352 24735 6354
rect 6821 6296 6826 6352
rect 6882 6296 24674 6352
rect 24730 6296 24735 6352
rect 6821 6294 24735 6296
rect 6821 6291 6887 6294
rect 24669 6291 24735 6294
rect 7189 6218 7255 6221
rect 24393 6218 24459 6221
rect 7189 6216 24459 6218
rect 7189 6160 7194 6216
rect 7250 6160 24398 6216
rect 24454 6160 24459 6216
rect 7189 6158 24459 6160
rect 7189 6155 7255 6158
rect 24393 6155 24459 6158
rect 6247 6016 6563 6017
rect 6247 5952 6253 6016
rect 6317 5952 6333 6016
rect 6397 5952 6413 6016
rect 6477 5952 6493 6016
rect 6557 5952 6563 6016
rect 6247 5951 6563 5952
rect 16850 6016 17166 6017
rect 16850 5952 16856 6016
rect 16920 5952 16936 6016
rect 17000 5952 17016 6016
rect 17080 5952 17096 6016
rect 17160 5952 17166 6016
rect 16850 5951 17166 5952
rect 27453 6016 27769 6017
rect 27453 5952 27459 6016
rect 27523 5952 27539 6016
rect 27603 5952 27619 6016
rect 27683 5952 27699 6016
rect 27763 5952 27769 6016
rect 27453 5951 27769 5952
rect 38056 6016 38372 6017
rect 38056 5952 38062 6016
rect 38126 5952 38142 6016
rect 38206 5952 38222 6016
rect 38286 5952 38302 6016
rect 38366 5952 38372 6016
rect 38056 5951 38372 5952
rect 12341 5810 12407 5813
rect 22829 5810 22895 5813
rect 12341 5808 22895 5810
rect 12341 5752 12346 5808
rect 12402 5752 22834 5808
rect 22890 5752 22895 5808
rect 12341 5750 22895 5752
rect 12341 5747 12407 5750
rect 22829 5747 22895 5750
rect 11548 5472 11864 5473
rect 11548 5408 11554 5472
rect 11618 5408 11634 5472
rect 11698 5408 11714 5472
rect 11778 5408 11794 5472
rect 11858 5408 11864 5472
rect 11548 5407 11864 5408
rect 22151 5472 22467 5473
rect 22151 5408 22157 5472
rect 22221 5408 22237 5472
rect 22301 5408 22317 5472
rect 22381 5408 22397 5472
rect 22461 5408 22467 5472
rect 22151 5407 22467 5408
rect 32754 5472 33070 5473
rect 32754 5408 32760 5472
rect 32824 5408 32840 5472
rect 32904 5408 32920 5472
rect 32984 5408 33000 5472
rect 33064 5408 33070 5472
rect 32754 5407 33070 5408
rect 43357 5472 43673 5473
rect 43357 5408 43363 5472
rect 43427 5408 43443 5472
rect 43507 5408 43523 5472
rect 43587 5408 43603 5472
rect 43667 5408 43673 5472
rect 43357 5407 43673 5408
rect 6247 4928 6563 4929
rect 6247 4864 6253 4928
rect 6317 4864 6333 4928
rect 6397 4864 6413 4928
rect 6477 4864 6493 4928
rect 6557 4864 6563 4928
rect 6247 4863 6563 4864
rect 16850 4928 17166 4929
rect 16850 4864 16856 4928
rect 16920 4864 16936 4928
rect 17000 4864 17016 4928
rect 17080 4864 17096 4928
rect 17160 4864 17166 4928
rect 16850 4863 17166 4864
rect 27453 4928 27769 4929
rect 27453 4864 27459 4928
rect 27523 4864 27539 4928
rect 27603 4864 27619 4928
rect 27683 4864 27699 4928
rect 27763 4864 27769 4928
rect 27453 4863 27769 4864
rect 38056 4928 38372 4929
rect 38056 4864 38062 4928
rect 38126 4864 38142 4928
rect 38206 4864 38222 4928
rect 38286 4864 38302 4928
rect 38366 4864 38372 4928
rect 38056 4863 38372 4864
rect 11548 4384 11864 4385
rect 11548 4320 11554 4384
rect 11618 4320 11634 4384
rect 11698 4320 11714 4384
rect 11778 4320 11794 4384
rect 11858 4320 11864 4384
rect 11548 4319 11864 4320
rect 22151 4384 22467 4385
rect 22151 4320 22157 4384
rect 22221 4320 22237 4384
rect 22301 4320 22317 4384
rect 22381 4320 22397 4384
rect 22461 4320 22467 4384
rect 22151 4319 22467 4320
rect 32754 4384 33070 4385
rect 32754 4320 32760 4384
rect 32824 4320 32840 4384
rect 32904 4320 32920 4384
rect 32984 4320 33000 4384
rect 33064 4320 33070 4384
rect 32754 4319 33070 4320
rect 43357 4384 43673 4385
rect 43357 4320 43363 4384
rect 43427 4320 43443 4384
rect 43507 4320 43523 4384
rect 43587 4320 43603 4384
rect 43667 4320 43673 4384
rect 43357 4319 43673 4320
rect 6247 3840 6563 3841
rect 6247 3776 6253 3840
rect 6317 3776 6333 3840
rect 6397 3776 6413 3840
rect 6477 3776 6493 3840
rect 6557 3776 6563 3840
rect 6247 3775 6563 3776
rect 16850 3840 17166 3841
rect 16850 3776 16856 3840
rect 16920 3776 16936 3840
rect 17000 3776 17016 3840
rect 17080 3776 17096 3840
rect 17160 3776 17166 3840
rect 16850 3775 17166 3776
rect 27453 3840 27769 3841
rect 27453 3776 27459 3840
rect 27523 3776 27539 3840
rect 27603 3776 27619 3840
rect 27683 3776 27699 3840
rect 27763 3776 27769 3840
rect 27453 3775 27769 3776
rect 38056 3840 38372 3841
rect 38056 3776 38062 3840
rect 38126 3776 38142 3840
rect 38206 3776 38222 3840
rect 38286 3776 38302 3840
rect 38366 3776 38372 3840
rect 38056 3775 38372 3776
rect 11548 3296 11864 3297
rect 11548 3232 11554 3296
rect 11618 3232 11634 3296
rect 11698 3232 11714 3296
rect 11778 3232 11794 3296
rect 11858 3232 11864 3296
rect 11548 3231 11864 3232
rect 22151 3296 22467 3297
rect 22151 3232 22157 3296
rect 22221 3232 22237 3296
rect 22301 3232 22317 3296
rect 22381 3232 22397 3296
rect 22461 3232 22467 3296
rect 22151 3231 22467 3232
rect 32754 3296 33070 3297
rect 32754 3232 32760 3296
rect 32824 3232 32840 3296
rect 32904 3232 32920 3296
rect 32984 3232 33000 3296
rect 33064 3232 33070 3296
rect 32754 3231 33070 3232
rect 43357 3296 43673 3297
rect 43357 3232 43363 3296
rect 43427 3232 43443 3296
rect 43507 3232 43523 3296
rect 43587 3232 43603 3296
rect 43667 3232 43673 3296
rect 43357 3231 43673 3232
rect 23381 2954 23447 2957
rect 34462 2954 34468 2956
rect 23381 2952 34468 2954
rect 23381 2896 23386 2952
rect 23442 2896 34468 2952
rect 23381 2894 34468 2896
rect 23381 2891 23447 2894
rect 34462 2892 34468 2894
rect 34532 2892 34538 2956
rect 6247 2752 6563 2753
rect 6247 2688 6253 2752
rect 6317 2688 6333 2752
rect 6397 2688 6413 2752
rect 6477 2688 6493 2752
rect 6557 2688 6563 2752
rect 6247 2687 6563 2688
rect 16850 2752 17166 2753
rect 16850 2688 16856 2752
rect 16920 2688 16936 2752
rect 17000 2688 17016 2752
rect 17080 2688 17096 2752
rect 17160 2688 17166 2752
rect 16850 2687 17166 2688
rect 27453 2752 27769 2753
rect 27453 2688 27459 2752
rect 27523 2688 27539 2752
rect 27603 2688 27619 2752
rect 27683 2688 27699 2752
rect 27763 2688 27769 2752
rect 27453 2687 27769 2688
rect 38056 2752 38372 2753
rect 38056 2688 38062 2752
rect 38126 2688 38142 2752
rect 38206 2688 38222 2752
rect 38286 2688 38302 2752
rect 38366 2688 38372 2752
rect 38056 2687 38372 2688
rect 11548 2208 11864 2209
rect 11548 2144 11554 2208
rect 11618 2144 11634 2208
rect 11698 2144 11714 2208
rect 11778 2144 11794 2208
rect 11858 2144 11864 2208
rect 11548 2143 11864 2144
rect 22151 2208 22467 2209
rect 22151 2144 22157 2208
rect 22221 2144 22237 2208
rect 22301 2144 22317 2208
rect 22381 2144 22397 2208
rect 22461 2144 22467 2208
rect 22151 2143 22467 2144
rect 32754 2208 33070 2209
rect 32754 2144 32760 2208
rect 32824 2144 32840 2208
rect 32904 2144 32920 2208
rect 32984 2144 33000 2208
rect 33064 2144 33070 2208
rect 32754 2143 33070 2144
rect 43357 2208 43673 2209
rect 43357 2144 43363 2208
rect 43427 2144 43443 2208
rect 43507 2144 43523 2208
rect 43587 2144 43603 2208
rect 43667 2144 43673 2208
rect 43357 2143 43673 2144
rect 6247 1664 6563 1665
rect 6247 1600 6253 1664
rect 6317 1600 6333 1664
rect 6397 1600 6413 1664
rect 6477 1600 6493 1664
rect 6557 1600 6563 1664
rect 6247 1599 6563 1600
rect 16850 1664 17166 1665
rect 16850 1600 16856 1664
rect 16920 1600 16936 1664
rect 17000 1600 17016 1664
rect 17080 1600 17096 1664
rect 17160 1600 17166 1664
rect 16850 1599 17166 1600
rect 27453 1664 27769 1665
rect 27453 1600 27459 1664
rect 27523 1600 27539 1664
rect 27603 1600 27619 1664
rect 27683 1600 27699 1664
rect 27763 1600 27769 1664
rect 27453 1599 27769 1600
rect 38056 1664 38372 1665
rect 38056 1600 38062 1664
rect 38126 1600 38142 1664
rect 38206 1600 38222 1664
rect 38286 1600 38302 1664
rect 38366 1600 38372 1664
rect 38056 1599 38372 1600
rect 11548 1120 11864 1121
rect 11548 1056 11554 1120
rect 11618 1056 11634 1120
rect 11698 1056 11714 1120
rect 11778 1056 11794 1120
rect 11858 1056 11864 1120
rect 11548 1055 11864 1056
rect 22151 1120 22467 1121
rect 22151 1056 22157 1120
rect 22221 1056 22237 1120
rect 22301 1056 22317 1120
rect 22381 1056 22397 1120
rect 22461 1056 22467 1120
rect 22151 1055 22467 1056
rect 32754 1120 33070 1121
rect 32754 1056 32760 1120
rect 32824 1056 32840 1120
rect 32904 1056 32920 1120
rect 32984 1056 33000 1120
rect 33064 1056 33070 1120
rect 32754 1055 33070 1056
rect 43357 1120 43673 1121
rect 43357 1056 43363 1120
rect 43427 1056 43443 1120
rect 43507 1056 43523 1120
rect 43587 1056 43603 1120
rect 43667 1056 43673 1120
rect 43357 1055 43673 1056
<< via3 >>
rect 19564 9888 19628 9892
rect 19564 9832 19614 9888
rect 19614 9832 19628 9888
rect 19564 9828 19628 9832
rect 11554 8732 11618 8736
rect 11554 8676 11558 8732
rect 11558 8676 11614 8732
rect 11614 8676 11618 8732
rect 11554 8672 11618 8676
rect 11634 8732 11698 8736
rect 11634 8676 11638 8732
rect 11638 8676 11694 8732
rect 11694 8676 11698 8732
rect 11634 8672 11698 8676
rect 11714 8732 11778 8736
rect 11714 8676 11718 8732
rect 11718 8676 11774 8732
rect 11774 8676 11778 8732
rect 11714 8672 11778 8676
rect 11794 8732 11858 8736
rect 11794 8676 11798 8732
rect 11798 8676 11854 8732
rect 11854 8676 11858 8732
rect 11794 8672 11858 8676
rect 22157 8732 22221 8736
rect 22157 8676 22161 8732
rect 22161 8676 22217 8732
rect 22217 8676 22221 8732
rect 22157 8672 22221 8676
rect 22237 8732 22301 8736
rect 22237 8676 22241 8732
rect 22241 8676 22297 8732
rect 22297 8676 22301 8732
rect 22237 8672 22301 8676
rect 22317 8732 22381 8736
rect 22317 8676 22321 8732
rect 22321 8676 22377 8732
rect 22377 8676 22381 8732
rect 22317 8672 22381 8676
rect 22397 8732 22461 8736
rect 22397 8676 22401 8732
rect 22401 8676 22457 8732
rect 22457 8676 22461 8732
rect 22397 8672 22461 8676
rect 32760 8732 32824 8736
rect 32760 8676 32764 8732
rect 32764 8676 32820 8732
rect 32820 8676 32824 8732
rect 32760 8672 32824 8676
rect 32840 8732 32904 8736
rect 32840 8676 32844 8732
rect 32844 8676 32900 8732
rect 32900 8676 32904 8732
rect 32840 8672 32904 8676
rect 32920 8732 32984 8736
rect 32920 8676 32924 8732
rect 32924 8676 32980 8732
rect 32980 8676 32984 8732
rect 32920 8672 32984 8676
rect 33000 8732 33064 8736
rect 33000 8676 33004 8732
rect 33004 8676 33060 8732
rect 33060 8676 33064 8732
rect 33000 8672 33064 8676
rect 43363 8732 43427 8736
rect 43363 8676 43367 8732
rect 43367 8676 43423 8732
rect 43423 8676 43427 8732
rect 43363 8672 43427 8676
rect 43443 8732 43507 8736
rect 43443 8676 43447 8732
rect 43447 8676 43503 8732
rect 43503 8676 43507 8732
rect 43443 8672 43507 8676
rect 43523 8732 43587 8736
rect 43523 8676 43527 8732
rect 43527 8676 43583 8732
rect 43583 8676 43587 8732
rect 43523 8672 43587 8676
rect 43603 8732 43667 8736
rect 43603 8676 43607 8732
rect 43607 8676 43663 8732
rect 43663 8676 43667 8732
rect 43603 8672 43667 8676
rect 19380 8392 19444 8396
rect 19380 8336 19394 8392
rect 19394 8336 19444 8392
rect 19380 8332 19444 8336
rect 34468 8332 34532 8396
rect 6253 8188 6317 8192
rect 6253 8132 6257 8188
rect 6257 8132 6313 8188
rect 6313 8132 6317 8188
rect 6253 8128 6317 8132
rect 6333 8188 6397 8192
rect 6333 8132 6337 8188
rect 6337 8132 6393 8188
rect 6393 8132 6397 8188
rect 6333 8128 6397 8132
rect 6413 8188 6477 8192
rect 6413 8132 6417 8188
rect 6417 8132 6473 8188
rect 6473 8132 6477 8188
rect 6413 8128 6477 8132
rect 6493 8188 6557 8192
rect 6493 8132 6497 8188
rect 6497 8132 6553 8188
rect 6553 8132 6557 8188
rect 6493 8128 6557 8132
rect 16856 8188 16920 8192
rect 16856 8132 16860 8188
rect 16860 8132 16916 8188
rect 16916 8132 16920 8188
rect 16856 8128 16920 8132
rect 16936 8188 17000 8192
rect 16936 8132 16940 8188
rect 16940 8132 16996 8188
rect 16996 8132 17000 8188
rect 16936 8128 17000 8132
rect 17016 8188 17080 8192
rect 17016 8132 17020 8188
rect 17020 8132 17076 8188
rect 17076 8132 17080 8188
rect 17016 8128 17080 8132
rect 17096 8188 17160 8192
rect 17096 8132 17100 8188
rect 17100 8132 17156 8188
rect 17156 8132 17160 8188
rect 17096 8128 17160 8132
rect 27459 8188 27523 8192
rect 27459 8132 27463 8188
rect 27463 8132 27519 8188
rect 27519 8132 27523 8188
rect 27459 8128 27523 8132
rect 27539 8188 27603 8192
rect 27539 8132 27543 8188
rect 27543 8132 27599 8188
rect 27599 8132 27603 8188
rect 27539 8128 27603 8132
rect 27619 8188 27683 8192
rect 27619 8132 27623 8188
rect 27623 8132 27679 8188
rect 27679 8132 27683 8188
rect 27619 8128 27683 8132
rect 27699 8188 27763 8192
rect 27699 8132 27703 8188
rect 27703 8132 27759 8188
rect 27759 8132 27763 8188
rect 27699 8128 27763 8132
rect 38062 8188 38126 8192
rect 38062 8132 38066 8188
rect 38066 8132 38122 8188
rect 38122 8132 38126 8188
rect 38062 8128 38126 8132
rect 38142 8188 38206 8192
rect 38142 8132 38146 8188
rect 38146 8132 38202 8188
rect 38202 8132 38206 8188
rect 38142 8128 38206 8132
rect 38222 8188 38286 8192
rect 38222 8132 38226 8188
rect 38226 8132 38282 8188
rect 38282 8132 38286 8188
rect 38222 8128 38286 8132
rect 38302 8188 38366 8192
rect 38302 8132 38306 8188
rect 38306 8132 38362 8188
rect 38362 8132 38366 8188
rect 38302 8128 38366 8132
rect 19380 7712 19444 7716
rect 19380 7656 19394 7712
rect 19394 7656 19444 7712
rect 19380 7652 19444 7656
rect 11554 7644 11618 7648
rect 11554 7588 11558 7644
rect 11558 7588 11614 7644
rect 11614 7588 11618 7644
rect 11554 7584 11618 7588
rect 11634 7644 11698 7648
rect 11634 7588 11638 7644
rect 11638 7588 11694 7644
rect 11694 7588 11698 7644
rect 11634 7584 11698 7588
rect 11714 7644 11778 7648
rect 11714 7588 11718 7644
rect 11718 7588 11774 7644
rect 11774 7588 11778 7644
rect 11714 7584 11778 7588
rect 11794 7644 11858 7648
rect 11794 7588 11798 7644
rect 11798 7588 11854 7644
rect 11854 7588 11858 7644
rect 11794 7584 11858 7588
rect 19564 7440 19628 7444
rect 19564 7384 19614 7440
rect 19614 7384 19628 7440
rect 19564 7380 19628 7384
rect 22157 7644 22221 7648
rect 22157 7588 22161 7644
rect 22161 7588 22217 7644
rect 22217 7588 22221 7644
rect 22157 7584 22221 7588
rect 22237 7644 22301 7648
rect 22237 7588 22241 7644
rect 22241 7588 22297 7644
rect 22297 7588 22301 7644
rect 22237 7584 22301 7588
rect 22317 7644 22381 7648
rect 22317 7588 22321 7644
rect 22321 7588 22377 7644
rect 22377 7588 22381 7644
rect 22317 7584 22381 7588
rect 22397 7644 22461 7648
rect 22397 7588 22401 7644
rect 22401 7588 22457 7644
rect 22457 7588 22461 7644
rect 22397 7584 22461 7588
rect 32760 7644 32824 7648
rect 32760 7588 32764 7644
rect 32764 7588 32820 7644
rect 32820 7588 32824 7644
rect 32760 7584 32824 7588
rect 32840 7644 32904 7648
rect 32840 7588 32844 7644
rect 32844 7588 32900 7644
rect 32900 7588 32904 7644
rect 32840 7584 32904 7588
rect 32920 7644 32984 7648
rect 32920 7588 32924 7644
rect 32924 7588 32980 7644
rect 32980 7588 32984 7644
rect 32920 7584 32984 7588
rect 33000 7644 33064 7648
rect 33000 7588 33004 7644
rect 33004 7588 33060 7644
rect 33060 7588 33064 7644
rect 33000 7584 33064 7588
rect 43363 7644 43427 7648
rect 43363 7588 43367 7644
rect 43367 7588 43423 7644
rect 43423 7588 43427 7644
rect 43363 7584 43427 7588
rect 43443 7644 43507 7648
rect 43443 7588 43447 7644
rect 43447 7588 43503 7644
rect 43503 7588 43507 7644
rect 43443 7584 43507 7588
rect 43523 7644 43587 7648
rect 43523 7588 43527 7644
rect 43527 7588 43583 7644
rect 43583 7588 43587 7644
rect 43523 7584 43587 7588
rect 43603 7644 43667 7648
rect 43603 7588 43607 7644
rect 43607 7588 43663 7644
rect 43663 7588 43667 7644
rect 43603 7584 43667 7588
rect 6253 7100 6317 7104
rect 6253 7044 6257 7100
rect 6257 7044 6313 7100
rect 6313 7044 6317 7100
rect 6253 7040 6317 7044
rect 6333 7100 6397 7104
rect 6333 7044 6337 7100
rect 6337 7044 6393 7100
rect 6393 7044 6397 7100
rect 6333 7040 6397 7044
rect 6413 7100 6477 7104
rect 6413 7044 6417 7100
rect 6417 7044 6473 7100
rect 6473 7044 6477 7100
rect 6413 7040 6477 7044
rect 6493 7100 6557 7104
rect 6493 7044 6497 7100
rect 6497 7044 6553 7100
rect 6553 7044 6557 7100
rect 6493 7040 6557 7044
rect 16856 7100 16920 7104
rect 16856 7044 16860 7100
rect 16860 7044 16916 7100
rect 16916 7044 16920 7100
rect 16856 7040 16920 7044
rect 16936 7100 17000 7104
rect 16936 7044 16940 7100
rect 16940 7044 16996 7100
rect 16996 7044 17000 7100
rect 16936 7040 17000 7044
rect 17016 7100 17080 7104
rect 17016 7044 17020 7100
rect 17020 7044 17076 7100
rect 17076 7044 17080 7100
rect 17016 7040 17080 7044
rect 17096 7100 17160 7104
rect 17096 7044 17100 7100
rect 17100 7044 17156 7100
rect 17156 7044 17160 7100
rect 17096 7040 17160 7044
rect 27459 7100 27523 7104
rect 27459 7044 27463 7100
rect 27463 7044 27519 7100
rect 27519 7044 27523 7100
rect 27459 7040 27523 7044
rect 27539 7100 27603 7104
rect 27539 7044 27543 7100
rect 27543 7044 27599 7100
rect 27599 7044 27603 7100
rect 27539 7040 27603 7044
rect 27619 7100 27683 7104
rect 27619 7044 27623 7100
rect 27623 7044 27679 7100
rect 27679 7044 27683 7100
rect 27619 7040 27683 7044
rect 27699 7100 27763 7104
rect 27699 7044 27703 7100
rect 27703 7044 27759 7100
rect 27759 7044 27763 7100
rect 27699 7040 27763 7044
rect 38062 7100 38126 7104
rect 38062 7044 38066 7100
rect 38066 7044 38122 7100
rect 38122 7044 38126 7100
rect 38062 7040 38126 7044
rect 38142 7100 38206 7104
rect 38142 7044 38146 7100
rect 38146 7044 38202 7100
rect 38202 7044 38206 7100
rect 38142 7040 38206 7044
rect 38222 7100 38286 7104
rect 38222 7044 38226 7100
rect 38226 7044 38282 7100
rect 38282 7044 38286 7100
rect 38222 7040 38286 7044
rect 38302 7100 38366 7104
rect 38302 7044 38306 7100
rect 38306 7044 38362 7100
rect 38362 7044 38366 7100
rect 38302 7040 38366 7044
rect 11554 6556 11618 6560
rect 11554 6500 11558 6556
rect 11558 6500 11614 6556
rect 11614 6500 11618 6556
rect 11554 6496 11618 6500
rect 11634 6556 11698 6560
rect 11634 6500 11638 6556
rect 11638 6500 11694 6556
rect 11694 6500 11698 6556
rect 11634 6496 11698 6500
rect 11714 6556 11778 6560
rect 11714 6500 11718 6556
rect 11718 6500 11774 6556
rect 11774 6500 11778 6556
rect 11714 6496 11778 6500
rect 11794 6556 11858 6560
rect 11794 6500 11798 6556
rect 11798 6500 11854 6556
rect 11854 6500 11858 6556
rect 11794 6496 11858 6500
rect 22157 6556 22221 6560
rect 22157 6500 22161 6556
rect 22161 6500 22217 6556
rect 22217 6500 22221 6556
rect 22157 6496 22221 6500
rect 22237 6556 22301 6560
rect 22237 6500 22241 6556
rect 22241 6500 22297 6556
rect 22297 6500 22301 6556
rect 22237 6496 22301 6500
rect 22317 6556 22381 6560
rect 22317 6500 22321 6556
rect 22321 6500 22377 6556
rect 22377 6500 22381 6556
rect 22317 6496 22381 6500
rect 22397 6556 22461 6560
rect 22397 6500 22401 6556
rect 22401 6500 22457 6556
rect 22457 6500 22461 6556
rect 22397 6496 22461 6500
rect 32760 6556 32824 6560
rect 32760 6500 32764 6556
rect 32764 6500 32820 6556
rect 32820 6500 32824 6556
rect 32760 6496 32824 6500
rect 32840 6556 32904 6560
rect 32840 6500 32844 6556
rect 32844 6500 32900 6556
rect 32900 6500 32904 6556
rect 32840 6496 32904 6500
rect 32920 6556 32984 6560
rect 32920 6500 32924 6556
rect 32924 6500 32980 6556
rect 32980 6500 32984 6556
rect 32920 6496 32984 6500
rect 33000 6556 33064 6560
rect 33000 6500 33004 6556
rect 33004 6500 33060 6556
rect 33060 6500 33064 6556
rect 33000 6496 33064 6500
rect 43363 6556 43427 6560
rect 43363 6500 43367 6556
rect 43367 6500 43423 6556
rect 43423 6500 43427 6556
rect 43363 6496 43427 6500
rect 43443 6556 43507 6560
rect 43443 6500 43447 6556
rect 43447 6500 43503 6556
rect 43503 6500 43507 6556
rect 43443 6496 43507 6500
rect 43523 6556 43587 6560
rect 43523 6500 43527 6556
rect 43527 6500 43583 6556
rect 43583 6500 43587 6556
rect 43523 6496 43587 6500
rect 43603 6556 43667 6560
rect 43603 6500 43607 6556
rect 43607 6500 43663 6556
rect 43663 6500 43667 6556
rect 43603 6496 43667 6500
rect 6253 6012 6317 6016
rect 6253 5956 6257 6012
rect 6257 5956 6313 6012
rect 6313 5956 6317 6012
rect 6253 5952 6317 5956
rect 6333 6012 6397 6016
rect 6333 5956 6337 6012
rect 6337 5956 6393 6012
rect 6393 5956 6397 6012
rect 6333 5952 6397 5956
rect 6413 6012 6477 6016
rect 6413 5956 6417 6012
rect 6417 5956 6473 6012
rect 6473 5956 6477 6012
rect 6413 5952 6477 5956
rect 6493 6012 6557 6016
rect 6493 5956 6497 6012
rect 6497 5956 6553 6012
rect 6553 5956 6557 6012
rect 6493 5952 6557 5956
rect 16856 6012 16920 6016
rect 16856 5956 16860 6012
rect 16860 5956 16916 6012
rect 16916 5956 16920 6012
rect 16856 5952 16920 5956
rect 16936 6012 17000 6016
rect 16936 5956 16940 6012
rect 16940 5956 16996 6012
rect 16996 5956 17000 6012
rect 16936 5952 17000 5956
rect 17016 6012 17080 6016
rect 17016 5956 17020 6012
rect 17020 5956 17076 6012
rect 17076 5956 17080 6012
rect 17016 5952 17080 5956
rect 17096 6012 17160 6016
rect 17096 5956 17100 6012
rect 17100 5956 17156 6012
rect 17156 5956 17160 6012
rect 17096 5952 17160 5956
rect 27459 6012 27523 6016
rect 27459 5956 27463 6012
rect 27463 5956 27519 6012
rect 27519 5956 27523 6012
rect 27459 5952 27523 5956
rect 27539 6012 27603 6016
rect 27539 5956 27543 6012
rect 27543 5956 27599 6012
rect 27599 5956 27603 6012
rect 27539 5952 27603 5956
rect 27619 6012 27683 6016
rect 27619 5956 27623 6012
rect 27623 5956 27679 6012
rect 27679 5956 27683 6012
rect 27619 5952 27683 5956
rect 27699 6012 27763 6016
rect 27699 5956 27703 6012
rect 27703 5956 27759 6012
rect 27759 5956 27763 6012
rect 27699 5952 27763 5956
rect 38062 6012 38126 6016
rect 38062 5956 38066 6012
rect 38066 5956 38122 6012
rect 38122 5956 38126 6012
rect 38062 5952 38126 5956
rect 38142 6012 38206 6016
rect 38142 5956 38146 6012
rect 38146 5956 38202 6012
rect 38202 5956 38206 6012
rect 38142 5952 38206 5956
rect 38222 6012 38286 6016
rect 38222 5956 38226 6012
rect 38226 5956 38282 6012
rect 38282 5956 38286 6012
rect 38222 5952 38286 5956
rect 38302 6012 38366 6016
rect 38302 5956 38306 6012
rect 38306 5956 38362 6012
rect 38362 5956 38366 6012
rect 38302 5952 38366 5956
rect 11554 5468 11618 5472
rect 11554 5412 11558 5468
rect 11558 5412 11614 5468
rect 11614 5412 11618 5468
rect 11554 5408 11618 5412
rect 11634 5468 11698 5472
rect 11634 5412 11638 5468
rect 11638 5412 11694 5468
rect 11694 5412 11698 5468
rect 11634 5408 11698 5412
rect 11714 5468 11778 5472
rect 11714 5412 11718 5468
rect 11718 5412 11774 5468
rect 11774 5412 11778 5468
rect 11714 5408 11778 5412
rect 11794 5468 11858 5472
rect 11794 5412 11798 5468
rect 11798 5412 11854 5468
rect 11854 5412 11858 5468
rect 11794 5408 11858 5412
rect 22157 5468 22221 5472
rect 22157 5412 22161 5468
rect 22161 5412 22217 5468
rect 22217 5412 22221 5468
rect 22157 5408 22221 5412
rect 22237 5468 22301 5472
rect 22237 5412 22241 5468
rect 22241 5412 22297 5468
rect 22297 5412 22301 5468
rect 22237 5408 22301 5412
rect 22317 5468 22381 5472
rect 22317 5412 22321 5468
rect 22321 5412 22377 5468
rect 22377 5412 22381 5468
rect 22317 5408 22381 5412
rect 22397 5468 22461 5472
rect 22397 5412 22401 5468
rect 22401 5412 22457 5468
rect 22457 5412 22461 5468
rect 22397 5408 22461 5412
rect 32760 5468 32824 5472
rect 32760 5412 32764 5468
rect 32764 5412 32820 5468
rect 32820 5412 32824 5468
rect 32760 5408 32824 5412
rect 32840 5468 32904 5472
rect 32840 5412 32844 5468
rect 32844 5412 32900 5468
rect 32900 5412 32904 5468
rect 32840 5408 32904 5412
rect 32920 5468 32984 5472
rect 32920 5412 32924 5468
rect 32924 5412 32980 5468
rect 32980 5412 32984 5468
rect 32920 5408 32984 5412
rect 33000 5468 33064 5472
rect 33000 5412 33004 5468
rect 33004 5412 33060 5468
rect 33060 5412 33064 5468
rect 33000 5408 33064 5412
rect 43363 5468 43427 5472
rect 43363 5412 43367 5468
rect 43367 5412 43423 5468
rect 43423 5412 43427 5468
rect 43363 5408 43427 5412
rect 43443 5468 43507 5472
rect 43443 5412 43447 5468
rect 43447 5412 43503 5468
rect 43503 5412 43507 5468
rect 43443 5408 43507 5412
rect 43523 5468 43587 5472
rect 43523 5412 43527 5468
rect 43527 5412 43583 5468
rect 43583 5412 43587 5468
rect 43523 5408 43587 5412
rect 43603 5468 43667 5472
rect 43603 5412 43607 5468
rect 43607 5412 43663 5468
rect 43663 5412 43667 5468
rect 43603 5408 43667 5412
rect 6253 4924 6317 4928
rect 6253 4868 6257 4924
rect 6257 4868 6313 4924
rect 6313 4868 6317 4924
rect 6253 4864 6317 4868
rect 6333 4924 6397 4928
rect 6333 4868 6337 4924
rect 6337 4868 6393 4924
rect 6393 4868 6397 4924
rect 6333 4864 6397 4868
rect 6413 4924 6477 4928
rect 6413 4868 6417 4924
rect 6417 4868 6473 4924
rect 6473 4868 6477 4924
rect 6413 4864 6477 4868
rect 6493 4924 6557 4928
rect 6493 4868 6497 4924
rect 6497 4868 6553 4924
rect 6553 4868 6557 4924
rect 6493 4864 6557 4868
rect 16856 4924 16920 4928
rect 16856 4868 16860 4924
rect 16860 4868 16916 4924
rect 16916 4868 16920 4924
rect 16856 4864 16920 4868
rect 16936 4924 17000 4928
rect 16936 4868 16940 4924
rect 16940 4868 16996 4924
rect 16996 4868 17000 4924
rect 16936 4864 17000 4868
rect 17016 4924 17080 4928
rect 17016 4868 17020 4924
rect 17020 4868 17076 4924
rect 17076 4868 17080 4924
rect 17016 4864 17080 4868
rect 17096 4924 17160 4928
rect 17096 4868 17100 4924
rect 17100 4868 17156 4924
rect 17156 4868 17160 4924
rect 17096 4864 17160 4868
rect 27459 4924 27523 4928
rect 27459 4868 27463 4924
rect 27463 4868 27519 4924
rect 27519 4868 27523 4924
rect 27459 4864 27523 4868
rect 27539 4924 27603 4928
rect 27539 4868 27543 4924
rect 27543 4868 27599 4924
rect 27599 4868 27603 4924
rect 27539 4864 27603 4868
rect 27619 4924 27683 4928
rect 27619 4868 27623 4924
rect 27623 4868 27679 4924
rect 27679 4868 27683 4924
rect 27619 4864 27683 4868
rect 27699 4924 27763 4928
rect 27699 4868 27703 4924
rect 27703 4868 27759 4924
rect 27759 4868 27763 4924
rect 27699 4864 27763 4868
rect 38062 4924 38126 4928
rect 38062 4868 38066 4924
rect 38066 4868 38122 4924
rect 38122 4868 38126 4924
rect 38062 4864 38126 4868
rect 38142 4924 38206 4928
rect 38142 4868 38146 4924
rect 38146 4868 38202 4924
rect 38202 4868 38206 4924
rect 38142 4864 38206 4868
rect 38222 4924 38286 4928
rect 38222 4868 38226 4924
rect 38226 4868 38282 4924
rect 38282 4868 38286 4924
rect 38222 4864 38286 4868
rect 38302 4924 38366 4928
rect 38302 4868 38306 4924
rect 38306 4868 38362 4924
rect 38362 4868 38366 4924
rect 38302 4864 38366 4868
rect 11554 4380 11618 4384
rect 11554 4324 11558 4380
rect 11558 4324 11614 4380
rect 11614 4324 11618 4380
rect 11554 4320 11618 4324
rect 11634 4380 11698 4384
rect 11634 4324 11638 4380
rect 11638 4324 11694 4380
rect 11694 4324 11698 4380
rect 11634 4320 11698 4324
rect 11714 4380 11778 4384
rect 11714 4324 11718 4380
rect 11718 4324 11774 4380
rect 11774 4324 11778 4380
rect 11714 4320 11778 4324
rect 11794 4380 11858 4384
rect 11794 4324 11798 4380
rect 11798 4324 11854 4380
rect 11854 4324 11858 4380
rect 11794 4320 11858 4324
rect 22157 4380 22221 4384
rect 22157 4324 22161 4380
rect 22161 4324 22217 4380
rect 22217 4324 22221 4380
rect 22157 4320 22221 4324
rect 22237 4380 22301 4384
rect 22237 4324 22241 4380
rect 22241 4324 22297 4380
rect 22297 4324 22301 4380
rect 22237 4320 22301 4324
rect 22317 4380 22381 4384
rect 22317 4324 22321 4380
rect 22321 4324 22377 4380
rect 22377 4324 22381 4380
rect 22317 4320 22381 4324
rect 22397 4380 22461 4384
rect 22397 4324 22401 4380
rect 22401 4324 22457 4380
rect 22457 4324 22461 4380
rect 22397 4320 22461 4324
rect 32760 4380 32824 4384
rect 32760 4324 32764 4380
rect 32764 4324 32820 4380
rect 32820 4324 32824 4380
rect 32760 4320 32824 4324
rect 32840 4380 32904 4384
rect 32840 4324 32844 4380
rect 32844 4324 32900 4380
rect 32900 4324 32904 4380
rect 32840 4320 32904 4324
rect 32920 4380 32984 4384
rect 32920 4324 32924 4380
rect 32924 4324 32980 4380
rect 32980 4324 32984 4380
rect 32920 4320 32984 4324
rect 33000 4380 33064 4384
rect 33000 4324 33004 4380
rect 33004 4324 33060 4380
rect 33060 4324 33064 4380
rect 33000 4320 33064 4324
rect 43363 4380 43427 4384
rect 43363 4324 43367 4380
rect 43367 4324 43423 4380
rect 43423 4324 43427 4380
rect 43363 4320 43427 4324
rect 43443 4380 43507 4384
rect 43443 4324 43447 4380
rect 43447 4324 43503 4380
rect 43503 4324 43507 4380
rect 43443 4320 43507 4324
rect 43523 4380 43587 4384
rect 43523 4324 43527 4380
rect 43527 4324 43583 4380
rect 43583 4324 43587 4380
rect 43523 4320 43587 4324
rect 43603 4380 43667 4384
rect 43603 4324 43607 4380
rect 43607 4324 43663 4380
rect 43663 4324 43667 4380
rect 43603 4320 43667 4324
rect 6253 3836 6317 3840
rect 6253 3780 6257 3836
rect 6257 3780 6313 3836
rect 6313 3780 6317 3836
rect 6253 3776 6317 3780
rect 6333 3836 6397 3840
rect 6333 3780 6337 3836
rect 6337 3780 6393 3836
rect 6393 3780 6397 3836
rect 6333 3776 6397 3780
rect 6413 3836 6477 3840
rect 6413 3780 6417 3836
rect 6417 3780 6473 3836
rect 6473 3780 6477 3836
rect 6413 3776 6477 3780
rect 6493 3836 6557 3840
rect 6493 3780 6497 3836
rect 6497 3780 6553 3836
rect 6553 3780 6557 3836
rect 6493 3776 6557 3780
rect 16856 3836 16920 3840
rect 16856 3780 16860 3836
rect 16860 3780 16916 3836
rect 16916 3780 16920 3836
rect 16856 3776 16920 3780
rect 16936 3836 17000 3840
rect 16936 3780 16940 3836
rect 16940 3780 16996 3836
rect 16996 3780 17000 3836
rect 16936 3776 17000 3780
rect 17016 3836 17080 3840
rect 17016 3780 17020 3836
rect 17020 3780 17076 3836
rect 17076 3780 17080 3836
rect 17016 3776 17080 3780
rect 17096 3836 17160 3840
rect 17096 3780 17100 3836
rect 17100 3780 17156 3836
rect 17156 3780 17160 3836
rect 17096 3776 17160 3780
rect 27459 3836 27523 3840
rect 27459 3780 27463 3836
rect 27463 3780 27519 3836
rect 27519 3780 27523 3836
rect 27459 3776 27523 3780
rect 27539 3836 27603 3840
rect 27539 3780 27543 3836
rect 27543 3780 27599 3836
rect 27599 3780 27603 3836
rect 27539 3776 27603 3780
rect 27619 3836 27683 3840
rect 27619 3780 27623 3836
rect 27623 3780 27679 3836
rect 27679 3780 27683 3836
rect 27619 3776 27683 3780
rect 27699 3836 27763 3840
rect 27699 3780 27703 3836
rect 27703 3780 27759 3836
rect 27759 3780 27763 3836
rect 27699 3776 27763 3780
rect 38062 3836 38126 3840
rect 38062 3780 38066 3836
rect 38066 3780 38122 3836
rect 38122 3780 38126 3836
rect 38062 3776 38126 3780
rect 38142 3836 38206 3840
rect 38142 3780 38146 3836
rect 38146 3780 38202 3836
rect 38202 3780 38206 3836
rect 38142 3776 38206 3780
rect 38222 3836 38286 3840
rect 38222 3780 38226 3836
rect 38226 3780 38282 3836
rect 38282 3780 38286 3836
rect 38222 3776 38286 3780
rect 38302 3836 38366 3840
rect 38302 3780 38306 3836
rect 38306 3780 38362 3836
rect 38362 3780 38366 3836
rect 38302 3776 38366 3780
rect 11554 3292 11618 3296
rect 11554 3236 11558 3292
rect 11558 3236 11614 3292
rect 11614 3236 11618 3292
rect 11554 3232 11618 3236
rect 11634 3292 11698 3296
rect 11634 3236 11638 3292
rect 11638 3236 11694 3292
rect 11694 3236 11698 3292
rect 11634 3232 11698 3236
rect 11714 3292 11778 3296
rect 11714 3236 11718 3292
rect 11718 3236 11774 3292
rect 11774 3236 11778 3292
rect 11714 3232 11778 3236
rect 11794 3292 11858 3296
rect 11794 3236 11798 3292
rect 11798 3236 11854 3292
rect 11854 3236 11858 3292
rect 11794 3232 11858 3236
rect 22157 3292 22221 3296
rect 22157 3236 22161 3292
rect 22161 3236 22217 3292
rect 22217 3236 22221 3292
rect 22157 3232 22221 3236
rect 22237 3292 22301 3296
rect 22237 3236 22241 3292
rect 22241 3236 22297 3292
rect 22297 3236 22301 3292
rect 22237 3232 22301 3236
rect 22317 3292 22381 3296
rect 22317 3236 22321 3292
rect 22321 3236 22377 3292
rect 22377 3236 22381 3292
rect 22317 3232 22381 3236
rect 22397 3292 22461 3296
rect 22397 3236 22401 3292
rect 22401 3236 22457 3292
rect 22457 3236 22461 3292
rect 22397 3232 22461 3236
rect 32760 3292 32824 3296
rect 32760 3236 32764 3292
rect 32764 3236 32820 3292
rect 32820 3236 32824 3292
rect 32760 3232 32824 3236
rect 32840 3292 32904 3296
rect 32840 3236 32844 3292
rect 32844 3236 32900 3292
rect 32900 3236 32904 3292
rect 32840 3232 32904 3236
rect 32920 3292 32984 3296
rect 32920 3236 32924 3292
rect 32924 3236 32980 3292
rect 32980 3236 32984 3292
rect 32920 3232 32984 3236
rect 33000 3292 33064 3296
rect 33000 3236 33004 3292
rect 33004 3236 33060 3292
rect 33060 3236 33064 3292
rect 33000 3232 33064 3236
rect 43363 3292 43427 3296
rect 43363 3236 43367 3292
rect 43367 3236 43423 3292
rect 43423 3236 43427 3292
rect 43363 3232 43427 3236
rect 43443 3292 43507 3296
rect 43443 3236 43447 3292
rect 43447 3236 43503 3292
rect 43503 3236 43507 3292
rect 43443 3232 43507 3236
rect 43523 3292 43587 3296
rect 43523 3236 43527 3292
rect 43527 3236 43583 3292
rect 43583 3236 43587 3292
rect 43523 3232 43587 3236
rect 43603 3292 43667 3296
rect 43603 3236 43607 3292
rect 43607 3236 43663 3292
rect 43663 3236 43667 3292
rect 43603 3232 43667 3236
rect 34468 2892 34532 2956
rect 6253 2748 6317 2752
rect 6253 2692 6257 2748
rect 6257 2692 6313 2748
rect 6313 2692 6317 2748
rect 6253 2688 6317 2692
rect 6333 2748 6397 2752
rect 6333 2692 6337 2748
rect 6337 2692 6393 2748
rect 6393 2692 6397 2748
rect 6333 2688 6397 2692
rect 6413 2748 6477 2752
rect 6413 2692 6417 2748
rect 6417 2692 6473 2748
rect 6473 2692 6477 2748
rect 6413 2688 6477 2692
rect 6493 2748 6557 2752
rect 6493 2692 6497 2748
rect 6497 2692 6553 2748
rect 6553 2692 6557 2748
rect 6493 2688 6557 2692
rect 16856 2748 16920 2752
rect 16856 2692 16860 2748
rect 16860 2692 16916 2748
rect 16916 2692 16920 2748
rect 16856 2688 16920 2692
rect 16936 2748 17000 2752
rect 16936 2692 16940 2748
rect 16940 2692 16996 2748
rect 16996 2692 17000 2748
rect 16936 2688 17000 2692
rect 17016 2748 17080 2752
rect 17016 2692 17020 2748
rect 17020 2692 17076 2748
rect 17076 2692 17080 2748
rect 17016 2688 17080 2692
rect 17096 2748 17160 2752
rect 17096 2692 17100 2748
rect 17100 2692 17156 2748
rect 17156 2692 17160 2748
rect 17096 2688 17160 2692
rect 27459 2748 27523 2752
rect 27459 2692 27463 2748
rect 27463 2692 27519 2748
rect 27519 2692 27523 2748
rect 27459 2688 27523 2692
rect 27539 2748 27603 2752
rect 27539 2692 27543 2748
rect 27543 2692 27599 2748
rect 27599 2692 27603 2748
rect 27539 2688 27603 2692
rect 27619 2748 27683 2752
rect 27619 2692 27623 2748
rect 27623 2692 27679 2748
rect 27679 2692 27683 2748
rect 27619 2688 27683 2692
rect 27699 2748 27763 2752
rect 27699 2692 27703 2748
rect 27703 2692 27759 2748
rect 27759 2692 27763 2748
rect 27699 2688 27763 2692
rect 38062 2748 38126 2752
rect 38062 2692 38066 2748
rect 38066 2692 38122 2748
rect 38122 2692 38126 2748
rect 38062 2688 38126 2692
rect 38142 2748 38206 2752
rect 38142 2692 38146 2748
rect 38146 2692 38202 2748
rect 38202 2692 38206 2748
rect 38142 2688 38206 2692
rect 38222 2748 38286 2752
rect 38222 2692 38226 2748
rect 38226 2692 38282 2748
rect 38282 2692 38286 2748
rect 38222 2688 38286 2692
rect 38302 2748 38366 2752
rect 38302 2692 38306 2748
rect 38306 2692 38362 2748
rect 38362 2692 38366 2748
rect 38302 2688 38366 2692
rect 11554 2204 11618 2208
rect 11554 2148 11558 2204
rect 11558 2148 11614 2204
rect 11614 2148 11618 2204
rect 11554 2144 11618 2148
rect 11634 2204 11698 2208
rect 11634 2148 11638 2204
rect 11638 2148 11694 2204
rect 11694 2148 11698 2204
rect 11634 2144 11698 2148
rect 11714 2204 11778 2208
rect 11714 2148 11718 2204
rect 11718 2148 11774 2204
rect 11774 2148 11778 2204
rect 11714 2144 11778 2148
rect 11794 2204 11858 2208
rect 11794 2148 11798 2204
rect 11798 2148 11854 2204
rect 11854 2148 11858 2204
rect 11794 2144 11858 2148
rect 22157 2204 22221 2208
rect 22157 2148 22161 2204
rect 22161 2148 22217 2204
rect 22217 2148 22221 2204
rect 22157 2144 22221 2148
rect 22237 2204 22301 2208
rect 22237 2148 22241 2204
rect 22241 2148 22297 2204
rect 22297 2148 22301 2204
rect 22237 2144 22301 2148
rect 22317 2204 22381 2208
rect 22317 2148 22321 2204
rect 22321 2148 22377 2204
rect 22377 2148 22381 2204
rect 22317 2144 22381 2148
rect 22397 2204 22461 2208
rect 22397 2148 22401 2204
rect 22401 2148 22457 2204
rect 22457 2148 22461 2204
rect 22397 2144 22461 2148
rect 32760 2204 32824 2208
rect 32760 2148 32764 2204
rect 32764 2148 32820 2204
rect 32820 2148 32824 2204
rect 32760 2144 32824 2148
rect 32840 2204 32904 2208
rect 32840 2148 32844 2204
rect 32844 2148 32900 2204
rect 32900 2148 32904 2204
rect 32840 2144 32904 2148
rect 32920 2204 32984 2208
rect 32920 2148 32924 2204
rect 32924 2148 32980 2204
rect 32980 2148 32984 2204
rect 32920 2144 32984 2148
rect 33000 2204 33064 2208
rect 33000 2148 33004 2204
rect 33004 2148 33060 2204
rect 33060 2148 33064 2204
rect 33000 2144 33064 2148
rect 43363 2204 43427 2208
rect 43363 2148 43367 2204
rect 43367 2148 43423 2204
rect 43423 2148 43427 2204
rect 43363 2144 43427 2148
rect 43443 2204 43507 2208
rect 43443 2148 43447 2204
rect 43447 2148 43503 2204
rect 43503 2148 43507 2204
rect 43443 2144 43507 2148
rect 43523 2204 43587 2208
rect 43523 2148 43527 2204
rect 43527 2148 43583 2204
rect 43583 2148 43587 2204
rect 43523 2144 43587 2148
rect 43603 2204 43667 2208
rect 43603 2148 43607 2204
rect 43607 2148 43663 2204
rect 43663 2148 43667 2204
rect 43603 2144 43667 2148
rect 6253 1660 6317 1664
rect 6253 1604 6257 1660
rect 6257 1604 6313 1660
rect 6313 1604 6317 1660
rect 6253 1600 6317 1604
rect 6333 1660 6397 1664
rect 6333 1604 6337 1660
rect 6337 1604 6393 1660
rect 6393 1604 6397 1660
rect 6333 1600 6397 1604
rect 6413 1660 6477 1664
rect 6413 1604 6417 1660
rect 6417 1604 6473 1660
rect 6473 1604 6477 1660
rect 6413 1600 6477 1604
rect 6493 1660 6557 1664
rect 6493 1604 6497 1660
rect 6497 1604 6553 1660
rect 6553 1604 6557 1660
rect 6493 1600 6557 1604
rect 16856 1660 16920 1664
rect 16856 1604 16860 1660
rect 16860 1604 16916 1660
rect 16916 1604 16920 1660
rect 16856 1600 16920 1604
rect 16936 1660 17000 1664
rect 16936 1604 16940 1660
rect 16940 1604 16996 1660
rect 16996 1604 17000 1660
rect 16936 1600 17000 1604
rect 17016 1660 17080 1664
rect 17016 1604 17020 1660
rect 17020 1604 17076 1660
rect 17076 1604 17080 1660
rect 17016 1600 17080 1604
rect 17096 1660 17160 1664
rect 17096 1604 17100 1660
rect 17100 1604 17156 1660
rect 17156 1604 17160 1660
rect 17096 1600 17160 1604
rect 27459 1660 27523 1664
rect 27459 1604 27463 1660
rect 27463 1604 27519 1660
rect 27519 1604 27523 1660
rect 27459 1600 27523 1604
rect 27539 1660 27603 1664
rect 27539 1604 27543 1660
rect 27543 1604 27599 1660
rect 27599 1604 27603 1660
rect 27539 1600 27603 1604
rect 27619 1660 27683 1664
rect 27619 1604 27623 1660
rect 27623 1604 27679 1660
rect 27679 1604 27683 1660
rect 27619 1600 27683 1604
rect 27699 1660 27763 1664
rect 27699 1604 27703 1660
rect 27703 1604 27759 1660
rect 27759 1604 27763 1660
rect 27699 1600 27763 1604
rect 38062 1660 38126 1664
rect 38062 1604 38066 1660
rect 38066 1604 38122 1660
rect 38122 1604 38126 1660
rect 38062 1600 38126 1604
rect 38142 1660 38206 1664
rect 38142 1604 38146 1660
rect 38146 1604 38202 1660
rect 38202 1604 38206 1660
rect 38142 1600 38206 1604
rect 38222 1660 38286 1664
rect 38222 1604 38226 1660
rect 38226 1604 38282 1660
rect 38282 1604 38286 1660
rect 38222 1600 38286 1604
rect 38302 1660 38366 1664
rect 38302 1604 38306 1660
rect 38306 1604 38362 1660
rect 38362 1604 38366 1660
rect 38302 1600 38366 1604
rect 11554 1116 11618 1120
rect 11554 1060 11558 1116
rect 11558 1060 11614 1116
rect 11614 1060 11618 1116
rect 11554 1056 11618 1060
rect 11634 1116 11698 1120
rect 11634 1060 11638 1116
rect 11638 1060 11694 1116
rect 11694 1060 11698 1116
rect 11634 1056 11698 1060
rect 11714 1116 11778 1120
rect 11714 1060 11718 1116
rect 11718 1060 11774 1116
rect 11774 1060 11778 1116
rect 11714 1056 11778 1060
rect 11794 1116 11858 1120
rect 11794 1060 11798 1116
rect 11798 1060 11854 1116
rect 11854 1060 11858 1116
rect 11794 1056 11858 1060
rect 22157 1116 22221 1120
rect 22157 1060 22161 1116
rect 22161 1060 22217 1116
rect 22217 1060 22221 1116
rect 22157 1056 22221 1060
rect 22237 1116 22301 1120
rect 22237 1060 22241 1116
rect 22241 1060 22297 1116
rect 22297 1060 22301 1116
rect 22237 1056 22301 1060
rect 22317 1116 22381 1120
rect 22317 1060 22321 1116
rect 22321 1060 22377 1116
rect 22377 1060 22381 1116
rect 22317 1056 22381 1060
rect 22397 1116 22461 1120
rect 22397 1060 22401 1116
rect 22401 1060 22457 1116
rect 22457 1060 22461 1116
rect 22397 1056 22461 1060
rect 32760 1116 32824 1120
rect 32760 1060 32764 1116
rect 32764 1060 32820 1116
rect 32820 1060 32824 1116
rect 32760 1056 32824 1060
rect 32840 1116 32904 1120
rect 32840 1060 32844 1116
rect 32844 1060 32900 1116
rect 32900 1060 32904 1116
rect 32840 1056 32904 1060
rect 32920 1116 32984 1120
rect 32920 1060 32924 1116
rect 32924 1060 32980 1116
rect 32980 1060 32984 1116
rect 32920 1056 32984 1060
rect 33000 1116 33064 1120
rect 33000 1060 33004 1116
rect 33004 1060 33060 1116
rect 33060 1060 33064 1116
rect 33000 1056 33064 1060
rect 43363 1116 43427 1120
rect 43363 1060 43367 1116
rect 43367 1060 43423 1116
rect 43423 1060 43427 1116
rect 43363 1056 43427 1060
rect 43443 1116 43507 1120
rect 43443 1060 43447 1116
rect 43447 1060 43503 1116
rect 43503 1060 43507 1116
rect 43443 1056 43507 1060
rect 43523 1116 43587 1120
rect 43523 1060 43527 1116
rect 43527 1060 43583 1116
rect 43583 1060 43587 1116
rect 43523 1056 43587 1060
rect 43603 1116 43667 1120
rect 43603 1060 43607 1116
rect 43607 1060 43663 1116
rect 43663 1060 43667 1116
rect 43603 1056 43667 1060
<< metal4 >>
rect 19563 9892 19629 9893
rect 19563 9828 19564 9892
rect 19628 9828 19629 9892
rect 19563 9827 19629 9828
rect 6245 8192 6565 8752
rect 6245 8128 6253 8192
rect 6317 8128 6333 8192
rect 6397 8128 6413 8192
rect 6477 8128 6493 8192
rect 6557 8128 6565 8192
rect 6245 7104 6565 8128
rect 6245 7040 6253 7104
rect 6317 7040 6333 7104
rect 6397 7040 6413 7104
rect 6477 7040 6493 7104
rect 6557 7040 6565 7104
rect 6245 6016 6565 7040
rect 6245 5952 6253 6016
rect 6317 5952 6333 6016
rect 6397 5952 6413 6016
rect 6477 5952 6493 6016
rect 6557 5952 6565 6016
rect 6245 4928 6565 5952
rect 6245 4864 6253 4928
rect 6317 4864 6333 4928
rect 6397 4864 6413 4928
rect 6477 4864 6493 4928
rect 6557 4864 6565 4928
rect 6245 3840 6565 4864
rect 6245 3776 6253 3840
rect 6317 3776 6333 3840
rect 6397 3776 6413 3840
rect 6477 3776 6493 3840
rect 6557 3776 6565 3840
rect 6245 2752 6565 3776
rect 6245 2688 6253 2752
rect 6317 2688 6333 2752
rect 6397 2688 6413 2752
rect 6477 2688 6493 2752
rect 6557 2688 6565 2752
rect 6245 1664 6565 2688
rect 6245 1600 6253 1664
rect 6317 1600 6333 1664
rect 6397 1600 6413 1664
rect 6477 1600 6493 1664
rect 6557 1600 6565 1664
rect 6245 1040 6565 1600
rect 11546 8736 11866 8752
rect 11546 8672 11554 8736
rect 11618 8672 11634 8736
rect 11698 8672 11714 8736
rect 11778 8672 11794 8736
rect 11858 8672 11866 8736
rect 11546 7648 11866 8672
rect 11546 7584 11554 7648
rect 11618 7584 11634 7648
rect 11698 7584 11714 7648
rect 11778 7584 11794 7648
rect 11858 7584 11866 7648
rect 11546 6560 11866 7584
rect 11546 6496 11554 6560
rect 11618 6496 11634 6560
rect 11698 6496 11714 6560
rect 11778 6496 11794 6560
rect 11858 6496 11866 6560
rect 11546 5472 11866 6496
rect 11546 5408 11554 5472
rect 11618 5408 11634 5472
rect 11698 5408 11714 5472
rect 11778 5408 11794 5472
rect 11858 5408 11866 5472
rect 11546 4384 11866 5408
rect 11546 4320 11554 4384
rect 11618 4320 11634 4384
rect 11698 4320 11714 4384
rect 11778 4320 11794 4384
rect 11858 4320 11866 4384
rect 11546 3296 11866 4320
rect 11546 3232 11554 3296
rect 11618 3232 11634 3296
rect 11698 3232 11714 3296
rect 11778 3232 11794 3296
rect 11858 3232 11866 3296
rect 11546 2208 11866 3232
rect 11546 2144 11554 2208
rect 11618 2144 11634 2208
rect 11698 2144 11714 2208
rect 11778 2144 11794 2208
rect 11858 2144 11866 2208
rect 11546 1120 11866 2144
rect 11546 1056 11554 1120
rect 11618 1056 11634 1120
rect 11698 1056 11714 1120
rect 11778 1056 11794 1120
rect 11858 1056 11866 1120
rect 11546 1040 11866 1056
rect 16848 8192 17168 8752
rect 19379 8396 19445 8397
rect 19379 8332 19380 8396
rect 19444 8332 19445 8396
rect 19379 8331 19445 8332
rect 16848 8128 16856 8192
rect 16920 8128 16936 8192
rect 17000 8128 17016 8192
rect 17080 8128 17096 8192
rect 17160 8128 17168 8192
rect 16848 7104 17168 8128
rect 19382 7717 19442 8331
rect 19379 7716 19445 7717
rect 19379 7652 19380 7716
rect 19444 7652 19445 7716
rect 19379 7651 19445 7652
rect 19566 7445 19626 9827
rect 22149 8736 22469 8752
rect 22149 8672 22157 8736
rect 22221 8672 22237 8736
rect 22301 8672 22317 8736
rect 22381 8672 22397 8736
rect 22461 8672 22469 8736
rect 22149 7648 22469 8672
rect 22149 7584 22157 7648
rect 22221 7584 22237 7648
rect 22301 7584 22317 7648
rect 22381 7584 22397 7648
rect 22461 7584 22469 7648
rect 19563 7444 19629 7445
rect 19563 7380 19564 7444
rect 19628 7380 19629 7444
rect 19563 7379 19629 7380
rect 16848 7040 16856 7104
rect 16920 7040 16936 7104
rect 17000 7040 17016 7104
rect 17080 7040 17096 7104
rect 17160 7040 17168 7104
rect 16848 6016 17168 7040
rect 16848 5952 16856 6016
rect 16920 5952 16936 6016
rect 17000 5952 17016 6016
rect 17080 5952 17096 6016
rect 17160 5952 17168 6016
rect 16848 4928 17168 5952
rect 16848 4864 16856 4928
rect 16920 4864 16936 4928
rect 17000 4864 17016 4928
rect 17080 4864 17096 4928
rect 17160 4864 17168 4928
rect 16848 3840 17168 4864
rect 16848 3776 16856 3840
rect 16920 3776 16936 3840
rect 17000 3776 17016 3840
rect 17080 3776 17096 3840
rect 17160 3776 17168 3840
rect 16848 2752 17168 3776
rect 16848 2688 16856 2752
rect 16920 2688 16936 2752
rect 17000 2688 17016 2752
rect 17080 2688 17096 2752
rect 17160 2688 17168 2752
rect 16848 1664 17168 2688
rect 16848 1600 16856 1664
rect 16920 1600 16936 1664
rect 17000 1600 17016 1664
rect 17080 1600 17096 1664
rect 17160 1600 17168 1664
rect 16848 1040 17168 1600
rect 22149 6560 22469 7584
rect 22149 6496 22157 6560
rect 22221 6496 22237 6560
rect 22301 6496 22317 6560
rect 22381 6496 22397 6560
rect 22461 6496 22469 6560
rect 22149 5472 22469 6496
rect 22149 5408 22157 5472
rect 22221 5408 22237 5472
rect 22301 5408 22317 5472
rect 22381 5408 22397 5472
rect 22461 5408 22469 5472
rect 22149 4384 22469 5408
rect 22149 4320 22157 4384
rect 22221 4320 22237 4384
rect 22301 4320 22317 4384
rect 22381 4320 22397 4384
rect 22461 4320 22469 4384
rect 22149 3296 22469 4320
rect 22149 3232 22157 3296
rect 22221 3232 22237 3296
rect 22301 3232 22317 3296
rect 22381 3232 22397 3296
rect 22461 3232 22469 3296
rect 22149 2208 22469 3232
rect 22149 2144 22157 2208
rect 22221 2144 22237 2208
rect 22301 2144 22317 2208
rect 22381 2144 22397 2208
rect 22461 2144 22469 2208
rect 22149 1120 22469 2144
rect 22149 1056 22157 1120
rect 22221 1056 22237 1120
rect 22301 1056 22317 1120
rect 22381 1056 22397 1120
rect 22461 1056 22469 1120
rect 22149 1040 22469 1056
rect 27451 8192 27771 8752
rect 27451 8128 27459 8192
rect 27523 8128 27539 8192
rect 27603 8128 27619 8192
rect 27683 8128 27699 8192
rect 27763 8128 27771 8192
rect 27451 7104 27771 8128
rect 27451 7040 27459 7104
rect 27523 7040 27539 7104
rect 27603 7040 27619 7104
rect 27683 7040 27699 7104
rect 27763 7040 27771 7104
rect 27451 6016 27771 7040
rect 27451 5952 27459 6016
rect 27523 5952 27539 6016
rect 27603 5952 27619 6016
rect 27683 5952 27699 6016
rect 27763 5952 27771 6016
rect 27451 4928 27771 5952
rect 27451 4864 27459 4928
rect 27523 4864 27539 4928
rect 27603 4864 27619 4928
rect 27683 4864 27699 4928
rect 27763 4864 27771 4928
rect 27451 3840 27771 4864
rect 27451 3776 27459 3840
rect 27523 3776 27539 3840
rect 27603 3776 27619 3840
rect 27683 3776 27699 3840
rect 27763 3776 27771 3840
rect 27451 2752 27771 3776
rect 27451 2688 27459 2752
rect 27523 2688 27539 2752
rect 27603 2688 27619 2752
rect 27683 2688 27699 2752
rect 27763 2688 27771 2752
rect 27451 1664 27771 2688
rect 27451 1600 27459 1664
rect 27523 1600 27539 1664
rect 27603 1600 27619 1664
rect 27683 1600 27699 1664
rect 27763 1600 27771 1664
rect 27451 1040 27771 1600
rect 32752 8736 33072 8752
rect 32752 8672 32760 8736
rect 32824 8672 32840 8736
rect 32904 8672 32920 8736
rect 32984 8672 33000 8736
rect 33064 8672 33072 8736
rect 32752 7648 33072 8672
rect 34467 8396 34533 8397
rect 34467 8332 34468 8396
rect 34532 8332 34533 8396
rect 34467 8331 34533 8332
rect 32752 7584 32760 7648
rect 32824 7584 32840 7648
rect 32904 7584 32920 7648
rect 32984 7584 33000 7648
rect 33064 7584 33072 7648
rect 32752 6560 33072 7584
rect 32752 6496 32760 6560
rect 32824 6496 32840 6560
rect 32904 6496 32920 6560
rect 32984 6496 33000 6560
rect 33064 6496 33072 6560
rect 32752 5472 33072 6496
rect 32752 5408 32760 5472
rect 32824 5408 32840 5472
rect 32904 5408 32920 5472
rect 32984 5408 33000 5472
rect 33064 5408 33072 5472
rect 32752 4384 33072 5408
rect 32752 4320 32760 4384
rect 32824 4320 32840 4384
rect 32904 4320 32920 4384
rect 32984 4320 33000 4384
rect 33064 4320 33072 4384
rect 32752 3296 33072 4320
rect 32752 3232 32760 3296
rect 32824 3232 32840 3296
rect 32904 3232 32920 3296
rect 32984 3232 33000 3296
rect 33064 3232 33072 3296
rect 32752 2208 33072 3232
rect 34470 2957 34530 8331
rect 38054 8192 38374 8752
rect 38054 8128 38062 8192
rect 38126 8128 38142 8192
rect 38206 8128 38222 8192
rect 38286 8128 38302 8192
rect 38366 8128 38374 8192
rect 38054 7104 38374 8128
rect 38054 7040 38062 7104
rect 38126 7040 38142 7104
rect 38206 7040 38222 7104
rect 38286 7040 38302 7104
rect 38366 7040 38374 7104
rect 38054 6016 38374 7040
rect 38054 5952 38062 6016
rect 38126 5952 38142 6016
rect 38206 5952 38222 6016
rect 38286 5952 38302 6016
rect 38366 5952 38374 6016
rect 38054 4928 38374 5952
rect 38054 4864 38062 4928
rect 38126 4864 38142 4928
rect 38206 4864 38222 4928
rect 38286 4864 38302 4928
rect 38366 4864 38374 4928
rect 38054 3840 38374 4864
rect 38054 3776 38062 3840
rect 38126 3776 38142 3840
rect 38206 3776 38222 3840
rect 38286 3776 38302 3840
rect 38366 3776 38374 3840
rect 34467 2956 34533 2957
rect 34467 2892 34468 2956
rect 34532 2892 34533 2956
rect 34467 2891 34533 2892
rect 32752 2144 32760 2208
rect 32824 2144 32840 2208
rect 32904 2144 32920 2208
rect 32984 2144 33000 2208
rect 33064 2144 33072 2208
rect 32752 1120 33072 2144
rect 32752 1056 32760 1120
rect 32824 1056 32840 1120
rect 32904 1056 32920 1120
rect 32984 1056 33000 1120
rect 33064 1056 33072 1120
rect 32752 1040 33072 1056
rect 38054 2752 38374 3776
rect 38054 2688 38062 2752
rect 38126 2688 38142 2752
rect 38206 2688 38222 2752
rect 38286 2688 38302 2752
rect 38366 2688 38374 2752
rect 38054 1664 38374 2688
rect 38054 1600 38062 1664
rect 38126 1600 38142 1664
rect 38206 1600 38222 1664
rect 38286 1600 38302 1664
rect 38366 1600 38374 1664
rect 38054 1040 38374 1600
rect 43355 8736 43675 8752
rect 43355 8672 43363 8736
rect 43427 8672 43443 8736
rect 43507 8672 43523 8736
rect 43587 8672 43603 8736
rect 43667 8672 43675 8736
rect 43355 7648 43675 8672
rect 43355 7584 43363 7648
rect 43427 7584 43443 7648
rect 43507 7584 43523 7648
rect 43587 7584 43603 7648
rect 43667 7584 43675 7648
rect 43355 6560 43675 7584
rect 43355 6496 43363 6560
rect 43427 6496 43443 6560
rect 43507 6496 43523 6560
rect 43587 6496 43603 6560
rect 43667 6496 43675 6560
rect 43355 5472 43675 6496
rect 43355 5408 43363 5472
rect 43427 5408 43443 5472
rect 43507 5408 43523 5472
rect 43587 5408 43603 5472
rect 43667 5408 43675 5472
rect 43355 4384 43675 5408
rect 43355 4320 43363 4384
rect 43427 4320 43443 4384
rect 43507 4320 43523 4384
rect 43587 4320 43603 4384
rect 43667 4320 43675 4384
rect 43355 3296 43675 4320
rect 43355 3232 43363 3296
rect 43427 3232 43443 3296
rect 43507 3232 43523 3296
rect 43587 3232 43603 3296
rect 43667 3232 43675 3296
rect 43355 2208 43675 3232
rect 43355 2144 43363 2208
rect 43427 2144 43443 2208
rect 43507 2144 43523 2208
rect 43587 2144 43603 2208
rect 43667 2144 43675 2208
rect 43355 1120 43675 2144
rect 43355 1056 43363 1120
rect 43427 1056 43443 1120
rect 43507 1056 43523 1120
rect 43587 1056 43603 1120
rect 43667 1056 43675 1120
rect 43355 1040 43675 1056
use sky130_ef_sc_hd__decap_12  FILLER_0_0_6 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1656 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_18 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 2760 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3588 0 1 1088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_29
timestamp 1688980957
transform 1 0 3772 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_41
timestamp 1688980957
transform 1 0 4876 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_50
timestamp 1688980957
transform 1 0 5704 0 1 1088
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_57
timestamp 1688980957
transform 1 0 6348 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_69
timestamp 1688980957
transform 1 0 7452 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_73 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 7820 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_81 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 8556 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_85
timestamp 1688980957
transform 1 0 8924 0 1 1088
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_96
timestamp 1688980957
transform 1 0 9936 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_108 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 11040 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_113
timestamp 1688980957
transform 1 0 11500 0 1 1088
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_119
timestamp 1688980957
transform 1 0 12052 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_131
timestamp 1688980957
transform 1 0 13156 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_139
timestamp 1688980957
transform 1 0 13892 0 1 1088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_144
timestamp 1688980957
transform 1 0 14352 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_156
timestamp 1688980957
transform 1 0 15456 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_165
timestamp 1688980957
transform 1 0 16284 0 1 1088
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_169
timestamp 1688980957
transform 1 0 16652 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_181
timestamp 1688980957
transform 1 0 17756 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_188
timestamp 1688980957
transform 1 0 18400 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_197
timestamp 1688980957
transform 1 0 19228 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_205
timestamp 1688980957
transform 1 0 19964 0 1 1088
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_211
timestamp 1688980957
transform 1 0 20516 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_223
timestamp 1688980957
transform 1 0 21620 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_225
timestamp 1688980957
transform 1 0 21804 0 1 1088
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_234
timestamp 1688980957
transform 1 0 22632 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_246
timestamp 1688980957
transform 1 0 23736 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_253
timestamp 1688980957
transform 1 0 24380 0 1 1088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_257
timestamp 1688980957
transform 1 0 24748 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_269
timestamp 1688980957
transform 1 0 25852 0 1 1088
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_281
timestamp 1688980957
transform 1 0 26956 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_293
timestamp 1688980957
transform 1 0 28060 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_299
timestamp 1688980957
transform 1 0 28612 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_303
timestamp 1688980957
transform 1 0 28980 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_307
timestamp 1688980957
transform 1 0 29348 0 1 1088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_309
timestamp 1688980957
transform 1 0 29532 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_321 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 30636 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_326
timestamp 1688980957
transform 1 0 31096 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_334
timestamp 1688980957
transform 1 0 31832 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_337
timestamp 1688980957
transform 1 0 32108 0 1 1088
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_345
timestamp 1688980957
transform 1 0 32844 0 1 1088
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_349
timestamp 1688980957
transform 1 0 33212 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_361
timestamp 1688980957
transform 1 0 34316 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_365
timestamp 1688980957
transform 1 0 34684 0 1 1088
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_372
timestamp 1688980957
transform 1 0 35328 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_0_384
timestamp 1688980957
transform 1 0 36432 0 1 1088
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_396
timestamp 1688980957
transform 1 0 37536 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_408
timestamp 1688980957
transform 1 0 38640 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_414
timestamp 1688980957
transform 1 0 39192 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_418
timestamp 1688980957
transform 1 0 39560 0 1 1088
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_421
timestamp 1688980957
transform 1 0 39836 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_0_433
timestamp 1688980957
transform 1 0 40940 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_437
timestamp 1688980957
transform 1 0 41308 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_441
timestamp 1688980957
transform 1 0 41676 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_447
timestamp 1688980957
transform 1 0 42228 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_449
timestamp 1688980957
transform 1 0 42412 0 1 1088
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 1688980957
transform 1 0 1380 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 1688980957
transform 1 0 2484 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_27
timestamp 1688980957
transform 1 0 3588 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_39
timestamp 1688980957
transform 1 0 4692 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_51
timestamp 1688980957
transform 1 0 5796 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 1688980957
transform 1 0 6164 0 -1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_57
timestamp 1688980957
transform 1 0 6348 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_69
timestamp 1688980957
transform 1 0 7452 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_81
timestamp 1688980957
transform 1 0 8556 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_93
timestamp 1688980957
transform 1 0 9660 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_105
timestamp 1688980957
transform 1 0 10764 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_111
timestamp 1688980957
transform 1 0 11316 0 -1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_113
timestamp 1688980957
transform 1 0 11500 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_125
timestamp 1688980957
transform 1 0 12604 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_137
timestamp 1688980957
transform 1 0 13708 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_149
timestamp 1688980957
transform 1 0 14812 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_161
timestamp 1688980957
transform 1 0 15916 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_167
timestamp 1688980957
transform 1 0 16468 0 -1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_169
timestamp 1688980957
transform 1 0 16652 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_181
timestamp 1688980957
transform 1 0 17756 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_193
timestamp 1688980957
transform 1 0 18860 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_205
timestamp 1688980957
transform 1 0 19964 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_217
timestamp 1688980957
transform 1 0 21068 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_223
timestamp 1688980957
transform 1 0 21620 0 -1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_225
timestamp 1688980957
transform 1 0 21804 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_237
timestamp 1688980957
transform 1 0 22908 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_249
timestamp 1688980957
transform 1 0 24012 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_261
timestamp 1688980957
transform 1 0 25116 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_273
timestamp 1688980957
transform 1 0 26220 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_279
timestamp 1688980957
transform 1 0 26772 0 -1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_281
timestamp 1688980957
transform 1 0 26956 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_293
timestamp 1688980957
transform 1 0 28060 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_305
timestamp 1688980957
transform 1 0 29164 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_317
timestamp 1688980957
transform 1 0 30268 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_329
timestamp 1688980957
transform 1 0 31372 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_335
timestamp 1688980957
transform 1 0 31924 0 -1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_337
timestamp 1688980957
transform 1 0 32108 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_349
timestamp 1688980957
transform 1 0 33212 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_361
timestamp 1688980957
transform 1 0 34316 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_373
timestamp 1688980957
transform 1 0 35420 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_385
timestamp 1688980957
transform 1 0 36524 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_391
timestamp 1688980957
transform 1 0 37076 0 -1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_393
timestamp 1688980957
transform 1 0 37260 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_405
timestamp 1688980957
transform 1 0 38364 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_409
timestamp 1688980957
transform 1 0 38732 0 -1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_413
timestamp 1688980957
transform 1 0 39100 0 -1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_425
timestamp 1688980957
transform 1 0 40204 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_437
timestamp 1688980957
transform 1 0 41308 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_445
timestamp 1688980957
transform 1 0 42044 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_1_449
timestamp 1688980957
transform 1 0 42412 0 -1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_457
timestamp 1688980957
transform 1 0 43148 0 -1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1688980957
transform 1 0 1380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 1688980957
transform 1 0 2484 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1688980957
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_29
timestamp 1688980957
transform 1 0 3772 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_41
timestamp 1688980957
transform 1 0 4876 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_53
timestamp 1688980957
transform 1 0 5980 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_65
timestamp 1688980957
transform 1 0 7084 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_77
timestamp 1688980957
transform 1 0 8188 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_83
timestamp 1688980957
transform 1 0 8740 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_85
timestamp 1688980957
transform 1 0 8924 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_97
timestamp 1688980957
transform 1 0 10028 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_109
timestamp 1688980957
transform 1 0 11132 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_121
timestamp 1688980957
transform 1 0 12236 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_133
timestamp 1688980957
transform 1 0 13340 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_139
timestamp 1688980957
transform 1 0 13892 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_141
timestamp 1688980957
transform 1 0 14076 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_153
timestamp 1688980957
transform 1 0 15180 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_165
timestamp 1688980957
transform 1 0 16284 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_177
timestamp 1688980957
transform 1 0 17388 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_189
timestamp 1688980957
transform 1 0 18492 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_195
timestamp 1688980957
transform 1 0 19044 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_197
timestamp 1688980957
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_209
timestamp 1688980957
transform 1 0 20332 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_221
timestamp 1688980957
transform 1 0 21436 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_225
timestamp 1688980957
transform 1 0 21804 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_229
timestamp 1688980957
transform 1 0 22172 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_241
timestamp 1688980957
transform 1 0 23276 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_249
timestamp 1688980957
transform 1 0 24012 0 1 2176
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_253
timestamp 1688980957
transform 1 0 24380 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_265
timestamp 1688980957
transform 1 0 25484 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_277
timestamp 1688980957
transform 1 0 26588 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_289
timestamp 1688980957
transform 1 0 27692 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_301
timestamp 1688980957
transform 1 0 28796 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_307
timestamp 1688980957
transform 1 0 29348 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_309
timestamp 1688980957
transform 1 0 29532 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_321
timestamp 1688980957
transform 1 0 30636 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_333
timestamp 1688980957
transform 1 0 31740 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_345
timestamp 1688980957
transform 1 0 32844 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_357
timestamp 1688980957
transform 1 0 33948 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_363
timestamp 1688980957
transform 1 0 34500 0 1 2176
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_365
timestamp 1688980957
transform 1 0 34684 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_377
timestamp 1688980957
transform 1 0 35788 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_389
timestamp 1688980957
transform 1 0 36892 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_401
timestamp 1688980957
transform 1 0 37996 0 1 2176
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_409
timestamp 1688980957
transform 1 0 38732 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_415
timestamp 1688980957
transform 1 0 39284 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_419
timestamp 1688980957
transform 1 0 39652 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_421
timestamp 1688980957
transform 1 0 39836 0 1 2176
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_428
timestamp 1688980957
transform 1 0 40480 0 1 2176
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_440
timestamp 1688980957
transform 1 0 41584 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_2_452
timestamp 1688980957
transform 1 0 42688 0 1 2176
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_3
timestamp 1688980957
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_15
timestamp 1688980957
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_27
timestamp 1688980957
transform 1 0 3588 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_39
timestamp 1688980957
transform 1 0 4692 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_51
timestamp 1688980957
transform 1 0 5796 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_55
timestamp 1688980957
transform 1 0 6164 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_57
timestamp 1688980957
transform 1 0 6348 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_69
timestamp 1688980957
transform 1 0 7452 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_81
timestamp 1688980957
transform 1 0 8556 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_93
timestamp 1688980957
transform 1 0 9660 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_105
timestamp 1688980957
transform 1 0 10764 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_111
timestamp 1688980957
transform 1 0 11316 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_113
timestamp 1688980957
transform 1 0 11500 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_125
timestamp 1688980957
transform 1 0 12604 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_137
timestamp 1688980957
transform 1 0 13708 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_149
timestamp 1688980957
transform 1 0 14812 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_161
timestamp 1688980957
transform 1 0 15916 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_167
timestamp 1688980957
transform 1 0 16468 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_169
timestamp 1688980957
transform 1 0 16652 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_181
timestamp 1688980957
transform 1 0 17756 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_189
timestamp 1688980957
transform 1 0 18492 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_193
timestamp 1688980957
transform 1 0 18860 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_205
timestamp 1688980957
transform 1 0 19964 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_223
timestamp 1688980957
transform 1 0 21620 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_225
timestamp 1688980957
transform 1 0 21804 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_233
timestamp 1688980957
transform 1 0 22540 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_237
timestamp 1688980957
transform 1 0 22908 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_249
timestamp 1688980957
transform 1 0 24012 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_261
timestamp 1688980957
transform 1 0 25116 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_273
timestamp 1688980957
transform 1 0 26220 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_279
timestamp 1688980957
transform 1 0 26772 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_281
timestamp 1688980957
transform 1 0 26956 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_293
timestamp 1688980957
transform 1 0 28060 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_308
timestamp 1688980957
transform 1 0 29440 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_320
timestamp 1688980957
transform 1 0 30544 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_3_332
timestamp 1688980957
transform 1 0 31648 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_337
timestamp 1688980957
transform 1 0 32108 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_349
timestamp 1688980957
transform 1 0 33212 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_361
timestamp 1688980957
transform 1 0 34316 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_373
timestamp 1688980957
transform 1 0 35420 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_382
timestamp 1688980957
transform 1 0 36248 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_390
timestamp 1688980957
transform 1 0 36984 0 -1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_393
timestamp 1688980957
transform 1 0 37260 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_405
timestamp 1688980957
transform 1 0 38364 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_417
timestamp 1688980957
transform 1 0 39468 0 -1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_423
timestamp 1688980957
transform 1 0 40020 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_435
timestamp 1688980957
transform 1 0 41124 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_447
timestamp 1688980957
transform 1 0 42228 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_449
timestamp 1688980957
transform 1 0 42412 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_457
timestamp 1688980957
transform 1 0 43148 0 -1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1688980957
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 1688980957
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1688980957
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 1688980957
transform 1 0 3772 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_41
timestamp 1688980957
transform 1 0 4876 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_53
timestamp 1688980957
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_65
timestamp 1688980957
transform 1 0 7084 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_77
timestamp 1688980957
transform 1 0 8188 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_83
timestamp 1688980957
transform 1 0 8740 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_85
timestamp 1688980957
transform 1 0 8924 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_97
timestamp 1688980957
transform 1 0 10028 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_109
timestamp 1688980957
transform 1 0 11132 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_121
timestamp 1688980957
transform 1 0 12236 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_133
timestamp 1688980957
transform 1 0 13340 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_139
timestamp 1688980957
transform 1 0 13892 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_141
timestamp 1688980957
transform 1 0 14076 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_153
timestamp 1688980957
transform 1 0 15180 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_165
timestamp 1688980957
transform 1 0 16284 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_177
timestamp 1688980957
transform 1 0 17388 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_189
timestamp 1688980957
transform 1 0 18492 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_195
timestamp 1688980957
transform 1 0 19044 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_197
timestamp 1688980957
transform 1 0 19228 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_202
timestamp 1688980957
transform 1 0 19688 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_214
timestamp 1688980957
transform 1 0 20792 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_235
timestamp 1688980957
transform 1 0 22724 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_239
timestamp 1688980957
transform 1 0 23092 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_251
timestamp 1688980957
transform 1 0 24196 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_253
timestamp 1688980957
transform 1 0 24380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_265
timestamp 1688980957
transform 1 0 25484 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_277
timestamp 1688980957
transform 1 0 26588 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_289
timestamp 1688980957
transform 1 0 27692 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_301
timestamp 1688980957
transform 1 0 28796 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_307
timestamp 1688980957
transform 1 0 29348 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_309
timestamp 1688980957
transform 1 0 29532 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_313
timestamp 1688980957
transform 1 0 29900 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_317
timestamp 1688980957
transform 1 0 30268 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_329
timestamp 1688980957
transform 1 0 31372 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_341
timestamp 1688980957
transform 1 0 32476 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_4_353
timestamp 1688980957
transform 1 0 33580 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_361
timestamp 1688980957
transform 1 0 34316 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_365
timestamp 1688980957
transform 1 0 34684 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_377
timestamp 1688980957
transform 1 0 35788 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_389
timestamp 1688980957
transform 1 0 36892 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_394
timestamp 1688980957
transform 1 0 37352 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_406
timestamp 1688980957
transform 1 0 38456 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_418
timestamp 1688980957
transform 1 0 39560 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_421
timestamp 1688980957
transform 1 0 39836 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_427
timestamp 1688980957
transform 1 0 40388 0 1 3264
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_431
timestamp 1688980957
transform 1 0 40756 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_443
timestamp 1688980957
transform 1 0 41860 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_4_455
timestamp 1688980957
transform 1 0 42964 0 1 3264
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_3
timestamp 1688980957
transform 1 0 1380 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_15
timestamp 1688980957
transform 1 0 2484 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_27
timestamp 1688980957
transform 1 0 3588 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_39
timestamp 1688980957
transform 1 0 4692 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_51
timestamp 1688980957
transform 1 0 5796 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_55
timestamp 1688980957
transform 1 0 6164 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_57
timestamp 1688980957
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_69
timestamp 1688980957
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_81
timestamp 1688980957
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_93
timestamp 1688980957
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_105
timestamp 1688980957
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_111
timestamp 1688980957
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_113
timestamp 1688980957
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_125
timestamp 1688980957
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_137
timestamp 1688980957
transform 1 0 13708 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_149
timestamp 1688980957
transform 1 0 14812 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_161
timestamp 1688980957
transform 1 0 15916 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_167
timestamp 1688980957
transform 1 0 16468 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_169
timestamp 1688980957
transform 1 0 16652 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_181
timestamp 1688980957
transform 1 0 17756 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_193
timestamp 1688980957
transform 1 0 18860 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_205
timestamp 1688980957
transform 1 0 19964 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_216
timestamp 1688980957
transform 1 0 20976 0 -1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_237
timestamp 1688980957
transform 1 0 22908 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_249
timestamp 1688980957
transform 1 0 24012 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_257
timestamp 1688980957
transform 1 0 24748 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_262
timestamp 1688980957
transform 1 0 25208 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_274
timestamp 1688980957
transform 1 0 26312 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_281
timestamp 1688980957
transform 1 0 26956 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_285
timestamp 1688980957
transform 1 0 27324 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_297
timestamp 1688980957
transform 1 0 28428 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_309
timestamp 1688980957
transform 1 0 29532 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_321
timestamp 1688980957
transform 1 0 30636 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_327
timestamp 1688980957
transform 1 0 31188 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_331
timestamp 1688980957
transform 1 0 31556 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_335
timestamp 1688980957
transform 1 0 31924 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_337
timestamp 1688980957
transform 1 0 32108 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_349
timestamp 1688980957
transform 1 0 33212 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_361
timestamp 1688980957
transform 1 0 34316 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_373
timestamp 1688980957
transform 1 0 35420 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_385
timestamp 1688980957
transform 1 0 36524 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_391
timestamp 1688980957
transform 1 0 37076 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_393
timestamp 1688980957
transform 1 0 37260 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_398
timestamp 1688980957
transform 1 0 37720 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_410
timestamp 1688980957
transform 1 0 38824 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_418
timestamp 1688980957
transform 1 0 39560 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_423
timestamp 1688980957
transform 1 0 40020 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_435
timestamp 1688980957
transform 1 0 41124 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_447
timestamp 1688980957
transform 1 0 42228 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_5_449
timestamp 1688980957
transform 1 0 42412 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_457
timestamp 1688980957
transform 1 0 43148 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_3
timestamp 1688980957
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_15
timestamp 1688980957
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_27
timestamp 1688980957
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_29
timestamp 1688980957
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_41
timestamp 1688980957
transform 1 0 4876 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_53
timestamp 1688980957
transform 1 0 5980 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_65
timestamp 1688980957
transform 1 0 7084 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_77
timestamp 1688980957
transform 1 0 8188 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_83
timestamp 1688980957
transform 1 0 8740 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_85
timestamp 1688980957
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_97
timestamp 1688980957
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_109
timestamp 1688980957
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_121
timestamp 1688980957
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_133
timestamp 1688980957
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_139
timestamp 1688980957
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_141
timestamp 1688980957
transform 1 0 14076 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_153
timestamp 1688980957
transform 1 0 15180 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_165
timestamp 1688980957
transform 1 0 16284 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_177
timestamp 1688980957
transform 1 0 17388 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_189
timestamp 1688980957
transform 1 0 18492 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_195
timestamp 1688980957
transform 1 0 19044 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_197
timestamp 1688980957
transform 1 0 19228 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_209
timestamp 1688980957
transform 1 0 20332 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_221
timestamp 1688980957
transform 1 0 21436 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_225
timestamp 1688980957
transform 1 0 21804 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_242
timestamp 1688980957
transform 1 0 23368 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_248
timestamp 1688980957
transform 1 0 23920 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_253
timestamp 1688980957
transform 1 0 24380 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_265
timestamp 1688980957
transform 1 0 25484 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_271
timestamp 1688980957
transform 1 0 26036 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_283
timestamp 1688980957
transform 1 0 27140 0 1 4352
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_294
timestamp 1688980957
transform 1 0 28152 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_306
timestamp 1688980957
transform 1 0 29256 0 1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_309
timestamp 1688980957
transform 1 0 29532 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_321
timestamp 1688980957
transform 1 0 30636 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_333
timestamp 1688980957
transform 1 0 31740 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_340
timestamp 1688980957
transform 1 0 32384 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_352
timestamp 1688980957
transform 1 0 33488 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_365
timestamp 1688980957
transform 1 0 34684 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_377
timestamp 1688980957
transform 1 0 35788 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_385
timestamp 1688980957
transform 1 0 36524 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_390
timestamp 1688980957
transform 1 0 36984 0 1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_6_398
timestamp 1688980957
transform 1 0 37720 0 1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_404
timestamp 1688980957
transform 1 0 38272 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_416
timestamp 1688980957
transform 1 0 39376 0 1 4352
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_421
timestamp 1688980957
transform 1 0 39836 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_433
timestamp 1688980957
transform 1 0 40940 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_445
timestamp 1688980957
transform 1 0 42044 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_457
timestamp 1688980957
transform 1 0 43148 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 1688980957
transform 1 0 1380 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 1688980957
transform 1 0 2484 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_27
timestamp 1688980957
transform 1 0 3588 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_39
timestamp 1688980957
transform 1 0 4692 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_51
timestamp 1688980957
transform 1 0 5796 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_55
timestamp 1688980957
transform 1 0 6164 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_57
timestamp 1688980957
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_69
timestamp 1688980957
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_81
timestamp 1688980957
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_93
timestamp 1688980957
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_105
timestamp 1688980957
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_111
timestamp 1688980957
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_113
timestamp 1688980957
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_125
timestamp 1688980957
transform 1 0 12604 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_137
timestamp 1688980957
transform 1 0 13708 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_149
timestamp 1688980957
transform 1 0 14812 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_161
timestamp 1688980957
transform 1 0 15916 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_167
timestamp 1688980957
transform 1 0 16468 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_169
timestamp 1688980957
transform 1 0 16652 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_181
timestamp 1688980957
transform 1 0 17756 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_193
timestamp 1688980957
transform 1 0 18860 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_205
timestamp 1688980957
transform 1 0 19964 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_217
timestamp 1688980957
transform 1 0 21068 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_223
timestamp 1688980957
transform 1 0 21620 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_225
timestamp 1688980957
transform 1 0 21804 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_237
timestamp 1688980957
transform 1 0 22908 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_249
timestamp 1688980957
transform 1 0 24012 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_261
timestamp 1688980957
transform 1 0 25116 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_273
timestamp 1688980957
transform 1 0 26220 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_279
timestamp 1688980957
transform 1 0 26772 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_281
timestamp 1688980957
transform 1 0 26956 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_293
timestamp 1688980957
transform 1 0 28060 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_305
timestamp 1688980957
transform 1 0 29164 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_317
timestamp 1688980957
transform 1 0 30268 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_329
timestamp 1688980957
transform 1 0 31372 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_335
timestamp 1688980957
transform 1 0 31924 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_337
timestamp 1688980957
transform 1 0 32108 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_349
timestamp 1688980957
transform 1 0 33212 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_361
timestamp 1688980957
transform 1 0 34316 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_373
timestamp 1688980957
transform 1 0 35420 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_385
timestamp 1688980957
transform 1 0 36524 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_391
timestamp 1688980957
transform 1 0 37076 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_393
timestamp 1688980957
transform 1 0 37260 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_397
timestamp 1688980957
transform 1 0 37628 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_409
timestamp 1688980957
transform 1 0 38732 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_421
timestamp 1688980957
transform 1 0 39836 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_433
timestamp 1688980957
transform 1 0 40940 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_445
timestamp 1688980957
transform 1 0 42044 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_7_449
timestamp 1688980957
transform 1 0 42412 0 -1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_457
timestamp 1688980957
transform 1 0 43148 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_3
timestamp 1688980957
transform 1 0 1380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_15
timestamp 1688980957
transform 1 0 2484 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_27
timestamp 1688980957
transform 1 0 3588 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_29
timestamp 1688980957
transform 1 0 3772 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_41
timestamp 1688980957
transform 1 0 4876 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_53
timestamp 1688980957
transform 1 0 5980 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_65
timestamp 1688980957
transform 1 0 7084 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_77
timestamp 1688980957
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_83
timestamp 1688980957
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_85
timestamp 1688980957
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_97
timestamp 1688980957
transform 1 0 10028 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_109
timestamp 1688980957
transform 1 0 11132 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_121
timestamp 1688980957
transform 1 0 12236 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_133
timestamp 1688980957
transform 1 0 13340 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_139
timestamp 1688980957
transform 1 0 13892 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_141
timestamp 1688980957
transform 1 0 14076 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_153
timestamp 1688980957
transform 1 0 15180 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_165
timestamp 1688980957
transform 1 0 16284 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_177
timestamp 1688980957
transform 1 0 17388 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_189
timestamp 1688980957
transform 1 0 18492 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_195
timestamp 1688980957
transform 1 0 19044 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_197
timestamp 1688980957
transform 1 0 19228 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_209
timestamp 1688980957
transform 1 0 20332 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_221
timestamp 1688980957
transform 1 0 21436 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_233
timestamp 1688980957
transform 1 0 22540 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_245
timestamp 1688980957
transform 1 0 23644 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_251
timestamp 1688980957
transform 1 0 24196 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_253
timestamp 1688980957
transform 1 0 24380 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_265
timestamp 1688980957
transform 1 0 25484 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_277
timestamp 1688980957
transform 1 0 26588 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_289
timestamp 1688980957
transform 1 0 27692 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_301
timestamp 1688980957
transform 1 0 28796 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_307
timestamp 1688980957
transform 1 0 29348 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_309
timestamp 1688980957
transform 1 0 29532 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_321
timestamp 1688980957
transform 1 0 30636 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_333
timestamp 1688980957
transform 1 0 31740 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_345
timestamp 1688980957
transform 1 0 32844 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_357
timestamp 1688980957
transform 1 0 33948 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_363
timestamp 1688980957
transform 1 0 34500 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_365
timestamp 1688980957
transform 1 0 34684 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_377
timestamp 1688980957
transform 1 0 35788 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_389
timestamp 1688980957
transform 1 0 36892 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_401
timestamp 1688980957
transform 1 0 37996 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_413
timestamp 1688980957
transform 1 0 39100 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_419
timestamp 1688980957
transform 1 0 39652 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_421
timestamp 1688980957
transform 1 0 39836 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_433
timestamp 1688980957
transform 1 0 40940 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_445
timestamp 1688980957
transform 1 0 42044 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_457
timestamp 1688980957
transform 1 0 43148 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 1688980957
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_15
timestamp 1688980957
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_27
timestamp 1688980957
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_39
timestamp 1688980957
transform 1 0 4692 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_9_51
timestamp 1688980957
transform 1 0 5796 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_55
timestamp 1688980957
transform 1 0 6164 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_57
timestamp 1688980957
transform 1 0 6348 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_69
timestamp 1688980957
transform 1 0 7452 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_81
timestamp 1688980957
transform 1 0 8556 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_93
timestamp 1688980957
transform 1 0 9660 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_105
timestamp 1688980957
transform 1 0 10764 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_111
timestamp 1688980957
transform 1 0 11316 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_113
timestamp 1688980957
transform 1 0 11500 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_125
timestamp 1688980957
transform 1 0 12604 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_137
timestamp 1688980957
transform 1 0 13708 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_149
timestamp 1688980957
transform 1 0 14812 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_161
timestamp 1688980957
transform 1 0 15916 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_167
timestamp 1688980957
transform 1 0 16468 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_169
timestamp 1688980957
transform 1 0 16652 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_181
timestamp 1688980957
transform 1 0 17756 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_193
timestamp 1688980957
transform 1 0 18860 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_205
timestamp 1688980957
transform 1 0 19964 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_217
timestamp 1688980957
transform 1 0 21068 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_223
timestamp 1688980957
transform 1 0 21620 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_225
timestamp 1688980957
transform 1 0 21804 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_237
timestamp 1688980957
transform 1 0 22908 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_249
timestamp 1688980957
transform 1 0 24012 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_261
timestamp 1688980957
transform 1 0 25116 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_273
timestamp 1688980957
transform 1 0 26220 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_279
timestamp 1688980957
transform 1 0 26772 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_281
timestamp 1688980957
transform 1 0 26956 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_293
timestamp 1688980957
transform 1 0 28060 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_305
timestamp 1688980957
transform 1 0 29164 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_317
timestamp 1688980957
transform 1 0 30268 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_329
timestamp 1688980957
transform 1 0 31372 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_335
timestamp 1688980957
transform 1 0 31924 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_337
timestamp 1688980957
transform 1 0 32108 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_349
timestamp 1688980957
transform 1 0 33212 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_361
timestamp 1688980957
transform 1 0 34316 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_373
timestamp 1688980957
transform 1 0 35420 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_385
timestamp 1688980957
transform 1 0 36524 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_391
timestamp 1688980957
transform 1 0 37076 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_393
timestamp 1688980957
transform 1 0 37260 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_405
timestamp 1688980957
transform 1 0 38364 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_417
timestamp 1688980957
transform 1 0 39468 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_429
timestamp 1688980957
transform 1 0 40572 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_441
timestamp 1688980957
transform 1 0 41676 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_447
timestamp 1688980957
transform 1 0 42228 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_449
timestamp 1688980957
transform 1 0 42412 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_457
timestamp 1688980957
transform 1 0 43148 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_3
timestamp 1688980957
transform 1 0 1380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_15
timestamp 1688980957
transform 1 0 2484 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 1688980957
transform 1 0 3588 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_29
timestamp 1688980957
transform 1 0 3772 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_41
timestamp 1688980957
transform 1 0 4876 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_53
timestamp 1688980957
transform 1 0 5980 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_65
timestamp 1688980957
transform 1 0 7084 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_77
timestamp 1688980957
transform 1 0 8188 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_83
timestamp 1688980957
transform 1 0 8740 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_85
timestamp 1688980957
transform 1 0 8924 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_97
timestamp 1688980957
transform 1 0 10028 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_109
timestamp 1688980957
transform 1 0 11132 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_121
timestamp 1688980957
transform 1 0 12236 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_133
timestamp 1688980957
transform 1 0 13340 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_139
timestamp 1688980957
transform 1 0 13892 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_141
timestamp 1688980957
transform 1 0 14076 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_153
timestamp 1688980957
transform 1 0 15180 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_165
timestamp 1688980957
transform 1 0 16284 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_177
timestamp 1688980957
transform 1 0 17388 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_189
timestamp 1688980957
transform 1 0 18492 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_195
timestamp 1688980957
transform 1 0 19044 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_197
timestamp 1688980957
transform 1 0 19228 0 1 6528
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_207
timestamp 1688980957
transform 1 0 20148 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_219
timestamp 1688980957
transform 1 0 21252 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_231
timestamp 1688980957
transform 1 0 22356 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_243
timestamp 1688980957
transform 1 0 23460 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_251
timestamp 1688980957
transform 1 0 24196 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_253
timestamp 1688980957
transform 1 0 24380 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_265
timestamp 1688980957
transform 1 0 25484 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_277
timestamp 1688980957
transform 1 0 26588 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_289
timestamp 1688980957
transform 1 0 27692 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_301
timestamp 1688980957
transform 1 0 28796 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_307
timestamp 1688980957
transform 1 0 29348 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_309
timestamp 1688980957
transform 1 0 29532 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_321
timestamp 1688980957
transform 1 0 30636 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_333
timestamp 1688980957
transform 1 0 31740 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_345
timestamp 1688980957
transform 1 0 32844 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_357
timestamp 1688980957
transform 1 0 33948 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_363
timestamp 1688980957
transform 1 0 34500 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_365
timestamp 1688980957
transform 1 0 34684 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_377
timestamp 1688980957
transform 1 0 35788 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_389
timestamp 1688980957
transform 1 0 36892 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_401
timestamp 1688980957
transform 1 0 37996 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_413
timestamp 1688980957
transform 1 0 39100 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_419
timestamp 1688980957
transform 1 0 39652 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_421
timestamp 1688980957
transform 1 0 39836 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_433
timestamp 1688980957
transform 1 0 40940 0 1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_445
timestamp 1688980957
transform 1 0 42044 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_457
timestamp 1688980957
transform 1 0 43148 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_3
timestamp 1688980957
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_15
timestamp 1688980957
transform 1 0 2484 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_27
timestamp 1688980957
transform 1 0 3588 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_39
timestamp 1688980957
transform 1 0 4692 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_51
timestamp 1688980957
transform 1 0 5796 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_55
timestamp 1688980957
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_57
timestamp 1688980957
transform 1 0 6348 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_63
timestamp 1688980957
transform 1 0 6900 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_68
timestamp 1688980957
transform 1 0 7360 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_84
timestamp 1688980957
transform 1 0 8832 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_96
timestamp 1688980957
transform 1 0 9936 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_108
timestamp 1688980957
transform 1 0 11040 0 -1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_113
timestamp 1688980957
transform 1 0 11500 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_125
timestamp 1688980957
transform 1 0 12604 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_137
timestamp 1688980957
transform 1 0 13708 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_143
timestamp 1688980957
transform 1 0 14260 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_148
timestamp 1688980957
transform 1 0 14720 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_160
timestamp 1688980957
transform 1 0 15824 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_169
timestamp 1688980957
transform 1 0 16652 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_11_189
timestamp 1688980957
transform 1 0 18492 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_204
timestamp 1688980957
transform 1 0 19872 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_211
timestamp 1688980957
transform 1 0 20516 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_228
timestamp 1688980957
transform 1 0 22080 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_232
timestamp 1688980957
transform 1 0 22448 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_236
timestamp 1688980957
transform 1 0 22816 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_248
timestamp 1688980957
transform 1 0 23920 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_256
timestamp 1688980957
transform 1 0 24656 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_260
timestamp 1688980957
transform 1 0 25024 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_275
timestamp 1688980957
transform 1 0 26404 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_279
timestamp 1688980957
transform 1 0 26772 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_281
timestamp 1688980957
transform 1 0 26956 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_293
timestamp 1688980957
transform 1 0 28060 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_305
timestamp 1688980957
transform 1 0 29164 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_317
timestamp 1688980957
transform 1 0 30268 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_329
timestamp 1688980957
transform 1 0 31372 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_335
timestamp 1688980957
transform 1 0 31924 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_337
timestamp 1688980957
transform 1 0 32108 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_349
timestamp 1688980957
transform 1 0 33212 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_361
timestamp 1688980957
transform 1 0 34316 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_373
timestamp 1688980957
transform 1 0 35420 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_385
timestamp 1688980957
transform 1 0 36524 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_391
timestamp 1688980957
transform 1 0 37076 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_393
timestamp 1688980957
transform 1 0 37260 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_405
timestamp 1688980957
transform 1 0 38364 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_417
timestamp 1688980957
transform 1 0 39468 0 -1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_429
timestamp 1688980957
transform 1 0 40572 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_11_441
timestamp 1688980957
transform 1 0 41676 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_447
timestamp 1688980957
transform 1 0 42228 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_449
timestamp 1688980957
transform 1 0 42412 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_457
timestamp 1688980957
transform 1 0 43148 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_3
timestamp 1688980957
transform 1 0 1380 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_15
timestamp 1688980957
transform 1 0 2484 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_27
timestamp 1688980957
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_29
timestamp 1688980957
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_41
timestamp 1688980957
transform 1 0 4876 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_49
timestamp 1688980957
transform 1 0 5612 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_70
timestamp 1688980957
transform 1 0 7544 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_85
timestamp 1688980957
transform 1 0 8924 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_94
timestamp 1688980957
transform 1 0 9752 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_106
timestamp 1688980957
transform 1 0 10856 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_121
timestamp 1688980957
transform 1 0 12236 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_130
timestamp 1688980957
transform 1 0 13064 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_139
timestamp 1688980957
transform 1 0 13892 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_141
timestamp 1688980957
transform 1 0 14076 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_154
timestamp 1688980957
transform 1 0 15272 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_178
timestamp 1688980957
transform 1 0 17480 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_192
timestamp 1688980957
transform 1 0 18768 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_251
timestamp 1688980957
transform 1 0 24196 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_292
timestamp 1688980957
transform 1 0 27968 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_304
timestamp 1688980957
transform 1 0 29072 0 1 7616
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_309
timestamp 1688980957
transform 1 0 29532 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_321
timestamp 1688980957
transform 1 0 30636 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_333
timestamp 1688980957
transform 1 0 31740 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_345
timestamp 1688980957
transform 1 0 32844 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_354
timestamp 1688980957
transform 1 0 33672 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_362
timestamp 1688980957
transform 1 0 34408 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_365
timestamp 1688980957
transform 1 0 34684 0 1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_373
timestamp 1688980957
transform 1 0 35420 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_417
timestamp 1688980957
transform 1 0 39468 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_433
timestamp 1688980957
transform 1 0 40940 0 1 7616
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_12_445
timestamp 1688980957
transform 1 0 42044 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_457
timestamp 1688980957
transform 1 0 43148 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_3
timestamp 1688980957
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_13_15
timestamp 1688980957
transform 1 0 2484 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_27
timestamp 1688980957
transform 1 0 3588 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_13_29
timestamp 1688980957
transform 1 0 3772 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_35
timestamp 1688980957
transform 1 0 4324 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_57
timestamp 1688980957
transform 1 0 6348 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_85
timestamp 1688980957
transform 1 0 8924 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_96
timestamp 1688980957
transform 1 0 9936 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_113
timestamp 1688980957
transform 1 0 11500 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_124
timestamp 1688980957
transform 1 0 12512 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_141
timestamp 1688980957
transform 1 0 14076 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_156
timestamp 1688980957
transform 1 0 15456 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_169
timestamp 1688980957
transform 1 0 16652 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_201
timestamp 1688980957
transform 1 0 19596 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_223
timestamp 1688980957
transform 1 0 21620 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_355
timestamp 1688980957
transform 1 0 33764 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_389
timestamp 1688980957
transform 1 0 36892 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_13_417
timestamp 1688980957
transform 1 0 39468 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_439
timestamp 1688980957
transform 1 0 41492 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_447
timestamp 1688980957
transform 1 0 42228 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_449
timestamp 1688980957
transform 1 0 42412 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_457
timestamp 1688980957
transform 1 0 43148 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  input1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3312 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input2 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 24748 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input3
timestamp 1688980957
transform -1 0 26864 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input4
timestamp 1688980957
transform -1 0 28980 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input5
timestamp 1688980957
transform -1 0 31096 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input6
timestamp 1688980957
transform -1 0 33212 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input7
timestamp 1688980957
transform -1 0 35328 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1688980957
transform -1 0 37536 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input9
timestamp 1688980957
transform 1 0 39284 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input10
timestamp 1688980957
transform 1 0 41400 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input11
timestamp 1688980957
transform 1 0 42964 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input12
timestamp 1688980957
transform 1 0 5428 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input13
timestamp 1688980957
transform 1 0 7544 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input14
timestamp 1688980957
transform 1 0 9660 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input15
timestamp 1688980957
transform 1 0 11776 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input16
timestamp 1688980957
transform -1 0 14352 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input17
timestamp 1688980957
transform -1 0 16284 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input18
timestamp 1688980957
transform -1 0 18400 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input19
timestamp 1688980957
transform -1 0 20516 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input20
timestamp 1688980957
transform -1 0 22632 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input21
timestamp 1688980957
transform 1 0 19596 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input22
timestamp 1688980957
transform 1 0 19872 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input23
timestamp 1688980957
transform 1 0 20240 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input24
timestamp 1688980957
transform 1 0 19504 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input25
timestamp 1688980957
transform 1 0 20240 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input26
timestamp 1688980957
transform 1 0 20516 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input27
timestamp 1688980957
transform 1 0 20792 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input28
timestamp 1688980957
transform 1 0 21068 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input29
timestamp 1688980957
transform 1 0 21804 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input30
timestamp 1688980957
transform 1 0 22080 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input31
timestamp 1688980957
transform 1 0 22356 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input32
timestamp 1688980957
transform 1 0 22632 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input33
timestamp 1688980957
transform 1 0 22908 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input34
timestamp 1688980957
transform 1 0 23184 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input35
timestamp 1688980957
transform 1 0 23460 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input36
timestamp 1688980957
transform 1 0 23736 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input37
timestamp 1688980957
transform 1 0 24012 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input38
timestamp 1688980957
transform -1 0 24656 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input39
timestamp 1688980957
transform -1 0 24932 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input40
timestamp 1688980957
transform -1 0 25208 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input41
timestamp 1688980957
transform -1 0 25484 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input42
timestamp 1688980957
transform 1 0 28060 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input43
timestamp 1688980957
transform 1 0 28336 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input44
timestamp 1688980957
transform 1 0 28612 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input45
timestamp 1688980957
transform 1 0 28888 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input46
timestamp 1688980957
transform 1 0 29164 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input47
timestamp 1688980957
transform 1 0 29532 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input48
timestamp 1688980957
transform 1 0 25484 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input49
timestamp 1688980957
transform -1 0 26036 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input50
timestamp 1688980957
transform -1 0 26312 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input51
timestamp 1688980957
transform -1 0 26588 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input52
timestamp 1688980957
transform -1 0 26864 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input53
timestamp 1688980957
transform 1 0 26956 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input54
timestamp 1688980957
transform -1 0 27508 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input55
timestamp 1688980957
transform -1 0 27784 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input56
timestamp 1688980957
transform -1 0 28060 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input57
timestamp 1688980957
transform -1 0 30084 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input58
timestamp 1688980957
transform -1 0 32936 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input59
timestamp 1688980957
transform -1 0 33212 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input60
timestamp 1688980957
transform -1 0 33488 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input61
timestamp 1688980957
transform -1 0 33764 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input62
timestamp 1688980957
transform -1 0 33672 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input63
timestamp 1688980957
transform -1 0 34592 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input64
timestamp 1688980957
transform -1 0 30360 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input65
timestamp 1688980957
transform -1 0 30636 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input66
timestamp 1688980957
transform -1 0 30912 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input67
timestamp 1688980957
transform -1 0 31188 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input68
timestamp 1688980957
transform -1 0 31464 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input69
timestamp 1688980957
transform -1 0 31740 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input70
timestamp 1688980957
transform -1 0 32016 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input71
timestamp 1688980957
transform -1 0 32384 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input72
timestamp 1688980957
transform -1 0 32660 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input73
timestamp 1688980957
transform 1 0 1380 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  inst_clk_buf
timestamp 1688980957
transform 1 0 21344 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_DSP_switch_matrix__00_
timestamp 1688980957
transform -1 0 25208 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_DSP_switch_matrix__01_
timestamp 1688980957
transform -1 0 24932 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_DSP_switch_matrix__02_
timestamp 1688980957
transform -1 0 24656 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_DSP_switch_matrix__03_
timestamp 1688980957
transform -1 0 23644 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_DSP_switch_matrix__04_
timestamp 1688980957
transform -1 0 23092 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_DSP_switch_matrix__05_
timestamp 1688980957
transform -1 0 22816 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_DSP_switch_matrix__06_
timestamp 1688980957
transform -1 0 22816 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_DSP_switch_matrix__07_
timestamp 1688980957
transform -1 0 22264 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_DSP_switch_matrix__08_
timestamp 1688980957
transform -1 0 21988 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_DSP_switch_matrix__09_
timestamp 1688980957
transform -1 0 21712 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_DSP_switch_matrix__10_
timestamp 1688980957
transform -1 0 21712 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_DSP_switch_matrix__11_
timestamp 1688980957
transform -1 0 21436 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_DSP_switch_matrix__12_
timestamp 1688980957
transform -1 0 20608 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_DSP_switch_matrix__13_
timestamp 1688980957
transform -1 0 20884 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_DSP_switch_matrix__14_
timestamp 1688980957
transform -1 0 20332 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_DSP_switch_matrix__15_
timestamp 1688980957
transform 1 0 19780 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_DSP_switch_matrix__16_
timestamp 1688980957
transform -1 0 22540 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_DSP_switch_matrix__17_
timestamp 1688980957
transform -1 0 23368 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_DSP_switch_matrix__18_
timestamp 1688980957
transform -1 0 26864 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_DSP_switch_matrix__19_
timestamp 1688980957
transform -1 0 26588 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_DSP_switch_matrix__20_
timestamp 1688980957
transform -1 0 26312 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_DSP_switch_matrix__21_
timestamp 1688980957
transform -1 0 26036 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_DSP_switch_matrix__22_
timestamp 1688980957
transform -1 0 25024 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_DSP_switch_matrix__23_
timestamp 1688980957
transform -1 0 25484 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_DSP_switch_matrix__24_
timestamp 1688980957
transform -1 0 24196 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_DSP_switch_matrix__25_
timestamp 1688980957
transform -1 0 23920 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_DSP_switch_matrix__26_
timestamp 1688980957
transform -1 0 25760 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_DSP_switch_matrix__27_
timestamp 1688980957
transform -1 0 27140 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_DSP_switch_matrix__28_
timestamp 1688980957
transform -1 0 27968 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_DSP_switch_matrix__29_
timestamp 1688980957
transform -1 0 27692 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_DSP_switch_matrix__30_
timestamp 1688980957
transform -1 0 27416 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_DSP_switch_matrix__31_
timestamp 1688980957
transform -1 0 26404 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_DSP_switch_matrix__32_
timestamp 1688980957
transform -1 0 21436 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_DSP_switch_matrix__33_
timestamp 1688980957
transform 1 0 20884 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_DSP_switch_matrix__34_
timestamp 1688980957
transform 1 0 18216 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_DSP_switch_matrix__35_
timestamp 1688980957
transform -1 0 17848 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_DSP_switch_matrix__36_
timestamp 1688980957
transform 1 0 18768 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_DSP_switch_matrix__37_
timestamp 1688980957
transform -1 0 19320 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_DSP_switch_matrix__38_
timestamp 1688980957
transform -1 0 19596 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_DSP_switch_matrix__39_
timestamp 1688980957
transform 1 0 19596 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_DSP_switch_matrix__40_
timestamp 1688980957
transform 1 0 21804 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_DSP_switch_matrix__41_
timestamp 1688980957
transform 1 0 21344 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_DSP_switch_matrix__42_
timestamp 1688980957
transform 1 0 20884 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_DSP_switch_matrix__43_
timestamp 1688980957
transform 1 0 20608 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_DSP_switch_matrix__44_
timestamp 1688980957
transform 1 0 19964 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_DSP_switch_matrix__45_
timestamp 1688980957
transform 1 0 17940 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_DSP_switch_matrix__46_
timestamp 1688980957
transform 1 0 17664 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_S_term_DSP_switch_matrix__47_
timestamp 1688980957
transform 1 0 17388 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_DSP_switch_matrix__48_
timestamp 1688980957
transform -1 0 19504 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_DSP_switch_matrix__49_
timestamp 1688980957
transform -1 0 19136 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_DSP_switch_matrix__50_
timestamp 1688980957
transform -1 0 18400 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  Inst_S_term_DSP_switch_matrix__51_
timestamp 1688980957
transform -1 0 18124 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  output74 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 34684 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output75
timestamp 1688980957
transform 1 0 38364 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output76
timestamp 1688980957
transform 1 0 38364 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output77
timestamp 1688980957
transform 1 0 38916 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output78
timestamp 1688980957
transform 1 0 37812 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output79
timestamp 1688980957
transform 1 0 39836 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output80
timestamp 1688980957
transform 1 0 40388 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output81
timestamp 1688980957
transform 1 0 38916 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output82
timestamp 1688980957
transform 1 0 39836 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output83
timestamp 1688980957
transform 1 0 40388 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output84
timestamp 1688980957
transform 1 0 40940 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output85
timestamp 1688980957
transform 1 0 35236 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output86
timestamp 1688980957
transform 1 0 35788 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output87
timestamp 1688980957
transform 1 0 36340 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output88
timestamp 1688980957
transform 1 0 36708 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output89
timestamp 1688980957
transform 1 0 35604 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output90
timestamp 1688980957
transform 1 0 37260 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output91
timestamp 1688980957
transform 1 0 36156 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output92
timestamp 1688980957
transform 1 0 37812 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output93
timestamp 1688980957
transform 1 0 37260 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output94 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform -1 0 4784 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output95
timestamp 1688980957
transform -1 0 5336 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output96
timestamp 1688980957
transform -1 0 5888 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output97
timestamp 1688980957
transform -1 0 6440 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output98
timestamp 1688980957
transform -1 0 6256 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output99
timestamp 1688980957
transform -1 0 6992 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output100
timestamp 1688980957
transform -1 0 6992 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output101
timestamp 1688980957
transform -1 0 7544 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output102
timestamp 1688980957
transform -1 0 7360 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output103
timestamp 1688980957
transform -1 0 7360 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output104
timestamp 1688980957
transform -1 0 7728 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output105
timestamp 1688980957
transform -1 0 8280 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output106
timestamp 1688980957
transform -1 0 8280 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output107
timestamp 1688980957
transform -1 0 8832 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output108
timestamp 1688980957
transform -1 0 8832 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output109
timestamp 1688980957
transform -1 0 9752 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output110
timestamp 1688980957
transform -1 0 8832 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output111
timestamp 1688980957
transform -1 0 9936 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output112
timestamp 1688980957
transform -1 0 9384 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output113
timestamp 1688980957
transform -1 0 10856 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output114
timestamp 1688980957
transform -1 0 10304 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output115
timestamp 1688980957
transform -1 0 13892 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output116
timestamp 1688980957
transform -1 0 13432 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output117
timestamp 1688980957
transform -1 0 13984 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output118
timestamp 1688980957
transform -1 0 14720 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output119
timestamp 1688980957
transform -1 0 14720 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output120
timestamp 1688980957
transform -1 0 15272 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output121
timestamp 1688980957
transform -1 0 11040 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output122
timestamp 1688980957
transform -1 0 11684 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output123
timestamp 1688980957
transform -1 0 10488 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output124
timestamp 1688980957
transform -1 0 12236 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output125
timestamp 1688980957
transform -1 0 11408 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output126
timestamp 1688980957
transform -1 0 12512 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output127
timestamp 1688980957
transform -1 0 13064 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output128
timestamp 1688980957
transform -1 0 11960 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output129
timestamp 1688980957
transform -1 0 13064 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output130
timestamp 1688980957
transform -1 0 14904 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output131
timestamp 1688980957
transform -1 0 18032 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output132
timestamp 1688980957
transform 1 0 18032 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output133
timestamp 1688980957
transform -1 0 18768 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output134
timestamp 1688980957
transform 1 0 19228 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output135
timestamp 1688980957
transform 1 0 19688 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output136
timestamp 1688980957
transform -1 0 19136 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output137
timestamp 1688980957
transform -1 0 15456 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output138
timestamp 1688980957
transform -1 0 15824 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output139
timestamp 1688980957
transform -1 0 16376 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output140
timestamp 1688980957
transform -1 0 16008 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output141
timestamp 1688980957
transform -1 0 16928 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output142
timestamp 1688980957
transform -1 0 16560 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output143
timestamp 1688980957
transform -1 0 17480 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output144
timestamp 1688980957
transform -1 0 17112 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output145
timestamp 1688980957
transform -1 0 17480 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output146
timestamp 1688980957
transform 1 0 33948 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1688980957
transform 1 0 1104 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1688980957
transform -1 0 43516 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1688980957
transform 1 0 1104 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1688980957
transform -1 0 43516 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1688980957
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1688980957
transform -1 0 43516 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1688980957
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1688980957
transform -1 0 43516 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1688980957
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1688980957
transform -1 0 43516 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1688980957
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1688980957
transform -1 0 43516 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1688980957
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1688980957
transform -1 0 43516 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1688980957
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1688980957
transform -1 0 43516 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1688980957
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1688980957
transform -1 0 43516 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1688980957
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1688980957
transform -1 0 43516 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1688980957
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1688980957
transform -1 0 43516 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1688980957
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1688980957
transform -1 0 43516 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1688980957
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1688980957
transform -1 0 43516 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1688980957
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1688980957
transform -1 0 43516 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_0__0_
timestamp 1688980957
transform -1 0 22172 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_1__0_
timestamp 1688980957
transform -1 0 22356 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_2__0_
timestamp 1688980957
transform -1 0 22080 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_3__0_
timestamp 1688980957
transform -1 0 22172 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_4__0_
timestamp 1688980957
transform -1 0 22632 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_5__0_
timestamp 1688980957
transform -1 0 21620 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_6__0_
timestamp 1688980957
transform -1 0 21344 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_7__0_
timestamp 1688980957
transform -1 0 18860 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_8__0_
timestamp 1688980957
transform -1 0 20976 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_9__0_
timestamp 1688980957
transform -1 0 23092 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_10__0_
timestamp 1688980957
transform -1 0 25208 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_11__0_
timestamp 1688980957
transform -1 0 27324 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_12__0_
timestamp 1688980957
transform -1 0 29440 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_13__0_
timestamp 1688980957
transform -1 0 31556 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_14__0_
timestamp 1688980957
transform -1 0 36984 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_15__0_
timestamp 1688980957
transform -1 0 36248 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_16__0_
timestamp 1688980957
transform -1 0 37720 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_17__0_
timestamp 1688980957
transform -1 0 39100 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_18__0_
timestamp 1688980957
transform 1 0 40480 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_19__0_
timestamp 1688980957
transform 1 0 40204 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  strobe_outbuf_0__0_
timestamp 1688980957
transform 1 0 22632 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  strobe_outbuf_1__0_
timestamp 1688980957
transform 1 0 22816 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  strobe_outbuf_2__0_
timestamp 1688980957
transform 1 0 22540 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  strobe_outbuf_3__0_
timestamp 1688980957
transform 1 0 22632 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  strobe_outbuf_4__0_
timestamp 1688980957
transform 1 0 23092 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  strobe_outbuf_5__0_
timestamp 1688980957
transform 1 0 22172 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  strobe_outbuf_6__0_
timestamp 1688980957
transform 1 0 22448 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  strobe_outbuf_7__0_
timestamp 1688980957
transform 1 0 19412 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  strobe_outbuf_8__0_
timestamp 1688980957
transform 1 0 21528 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  strobe_outbuf_9__0_
timestamp 1688980957
transform 1 0 23644 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  strobe_outbuf_10__0_
timestamp 1688980957
transform 1 0 25760 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  strobe_outbuf_11__0_
timestamp 1688980957
transform 1 0 27876 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  strobe_outbuf_12__0_
timestamp 1688980957
transform 1 0 29992 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_13__0_
timestamp 1688980957
transform -1 0 32384 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_14__0_
timestamp 1688980957
transform -1 0 37628 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_15__0_
timestamp 1688980957
transform -1 0 37352 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_16__0_
timestamp 1688980957
transform -1 0 38272 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_17__0_
timestamp 1688980957
transform -1 0 39284 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_18__0_
timestamp 1688980957
transform -1 0 40020 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_19__0_
timestamp 1688980957
transform -1 0 40020 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_28 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3680 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_29
timestamp 1688980957
transform 1 0 6256 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_30
timestamp 1688980957
transform 1 0 8832 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_31
timestamp 1688980957
transform 1 0 11408 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_32
timestamp 1688980957
transform 1 0 13984 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_33
timestamp 1688980957
transform 1 0 16560 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_34
timestamp 1688980957
transform 1 0 19136 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_35
timestamp 1688980957
transform 1 0 21712 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_36
timestamp 1688980957
transform 1 0 24288 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_37
timestamp 1688980957
transform 1 0 26864 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_38
timestamp 1688980957
transform 1 0 29440 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_39
timestamp 1688980957
transform 1 0 32016 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_40
timestamp 1688980957
transform 1 0 34592 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_41
timestamp 1688980957
transform 1 0 37168 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_42
timestamp 1688980957
transform 1 0 39744 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_43
timestamp 1688980957
transform 1 0 42320 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_44
timestamp 1688980957
transform 1 0 6256 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_45
timestamp 1688980957
transform 1 0 11408 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_46
timestamp 1688980957
transform 1 0 16560 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_47
timestamp 1688980957
transform 1 0 21712 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_48
timestamp 1688980957
transform 1 0 26864 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_49
timestamp 1688980957
transform 1 0 32016 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_50
timestamp 1688980957
transform 1 0 37168 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_51
timestamp 1688980957
transform 1 0 42320 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_52
timestamp 1688980957
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_53
timestamp 1688980957
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_54
timestamp 1688980957
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_55
timestamp 1688980957
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_56
timestamp 1688980957
transform 1 0 24288 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_57
timestamp 1688980957
transform 1 0 29440 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_58
timestamp 1688980957
transform 1 0 34592 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_59
timestamp 1688980957
transform 1 0 39744 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_60
timestamp 1688980957
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_61
timestamp 1688980957
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_62
timestamp 1688980957
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_63
timestamp 1688980957
transform 1 0 21712 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_64
timestamp 1688980957
transform 1 0 26864 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_65
timestamp 1688980957
transform 1 0 32016 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_66
timestamp 1688980957
transform 1 0 37168 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_67
timestamp 1688980957
transform 1 0 42320 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_68
timestamp 1688980957
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_69
timestamp 1688980957
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_70
timestamp 1688980957
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_71
timestamp 1688980957
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_72
timestamp 1688980957
transform 1 0 24288 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_73
timestamp 1688980957
transform 1 0 29440 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_74
timestamp 1688980957
transform 1 0 34592 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_75
timestamp 1688980957
transform 1 0 39744 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_76
timestamp 1688980957
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_77
timestamp 1688980957
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_78
timestamp 1688980957
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_79
timestamp 1688980957
transform 1 0 21712 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_80
timestamp 1688980957
transform 1 0 26864 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_81
timestamp 1688980957
transform 1 0 32016 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_82
timestamp 1688980957
transform 1 0 37168 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_83
timestamp 1688980957
transform 1 0 42320 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_84
timestamp 1688980957
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_85
timestamp 1688980957
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_86
timestamp 1688980957
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_87
timestamp 1688980957
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_88
timestamp 1688980957
transform 1 0 24288 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_89
timestamp 1688980957
transform 1 0 29440 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_90
timestamp 1688980957
transform 1 0 34592 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_91
timestamp 1688980957
transform 1 0 39744 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_92
timestamp 1688980957
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_93
timestamp 1688980957
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_94
timestamp 1688980957
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_95
timestamp 1688980957
transform 1 0 21712 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_96
timestamp 1688980957
transform 1 0 26864 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_97
timestamp 1688980957
transform 1 0 32016 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_98
timestamp 1688980957
transform 1 0 37168 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_99
timestamp 1688980957
transform 1 0 42320 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_100
timestamp 1688980957
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_101
timestamp 1688980957
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_102
timestamp 1688980957
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_103
timestamp 1688980957
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_104
timestamp 1688980957
transform 1 0 24288 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_105
timestamp 1688980957
transform 1 0 29440 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_106
timestamp 1688980957
transform 1 0 34592 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_107
timestamp 1688980957
transform 1 0 39744 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_108
timestamp 1688980957
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_109
timestamp 1688980957
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_110
timestamp 1688980957
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_111
timestamp 1688980957
transform 1 0 21712 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_112
timestamp 1688980957
transform 1 0 26864 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_113
timestamp 1688980957
transform 1 0 32016 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_114
timestamp 1688980957
transform 1 0 37168 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_115
timestamp 1688980957
transform 1 0 42320 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_116
timestamp 1688980957
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_117
timestamp 1688980957
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_118
timestamp 1688980957
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_119
timestamp 1688980957
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_120
timestamp 1688980957
transform 1 0 24288 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_121
timestamp 1688980957
transform 1 0 29440 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_122
timestamp 1688980957
transform 1 0 34592 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_123
timestamp 1688980957
transform 1 0 39744 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_124
timestamp 1688980957
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_125
timestamp 1688980957
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_126
timestamp 1688980957
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_127
timestamp 1688980957
transform 1 0 21712 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_128
timestamp 1688980957
transform 1 0 26864 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_129
timestamp 1688980957
transform 1 0 32016 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_130
timestamp 1688980957
transform 1 0 37168 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_131
timestamp 1688980957
transform 1 0 42320 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_132
timestamp 1688980957
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_133
timestamp 1688980957
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_134
timestamp 1688980957
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_135
timestamp 1688980957
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_136
timestamp 1688980957
transform 1 0 24288 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_137
timestamp 1688980957
transform 1 0 29440 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_138
timestamp 1688980957
transform 1 0 34592 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_139
timestamp 1688980957
transform 1 0 39744 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_140
timestamp 1688980957
transform 1 0 3680 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_141
timestamp 1688980957
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_142
timestamp 1688980957
transform 1 0 8832 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_143
timestamp 1688980957
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_144
timestamp 1688980957
transform 1 0 13984 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_145
timestamp 1688980957
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_146
timestamp 1688980957
transform 1 0 19136 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_147
timestamp 1688980957
transform 1 0 21712 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_148
timestamp 1688980957
transform 1 0 24288 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_149
timestamp 1688980957
transform 1 0 26864 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_150
timestamp 1688980957
transform 1 0 29440 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_151
timestamp 1688980957
transform 1 0 32016 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_152
timestamp 1688980957
transform 1 0 34592 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_153
timestamp 1688980957
transform 1 0 37168 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_154
timestamp 1688980957
transform 1 0 39744 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_155
timestamp 1688980957
transform 1 0 42320 0 -1 8704
box -38 -48 130 592
<< labels >>
flabel metal2 s 3238 -300 3294 160 0 FreeSans 224 90 0 0 FrameStrobe[0]
port 0 nsew signal input
flabel metal2 s 24398 -300 24454 160 0 FreeSans 224 90 0 0 FrameStrobe[10]
port 1 nsew signal input
flabel metal2 s 26514 -300 26570 160 0 FreeSans 224 90 0 0 FrameStrobe[11]
port 2 nsew signal input
flabel metal2 s 28630 -300 28686 160 0 FreeSans 224 90 0 0 FrameStrobe[12]
port 3 nsew signal input
flabel metal2 s 30746 -300 30802 160 0 FreeSans 224 90 0 0 FrameStrobe[13]
port 4 nsew signal input
flabel metal2 s 32862 -300 32918 160 0 FreeSans 224 90 0 0 FrameStrobe[14]
port 5 nsew signal input
flabel metal2 s 34978 -300 35034 160 0 FreeSans 224 90 0 0 FrameStrobe[15]
port 6 nsew signal input
flabel metal2 s 37094 -300 37150 160 0 FreeSans 224 90 0 0 FrameStrobe[16]
port 7 nsew signal input
flabel metal2 s 39210 -300 39266 160 0 FreeSans 224 90 0 0 FrameStrobe[17]
port 8 nsew signal input
flabel metal2 s 41326 -300 41382 160 0 FreeSans 224 90 0 0 FrameStrobe[18]
port 9 nsew signal input
flabel metal2 s 43442 -300 43498 160 0 FreeSans 224 90 0 0 FrameStrobe[19]
port 10 nsew signal input
flabel metal2 s 5354 -300 5410 160 0 FreeSans 224 90 0 0 FrameStrobe[1]
port 11 nsew signal input
flabel metal2 s 7470 -300 7526 160 0 FreeSans 224 90 0 0 FrameStrobe[2]
port 12 nsew signal input
flabel metal2 s 9586 -300 9642 160 0 FreeSans 224 90 0 0 FrameStrobe[3]
port 13 nsew signal input
flabel metal2 s 11702 -300 11758 160 0 FreeSans 224 90 0 0 FrameStrobe[4]
port 14 nsew signal input
flabel metal2 s 13818 -300 13874 160 0 FreeSans 224 90 0 0 FrameStrobe[5]
port 15 nsew signal input
flabel metal2 s 15934 -300 15990 160 0 FreeSans 224 90 0 0 FrameStrobe[6]
port 16 nsew signal input
flabel metal2 s 18050 -300 18106 160 0 FreeSans 224 90 0 0 FrameStrobe[7]
port 17 nsew signal input
flabel metal2 s 20166 -300 20222 160 0 FreeSans 224 90 0 0 FrameStrobe[8]
port 18 nsew signal input
flabel metal2 s 22282 -300 22338 160 0 FreeSans 224 90 0 0 FrameStrobe[9]
port 19 nsew signal input
flabel metal2 s 34150 9840 34206 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[0]
port 20 nsew signal tristate
flabel metal2 s 36910 9840 36966 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[10]
port 21 nsew signal tristate
flabel metal2 s 37186 9840 37242 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[11]
port 22 nsew signal tristate
flabel metal2 s 37462 9840 37518 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[12]
port 23 nsew signal tristate
flabel metal2 s 37738 9840 37794 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[13]
port 24 nsew signal tristate
flabel metal2 s 38014 9840 38070 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[14]
port 25 nsew signal tristate
flabel metal2 s 38290 9840 38346 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[15]
port 26 nsew signal tristate
flabel metal2 s 38566 9840 38622 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[16]
port 27 nsew signal tristate
flabel metal2 s 38842 9840 38898 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[17]
port 28 nsew signal tristate
flabel metal2 s 39118 9840 39174 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[18]
port 29 nsew signal tristate
flabel metal2 s 39394 9840 39450 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[19]
port 30 nsew signal tristate
flabel metal2 s 34426 9840 34482 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[1]
port 31 nsew signal tristate
flabel metal2 s 34702 9840 34758 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[2]
port 32 nsew signal tristate
flabel metal2 s 34978 9840 35034 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[3]
port 33 nsew signal tristate
flabel metal2 s 35254 9840 35310 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[4]
port 34 nsew signal tristate
flabel metal2 s 35530 9840 35586 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[5]
port 35 nsew signal tristate
flabel metal2 s 35806 9840 35862 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[6]
port 36 nsew signal tristate
flabel metal2 s 36082 9840 36138 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[7]
port 37 nsew signal tristate
flabel metal2 s 36358 9840 36414 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[8]
port 38 nsew signal tristate
flabel metal2 s 36634 9840 36690 10300 0 FreeSans 224 90 0 0 FrameStrobe_O[9]
port 39 nsew signal tristate
flabel metal2 s 5170 9840 5226 10300 0 FreeSans 224 90 0 0 N1BEG[0]
port 40 nsew signal tristate
flabel metal2 s 5446 9840 5502 10300 0 FreeSans 224 90 0 0 N1BEG[1]
port 41 nsew signal tristate
flabel metal2 s 5722 9840 5778 10300 0 FreeSans 224 90 0 0 N1BEG[2]
port 42 nsew signal tristate
flabel metal2 s 5998 9840 6054 10300 0 FreeSans 224 90 0 0 N1BEG[3]
port 43 nsew signal tristate
flabel metal2 s 6274 9840 6330 10300 0 FreeSans 224 90 0 0 N2BEG[0]
port 44 nsew signal tristate
flabel metal2 s 6550 9840 6606 10300 0 FreeSans 224 90 0 0 N2BEG[1]
port 45 nsew signal tristate
flabel metal2 s 6826 9840 6882 10300 0 FreeSans 224 90 0 0 N2BEG[2]
port 46 nsew signal tristate
flabel metal2 s 7102 9840 7158 10300 0 FreeSans 224 90 0 0 N2BEG[3]
port 47 nsew signal tristate
flabel metal2 s 7378 9840 7434 10300 0 FreeSans 224 90 0 0 N2BEG[4]
port 48 nsew signal tristate
flabel metal2 s 7654 9840 7710 10300 0 FreeSans 224 90 0 0 N2BEG[5]
port 49 nsew signal tristate
flabel metal2 s 7930 9840 7986 10300 0 FreeSans 224 90 0 0 N2BEG[6]
port 50 nsew signal tristate
flabel metal2 s 8206 9840 8262 10300 0 FreeSans 224 90 0 0 N2BEG[7]
port 51 nsew signal tristate
flabel metal2 s 8482 9840 8538 10300 0 FreeSans 224 90 0 0 N2BEGb[0]
port 52 nsew signal tristate
flabel metal2 s 8758 9840 8814 10300 0 FreeSans 224 90 0 0 N2BEGb[1]
port 53 nsew signal tristate
flabel metal2 s 9034 9840 9090 10300 0 FreeSans 224 90 0 0 N2BEGb[2]
port 54 nsew signal tristate
flabel metal2 s 9310 9840 9366 10300 0 FreeSans 224 90 0 0 N2BEGb[3]
port 55 nsew signal tristate
flabel metal2 s 9586 9840 9642 10300 0 FreeSans 224 90 0 0 N2BEGb[4]
port 56 nsew signal tristate
flabel metal2 s 9862 9840 9918 10300 0 FreeSans 224 90 0 0 N2BEGb[5]
port 57 nsew signal tristate
flabel metal2 s 10138 9840 10194 10300 0 FreeSans 224 90 0 0 N2BEGb[6]
port 58 nsew signal tristate
flabel metal2 s 10414 9840 10470 10300 0 FreeSans 224 90 0 0 N2BEGb[7]
port 59 nsew signal tristate
flabel metal2 s 10690 9840 10746 10300 0 FreeSans 224 90 0 0 N4BEG[0]
port 60 nsew signal tristate
flabel metal2 s 13450 9840 13506 10300 0 FreeSans 224 90 0 0 N4BEG[10]
port 61 nsew signal tristate
flabel metal2 s 13726 9840 13782 10300 0 FreeSans 224 90 0 0 N4BEG[11]
port 62 nsew signal tristate
flabel metal2 s 14002 9840 14058 10300 0 FreeSans 224 90 0 0 N4BEG[12]
port 63 nsew signal tristate
flabel metal2 s 14278 9840 14334 10300 0 FreeSans 224 90 0 0 N4BEG[13]
port 64 nsew signal tristate
flabel metal2 s 14554 9840 14610 10300 0 FreeSans 224 90 0 0 N4BEG[14]
port 65 nsew signal tristate
flabel metal2 s 14830 9840 14886 10300 0 FreeSans 224 90 0 0 N4BEG[15]
port 66 nsew signal tristate
flabel metal2 s 10966 9840 11022 10300 0 FreeSans 224 90 0 0 N4BEG[1]
port 67 nsew signal tristate
flabel metal2 s 11242 9840 11298 10300 0 FreeSans 224 90 0 0 N4BEG[2]
port 68 nsew signal tristate
flabel metal2 s 11518 9840 11574 10300 0 FreeSans 224 90 0 0 N4BEG[3]
port 69 nsew signal tristate
flabel metal2 s 11794 9840 11850 10300 0 FreeSans 224 90 0 0 N4BEG[4]
port 70 nsew signal tristate
flabel metal2 s 12070 9840 12126 10300 0 FreeSans 224 90 0 0 N4BEG[5]
port 71 nsew signal tristate
flabel metal2 s 12346 9840 12402 10300 0 FreeSans 224 90 0 0 N4BEG[6]
port 72 nsew signal tristate
flabel metal2 s 12622 9840 12678 10300 0 FreeSans 224 90 0 0 N4BEG[7]
port 73 nsew signal tristate
flabel metal2 s 12898 9840 12954 10300 0 FreeSans 224 90 0 0 N4BEG[8]
port 74 nsew signal tristate
flabel metal2 s 13174 9840 13230 10300 0 FreeSans 224 90 0 0 N4BEG[9]
port 75 nsew signal tristate
flabel metal2 s 15106 9840 15162 10300 0 FreeSans 224 90 0 0 NN4BEG[0]
port 76 nsew signal tristate
flabel metal2 s 17866 9840 17922 10300 0 FreeSans 224 90 0 0 NN4BEG[10]
port 77 nsew signal tristate
flabel metal2 s 18142 9840 18198 10300 0 FreeSans 224 90 0 0 NN4BEG[11]
port 78 nsew signal tristate
flabel metal2 s 18418 9840 18474 10300 0 FreeSans 224 90 0 0 NN4BEG[12]
port 79 nsew signal tristate
flabel metal2 s 18694 9840 18750 10300 0 FreeSans 224 90 0 0 NN4BEG[13]
port 80 nsew signal tristate
flabel metal2 s 18970 9840 19026 10300 0 FreeSans 224 90 0 0 NN4BEG[14]
port 81 nsew signal tristate
flabel metal2 s 19246 9840 19302 10300 0 FreeSans 224 90 0 0 NN4BEG[15]
port 82 nsew signal tristate
flabel metal2 s 15382 9840 15438 10300 0 FreeSans 224 90 0 0 NN4BEG[1]
port 83 nsew signal tristate
flabel metal2 s 15658 9840 15714 10300 0 FreeSans 224 90 0 0 NN4BEG[2]
port 84 nsew signal tristate
flabel metal2 s 15934 9840 15990 10300 0 FreeSans 224 90 0 0 NN4BEG[3]
port 85 nsew signal tristate
flabel metal2 s 16210 9840 16266 10300 0 FreeSans 224 90 0 0 NN4BEG[4]
port 86 nsew signal tristate
flabel metal2 s 16486 9840 16542 10300 0 FreeSans 224 90 0 0 NN4BEG[5]
port 87 nsew signal tristate
flabel metal2 s 16762 9840 16818 10300 0 FreeSans 224 90 0 0 NN4BEG[6]
port 88 nsew signal tristate
flabel metal2 s 17038 9840 17094 10300 0 FreeSans 224 90 0 0 NN4BEG[7]
port 89 nsew signal tristate
flabel metal2 s 17314 9840 17370 10300 0 FreeSans 224 90 0 0 NN4BEG[8]
port 90 nsew signal tristate
flabel metal2 s 17590 9840 17646 10300 0 FreeSans 224 90 0 0 NN4BEG[9]
port 91 nsew signal tristate
flabel metal2 s 19522 9840 19578 10300 0 FreeSans 224 90 0 0 S1END[0]
port 92 nsew signal input
flabel metal2 s 19798 9840 19854 10300 0 FreeSans 224 90 0 0 S1END[1]
port 93 nsew signal input
flabel metal2 s 20074 9840 20130 10300 0 FreeSans 224 90 0 0 S1END[2]
port 94 nsew signal input
flabel metal2 s 20350 9840 20406 10300 0 FreeSans 224 90 0 0 S1END[3]
port 95 nsew signal input
flabel metal2 s 20626 9840 20682 10300 0 FreeSans 224 90 0 0 S2END[0]
port 96 nsew signal input
flabel metal2 s 20902 9840 20958 10300 0 FreeSans 224 90 0 0 S2END[1]
port 97 nsew signal input
flabel metal2 s 21178 9840 21234 10300 0 FreeSans 224 90 0 0 S2END[2]
port 98 nsew signal input
flabel metal2 s 21454 9840 21510 10300 0 FreeSans 224 90 0 0 S2END[3]
port 99 nsew signal input
flabel metal2 s 21730 9840 21786 10300 0 FreeSans 224 90 0 0 S2END[4]
port 100 nsew signal input
flabel metal2 s 22006 9840 22062 10300 0 FreeSans 224 90 0 0 S2END[5]
port 101 nsew signal input
flabel metal2 s 22282 9840 22338 10300 0 FreeSans 224 90 0 0 S2END[6]
port 102 nsew signal input
flabel metal2 s 22558 9840 22614 10300 0 FreeSans 224 90 0 0 S2END[7]
port 103 nsew signal input
flabel metal2 s 22834 9840 22890 10300 0 FreeSans 224 90 0 0 S2MID[0]
port 104 nsew signal input
flabel metal2 s 23110 9840 23166 10300 0 FreeSans 224 90 0 0 S2MID[1]
port 105 nsew signal input
flabel metal2 s 23386 9840 23442 10300 0 FreeSans 224 90 0 0 S2MID[2]
port 106 nsew signal input
flabel metal2 s 23662 9840 23718 10300 0 FreeSans 224 90 0 0 S2MID[3]
port 107 nsew signal input
flabel metal2 s 23938 9840 23994 10300 0 FreeSans 224 90 0 0 S2MID[4]
port 108 nsew signal input
flabel metal2 s 24214 9840 24270 10300 0 FreeSans 224 90 0 0 S2MID[5]
port 109 nsew signal input
flabel metal2 s 24490 9840 24546 10300 0 FreeSans 224 90 0 0 S2MID[6]
port 110 nsew signal input
flabel metal2 s 24766 9840 24822 10300 0 FreeSans 224 90 0 0 S2MID[7]
port 111 nsew signal input
flabel metal2 s 25042 9840 25098 10300 0 FreeSans 224 90 0 0 S4END[0]
port 112 nsew signal input
flabel metal2 s 27802 9840 27858 10300 0 FreeSans 224 90 0 0 S4END[10]
port 113 nsew signal input
flabel metal2 s 28078 9840 28134 10300 0 FreeSans 224 90 0 0 S4END[11]
port 114 nsew signal input
flabel metal2 s 28354 9840 28410 10300 0 FreeSans 224 90 0 0 S4END[12]
port 115 nsew signal input
flabel metal2 s 28630 9840 28686 10300 0 FreeSans 224 90 0 0 S4END[13]
port 116 nsew signal input
flabel metal2 s 28906 9840 28962 10300 0 FreeSans 224 90 0 0 S4END[14]
port 117 nsew signal input
flabel metal2 s 29182 9840 29238 10300 0 FreeSans 224 90 0 0 S4END[15]
port 118 nsew signal input
flabel metal2 s 25318 9840 25374 10300 0 FreeSans 224 90 0 0 S4END[1]
port 119 nsew signal input
flabel metal2 s 25594 9840 25650 10300 0 FreeSans 224 90 0 0 S4END[2]
port 120 nsew signal input
flabel metal2 s 25870 9840 25926 10300 0 FreeSans 224 90 0 0 S4END[3]
port 121 nsew signal input
flabel metal2 s 26146 9840 26202 10300 0 FreeSans 224 90 0 0 S4END[4]
port 122 nsew signal input
flabel metal2 s 26422 9840 26478 10300 0 FreeSans 224 90 0 0 S4END[5]
port 123 nsew signal input
flabel metal2 s 26698 9840 26754 10300 0 FreeSans 224 90 0 0 S4END[6]
port 124 nsew signal input
flabel metal2 s 26974 9840 27030 10300 0 FreeSans 224 90 0 0 S4END[7]
port 125 nsew signal input
flabel metal2 s 27250 9840 27306 10300 0 FreeSans 224 90 0 0 S4END[8]
port 126 nsew signal input
flabel metal2 s 27526 9840 27582 10300 0 FreeSans 224 90 0 0 S4END[9]
port 127 nsew signal input
flabel metal2 s 29458 9840 29514 10300 0 FreeSans 224 90 0 0 SS4END[0]
port 128 nsew signal input
flabel metal2 s 32218 9840 32274 10300 0 FreeSans 224 90 0 0 SS4END[10]
port 129 nsew signal input
flabel metal2 s 32494 9840 32550 10300 0 FreeSans 224 90 0 0 SS4END[11]
port 130 nsew signal input
flabel metal2 s 32770 9840 32826 10300 0 FreeSans 224 90 0 0 SS4END[12]
port 131 nsew signal input
flabel metal2 s 33046 9840 33102 10300 0 FreeSans 224 90 0 0 SS4END[13]
port 132 nsew signal input
flabel metal2 s 33322 9840 33378 10300 0 FreeSans 224 90 0 0 SS4END[14]
port 133 nsew signal input
flabel metal2 s 33598 9840 33654 10300 0 FreeSans 224 90 0 0 SS4END[15]
port 134 nsew signal input
flabel metal2 s 29734 9840 29790 10300 0 FreeSans 224 90 0 0 SS4END[1]
port 135 nsew signal input
flabel metal2 s 30010 9840 30066 10300 0 FreeSans 224 90 0 0 SS4END[2]
port 136 nsew signal input
flabel metal2 s 30286 9840 30342 10300 0 FreeSans 224 90 0 0 SS4END[3]
port 137 nsew signal input
flabel metal2 s 30562 9840 30618 10300 0 FreeSans 224 90 0 0 SS4END[4]
port 138 nsew signal input
flabel metal2 s 30838 9840 30894 10300 0 FreeSans 224 90 0 0 SS4END[5]
port 139 nsew signal input
flabel metal2 s 31114 9840 31170 10300 0 FreeSans 224 90 0 0 SS4END[6]
port 140 nsew signal input
flabel metal2 s 31390 9840 31446 10300 0 FreeSans 224 90 0 0 SS4END[7]
port 141 nsew signal input
flabel metal2 s 31666 9840 31722 10300 0 FreeSans 224 90 0 0 SS4END[8]
port 142 nsew signal input
flabel metal2 s 31942 9840 31998 10300 0 FreeSans 224 90 0 0 SS4END[9]
port 143 nsew signal input
flabel metal2 s 1122 -300 1178 160 0 FreeSans 224 90 0 0 UserCLK
port 144 nsew signal input
flabel metal2 s 33874 9840 33930 10300 0 FreeSans 224 90 0 0 UserCLKo
port 145 nsew signal tristate
flabel metal4 s 6245 1040 6565 8752 0 FreeSans 1920 90 0 0 vccd1
port 146 nsew power bidirectional
flabel metal4 s 16848 1040 17168 8752 0 FreeSans 1920 90 0 0 vccd1
port 146 nsew power bidirectional
flabel metal4 s 27451 1040 27771 8752 0 FreeSans 1920 90 0 0 vccd1
port 146 nsew power bidirectional
flabel metal4 s 38054 1040 38374 8752 0 FreeSans 1920 90 0 0 vccd1
port 146 nsew power bidirectional
flabel metal4 s 11546 1040 11866 8752 0 FreeSans 1920 90 0 0 vssd1
port 147 nsew ground bidirectional
flabel metal4 s 22149 1040 22469 8752 0 FreeSans 1920 90 0 0 vssd1
port 147 nsew ground bidirectional
flabel metal4 s 32752 1040 33072 8752 0 FreeSans 1920 90 0 0 vssd1
port 147 nsew ground bidirectional
flabel metal4 s 43355 1040 43675 8752 0 FreeSans 1920 90 0 0 vssd1
port 147 nsew ground bidirectional
rlabel metal1 22310 8160 22310 8160 0 vccd1
rlabel via1 22389 8704 22389 8704 0 vssd1
rlabel metal2 3319 68 3319 68 0 FrameStrobe[0]
rlabel metal2 24479 68 24479 68 0 FrameStrobe[10]
rlabel metal2 26595 68 26595 68 0 FrameStrobe[11]
rlabel metal2 28711 68 28711 68 0 FrameStrobe[12]
rlabel metal2 30827 68 30827 68 0 FrameStrobe[13]
rlabel metal2 32791 68 32791 68 0 FrameStrobe[14]
rlabel metal2 35059 68 35059 68 0 FrameStrobe[15]
rlabel metal2 37122 415 37122 415 0 FrameStrobe[16]
rlabel metal2 39383 68 39383 68 0 FrameStrobe[17]
rlabel metal2 41354 704 41354 704 0 FrameStrobe[18]
rlabel metal2 43325 68 43325 68 0 FrameStrobe[19]
rlabel metal2 5435 68 5435 68 0 FrameStrobe[1]
rlabel metal2 7551 68 7551 68 0 FrameStrobe[2]
rlabel metal2 9667 68 9667 68 0 FrameStrobe[3]
rlabel metal2 11829 68 11829 68 0 FrameStrobe[4]
rlabel metal2 13991 68 13991 68 0 FrameStrobe[5]
rlabel metal2 16015 68 16015 68 0 FrameStrobe[6]
rlabel metal2 18131 68 18131 68 0 FrameStrobe[7]
rlabel metal2 20247 68 20247 68 0 FrameStrobe[8]
rlabel metal2 22455 68 22455 68 0 FrameStrobe[9]
rlabel metal2 34178 9445 34178 9445 0 FrameStrobe_O[0]
rlabel metal1 37812 6766 37812 6766 0 FrameStrobe_O[10]
rlabel metal1 37996 6698 37996 6698 0 FrameStrobe_O[11]
rlabel metal2 37490 9717 37490 9717 0 FrameStrobe_O[12]
rlabel metal2 37766 8952 37766 8952 0 FrameStrobe_O[13]
rlabel metal2 38042 9649 38042 9649 0 FrameStrobe_O[14]
rlabel metal2 38318 9785 38318 9785 0 FrameStrobe_O[15]
rlabel metal1 38870 6834 38870 6834 0 FrameStrobe_O[16]
rlabel metal2 38870 8952 38870 8952 0 FrameStrobe_O[17]
rlabel metal2 39146 8918 39146 8918 0 FrameStrobe_O[18]
rlabel metal2 39422 9785 39422 9785 0 FrameStrobe_O[19]
rlabel metal2 34454 9088 34454 9088 0 FrameStrobe_O[1]
rlabel metal2 34730 9530 34730 9530 0 FrameStrobe_O[2]
rlabel metal1 36570 8568 36570 8568 0 FrameStrobe_O[3]
rlabel metal2 35282 8782 35282 8782 0 FrameStrobe_O[4]
rlabel metal2 35558 9037 35558 9037 0 FrameStrobe_O[5]
rlabel metal2 35834 9088 35834 9088 0 FrameStrobe_O[6]
rlabel metal2 36110 8952 36110 8952 0 FrameStrobe_O[7]
rlabel metal2 36386 9445 36386 9445 0 FrameStrobe_O[8]
rlabel metal2 36662 9513 36662 9513 0 FrameStrobe_O[9]
rlabel metal1 22402 2618 22402 2618 0 FrameStrobe_O_i\[0\]
rlabel metal1 25484 4250 25484 4250 0 FrameStrobe_O_i\[10\]
rlabel metal1 27278 4012 27278 4012 0 FrameStrobe_O_i\[11\]
rlabel metal1 29716 3162 29716 3162 0 FrameStrobe_O_i\[12\]
rlabel metal1 32154 4012 32154 4012 0 FrameStrobe_O_i\[13\]
rlabel metal1 37168 4794 37168 4794 0 FrameStrobe_O_i\[14\]
rlabel metal1 36662 3162 36662 3162 0 FrameStrobe_O_i\[15\]
rlabel metal1 37858 4250 37858 4250 0 FrameStrobe_O_i\[16\]
rlabel metal2 39054 2244 39054 2244 0 FrameStrobe_O_i\[17\]
rlabel metal1 40158 3706 40158 3706 0 FrameStrobe_O_i\[18\]
rlabel metal2 40250 2822 40250 2822 0 FrameStrobe_O_i\[19\]
rlabel metal1 22402 3910 22402 3910 0 FrameStrobe_O_i\[1\]
rlabel metal2 22586 4420 22586 4420 0 FrameStrobe_O_i\[2\]
rlabel metal1 22310 3706 22310 3706 0 FrameStrobe_O_i\[3\]
rlabel metal1 22632 3910 22632 3910 0 FrameStrobe_O_i\[4\]
rlabel metal1 21804 3162 21804 3162 0 FrameStrobe_O_i\[5\]
rlabel metal2 21298 3298 21298 3298 0 FrameStrobe_O_i\[6\]
rlabel metal1 19136 3162 19136 3162 0 FrameStrobe_O_i\[7\]
rlabel metal1 21252 4250 21252 4250 0 FrameStrobe_O_i\[8\]
rlabel metal1 23368 3706 23368 3706 0 FrameStrobe_O_i\[9\]
rlabel metal1 4876 8330 4876 8330 0 N1BEG[0]
rlabel metal1 5290 8602 5290 8602 0 N1BEG[1]
rlabel metal1 5704 8602 5704 8602 0 N1BEG[2]
rlabel metal2 6026 8952 6026 8952 0 N1BEG[3]
rlabel metal1 6164 8602 6164 8602 0 N2BEG[0]
rlabel metal2 6578 9326 6578 9326 0 N2BEG[1]
rlabel metal1 6808 8602 6808 8602 0 N2BEG[2]
rlabel metal2 7130 8952 7130 8952 0 N2BEG[3]
rlabel metal1 7268 7242 7268 7242 0 N2BEG[4]
rlabel metal1 7406 8330 7406 8330 0 N2BEG[5]
rlabel metal1 7728 8602 7728 8602 0 N2BEG[6]
rlabel metal2 8234 8952 8234 8952 0 N2BEG[7]
rlabel metal1 8280 8602 8280 8602 0 N2BEGb[0]
rlabel metal2 8786 8952 8786 8952 0 N2BEGb[1]
rlabel metal1 8648 7242 8648 7242 0 N2BEGb[2]
rlabel metal2 9338 8952 9338 8952 0 N2BEGb[3]
rlabel metal1 8602 8568 8602 8568 0 N2BEGb[4]
rlabel metal1 9706 8602 9706 8602 0 N2BEGb[5]
rlabel metal1 9706 6834 9706 6834 0 N2BEGb[6]
rlabel metal2 10442 8952 10442 8952 0 N2BEGb[7]
rlabel metal1 10396 7990 10396 7990 0 N4BEG[0]
rlabel metal2 13478 8952 13478 8952 0 N4BEG[10]
rlabel metal1 13386 8602 13386 8602 0 N4BEG[11]
rlabel metal1 13892 8602 13892 8602 0 N4BEG[12]
rlabel metal2 14306 8952 14306 8952 0 N4BEG[13]
rlabel metal1 14536 7514 14536 7514 0 N4BEG[14]
rlabel metal2 14858 8952 14858 8952 0 N4BEG[15]
rlabel metal1 10902 8602 10902 8602 0 N4BEG[1]
rlabel metal2 11270 8952 11270 8952 0 N4BEG[2]
rlabel metal1 10258 8568 10258 8568 0 N4BEG[3]
rlabel metal2 11822 9326 11822 9326 0 N4BEG[4]
rlabel metal1 11638 8602 11638 8602 0 N4BEG[5]
rlabel metal1 12328 8602 12328 8602 0 N4BEG[6]
rlabel metal2 12650 8952 12650 8952 0 N4BEG[7]
rlabel metal1 11730 8364 11730 8364 0 N4BEG[8]
rlabel metal1 12972 8602 12972 8602 0 N4BEG[9]
rlabel metal1 14674 8568 14674 8568 0 NN4BEG[0]
rlabel metal1 17848 8602 17848 8602 0 NN4BEG[10]
rlabel metal2 18170 9224 18170 9224 0 NN4BEG[11]
rlabel metal1 18492 8058 18492 8058 0 NN4BEG[12]
rlabel metal1 19090 8330 19090 8330 0 NN4BEG[13]
rlabel metal2 19366 8857 19366 8857 0 NN4BEG[14]
rlabel metal1 18998 8602 18998 8602 0 NN4BEG[15]
rlabel metal1 15226 8602 15226 8602 0 NN4BEG[1]
rlabel metal1 15640 8058 15640 8058 0 NN4BEG[2]
rlabel metal2 15962 8952 15962 8952 0 NN4BEG[3]
rlabel metal1 16008 8602 16008 8602 0 NN4BEG[4]
rlabel metal2 16514 8952 16514 8952 0 NN4BEG[5]
rlabel metal1 16560 8602 16560 8602 0 NN4BEG[6]
rlabel metal2 17066 9309 17066 9309 0 NN4BEG[7]
rlabel metal1 16882 8568 16882 8568 0 NN4BEG[8]
rlabel metal1 17434 8602 17434 8602 0 NN4BEG[9]
rlabel metal2 19550 9836 19550 9836 0 S1END[0]
rlabel metal2 19826 9224 19826 9224 0 S1END[1]
rlabel metal2 20102 9241 20102 9241 0 S1END[2]
rlabel metal2 20378 9360 20378 9360 0 S1END[3]
rlabel metal2 20654 9156 20654 9156 0 S2END[0]
rlabel metal2 20930 9156 20930 9156 0 S2END[1]
rlabel metal2 21206 9156 21206 9156 0 S2END[2]
rlabel metal2 21482 9156 21482 9156 0 S2END[3]
rlabel metal2 21758 9156 21758 9156 0 S2END[4]
rlabel metal2 22034 9156 22034 9156 0 S2END[5]
rlabel metal2 22310 9513 22310 9513 0 S2END[6]
rlabel metal2 22586 9564 22586 9564 0 S2END[7]
rlabel metal2 22862 9513 22862 9513 0 S2MID[0]
rlabel metal2 23138 9513 23138 9513 0 S2MID[1]
rlabel metal2 23414 9513 23414 9513 0 S2MID[2]
rlabel metal2 23690 9513 23690 9513 0 S2MID[3]
rlabel metal2 23966 9513 23966 9513 0 S2MID[4]
rlabel metal2 24242 9156 24242 9156 0 S2MID[5]
rlabel metal2 24518 9156 24518 9156 0 S2MID[6]
rlabel metal2 24794 9156 24794 9156 0 S2MID[7]
rlabel metal2 25070 9156 25070 9156 0 S4END[0]
rlabel metal2 27830 9156 27830 9156 0 S4END[10]
rlabel metal2 28106 9190 28106 9190 0 S4END[11]
rlabel metal2 28382 9836 28382 9836 0 S4END[12]
rlabel metal2 28658 9156 28658 9156 0 S4END[13]
rlabel metal2 28934 9513 28934 9513 0 S4END[14]
rlabel metal2 29210 9122 29210 9122 0 S4END[15]
rlabel metal2 25346 9156 25346 9156 0 S4END[1]
rlabel metal2 25622 9156 25622 9156 0 S4END[2]
rlabel metal2 25898 9513 25898 9513 0 S4END[3]
rlabel metal2 26174 9156 26174 9156 0 S4END[4]
rlabel metal2 26450 9156 26450 9156 0 S4END[5]
rlabel metal2 26726 9156 26726 9156 0 S4END[6]
rlabel metal2 27002 9190 27002 9190 0 S4END[7]
rlabel metal2 27278 9156 27278 9156 0 S4END[8]
rlabel metal2 27554 9224 27554 9224 0 S4END[9]
rlabel metal2 29486 9513 29486 9513 0 SS4END[0]
rlabel metal2 32246 9190 32246 9190 0 SS4END[10]
rlabel metal2 32522 9224 32522 9224 0 SS4END[11]
rlabel metal2 32798 9513 32798 9513 0 SS4END[12]
rlabel metal2 33074 9377 33074 9377 0 SS4END[13]
rlabel metal2 33350 8850 33350 8850 0 SS4END[14]
rlabel metal2 33626 9513 33626 9513 0 SS4END[15]
rlabel metal2 29762 9224 29762 9224 0 SS4END[1]
rlabel metal2 30038 9173 30038 9173 0 SS4END[2]
rlabel metal2 30314 9088 30314 9088 0 SS4END[3]
rlabel metal2 30590 9190 30590 9190 0 SS4END[4]
rlabel metal2 30866 9224 30866 9224 0 SS4END[5]
rlabel metal2 31142 9513 31142 9513 0 SS4END[6]
rlabel metal1 31970 8432 31970 8432 0 SS4END[7]
rlabel metal2 31786 8585 31786 8585 0 SS4END[8]
rlabel metal2 31970 9513 31970 9513 0 SS4END[9]
rlabel metal2 1150 704 1150 704 0 UserCLK
rlabel metal1 34040 8602 34040 8602 0 UserCLKo
rlabel metal2 3542 1972 3542 1972 0 net1
rlabel metal1 41078 1190 41078 1190 0 net10
rlabel metal1 7038 8466 7038 8466 0 net100
rlabel metal1 9706 7718 9706 7718 0 net101
rlabel metal1 9844 6970 9844 6970 0 net102
rlabel metal1 11822 8296 11822 8296 0 net103
rlabel metal1 8602 9724 8602 9724 0 net104
rlabel metal2 8142 7344 8142 7344 0 net105
rlabel metal1 8280 8534 8280 8534 0 net106
rlabel metal2 9522 7616 9522 7616 0 net107
rlabel metal1 8786 7276 8786 7276 0 net108
rlabel metal1 9614 7344 9614 7344 0 net109
rlabel metal2 43010 1972 43010 1972 0 net11
rlabel metal2 8694 8670 8694 8670 0 net110
rlabel metal1 11638 8466 11638 8466 0 net111
rlabel metal2 9706 8636 9706 8636 0 net112
rlabel metal2 17986 7242 17986 7242 0 net113
rlabel via2 11914 7803 11914 7803 0 net114
rlabel metal2 13754 7905 13754 7905 0 net115
rlabel metal3 21804 8976 21804 8976 0 net116
rlabel metal2 13846 8738 13846 8738 0 net117
rlabel metal2 19412 7854 19412 7854 0 net118
rlabel metal2 14674 7174 14674 7174 0 net119
rlabel metal1 5658 1258 5658 1258 0 net12
rlabel metal2 17526 7140 17526 7140 0 net120
rlabel metal1 11040 8466 11040 8466 0 net121
rlabel metal2 13662 7786 13662 7786 0 net122
rlabel metal2 10810 9044 10810 9044 0 net123
rlabel metal1 25254 8058 25254 8058 0 net124
rlabel metal1 11362 9248 11362 9248 0 net125
rlabel metal2 12558 8840 12558 8840 0 net126
rlabel metal3 21436 7412 21436 7412 0 net127
rlabel metal1 12282 9214 12282 9214 0 net128
rlabel via2 21850 9163 21850 9163 0 net129
rlabel metal2 7774 2618 7774 2618 0 net13
rlabel metal2 21206 8041 21206 8041 0 net130
rlabel metal1 18170 7514 18170 7514 0 net131
rlabel metal2 17802 8228 17802 8228 0 net132
rlabel metal1 18768 7514 18768 7514 0 net133
rlabel metal2 19274 8007 19274 8007 0 net134
rlabel metal1 19688 7514 19688 7514 0 net135
rlabel metal1 18998 8432 18998 8432 0 net136
rlabel metal2 20930 8177 20930 8177 0 net137
rlabel metal1 21666 7174 21666 7174 0 net138
rlabel metal1 16330 7854 16330 7854 0 net139
rlabel metal2 9890 1088 9890 1088 0 net14
rlabel metal1 20838 7174 20838 7174 0 net140
rlabel metal1 17158 7854 17158 7854 0 net141
rlabel metal1 19872 7174 19872 7174 0 net142
rlabel metal1 17940 7242 17940 7242 0 net143
rlabel metal1 17480 7514 17480 7514 0 net144
rlabel metal2 17434 7820 17434 7820 0 net145
rlabel metal1 27784 1734 27784 1734 0 net146
rlabel metal2 18262 1258 18262 1258 0 net15
rlabel metal1 18078 1360 18078 1360 0 net16
rlabel metal1 18676 2958 18676 2958 0 net17
rlabel metal1 18492 1190 18492 1190 0 net18
rlabel metal1 20608 4114 20608 4114 0 net19
rlabel metal1 24748 1190 24748 1190 0 net2
rlabel metal1 22678 1190 22678 1190 0 net20
rlabel metal1 18952 6630 18952 6630 0 net21
rlabel metal1 19918 6664 19918 6664 0 net22
rlabel metal1 20102 7514 20102 7514 0 net23
rlabel metal1 19504 7854 19504 7854 0 net24
rlabel metal1 20056 7854 20056 7854 0 net25
rlabel metal1 20332 7854 20332 7854 0 net26
rlabel metal1 20838 7446 20838 7446 0 net27
rlabel metal1 20562 7888 20562 7888 0 net28
rlabel metal1 21482 7378 21482 7378 0 net29
rlabel metal1 26956 1190 26956 1190 0 net3
rlabel metal2 22034 7667 22034 7667 0 net30
rlabel metal1 21850 7886 21850 7886 0 net31
rlabel metal1 22126 7786 22126 7786 0 net32
rlabel metal1 22218 7820 22218 7820 0 net33
rlabel metal1 23000 7378 23000 7378 0 net34
rlabel metal1 22770 7888 22770 7888 0 net35
rlabel metal1 23046 7820 23046 7820 0 net36
rlabel metal1 23598 7820 23598 7820 0 net37
rlabel metal2 24610 8058 24610 8058 0 net38
rlabel metal2 24886 8058 24886 8058 0 net39
rlabel metal1 28934 1258 28934 1258 0 net4
rlabel metal2 25162 8058 25162 8058 0 net40
rlabel metal2 25438 8058 25438 8058 0 net41
rlabel metal1 27094 7888 27094 7888 0 net42
rlabel metal1 25714 7922 25714 7922 0 net43
rlabel metal2 23874 7548 23874 7548 0 net44
rlabel metal1 24150 7888 24150 7888 0 net45
rlabel metal2 23322 7684 23322 7684 0 net46
rlabel metal1 28934 8568 28934 8568 0 net47
rlabel metal1 24978 7412 24978 7412 0 net48
rlabel metal2 25990 8058 25990 8058 0 net49
rlabel metal1 31188 1190 31188 1190 0 net5
rlabel metal2 26266 8058 26266 8058 0 net50
rlabel metal2 26542 8058 26542 8058 0 net51
rlabel metal2 26818 8058 26818 8058 0 net52
rlabel metal1 26358 7412 26358 7412 0 net53
rlabel metal2 27370 8058 27370 8058 0 net54
rlabel metal1 27738 7854 27738 7854 0 net55
rlabel metal1 27968 7854 27968 7854 0 net56
rlabel metal1 29026 8296 29026 8296 0 net57
rlabel metal1 32430 8262 32430 8262 0 net58
rlabel metal2 25438 8772 25438 8772 0 net59
rlabel metal1 33856 1190 33856 1190 0 net6
rlabel metal1 33350 8262 33350 8262 0 net60
rlabel metal2 24610 9044 24610 9044 0 net61
rlabel metal1 33442 7344 33442 7344 0 net62
rlabel metal2 33626 8143 33626 8143 0 net63
rlabel metal3 21988 8840 21988 8840 0 net64
rlabel metal2 18906 8279 18906 8279 0 net65
rlabel metal1 19458 8568 19458 8568 0 net66
rlabel metal2 30958 8670 30958 8670 0 net67
rlabel metal2 18630 8398 18630 8398 0 net68
rlabel metal2 21850 9435 21850 9435 0 net69
rlabel metal1 35282 1258 35282 1258 0 net7
rlabel metal1 17802 9724 17802 9724 0 net70
rlabel metal1 32016 8602 32016 8602 0 net71
rlabel metal3 21620 7548 21620 7548 0 net72
rlabel metal2 1610 1734 1610 1734 0 net73
rlabel metal3 34661 8364 34661 8364 0 net74
rlabel metal1 38272 8534 38272 8534 0 net75
rlabel metal1 37996 7854 37996 7854 0 net76
rlabel metal1 39054 8568 39054 8568 0 net77
rlabel metal2 37950 6256 37950 6256 0 net78
rlabel metal1 38456 5338 38456 5338 0 net79
rlabel metal1 37490 1258 37490 1258 0 net8
rlabel metal1 38456 3706 38456 3706 0 net80
rlabel metal1 38318 4794 38318 4794 0 net81
rlabel metal1 39606 2618 39606 2618 0 net82
rlabel metal1 39928 3910 39928 3910 0 net83
rlabel metal1 40526 3162 40526 3162 0 net84
rlabel metal2 23046 5202 23046 5202 0 net85
rlabel metal2 35926 8704 35926 8704 0 net86
rlabel metal1 36478 8432 36478 8432 0 net87
rlabel metal2 36846 6290 36846 6290 0 net88
rlabel metal1 35742 3468 35742 3468 0 net89
rlabel metal1 39100 1530 39100 1530 0 net9
rlabel metal2 36662 5916 36662 5916 0 net90
rlabel metal2 36294 5712 36294 5712 0 net91
rlabel metal1 37766 8534 37766 8534 0 net92
rlabel metal1 37398 7888 37398 7888 0 net93
rlabel metal1 4738 9384 4738 9384 0 net94
rlabel metal1 5382 8534 5382 8534 0 net95
rlabel metal1 5750 8500 5750 8500 0 net96
rlabel metal2 6302 7650 6302 7650 0 net97
rlabel metal2 6210 8636 6210 8636 0 net98
rlabel metal2 6854 7055 6854 7055 0 net99
<< properties >>
string FIXED_BBOX 0 0 44700 10000
<< end >>
