magic
tech sky130A
magscale 1 2
timestamp 1734828900
<< viali >>
rect 2237 43401 2271 43435
rect 3157 43401 3191 43435
rect 3985 43401 4019 43435
rect 5273 43401 5307 43435
rect 5825 43401 5859 43435
rect 6837 43401 6871 43435
rect 8309 43401 8343 43435
rect 8677 43401 8711 43435
rect 9137 43401 9171 43435
rect 12173 43401 12207 43435
rect 12449 43401 12483 43435
rect 13921 43401 13955 43435
rect 16865 43401 16899 43435
rect 17417 43401 17451 43435
rect 17785 43401 17819 43435
rect 18153 43401 18187 43435
rect 19441 43401 19475 43435
rect 2881 43333 2915 43367
rect 4997 43333 5031 43367
rect 7849 43333 7883 43367
rect 9781 43333 9815 43367
rect 10333 43333 10367 43367
rect 10885 43333 10919 43367
rect 12357 43333 12391 43367
rect 12909 43333 12943 43367
rect 20821 43333 20855 43367
rect 1961 43265 1995 43299
rect 2053 43265 2087 43299
rect 2513 43265 2547 43299
rect 3065 43265 3099 43299
rect 3801 43265 3835 43299
rect 4169 43265 4203 43299
rect 4629 43265 4663 43299
rect 5181 43265 5215 43299
rect 5733 43265 5767 43299
rect 6561 43265 6595 43299
rect 7021 43265 7055 43299
rect 7481 43265 7515 43299
rect 8033 43265 8067 43299
rect 8493 43265 8527 43299
rect 8953 43265 8987 43299
rect 9321 43265 9355 43299
rect 11345 43265 11379 43299
rect 11713 43265 11747 43299
rect 11989 43265 12023 43299
rect 13645 43265 13679 43299
rect 13737 43265 13771 43299
rect 14105 43265 14139 43299
rect 14473 43265 14507 43299
rect 15025 43265 15059 43299
rect 15301 43265 15335 43299
rect 15577 43265 15611 43299
rect 15853 43265 15887 43299
rect 16129 43265 16163 43299
rect 16405 43265 16439 43299
rect 16773 43265 16807 43299
rect 17233 43265 17267 43299
rect 17601 43265 17635 43299
rect 18061 43265 18095 43299
rect 18613 43265 18647 43299
rect 19349 43265 19383 43299
rect 19901 43265 19935 43299
rect 20453 43265 20487 43299
rect 21005 43265 21039 43299
rect 1777 43129 1811 43163
rect 11069 43129 11103 43163
rect 13093 43129 13127 43163
rect 13461 43129 13495 43163
rect 16221 43129 16255 43163
rect 4353 43061 4387 43095
rect 7205 43061 7239 43095
rect 9505 43061 9539 43095
rect 9873 43061 9907 43095
rect 10425 43061 10459 43095
rect 11161 43061 11195 43095
rect 11897 43061 11931 43095
rect 14289 43061 14323 43095
rect 14657 43061 14691 43095
rect 14841 43061 14875 43095
rect 15117 43061 15151 43095
rect 15393 43061 15427 43095
rect 15669 43061 15703 43095
rect 15945 43061 15979 43095
rect 18705 43061 18739 43095
rect 19993 43061 20027 43095
rect 21097 43061 21131 43095
rect 5365 42857 5399 42891
rect 11529 42857 11563 42891
rect 17233 42857 17267 42891
rect 17785 42857 17819 42891
rect 20545 42857 20579 42891
rect 2973 42789 3007 42823
rect 3525 42721 3559 42755
rect 4261 42721 4295 42755
rect 4813 42721 4847 42755
rect 6469 42721 6503 42755
rect 7021 42721 7055 42755
rect 7573 42721 7607 42755
rect 8125 42721 8159 42755
rect 8677 42721 8711 42755
rect 9689 42721 9723 42755
rect 18521 42721 18555 42755
rect 19625 42721 19659 42755
rect 21281 42721 21315 42755
rect 1961 42653 1995 42687
rect 2513 42653 2547 42687
rect 3249 42653 3283 42687
rect 6009 42653 6043 42687
rect 9137 42653 9171 42687
rect 9873 42653 9907 42687
rect 10517 42653 10551 42687
rect 10793 42653 10827 42687
rect 11069 42653 11103 42687
rect 11345 42653 11379 42687
rect 11713 42653 11747 42687
rect 11897 42653 11931 42687
rect 12173 42653 12207 42687
rect 12633 42653 12667 42687
rect 13093 42653 13127 42687
rect 13185 42653 13219 42687
rect 13645 42653 13679 42687
rect 14197 42653 14231 42687
rect 14657 42653 14691 42687
rect 14933 42653 14967 42687
rect 18889 42653 18923 42687
rect 2145 42585 2179 42619
rect 2697 42585 2731 42619
rect 3985 42585 4019 42619
rect 4537 42585 4571 42619
rect 5089 42585 5123 42619
rect 5641 42585 5675 42619
rect 6193 42585 6227 42619
rect 6745 42585 6779 42619
rect 7297 42585 7331 42619
rect 7849 42585 7883 42619
rect 8401 42585 8435 42619
rect 9413 42585 9447 42619
rect 15117 42585 15151 42619
rect 16865 42585 16899 42619
rect 17141 42585 17175 42619
rect 17693 42585 17727 42619
rect 18245 42585 18279 42619
rect 19349 42585 19383 42619
rect 19901 42585 19935 42619
rect 20453 42585 20487 42619
rect 21005 42585 21039 42619
rect 1777 42517 1811 42551
rect 8953 42517 8987 42551
rect 10057 42517 10091 42551
rect 10333 42517 10367 42551
rect 10609 42517 10643 42551
rect 10885 42517 10919 42551
rect 11161 42517 11195 42551
rect 12081 42517 12115 42551
rect 12357 42517 12391 42551
rect 12817 42517 12851 42551
rect 12909 42517 12943 42551
rect 13369 42517 13403 42551
rect 13737 42517 13771 42551
rect 14289 42517 14323 42551
rect 14473 42517 14507 42551
rect 14749 42517 14783 42551
rect 18705 42517 18739 42551
rect 19993 42517 20027 42551
rect 2513 42313 2547 42347
rect 2789 42313 2823 42347
rect 3065 42313 3099 42347
rect 3525 42313 3559 42347
rect 4169 42313 4203 42347
rect 4537 42313 4571 42347
rect 5089 42313 5123 42347
rect 5641 42313 5675 42347
rect 6009 42313 6043 42347
rect 6561 42313 6595 42347
rect 7481 42313 7515 42347
rect 10333 42313 10367 42347
rect 10609 42313 10643 42347
rect 17969 42313 18003 42347
rect 18337 42313 18371 42347
rect 18981 42313 19015 42347
rect 19625 42313 19659 42347
rect 20177 42313 20211 42347
rect 14197 42245 14231 42279
rect 15117 42245 15151 42279
rect 20821 42245 20855 42279
rect 21373 42245 21407 42279
rect 2697 42177 2731 42211
rect 2973 42177 3007 42211
rect 3249 42177 3283 42211
rect 3341 42177 3375 42211
rect 3893 42177 3927 42211
rect 4445 42177 4479 42211
rect 4905 42177 4939 42211
rect 5549 42177 5583 42211
rect 6193 42177 6227 42211
rect 6377 42177 6411 42211
rect 6929 42177 6963 42211
rect 7389 42177 7423 42211
rect 8309 42177 8343 42211
rect 9137 42177 9171 42211
rect 9413 42177 9447 42211
rect 9689 42177 9723 42211
rect 10517 42177 10551 42211
rect 10793 42177 10827 42211
rect 13553 42177 13587 42211
rect 14657 42177 14691 42211
rect 15393 42177 15427 42211
rect 15761 42177 15795 42211
rect 16221 42177 16255 42211
rect 16773 42177 16807 42211
rect 17233 42177 17267 42211
rect 17509 42177 17543 42211
rect 17785 42177 17819 42211
rect 18245 42177 18279 42211
rect 18889 42177 18923 42211
rect 19165 42177 19199 42211
rect 19533 42177 19567 42211
rect 19993 42177 20027 42211
rect 20453 42177 20487 42211
rect 21005 42177 21039 42211
rect 7113 42041 7147 42075
rect 8953 42041 8987 42075
rect 18705 42041 18739 42075
rect 8585 41973 8619 42007
rect 9229 41973 9263 42007
rect 9505 41973 9539 42007
rect 9965 41973 9999 42007
rect 13737 41973 13771 42007
rect 14289 41973 14323 42007
rect 14841 41973 14875 42007
rect 15209 41973 15243 42007
rect 15577 41973 15611 42007
rect 15945 41973 15979 42007
rect 16313 41973 16347 42007
rect 16865 41973 16899 42007
rect 17049 41973 17083 42007
rect 17325 41973 17359 42007
rect 3157 41769 3191 41803
rect 3801 41769 3835 41803
rect 4353 41769 4387 41803
rect 4629 41769 4663 41803
rect 4905 41769 4939 41803
rect 5457 41769 5491 41803
rect 5733 41769 5767 41803
rect 6009 41769 6043 41803
rect 6469 41769 6503 41803
rect 7757 41769 7791 41803
rect 8585 41769 8619 41803
rect 14197 41769 14231 41803
rect 15945 41769 15979 41803
rect 16221 41769 16255 41803
rect 18705 41769 18739 41803
rect 20545 41769 20579 41803
rect 20913 41769 20947 41803
rect 3433 41701 3467 41735
rect 4077 41701 4111 41735
rect 5181 41701 5215 41735
rect 6837 41701 6871 41735
rect 7205 41701 7239 41735
rect 8953 41701 8987 41735
rect 17049 41701 17083 41735
rect 17601 41701 17635 41735
rect 17877 41701 17911 41735
rect 20085 41701 20119 41735
rect 15117 41633 15151 41667
rect 1409 41565 1443 41599
rect 1961 41565 1995 41599
rect 3341 41565 3375 41599
rect 3617 41565 3651 41599
rect 3985 41565 4019 41599
rect 4261 41565 4295 41599
rect 4537 41565 4571 41599
rect 4813 41565 4847 41599
rect 5089 41565 5123 41599
rect 5365 41565 5399 41599
rect 5641 41565 5675 41599
rect 5917 41565 5951 41599
rect 6193 41565 6227 41599
rect 7021 41565 7055 41599
rect 7389 41565 7423 41599
rect 7665 41565 7699 41599
rect 7941 41565 7975 41599
rect 8769 41565 8803 41599
rect 9137 41565 9171 41599
rect 9421 41565 9455 41599
rect 9689 41565 9723 41599
rect 9965 41565 9999 41599
rect 14381 41565 14415 41599
rect 14565 41565 14599 41599
rect 15301 41565 15335 41599
rect 15669 41565 15703 41599
rect 16137 41561 16171 41595
rect 16405 41565 16439 41599
rect 16681 41565 16715 41599
rect 16957 41565 16991 41599
rect 17233 41565 17267 41599
rect 17509 41565 17543 41599
rect 17785 41565 17819 41599
rect 18061 41581 18095 41615
rect 18337 41565 18371 41599
rect 18613 41565 18647 41599
rect 18889 41565 18923 41599
rect 19441 41565 19475 41599
rect 20269 41565 20303 41599
rect 20361 41565 20395 41599
rect 20729 41565 20763 41599
rect 1685 41497 1719 41531
rect 2237 41497 2271 41531
rect 8125 41497 8159 41531
rect 14933 41497 14967 41531
rect 21189 41497 21223 41531
rect 21557 41497 21591 41531
rect 7481 41429 7515 41463
rect 8401 41429 8435 41463
rect 9229 41429 9263 41463
rect 9505 41429 9539 41463
rect 9781 41429 9815 41463
rect 14657 41429 14691 41463
rect 15393 41429 15427 41463
rect 15761 41429 15795 41463
rect 16497 41429 16531 41463
rect 16773 41429 16807 41463
rect 17325 41429 17359 41463
rect 18153 41429 18187 41463
rect 18429 41429 18463 41463
rect 19257 41429 19291 41463
rect 19809 41429 19843 41463
rect 3985 41225 4019 41259
rect 5181 41225 5215 41259
rect 5457 41225 5491 41259
rect 5733 41225 5767 41259
rect 6009 41225 6043 41259
rect 8125 41225 8159 41259
rect 8401 41225 8435 41259
rect 14657 41225 14691 41259
rect 14933 41225 14967 41259
rect 15209 41225 15243 41259
rect 15945 41225 15979 41259
rect 17417 41225 17451 41259
rect 17693 41225 17727 41259
rect 18245 41225 18279 41259
rect 19441 41225 19475 41259
rect 20269 41225 20303 41259
rect 20821 41225 20855 41259
rect 2237 41157 2271 41191
rect 1409 41089 1443 41123
rect 1961 41089 1995 41123
rect 2513 41089 2547 41123
rect 4169 41089 4203 41123
rect 4905 41089 4939 41123
rect 5365 41089 5399 41123
rect 5641 41089 5675 41123
rect 5917 41089 5951 41123
rect 6193 41089 6227 41123
rect 6561 41089 6595 41123
rect 6929 41089 6963 41123
rect 7205 41089 7239 41123
rect 7481 41089 7515 41123
rect 8309 41089 8343 41123
rect 8585 41089 8619 41123
rect 14841 41089 14875 41123
rect 15117 41089 15151 41123
rect 15393 41089 15427 41123
rect 15669 41089 15703 41123
rect 16129 41089 16163 41123
rect 16497 41089 16531 41123
rect 16865 41089 16899 41123
rect 17141 41089 17175 41123
rect 17233 41089 17267 41123
rect 17877 41089 17911 41123
rect 18153 41113 18187 41147
rect 18429 41089 18463 41123
rect 18797 41089 18831 41123
rect 19073 41089 19107 41123
rect 19349 41073 19383 41107
rect 19625 41089 19659 41123
rect 19901 41089 19935 41123
rect 20177 41089 20211 41123
rect 20453 41089 20487 41123
rect 20729 41089 20763 41123
rect 21005 41089 21039 41123
rect 21281 41089 21315 41123
rect 1593 41021 1627 41055
rect 2697 41021 2731 41055
rect 6377 40953 6411 40987
rect 7021 40953 7055 40987
rect 7297 40953 7331 40987
rect 15485 40953 15519 40987
rect 16681 40953 16715 40987
rect 19165 40953 19199 40987
rect 20545 40953 20579 40987
rect 7757 40885 7791 40919
rect 16313 40885 16347 40919
rect 16957 40885 16991 40919
rect 17969 40885 18003 40919
rect 18613 40885 18647 40919
rect 18889 40885 18923 40919
rect 19717 40885 19751 40919
rect 19993 40885 20027 40919
rect 21465 40885 21499 40919
rect 5457 40681 5491 40715
rect 7113 40681 7147 40715
rect 19073 40681 19107 40715
rect 19717 40681 19751 40715
rect 20821 40681 20855 40715
rect 17509 40613 17543 40647
rect 17785 40613 17819 40647
rect 18337 40613 18371 40647
rect 19993 40613 20027 40647
rect 1409 40477 1443 40511
rect 1961 40477 1995 40511
rect 2513 40477 2547 40511
rect 5641 40477 5675 40511
rect 6837 40477 6871 40511
rect 7297 40477 7331 40511
rect 17417 40477 17451 40511
rect 17693 40477 17727 40511
rect 17969 40477 18003 40511
rect 18245 40477 18279 40511
rect 18521 40477 18555 40511
rect 18797 40477 18831 40511
rect 18889 40477 18923 40511
rect 19625 40477 19659 40511
rect 19901 40477 19935 40511
rect 20177 40477 20211 40511
rect 20453 40477 20487 40511
rect 20729 40477 20763 40511
rect 21005 40477 21039 40511
rect 21281 40477 21315 40511
rect 1685 40409 1719 40443
rect 2237 40409 2271 40443
rect 2789 40409 2823 40443
rect 17233 40341 17267 40375
rect 18061 40341 18095 40375
rect 18613 40341 18647 40375
rect 19441 40341 19475 40375
rect 20269 40341 20303 40375
rect 20545 40341 20579 40375
rect 21465 40341 21499 40375
rect 16129 40137 16163 40171
rect 17509 40137 17543 40171
rect 17785 40137 17819 40171
rect 18061 40137 18095 40171
rect 18337 40137 18371 40171
rect 18613 40137 18647 40171
rect 19165 40137 19199 40171
rect 19441 40137 19475 40171
rect 20545 40137 20579 40171
rect 20821 40137 20855 40171
rect 2053 40069 2087 40103
rect 21189 40069 21223 40103
rect 1777 40001 1811 40035
rect 2329 40001 2363 40035
rect 3065 40001 3099 40035
rect 16313 40001 16347 40035
rect 17693 40001 17727 40035
rect 17969 40001 18003 40035
rect 18245 40001 18279 40035
rect 18521 40001 18555 40035
rect 18797 40001 18831 40035
rect 19073 40001 19107 40035
rect 19349 40001 19383 40035
rect 19625 40001 19659 40035
rect 19993 40001 20027 40035
rect 20453 40001 20487 40035
rect 20729 40001 20763 40035
rect 21005 40001 21039 40035
rect 2605 39933 2639 39967
rect 3341 39933 3375 39967
rect 18889 39865 18923 39899
rect 20269 39865 20303 39899
rect 19809 39797 19843 39831
rect 21465 39797 21499 39831
rect 6193 39593 6227 39627
rect 15945 39593 15979 39627
rect 17417 39593 17451 39627
rect 18061 39593 18095 39627
rect 18889 39593 18923 39627
rect 19809 39593 19843 39627
rect 19533 39525 19567 39559
rect 20085 39525 20119 39559
rect 4077 39457 4111 39491
rect 1501 39389 1535 39423
rect 1775 39389 1809 39423
rect 2881 39389 2915 39423
rect 3801 39389 3835 39423
rect 6377 39389 6411 39423
rect 16129 39389 16163 39423
rect 17601 39389 17635 39423
rect 17877 39389 17911 39423
rect 18245 39389 18279 39423
rect 19073 39389 19107 39423
rect 19441 39389 19475 39423
rect 19717 39389 19751 39423
rect 19993 39389 20027 39423
rect 20269 39389 20303 39423
rect 20545 39389 20579 39423
rect 21005 39389 21039 39423
rect 21281 39389 21315 39423
rect 3157 39321 3191 39355
rect 2513 39253 2547 39287
rect 17693 39253 17727 39287
rect 19257 39253 19291 39287
rect 20361 39253 20395 39287
rect 20821 39253 20855 39287
rect 21465 39253 21499 39287
rect 6009 39049 6043 39083
rect 15669 39049 15703 39083
rect 18797 39049 18831 39083
rect 19717 39049 19751 39083
rect 20085 39049 20119 39083
rect 20545 39049 20579 39083
rect 1685 38981 1719 39015
rect 21189 38981 21223 39015
rect 1409 38913 1443 38947
rect 2235 38913 2269 38947
rect 4059 38913 4093 38947
rect 6193 38913 6227 38947
rect 6377 38913 6411 38947
rect 6651 38913 6685 38947
rect 15853 38913 15887 38947
rect 18981 38913 19015 38947
rect 19901 38913 19935 38947
rect 20269 38913 20303 38947
rect 20729 38913 20763 38947
rect 21005 38913 21039 38947
rect 1961 38845 1995 38879
rect 3801 38845 3835 38879
rect 2973 38709 3007 38743
rect 4813 38709 4847 38743
rect 7389 38709 7423 38743
rect 20821 38709 20855 38743
rect 21465 38709 21499 38743
rect 16129 38505 16163 38539
rect 17325 38505 17359 38539
rect 17877 38505 17911 38539
rect 19717 38505 19751 38539
rect 19993 38437 20027 38471
rect 20269 38437 20303 38471
rect 1685 38369 1719 38403
rect 3893 38369 3927 38403
rect 5365 38369 5399 38403
rect 1959 38301 1993 38335
rect 3157 38301 3191 38335
rect 4167 38301 4201 38335
rect 5607 38301 5641 38335
rect 6745 38301 6779 38335
rect 7019 38301 7053 38335
rect 16313 38301 16347 38335
rect 17509 38301 17543 38335
rect 18061 38301 18095 38335
rect 19901 38301 19935 38335
rect 20177 38301 20211 38335
rect 20453 38301 20487 38335
rect 20729 38301 20763 38335
rect 21005 38301 21039 38335
rect 21281 38301 21315 38335
rect 3433 38233 3467 38267
rect 2697 38165 2731 38199
rect 4905 38165 4939 38199
rect 6377 38165 6411 38199
rect 7757 38165 7791 38199
rect 20545 38165 20579 38199
rect 20821 38165 20855 38199
rect 21465 38165 21499 38199
rect 3801 37961 3835 37995
rect 6009 37961 6043 37995
rect 8217 37961 8251 37995
rect 18613 37961 18647 37995
rect 19901 37961 19935 37995
rect 20545 37961 20579 37995
rect 7113 37893 7147 37927
rect 7389 37893 7423 37927
rect 7481 37893 7515 37927
rect 1409 37825 1443 37859
rect 3157 37825 3191 37859
rect 4903 37825 4937 37859
rect 6193 37825 6227 37859
rect 7849 37825 7883 37859
rect 9689 37825 9723 37859
rect 9963 37825 9997 37859
rect 13001 37825 13035 37859
rect 13275 37825 13309 37859
rect 14839 37835 14873 37869
rect 18797 37825 18831 37859
rect 20085 37825 20119 37859
rect 20453 37825 20487 37859
rect 20729 37825 20763 37859
rect 21005 37825 21039 37859
rect 21281 37825 21315 37859
rect 1685 37757 1719 37791
rect 1961 37757 1995 37791
rect 2145 37757 2179 37791
rect 2605 37757 2639 37791
rect 2881 37757 2915 37791
rect 3019 37757 3053 37791
rect 4629 37757 4663 37791
rect 14565 37757 14599 37791
rect 20269 37689 20303 37723
rect 4537 37621 4571 37655
rect 5641 37621 5675 37655
rect 6653 37621 6687 37655
rect 8401 37621 8435 37655
rect 10701 37621 10735 37655
rect 14013 37621 14047 37655
rect 15577 37621 15611 37655
rect 20821 37621 20855 37655
rect 21465 37621 21499 37655
rect 5733 37417 5767 37451
rect 11529 37417 11563 37451
rect 19717 37417 19751 37451
rect 19993 37417 20027 37451
rect 20269 37417 20303 37451
rect 20545 37417 20579 37451
rect 4445 37349 4479 37383
rect 4721 37281 4755 37315
rect 4997 37281 5031 37315
rect 5641 37281 5675 37315
rect 12357 37281 12391 37315
rect 1501 37213 1535 37247
rect 1775 37213 1809 37247
rect 3065 37213 3099 37247
rect 3801 37213 3835 37247
rect 3985 37213 4019 37247
rect 4859 37213 4893 37247
rect 5917 37213 5951 37247
rect 6469 37213 6503 37247
rect 10517 37213 10551 37247
rect 11713 37213 11747 37247
rect 12615 37183 12649 37217
rect 14289 37213 14323 37247
rect 15761 37213 15795 37247
rect 16037 37213 16071 37247
rect 16221 37213 16255 37247
rect 16497 37213 16531 37247
rect 17233 37213 17267 37247
rect 17877 37213 17911 37247
rect 17969 37213 18003 37247
rect 18153 37213 18187 37247
rect 18981 37213 19015 37247
rect 19901 37213 19935 37247
rect 20177 37213 20211 37247
rect 20453 37213 20487 37247
rect 20729 37213 20763 37247
rect 21005 37213 21039 37247
rect 21189 37213 21223 37247
rect 3341 37145 3375 37179
rect 6561 37145 6595 37179
rect 6929 37145 6963 37179
rect 10609 37145 10643 37179
rect 10977 37145 11011 37179
rect 14534 37145 14568 37179
rect 21557 37145 21591 37179
rect 2513 37077 2547 37111
rect 6193 37077 6227 37111
rect 7297 37077 7331 37111
rect 7481 37077 7515 37111
rect 9781 37077 9815 37111
rect 10241 37077 10275 37111
rect 11345 37077 11379 37111
rect 11897 37077 11931 37111
rect 13369 37077 13403 37111
rect 15669 37077 15703 37111
rect 15853 37077 15887 37111
rect 16129 37077 16163 37111
rect 16313 37077 16347 37111
rect 17325 37077 17359 37111
rect 17693 37077 17727 37111
rect 18153 37077 18187 37111
rect 18797 37077 18831 37111
rect 20821 37077 20855 37111
rect 6009 36873 6043 36907
rect 8309 36873 8343 36907
rect 11069 36873 11103 36907
rect 14841 36873 14875 36907
rect 16221 36873 16255 36907
rect 18061 36873 18095 36907
rect 19901 36873 19935 36907
rect 20913 36873 20947 36907
rect 11621 36805 11655 36839
rect 16037 36805 16071 36839
rect 18705 36805 18739 36839
rect 2939 36737 2973 36771
rect 4351 36737 4385 36771
rect 5733 36737 5767 36771
rect 6193 36737 6227 36771
rect 6377 36737 6411 36771
rect 7539 36737 7573 36771
rect 8677 36737 8711 36771
rect 8951 36737 8985 36771
rect 10057 36737 10091 36771
rect 10331 36737 10365 36771
rect 13967 36737 14001 36771
rect 15025 36737 15059 36771
rect 15669 36737 15703 36771
rect 15945 36737 15979 36771
rect 16405 36737 16439 36771
rect 16937 36737 16971 36771
rect 18337 36737 18371 36771
rect 19625 36737 19659 36771
rect 20085 36737 20119 36771
rect 20361 36737 20395 36771
rect 20545 36737 20579 36771
rect 20821 36737 20855 36771
rect 21097 36737 21131 36771
rect 21281 36737 21315 36771
rect 2697 36669 2731 36703
rect 4077 36669 4111 36703
rect 6561 36669 6595 36703
rect 7297 36669 7331 36703
rect 12909 36669 12943 36703
rect 13093 36669 13127 36703
rect 13553 36669 13587 36703
rect 13829 36669 13863 36703
rect 14105 36669 14139 36703
rect 15485 36669 15519 36703
rect 16681 36669 16715 36703
rect 18153 36669 18187 36703
rect 11805 36601 11839 36635
rect 18613 36601 18647 36635
rect 20637 36601 20671 36635
rect 3709 36533 3743 36567
rect 5089 36533 5123 36567
rect 9689 36533 9723 36567
rect 14749 36533 14783 36567
rect 20453 36533 20487 36567
rect 21465 36533 21499 36567
rect 3985 36329 4019 36363
rect 7113 36329 7147 36363
rect 14289 36329 14323 36363
rect 15945 36329 15979 36363
rect 16589 36329 16623 36363
rect 17877 36329 17911 36363
rect 19533 36329 19567 36363
rect 12265 36261 12299 36295
rect 19809 36261 19843 36295
rect 2237 36193 2271 36227
rect 8953 36193 8987 36227
rect 16865 36193 16899 36227
rect 1409 36125 1443 36159
rect 2511 36125 2545 36159
rect 4169 36125 4203 36159
rect 6101 36125 6135 36159
rect 6193 36125 6227 36159
rect 7481 36125 7515 36159
rect 7755 36125 7789 36159
rect 9195 36125 9229 36159
rect 10517 36125 10551 36159
rect 11253 36125 11287 36159
rect 11527 36125 11561 36159
rect 16129 36125 16163 36159
rect 16773 36125 16807 36159
rect 17139 36125 17173 36159
rect 19441 36125 19475 36159
rect 19717 36121 19751 36155
rect 19993 36101 20027 36135
rect 20261 36125 20295 36159
rect 20637 36125 20671 36159
rect 21005 36125 21039 36159
rect 1685 36057 1719 36091
rect 6561 36057 6595 36091
rect 21189 36057 21223 36091
rect 21557 36057 21591 36091
rect 3249 35989 3283 36023
rect 5273 35989 5307 36023
rect 5825 35989 5859 36023
rect 6929 35989 6963 36023
rect 8493 35989 8527 36023
rect 9965 35989 9999 36023
rect 10609 35989 10643 36023
rect 19257 35989 19291 36023
rect 20085 35989 20119 36023
rect 20453 35989 20487 36023
rect 20821 35989 20855 36023
rect 5917 35785 5951 35819
rect 20177 35785 20211 35819
rect 20545 35785 20579 35819
rect 18950 35717 18984 35751
rect 1685 35649 1719 35683
rect 1961 35649 1995 35683
rect 2973 35649 3007 35683
rect 3801 35649 3835 35683
rect 4261 35649 4295 35683
rect 5147 35649 5181 35683
rect 6377 35649 6411 35683
rect 6653 35649 6687 35683
rect 7295 35649 7329 35683
rect 8401 35649 8435 35683
rect 9321 35649 9355 35683
rect 12063 35679 12097 35713
rect 15485 35649 15519 35683
rect 16865 35649 16899 35683
rect 17233 35649 17267 35683
rect 18613 35649 18647 35683
rect 20361 35649 20395 35683
rect 20729 35649 20763 35683
rect 21005 35649 21039 35683
rect 21281 35649 21315 35683
rect 1777 35581 1811 35615
rect 2421 35581 2455 35615
rect 2697 35581 2731 35615
rect 2814 35581 2848 35615
rect 4537 35581 4571 35615
rect 4905 35581 4939 35615
rect 7021 35581 7055 35615
rect 8585 35581 8619 35615
rect 9045 35581 9079 35615
rect 9438 35581 9472 35615
rect 9597 35581 9631 35615
rect 11805 35581 11839 35615
rect 17049 35581 17083 35615
rect 18705 35581 18739 35615
rect 13369 35513 13403 35547
rect 18429 35513 18463 35547
rect 20085 35513 20119 35547
rect 3617 35445 3651 35479
rect 4077 35445 4111 35479
rect 8033 35445 8067 35479
rect 10241 35445 10275 35479
rect 12817 35445 12851 35479
rect 15301 35445 15335 35479
rect 17141 35445 17175 35479
rect 20821 35445 20855 35479
rect 21465 35445 21499 35479
rect 7297 35241 7331 35275
rect 17325 35241 17359 35275
rect 17785 35241 17819 35275
rect 20269 35241 20303 35275
rect 12265 35173 12299 35207
rect 4905 35105 4939 35139
rect 6285 35105 6319 35139
rect 12541 35105 12575 35139
rect 12817 35105 12851 35139
rect 14841 35105 14875 35139
rect 16313 35105 16347 35139
rect 19257 35105 19291 35139
rect 20637 35105 20671 35139
rect 1409 35037 1443 35071
rect 2513 35037 2547 35071
rect 2605 35037 2639 35071
rect 4261 35037 4295 35071
rect 5147 35037 5181 35071
rect 6543 35037 6577 35071
rect 9413 35037 9447 35071
rect 9505 35037 9539 35071
rect 11069 35037 11103 35071
rect 11621 35037 11655 35071
rect 11805 35037 11839 35071
rect 12658 35037 12692 35071
rect 16587 35037 16621 35071
rect 17693 35037 17727 35071
rect 17877 35037 17911 35071
rect 18889 35037 18923 35071
rect 19499 35037 19533 35071
rect 20821 35037 20855 35071
rect 21189 35037 21223 35071
rect 21281 35037 21315 35071
rect 1685 34969 1719 35003
rect 2973 34969 3007 35003
rect 3893 34969 3927 35003
rect 4445 34969 4479 35003
rect 9137 34969 9171 35003
rect 9873 34969 9907 35003
rect 10241 34969 10275 35003
rect 10793 34969 10827 35003
rect 11253 34969 11287 35003
rect 13461 34969 13495 35003
rect 15086 34969 15120 35003
rect 18981 34969 19015 35003
rect 21097 34969 21131 35003
rect 2237 34901 2271 34935
rect 3341 34901 3375 34935
rect 3525 34901 3559 34935
rect 4537 34901 4571 34935
rect 5917 34901 5951 34935
rect 10425 34901 10459 34935
rect 16221 34901 16255 34935
rect 21465 34901 21499 34935
rect 6377 34697 6411 34731
rect 9229 34697 9263 34731
rect 10885 34697 10919 34731
rect 16037 34697 16071 34731
rect 16313 34697 16347 34731
rect 16773 34697 16807 34731
rect 18889 34697 18923 34731
rect 19717 34697 19751 34731
rect 19993 34697 20027 34731
rect 20269 34697 20303 34731
rect 20545 34697 20579 34731
rect 4813 34629 4847 34663
rect 5089 34629 5123 34663
rect 5181 34629 5215 34663
rect 5917 34629 5951 34663
rect 9505 34629 9539 34663
rect 10333 34629 10367 34663
rect 10793 34629 10827 34663
rect 21189 34629 21223 34663
rect 1869 34561 1903 34595
rect 2143 34561 2177 34595
rect 3523 34561 3557 34595
rect 5549 34561 5583 34595
rect 6561 34561 6595 34595
rect 7665 34561 7699 34595
rect 7939 34561 7973 34595
rect 9597 34561 9631 34595
rect 9965 34561 9999 34595
rect 13001 34561 13035 34595
rect 13243 34561 13277 34595
rect 14381 34561 14415 34595
rect 14639 34591 14673 34625
rect 15945 34561 15979 34595
rect 16497 34561 16531 34595
rect 16957 34561 16991 34595
rect 17233 34561 17267 34595
rect 17491 34591 17525 34625
rect 19073 34561 19107 34595
rect 19625 34561 19659 34595
rect 19901 34561 19935 34595
rect 20177 34561 20211 34595
rect 20453 34561 20487 34595
rect 20729 34561 20763 34595
rect 21005 34561 21039 34595
rect 3249 34493 3283 34527
rect 6101 34425 6135 34459
rect 8677 34425 8711 34459
rect 10517 34425 10551 34459
rect 19441 34425 19475 34459
rect 2881 34357 2915 34391
rect 4261 34357 4295 34391
rect 14013 34357 14047 34391
rect 15393 34357 15427 34391
rect 18245 34357 18279 34391
rect 20821 34357 20855 34391
rect 21465 34357 21499 34391
rect 7941 34153 7975 34187
rect 10333 34153 10367 34187
rect 18061 34153 18095 34187
rect 19257 34153 19291 34187
rect 17969 34085 18003 34119
rect 18889 34085 18923 34119
rect 19993 34085 20027 34119
rect 6377 34017 6411 34051
rect 8033 34017 8067 34051
rect 9321 34017 9355 34051
rect 10701 34017 10735 34051
rect 16313 34017 16347 34051
rect 18153 34017 18187 34051
rect 1593 33949 1627 33983
rect 1851 33919 1885 33953
rect 2973 33949 3007 33983
rect 3249 33949 3283 33983
rect 3801 33949 3835 33983
rect 5181 33949 5215 33983
rect 5273 33949 5307 33983
rect 5641 33949 5675 33983
rect 6651 33949 6685 33983
rect 7757 33949 7791 33983
rect 7849 33949 7883 33983
rect 9563 33949 9597 33983
rect 10975 33949 11009 33983
rect 14933 33949 14967 33983
rect 15207 33949 15241 33983
rect 17877 33949 17911 33983
rect 18245 33949 18279 33983
rect 18705 33949 18739 33983
rect 18797 33949 18831 33983
rect 18981 33949 19015 33983
rect 19441 33949 19475 33983
rect 19901 33949 19935 33983
rect 20177 33949 20211 33983
rect 20361 33949 20395 33983
rect 20637 33949 20671 33983
rect 20821 33949 20855 33983
rect 21189 33949 21223 33983
rect 21281 33949 21315 33983
rect 4077 33881 4111 33915
rect 4905 33881 4939 33915
rect 16580 33881 16614 33915
rect 18337 33881 18371 33915
rect 2605 33813 2639 33847
rect 6009 33813 6043 33847
rect 6193 33813 6227 33847
rect 7389 33813 7423 33847
rect 11713 33813 11747 33847
rect 15945 33813 15979 33847
rect 17693 33813 17727 33847
rect 18521 33813 18555 33847
rect 19717 33813 19751 33847
rect 20453 33813 20487 33847
rect 20821 33813 20855 33847
rect 21005 33813 21039 33847
rect 21465 33813 21499 33847
rect 4169 33609 4203 33643
rect 16681 33609 16715 33643
rect 17049 33609 17083 33643
rect 19165 33609 19199 33643
rect 19993 33609 20027 33643
rect 2881 33541 2915 33575
rect 3157 33541 3191 33575
rect 3985 33541 4019 33575
rect 10701 33541 10735 33575
rect 11253 33541 11287 33575
rect 13185 33541 13219 33575
rect 13461 33541 13495 33575
rect 13553 33541 13587 33575
rect 13921 33541 13955 33575
rect 14289 33541 14323 33575
rect 20453 33541 20487 33575
rect 21005 33541 21039 33575
rect 1409 33473 1443 33507
rect 1961 33473 1995 33507
rect 3249 33473 3283 33507
rect 3617 33473 3651 33507
rect 4903 33473 4937 33507
rect 7479 33473 7513 33507
rect 9319 33473 9353 33507
rect 11771 33473 11805 33507
rect 14657 33473 14691 33507
rect 14931 33473 14965 33507
rect 16865 33473 16899 33507
rect 17233 33473 17267 33507
rect 17325 33473 17359 33507
rect 19349 33473 19383 33507
rect 19901 33473 19935 33507
rect 20177 33473 20211 33507
rect 1685 33405 1719 33439
rect 2237 33405 2271 33439
rect 4629 33405 4663 33439
rect 7205 33405 7239 33439
rect 9045 33405 9079 33439
rect 11529 33405 11563 33439
rect 19717 33337 19751 33371
rect 5641 33269 5675 33303
rect 8217 33269 8251 33303
rect 10057 33269 10091 33303
rect 10793 33269 10827 33303
rect 12541 33269 12575 33303
rect 14473 33269 14507 33303
rect 15669 33269 15703 33303
rect 17417 33269 17451 33303
rect 20729 33269 20763 33303
rect 21281 33269 21315 33303
rect 3341 33065 3375 33099
rect 7021 33065 7055 33099
rect 7297 33065 7331 33099
rect 12357 33065 12391 33099
rect 18061 33065 18095 33099
rect 18889 33065 18923 33099
rect 6745 32997 6779 33031
rect 15209 32997 15243 33031
rect 17877 32997 17911 33031
rect 18705 32997 18739 33031
rect 21097 32997 21131 33031
rect 2329 32929 2363 32963
rect 3801 32929 3835 32963
rect 7481 32929 7515 32963
rect 9045 32929 9079 32963
rect 12633 32929 12667 32963
rect 15602 32929 15636 32963
rect 15761 32929 15795 32963
rect 16497 32929 16531 32963
rect 18245 32929 18279 32963
rect 21005 32929 21039 32963
rect 2603 32861 2637 32895
rect 4059 32831 4093 32865
rect 5825 32861 5859 32895
rect 6929 32861 6963 32895
rect 7205 32861 7239 32895
rect 7389 32861 7423 32895
rect 7723 32861 7757 32895
rect 9303 32831 9337 32865
rect 10885 32861 10919 32895
rect 11727 32861 11761 32895
rect 12891 32831 12925 32865
rect 14565 32861 14599 32895
rect 14749 32861 14783 32895
rect 15485 32861 15519 32895
rect 16405 32861 16439 32895
rect 17969 32861 18003 32895
rect 18521 32861 18555 32895
rect 18613 32861 18647 32895
rect 18797 32861 18831 32895
rect 19073 32861 19107 32895
rect 19257 32861 19291 32895
rect 20729 32861 20763 32895
rect 20821 32861 20855 32895
rect 21281 32861 21315 32895
rect 21557 32861 21591 32895
rect 1501 32793 1535 32827
rect 1685 32793 1719 32827
rect 5733 32793 5767 32827
rect 6193 32793 6227 32827
rect 10977 32793 11011 32827
rect 11345 32793 11379 32827
rect 16764 32793 16798 32827
rect 19524 32793 19558 32827
rect 4813 32725 4847 32759
rect 5457 32725 5491 32759
rect 6561 32725 6595 32759
rect 8493 32725 8527 32759
rect 10057 32725 10091 32759
rect 10609 32725 10643 32759
rect 11897 32725 11931 32759
rect 13645 32725 13679 32759
rect 18245 32725 18279 32759
rect 18337 32725 18371 32759
rect 20637 32725 20671 32759
rect 21005 32725 21039 32759
rect 21373 32725 21407 32759
rect 6377 32521 6411 32555
rect 7021 32521 7055 32555
rect 11253 32521 11287 32555
rect 17877 32521 17911 32555
rect 18981 32521 19015 32555
rect 20637 32521 20671 32555
rect 3249 32453 3283 32487
rect 9137 32453 9171 32487
rect 9413 32453 9447 32487
rect 9505 32453 9539 32487
rect 10241 32453 10275 32487
rect 1835 32385 1869 32419
rect 2973 32385 3007 32419
rect 3709 32385 3743 32419
rect 5549 32385 5583 32419
rect 6561 32385 6595 32419
rect 7205 32385 7239 32419
rect 7297 32385 7331 32419
rect 7571 32385 7605 32419
rect 9873 32385 9907 32419
rect 11069 32385 11103 32419
rect 12633 32385 12667 32419
rect 12907 32385 12941 32419
rect 14255 32385 14289 32419
rect 15669 32385 15703 32419
rect 17139 32385 17173 32419
rect 19165 32385 19199 32419
rect 19441 32385 19475 32419
rect 19625 32385 19659 32419
rect 19899 32385 19933 32419
rect 21189 32385 21223 32419
rect 21281 32385 21315 32419
rect 1593 32317 1627 32351
rect 3893 32317 3927 32351
rect 4629 32317 4663 32351
rect 4767 32317 4801 32351
rect 4905 32317 4939 32351
rect 14013 32317 14047 32351
rect 16865 32317 16899 32351
rect 4353 32249 4387 32283
rect 10425 32249 10459 32283
rect 2605 32181 2639 32215
rect 8309 32181 8343 32215
rect 10977 32181 11011 32215
rect 13645 32181 13679 32215
rect 15025 32181 15059 32215
rect 19257 32181 19291 32215
rect 21005 32181 21039 32215
rect 21465 32181 21499 32215
rect 6837 31977 6871 32011
rect 17049 31977 17083 32011
rect 19257 31977 19291 32011
rect 19993 31977 20027 32011
rect 20269 31977 20303 32011
rect 10425 31909 10459 31943
rect 13829 31909 13863 31943
rect 14749 31909 14783 31943
rect 18153 31909 18187 31943
rect 18705 31909 18739 31943
rect 19625 31909 19659 31943
rect 1961 31841 1995 31875
rect 2421 31841 2455 31875
rect 2814 31841 2848 31875
rect 3617 31841 3651 31875
rect 4997 31841 5031 31875
rect 5641 31841 5675 31875
rect 5917 31841 5951 31875
rect 6034 31841 6068 31875
rect 7481 31841 7515 31875
rect 9781 31841 9815 31875
rect 10701 31841 10735 31875
rect 10839 31841 10873 31875
rect 14289 31841 14323 31875
rect 15025 31841 15059 31875
rect 15301 31841 15335 31875
rect 16037 31841 16071 31875
rect 20729 31841 20763 31875
rect 1409 31773 1443 31807
rect 1777 31773 1811 31807
rect 2697 31773 2731 31807
rect 2973 31773 3007 31807
rect 3801 31773 3835 31807
rect 4077 31773 4111 31807
rect 4721 31773 4755 31807
rect 5181 31773 5215 31807
rect 6193 31773 6227 31807
rect 7755 31773 7789 31807
rect 9965 31773 9999 31807
rect 10977 31773 11011 31807
rect 11621 31773 11655 31807
rect 12817 31773 12851 31807
rect 12909 31773 12943 31807
rect 14105 31773 14139 31807
rect 15142 31773 15176 31807
rect 15945 31773 15979 31807
rect 16311 31773 16345 31807
rect 18337 31773 18371 31807
rect 18429 31773 18463 31807
rect 18613 31773 18647 31807
rect 18889 31773 18923 31807
rect 19441 31773 19475 31807
rect 19809 31773 19843 31807
rect 20177 31773 20211 31807
rect 20453 31773 20487 31807
rect 20637 31773 20671 31807
rect 21189 31773 21223 31807
rect 13277 31705 13311 31739
rect 13645 31705 13679 31739
rect 1593 31637 1627 31671
rect 4537 31637 4571 31671
rect 8493 31637 8527 31671
rect 12541 31637 12575 31671
rect 18521 31637 18555 31671
rect 21465 31637 21499 31671
rect 2421 31433 2455 31467
rect 10793 31433 10827 31467
rect 18061 31433 18095 31467
rect 19625 31433 19659 31467
rect 19901 31433 19935 31467
rect 9137 31365 9171 31399
rect 1409 31297 1443 31331
rect 1683 31297 1717 31331
rect 3123 31297 3157 31331
rect 4261 31297 4295 31331
rect 4905 31297 4939 31331
rect 5179 31297 5213 31331
rect 6377 31297 6411 31331
rect 7481 31297 7515 31331
rect 8493 31297 8527 31331
rect 9781 31297 9815 31331
rect 10055 31297 10089 31331
rect 11787 31327 11821 31361
rect 12909 31297 12943 31331
rect 13093 31297 13127 31331
rect 14715 31297 14749 31331
rect 16681 31297 16715 31331
rect 16937 31297 16971 31331
rect 18153 31297 18187 31331
rect 18427 31297 18461 31331
rect 19809 31297 19843 31331
rect 20085 31297 20119 31331
rect 20545 31297 20579 31331
rect 21005 31297 21039 31331
rect 21281 31297 21315 31331
rect 2881 31229 2915 31263
rect 4445 31229 4479 31263
rect 7297 31229 7331 31263
rect 7941 31229 7975 31263
rect 8217 31229 8251 31263
rect 8355 31229 8389 31263
rect 11529 31229 11563 31263
rect 14473 31229 14507 31263
rect 20361 31161 20395 31195
rect 3893 31093 3927 31127
rect 5917 31093 5951 31127
rect 6561 31093 6595 31127
rect 12541 31093 12575 31127
rect 13001 31093 13035 31127
rect 15485 31093 15519 31127
rect 19165 31093 19199 31127
rect 20821 31093 20855 31127
rect 21465 31093 21499 31127
rect 8493 30889 8527 30923
rect 11897 30889 11931 30923
rect 20637 30889 20671 30923
rect 4445 30821 4479 30855
rect 12449 30821 12483 30855
rect 12725 30821 12759 30855
rect 17049 30821 17083 30855
rect 17417 30821 17451 30855
rect 1409 30753 1443 30787
rect 3985 30753 4019 30787
rect 4838 30753 4872 30787
rect 11989 30753 12023 30787
rect 14105 30753 14139 30787
rect 17877 30753 17911 30787
rect 18245 30753 18279 30787
rect 18429 30753 18463 30787
rect 1651 30685 1685 30719
rect 2789 30685 2823 30719
rect 3065 30685 3099 30719
rect 3801 30685 3835 30719
rect 4721 30685 4755 30719
rect 4997 30685 5031 30719
rect 11713 30685 11747 30719
rect 11805 30685 11839 30719
rect 12173 30685 12207 30719
rect 12633 30685 12667 30719
rect 12909 30685 12943 30719
rect 14347 30685 14381 30719
rect 15669 30685 15703 30719
rect 17325 30685 17359 30719
rect 17601 30685 17635 30719
rect 17785 30685 17819 30719
rect 18153 30685 18187 30719
rect 18705 30685 18739 30719
rect 19257 30685 19291 30719
rect 21005 30685 21039 30719
rect 21189 30685 21223 30719
rect 5641 30617 5675 30651
rect 6101 30617 6135 30651
rect 6377 30617 6411 30651
rect 6469 30617 6503 30651
rect 6837 30617 6871 30651
rect 12265 30617 12299 30651
rect 15936 30617 15970 30651
rect 19524 30617 19558 30651
rect 21557 30617 21591 30651
rect 2421 30549 2455 30583
rect 7205 30549 7239 30583
rect 7389 30549 7423 30583
rect 15117 30549 15151 30583
rect 17141 30549 17175 30583
rect 18429 30549 18463 30583
rect 18521 30549 18555 30583
rect 20821 30549 20855 30583
rect 3249 30345 3283 30379
rect 4353 30345 4387 30379
rect 7389 30345 7423 30379
rect 13369 30345 13403 30379
rect 19257 30345 19291 30379
rect 21189 30277 21223 30311
rect 1409 30209 1443 30243
rect 1685 30209 1719 30243
rect 1943 30239 1977 30273
rect 3065 30209 3099 30243
rect 3615 30209 3649 30243
rect 5179 30209 5213 30243
rect 6635 30209 6669 30243
rect 8585 30209 8619 30243
rect 8827 30219 8861 30253
rect 12449 30209 12483 30243
rect 13461 30209 13495 30243
rect 13735 30209 13769 30243
rect 15115 30209 15149 30243
rect 16313 30209 16347 30243
rect 16497 30209 16531 30243
rect 16681 30209 16715 30243
rect 16955 30209 16989 30243
rect 18981 30209 19015 30243
rect 19165 30209 19199 30243
rect 19441 30209 19475 30243
rect 19533 30209 19567 30243
rect 19807 30209 19841 30243
rect 3341 30141 3375 30175
rect 4905 30141 4939 30175
rect 6377 30141 6411 30175
rect 11529 30141 11563 30175
rect 11713 30141 11747 30175
rect 12566 30141 12600 30175
rect 12725 30141 12759 30175
rect 14841 30141 14875 30175
rect 1593 30073 1627 30107
rect 12173 30073 12207 30107
rect 2697 30005 2731 30039
rect 5917 30005 5951 30039
rect 9597 30005 9631 30039
rect 14473 30005 14507 30039
rect 15853 30005 15887 30039
rect 16405 30005 16439 30039
rect 17693 30005 17727 30039
rect 19073 30005 19107 30039
rect 20545 30005 20579 30039
rect 21465 30005 21499 30039
rect 13001 29801 13035 29835
rect 20085 29801 20119 29835
rect 21005 29801 21039 29835
rect 10793 29733 10827 29767
rect 11785 29733 11819 29767
rect 14749 29733 14783 29767
rect 16037 29733 16071 29767
rect 16681 29733 16715 29767
rect 16957 29733 16991 29767
rect 20361 29733 20395 29767
rect 4537 29665 4571 29699
rect 11345 29665 11379 29699
rect 12081 29665 12115 29699
rect 12219 29665 12253 29699
rect 14289 29665 14323 29699
rect 15301 29665 15335 29699
rect 17141 29665 17175 29699
rect 21189 29665 21223 29699
rect 1501 29597 1535 29631
rect 2421 29597 2455 29631
rect 2789 29597 2823 29631
rect 4261 29597 4295 29631
rect 7481 29597 7515 29631
rect 7723 29597 7757 29631
rect 9781 29597 9815 29631
rect 10055 29597 10089 29631
rect 11161 29597 11195 29631
rect 12357 29597 12391 29631
rect 14105 29597 14139 29631
rect 15025 29597 15059 29631
rect 15142 29597 15176 29631
rect 15945 29597 15979 29631
rect 16221 29597 16255 29631
rect 16589 29597 16623 29631
rect 16865 29597 16899 29631
rect 17417 29597 17451 29631
rect 18153 29597 18187 29631
rect 19993 29597 20027 29631
rect 20269 29597 20303 29631
rect 20545 29597 20579 29631
rect 20821 29597 20855 29631
rect 20913 29597 20947 29631
rect 21281 29597 21315 29631
rect 1685 29529 1719 29563
rect 2053 29529 2087 29563
rect 2329 29529 2363 29563
rect 5365 29529 5399 29563
rect 5641 29529 5675 29563
rect 5733 29529 5767 29563
rect 6101 29529 6135 29563
rect 3157 29461 3191 29495
rect 3341 29461 3375 29495
rect 6469 29461 6503 29495
rect 6653 29461 6687 29495
rect 8493 29461 8527 29495
rect 17141 29461 17175 29495
rect 17233 29461 17267 29495
rect 17969 29461 18003 29495
rect 19809 29461 19843 29495
rect 20637 29461 20671 29495
rect 21189 29461 21223 29495
rect 21465 29461 21499 29495
rect 3157 29257 3191 29291
rect 5917 29257 5951 29291
rect 12541 29257 12575 29291
rect 15117 29257 15151 29291
rect 18061 29257 18095 29291
rect 19993 29257 20027 29291
rect 20453 29257 20487 29291
rect 20729 29257 20763 29291
rect 9229 29189 9263 29223
rect 9459 29189 9493 29223
rect 9781 29189 9815 29223
rect 10609 29189 10643 29223
rect 21189 29189 21223 29223
rect 1867 29121 1901 29155
rect 2973 29121 3007 29155
rect 3523 29121 3557 29155
rect 4905 29121 4939 29155
rect 5179 29121 5213 29155
rect 7389 29121 7423 29155
rect 8447 29121 8481 29155
rect 8585 29121 8619 29155
rect 9873 29121 9907 29155
rect 10241 29121 10275 29155
rect 11529 29121 11563 29155
rect 11803 29121 11837 29155
rect 14314 29121 14348 29155
rect 14473 29121 14507 29155
rect 15209 29121 15243 29155
rect 15483 29121 15517 29155
rect 16681 29121 16715 29155
rect 16948 29121 16982 29155
rect 18337 29121 18371 29155
rect 18611 29121 18645 29155
rect 20177 29121 20211 29155
rect 20637 29121 20671 29155
rect 20913 29121 20947 29155
rect 1593 29053 1627 29087
rect 3249 29053 3283 29087
rect 7573 29053 7607 29087
rect 8033 29053 8067 29087
rect 8309 29053 8343 29087
rect 13277 29053 13311 29087
rect 13461 29053 13495 29087
rect 13921 29053 13955 29087
rect 14197 29053 14231 29087
rect 4261 28985 4295 29019
rect 10793 28985 10827 29019
rect 2605 28917 2639 28951
rect 16221 28917 16255 28951
rect 19349 28917 19383 28951
rect 21465 28917 21499 28951
rect 1593 28713 1627 28747
rect 10701 28713 10735 28747
rect 17049 28713 17083 28747
rect 19073 28713 19107 28747
rect 8125 28645 8159 28679
rect 2237 28577 2271 28611
rect 3893 28577 3927 28611
rect 5273 28577 5307 28611
rect 5549 28577 5583 28611
rect 9689 28577 9723 28611
rect 14289 28577 14323 28611
rect 14749 28577 14783 28611
rect 15142 28577 15176 28611
rect 15945 28577 15979 28611
rect 17693 28577 17727 28611
rect 19533 28577 19567 28611
rect 19993 28577 20027 28611
rect 1501 28509 1535 28543
rect 1777 28509 1811 28543
rect 2479 28509 2513 28543
rect 4135 28509 4169 28543
rect 7113 28509 7147 28543
rect 7387 28509 7421 28543
rect 9931 28509 9965 28543
rect 11437 28509 11471 28543
rect 11711 28509 11745 28543
rect 14105 28509 14139 28543
rect 15025 28509 15059 28543
rect 15301 28509 15335 28543
rect 16037 28509 16071 28543
rect 16311 28509 16345 28543
rect 17417 28509 17451 28543
rect 19257 28509 19291 28543
rect 19349 28509 19383 28543
rect 19809 28509 19843 28543
rect 19901 28509 19935 28543
rect 20085 28509 20119 28543
rect 20361 28509 20395 28543
rect 20637 28509 20671 28543
rect 20913 28509 20947 28543
rect 21189 28509 21223 28543
rect 21281 28509 21315 28543
rect 17938 28441 17972 28475
rect 1961 28373 1995 28407
rect 3249 28373 3283 28407
rect 4905 28373 4939 28407
rect 12449 28373 12483 28407
rect 17509 28373 17543 28407
rect 19533 28373 19567 28407
rect 19625 28373 19659 28407
rect 20177 28373 20211 28407
rect 20453 28373 20487 28407
rect 20729 28373 20763 28407
rect 21005 28373 21039 28407
rect 21465 28373 21499 28407
rect 2329 28169 2363 28203
rect 3617 28169 3651 28203
rect 5273 28169 5307 28203
rect 10057 28169 10091 28203
rect 17049 28169 17083 28203
rect 19257 28169 19291 28203
rect 19993 28169 20027 28203
rect 20361 28169 20395 28203
rect 2697 28101 2731 28135
rect 3433 28101 3467 28135
rect 3985 28101 4019 28135
rect 4353 28101 4387 28135
rect 5089 28101 5123 28135
rect 1501 28033 1535 28067
rect 1961 28033 1995 28067
rect 2605 28033 2639 28067
rect 3065 28033 3099 28067
rect 4261 28033 4295 28067
rect 4721 28033 4755 28067
rect 7923 28063 7957 28097
rect 9287 28043 9321 28077
rect 11895 28033 11929 28067
rect 14287 28033 14321 28067
rect 16405 28033 16439 28067
rect 16865 28033 16899 28067
rect 17383 28033 17417 28067
rect 18521 28033 18555 28067
rect 18613 28033 18647 28067
rect 18889 28033 18923 28067
rect 19073 28033 19107 28067
rect 19165 28033 19199 28067
rect 19625 28033 19659 28067
rect 19901 28033 19935 28067
rect 20177 28033 20211 28067
rect 20545 28033 20579 28067
rect 20821 28033 20855 28067
rect 20913 28033 20947 28067
rect 21281 28033 21315 28067
rect 7665 27965 7699 27999
rect 9045 27965 9079 27999
rect 11621 27965 11655 27999
rect 14013 27965 14047 27999
rect 17141 27965 17175 27999
rect 18797 27965 18831 27999
rect 18981 27965 19015 27999
rect 1685 27897 1719 27931
rect 18153 27897 18187 27931
rect 19441 27897 19475 27931
rect 1777 27829 1811 27863
rect 8677 27829 8711 27863
rect 12633 27829 12667 27863
rect 15025 27829 15059 27863
rect 16221 27829 16255 27863
rect 18705 27829 18739 27863
rect 19717 27829 19751 27863
rect 20637 27829 20671 27863
rect 21097 27829 21131 27863
rect 21465 27829 21499 27863
rect 17693 27625 17727 27659
rect 3985 27557 4019 27591
rect 8677 27557 8711 27591
rect 10977 27557 11011 27591
rect 20637 27557 20671 27591
rect 9965 27489 9999 27523
rect 14105 27489 14139 27523
rect 17601 27489 17635 27523
rect 19257 27489 19291 27523
rect 1593 27421 1627 27455
rect 1867 27421 1901 27455
rect 2973 27421 3007 27455
rect 3249 27421 3283 27455
rect 3801 27421 3835 27455
rect 4261 27421 4295 27455
rect 4503 27421 4537 27455
rect 5641 27421 5675 27455
rect 5883 27421 5917 27455
rect 10239 27421 10273 27455
rect 12657 27421 12691 27455
rect 14379 27421 14413 27455
rect 15853 27421 15887 27455
rect 17325 27421 17359 27455
rect 17417 27421 17451 27455
rect 17877 27421 17911 27455
rect 19513 27421 19547 27455
rect 21005 27421 21039 27455
rect 7665 27353 7699 27387
rect 7757 27353 7791 27387
rect 8125 27353 8159 27387
rect 11805 27353 11839 27387
rect 11897 27353 11931 27387
rect 12265 27353 12299 27387
rect 16098 27353 16132 27387
rect 21373 27353 21407 27387
rect 2605 27285 2639 27319
rect 3157 27285 3191 27319
rect 3433 27285 3467 27319
rect 5273 27285 5307 27319
rect 6653 27285 6687 27319
rect 7389 27285 7423 27319
rect 8493 27285 8527 27319
rect 11529 27285 11563 27319
rect 12817 27285 12851 27319
rect 15117 27285 15151 27319
rect 17233 27285 17267 27319
rect 17601 27285 17635 27319
rect 2789 27081 2823 27115
rect 11713 27081 11747 27115
rect 18153 27081 18187 27115
rect 19349 27081 19383 27115
rect 21373 27081 21407 27115
rect 3893 27013 3927 27047
rect 11989 27013 12023 27047
rect 12081 27013 12115 27047
rect 12449 27013 12483 27047
rect 12817 27013 12851 27047
rect 1409 26945 1443 26979
rect 2329 26945 2363 26979
rect 3065 26945 3099 26979
rect 3157 26945 3191 26979
rect 3525 26945 3559 26979
rect 4261 26945 4295 26979
rect 4905 26945 4939 26979
rect 5179 26945 5213 26979
rect 7414 26945 7448 26979
rect 7573 26945 7607 26979
rect 8583 26945 8617 26979
rect 9689 26945 9723 26979
rect 9873 26945 9907 26979
rect 10057 26945 10091 26979
rect 10299 26945 10333 26979
rect 14657 26945 14691 26979
rect 15577 26945 15611 26979
rect 15853 26945 15887 26979
rect 16129 26945 16163 26979
rect 16221 26945 16255 26979
rect 16955 26945 16989 26979
rect 18061 26945 18095 26979
rect 18245 26945 18279 26979
rect 19533 26945 19567 26979
rect 19883 26975 19917 27009
rect 21005 26945 21039 26979
rect 21557 26945 21591 26979
rect 1685 26877 1719 26911
rect 6377 26877 6411 26911
rect 6561 26877 6595 26911
rect 7021 26877 7055 26911
rect 7297 26877 7331 26911
rect 8297 26877 8331 26911
rect 13737 26877 13771 26911
rect 13921 26877 13955 26911
rect 14381 26877 14415 26911
rect 14774 26877 14808 26911
rect 14933 26877 14967 26911
rect 16681 26877 16715 26911
rect 19625 26877 19659 26911
rect 21281 26877 21315 26911
rect 2513 26809 2547 26843
rect 11069 26809 11103 26843
rect 15945 26809 15979 26843
rect 17693 26809 17727 26843
rect 20637 26809 20671 26843
rect 4077 26741 4111 26775
rect 4445 26741 4479 26775
rect 5917 26741 5951 26775
rect 8217 26741 8251 26775
rect 9321 26741 9355 26775
rect 9781 26741 9815 26775
rect 13001 26741 13035 26775
rect 15669 26741 15703 26775
rect 16313 26741 16347 26775
rect 21097 26741 21131 26775
rect 21189 26741 21223 26775
rect 2973 26537 3007 26571
rect 4813 26537 4847 26571
rect 9413 26537 9447 26571
rect 12633 26537 12667 26571
rect 15945 26537 15979 26571
rect 17509 26537 17543 26571
rect 20085 26537 20119 26571
rect 20453 26537 20487 26571
rect 20913 26537 20947 26571
rect 3249 26469 3283 26503
rect 3525 26469 3559 26503
rect 10793 26469 10827 26503
rect 14749 26469 14783 26503
rect 18337 26469 18371 26503
rect 1409 26401 1443 26435
rect 5549 26401 5583 26435
rect 6009 26401 6043 26435
rect 6402 26401 6436 26435
rect 6561 26401 6595 26435
rect 9321 26401 9355 26435
rect 15025 26401 15059 26435
rect 15163 26401 15197 26435
rect 15301 26401 15335 26435
rect 16037 26401 16071 26435
rect 1683 26333 1717 26367
rect 2789 26333 2823 26367
rect 3065 26333 3099 26367
rect 3341 26333 3375 26367
rect 3801 26333 3835 26367
rect 4075 26333 4109 26367
rect 5365 26333 5399 26367
rect 6285 26333 6319 26367
rect 7481 26333 7515 26367
rect 7755 26333 7789 26367
rect 9137 26333 9171 26367
rect 9505 26333 9539 26367
rect 9781 26333 9815 26367
rect 10055 26333 10089 26367
rect 11713 26333 11747 26367
rect 14105 26333 14139 26367
rect 14289 26333 14323 26367
rect 16295 26303 16329 26337
rect 17417 26333 17451 26367
rect 18521 26333 18555 26367
rect 19257 26333 19291 26367
rect 19349 26333 19383 26367
rect 19717 26333 19751 26367
rect 20269 26333 20303 26367
rect 20361 26333 20395 26367
rect 20821 26333 20855 26367
rect 21005 26333 21039 26367
rect 21189 26333 21223 26367
rect 11621 26265 11655 26299
rect 12081 26265 12115 26299
rect 12449 26265 12483 26299
rect 21557 26265 21591 26299
rect 2421 26197 2455 26231
rect 7205 26197 7239 26231
rect 8493 26197 8527 26231
rect 11345 26197 11379 26231
rect 17049 26197 17083 26231
rect 19533 26197 19567 26231
rect 1409 25993 1443 26027
rect 4353 25993 4387 26027
rect 8217 25993 8251 26027
rect 10701 25993 10735 26027
rect 13921 25993 13955 26027
rect 19165 25993 19199 26027
rect 3249 25925 3283 25959
rect 3617 25925 3651 25959
rect 3985 25925 4019 25959
rect 8493 25925 8527 25959
rect 8585 25925 8619 25959
rect 8953 25925 8987 25959
rect 9321 25925 9355 25959
rect 16037 25925 16071 25959
rect 16313 25925 16347 25959
rect 1593 25857 1627 25891
rect 1685 25857 1719 25891
rect 1959 25857 1993 25891
rect 3525 25857 3559 25891
rect 6561 25857 6595 25891
rect 6927 25857 6961 25891
rect 9689 25857 9723 25891
rect 9963 25857 9997 25891
rect 11529 25857 11563 25891
rect 11803 25857 11837 25891
rect 13183 25857 13217 25891
rect 15669 25857 15703 25891
rect 15853 25857 15887 25891
rect 16221 25857 16255 25891
rect 16405 25857 16439 25891
rect 17785 25857 17819 25891
rect 18041 25857 18075 25891
rect 19515 25887 19549 25921
rect 20913 25857 20947 25891
rect 21005 25857 21039 25891
rect 21281 25857 21315 25891
rect 6653 25789 6687 25823
rect 12909 25789 12943 25823
rect 19257 25789 19291 25823
rect 4537 25721 4571 25755
rect 7665 25721 7699 25755
rect 2697 25653 2731 25687
rect 6377 25653 6411 25687
rect 9505 25653 9539 25687
rect 12541 25653 12575 25687
rect 15945 25653 15979 25687
rect 20269 25653 20303 25687
rect 20729 25653 20763 25687
rect 21097 25653 21131 25687
rect 21465 25653 21499 25687
rect 3341 25449 3375 25483
rect 8125 25449 8159 25483
rect 10793 25449 10827 25483
rect 19533 25449 19567 25483
rect 19625 25449 19659 25483
rect 20085 25449 20119 25483
rect 3985 25381 4019 25415
rect 6377 25381 6411 25415
rect 9597 25381 9631 25415
rect 18705 25381 18739 25415
rect 1685 25313 1719 25347
rect 2329 25313 2363 25347
rect 5917 25313 5951 25347
rect 6653 25313 6687 25347
rect 6791 25313 6825 25347
rect 9137 25313 9171 25347
rect 9990 25313 10024 25347
rect 19717 25313 19751 25347
rect 19901 25313 19935 25347
rect 1409 25245 1443 25279
rect 2571 25245 2605 25279
rect 3801 25245 3835 25279
rect 4353 25245 4387 25279
rect 4627 25245 4661 25279
rect 5733 25245 5767 25279
rect 6929 25245 6963 25279
rect 7573 25245 7607 25279
rect 7941 25245 7975 25279
rect 8033 25245 8067 25279
rect 8953 25245 8987 25279
rect 9873 25245 9907 25279
rect 10149 25245 10183 25279
rect 11805 25245 11839 25279
rect 14105 25245 14139 25279
rect 15117 25245 15151 25279
rect 15391 25245 15425 25279
rect 16497 25245 16531 25279
rect 16755 25215 16789 25249
rect 18061 25245 18095 25279
rect 18429 25245 18463 25279
rect 18613 25245 18647 25279
rect 18889 25245 18923 25279
rect 19441 25245 19475 25279
rect 19809 25245 19843 25279
rect 19993 25245 20027 25279
rect 20269 25245 20303 25279
rect 20453 25245 20487 25279
rect 20637 25245 20671 25279
rect 20913 25245 20947 25279
rect 21189 25245 21223 25279
rect 11897 25177 11931 25211
rect 12265 25177 12299 25211
rect 21557 25177 21591 25211
rect 5365 25109 5399 25143
rect 7757 25109 7791 25143
rect 11529 25109 11563 25143
rect 12633 25109 12667 25143
rect 12817 25109 12851 25143
rect 14197 25109 14231 25143
rect 16129 25109 16163 25143
rect 17509 25109 17543 25143
rect 17877 25109 17911 25143
rect 18613 25109 18647 25143
rect 20637 25109 20671 25143
rect 20729 25109 20763 25143
rect 1409 24905 1443 24939
rect 10609 24905 10643 24939
rect 12541 24905 12575 24939
rect 18705 24905 18739 24939
rect 21005 24905 21039 24939
rect 1869 24837 1903 24871
rect 2145 24837 2179 24871
rect 2973 24837 3007 24871
rect 19892 24837 19926 24871
rect 1593 24769 1627 24803
rect 2237 24769 2271 24803
rect 2605 24769 2639 24803
rect 4719 24769 4753 24803
rect 7665 24769 7699 24803
rect 8723 24769 8757 24803
rect 9871 24769 9905 24803
rect 11803 24769 11837 24803
rect 13459 24779 13493 24813
rect 14565 24769 14599 24803
rect 14749 24769 14783 24803
rect 15025 24769 15059 24803
rect 15283 24799 15317 24833
rect 17325 24769 17359 24803
rect 17581 24769 17615 24803
rect 18797 24769 18831 24803
rect 19165 24769 19199 24803
rect 19625 24769 19659 24803
rect 21189 24769 21223 24803
rect 4445 24701 4479 24735
rect 7849 24701 7883 24735
rect 8585 24701 8619 24735
rect 8861 24701 8895 24735
rect 9597 24701 9631 24735
rect 11529 24701 11563 24735
rect 13185 24701 13219 24735
rect 19073 24701 19107 24735
rect 8309 24633 8343 24667
rect 14197 24633 14231 24667
rect 18889 24633 18923 24667
rect 19257 24633 19291 24667
rect 3157 24565 3191 24599
rect 5457 24565 5491 24599
rect 9505 24565 9539 24599
rect 14657 24565 14691 24599
rect 16037 24565 16071 24599
rect 18981 24565 19015 24599
rect 21465 24565 21499 24599
rect 1593 24361 1627 24395
rect 2697 24361 2731 24395
rect 8217 24361 8251 24395
rect 14749 24361 14783 24395
rect 17233 24361 17267 24395
rect 18613 24361 18647 24395
rect 20821 24361 20855 24395
rect 5365 24293 5399 24327
rect 16037 24293 16071 24327
rect 1685 24225 1719 24259
rect 5779 24225 5813 24259
rect 12449 24225 12483 24259
rect 14381 24225 14415 24259
rect 15577 24225 15611 24259
rect 16589 24225 16623 24259
rect 17601 24225 17635 24259
rect 19257 24225 19291 24259
rect 21005 24225 21039 24259
rect 1409 24157 1443 24191
rect 1943 24127 1977 24161
rect 4721 24157 4755 24191
rect 4905 24157 4939 24191
rect 5641 24157 5675 24191
rect 5917 24157 5951 24191
rect 7205 24157 7239 24191
rect 7463 24157 7497 24191
rect 10057 24157 10091 24191
rect 10149 24157 10183 24191
rect 10423 24157 10457 24191
rect 11529 24157 11563 24191
rect 11713 24157 11747 24191
rect 12723 24157 12757 24191
rect 14289 24157 14323 24191
rect 14657 24157 14691 24191
rect 14933 24157 14967 24191
rect 15393 24157 15427 24191
rect 16313 24157 16347 24191
rect 16430 24157 16464 24191
rect 17859 24127 17893 24161
rect 20729 24157 20763 24191
rect 21281 24157 21315 24191
rect 14565 24089 14599 24123
rect 19502 24089 19536 24123
rect 6561 24021 6595 24055
rect 9873 24021 9907 24055
rect 11161 24021 11195 24055
rect 11713 24021 11747 24055
rect 13461 24021 13495 24055
rect 20637 24021 20671 24055
rect 21005 24021 21039 24055
rect 21465 24021 21499 24055
rect 14749 23817 14783 23851
rect 19349 23817 19383 23851
rect 20637 23817 20671 23851
rect 11345 23749 11379 23783
rect 19165 23749 19199 23783
rect 1409 23681 1443 23715
rect 1683 23681 1717 23715
rect 4905 23681 4939 23715
rect 5179 23681 5213 23715
rect 7021 23681 7055 23715
rect 7389 23681 7423 23715
rect 7941 23681 7975 23715
rect 9597 23681 9631 23715
rect 10425 23681 10459 23715
rect 10517 23681 10551 23715
rect 10609 23681 10643 23715
rect 10977 23681 11011 23715
rect 11161 23681 11195 23715
rect 13829 23681 13863 23715
rect 15083 23681 15117 23715
rect 16923 23681 16957 23715
rect 19073 23681 19107 23715
rect 19257 23681 19291 23715
rect 19533 23681 19567 23715
rect 19899 23681 19933 23715
rect 21005 23681 21039 23715
rect 21373 23681 21407 23715
rect 2789 23613 2823 23647
rect 3065 23613 3099 23647
rect 7757 23613 7791 23647
rect 8401 23613 8435 23647
rect 8677 23613 8711 23647
rect 8794 23613 8828 23647
rect 8953 23613 8987 23647
rect 12909 23613 12943 23647
rect 13093 23613 13127 23647
rect 13553 23613 13587 23647
rect 13946 23613 13980 23647
rect 14105 23613 14139 23647
rect 14841 23613 14875 23647
rect 16681 23613 16715 23647
rect 19625 23613 19659 23647
rect 21281 23613 21315 23647
rect 6837 23545 6871 23579
rect 21097 23545 21131 23579
rect 21465 23545 21499 23579
rect 2421 23477 2455 23511
rect 5917 23477 5951 23511
rect 7481 23477 7515 23511
rect 10241 23477 10275 23511
rect 11253 23477 11287 23511
rect 15853 23477 15887 23511
rect 17693 23477 17727 23511
rect 21189 23477 21223 23511
rect 3525 23273 3559 23307
rect 8493 23273 8527 23307
rect 14657 23273 14691 23307
rect 20545 23273 20579 23307
rect 21465 23273 21499 23307
rect 3249 23205 3283 23239
rect 5917 23205 5951 23239
rect 16037 23205 16071 23239
rect 17233 23205 17267 23239
rect 19257 23205 19291 23239
rect 1685 23137 1719 23171
rect 6193 23137 6227 23171
rect 6310 23137 6344 23171
rect 6469 23137 6503 23171
rect 7481 23137 7515 23171
rect 11069 23137 11103 23171
rect 12449 23137 12483 23171
rect 15577 23137 15611 23171
rect 16313 23137 16347 23171
rect 16589 23137 16623 23171
rect 19533 23137 19567 23171
rect 1409 23069 1443 23103
rect 1959 23069 1993 23103
rect 3065 23069 3099 23103
rect 3341 23069 3375 23103
rect 3801 23069 3835 23103
rect 4075 23069 4109 23103
rect 5273 23069 5307 23103
rect 5457 23069 5491 23103
rect 7113 23069 7147 23103
rect 7389 23069 7423 23103
rect 7755 23069 7789 23103
rect 9689 23069 9723 23103
rect 9931 23069 9965 23103
rect 11343 23069 11377 23103
rect 12723 23069 12757 23103
rect 14841 23069 14875 23103
rect 15393 23069 15427 23103
rect 16430 23069 16464 23103
rect 18521 23069 18555 23103
rect 18889 23069 18923 23103
rect 19073 23069 19107 23103
rect 19441 23045 19475 23079
rect 19791 23039 19825 23073
rect 21189 23069 21223 23103
rect 1593 22933 1627 22967
rect 2697 22933 2731 22967
rect 4813 22933 4847 22967
rect 7205 22933 7239 22967
rect 10701 22933 10735 22967
rect 12081 22933 12115 22967
rect 13461 22933 13495 22967
rect 18337 22933 18371 22967
rect 19073 22933 19107 22967
rect 1685 22729 1719 22763
rect 2973 22729 3007 22763
rect 3341 22729 3375 22763
rect 9873 22729 9907 22763
rect 14749 22729 14783 22763
rect 19257 22729 19291 22763
rect 20361 22729 20395 22763
rect 21097 22729 21131 22763
rect 2053 22661 2087 22695
rect 2789 22661 2823 22695
rect 3617 22661 3651 22695
rect 3709 22661 3743 22695
rect 4077 22661 4111 22695
rect 4445 22661 4479 22695
rect 10241 22661 10275 22695
rect 10977 22661 11011 22695
rect 1961 22593 1995 22627
rect 2421 22593 2455 22627
rect 6837 22593 6871 22627
rect 7111 22593 7145 22627
rect 8585 22593 8619 22627
rect 9045 22593 9079 22627
rect 10149 22593 10183 22627
rect 10609 22593 10643 22627
rect 12909 22593 12943 22627
rect 13093 22593 13127 22627
rect 15191 22623 15225 22657
rect 17877 22593 17911 22627
rect 18144 22593 18178 22627
rect 19591 22593 19625 22627
rect 20913 22593 20947 22627
rect 21281 22593 21315 22627
rect 8309 22525 8343 22559
rect 13553 22525 13587 22559
rect 13829 22525 13863 22559
rect 13946 22525 13980 22559
rect 14105 22525 14139 22559
rect 14933 22525 14967 22559
rect 19349 22525 19383 22559
rect 21557 22525 21591 22559
rect 4629 22457 4663 22491
rect 7849 22457 7883 22491
rect 9045 22457 9079 22491
rect 11161 22389 11195 22423
rect 15945 22389 15979 22423
rect 21373 22389 21407 22423
rect 21465 22389 21499 22423
rect 10149 22185 10183 22219
rect 21465 22185 21499 22219
rect 2789 22117 2823 22151
rect 3433 22117 3467 22151
rect 6377 22117 6411 22151
rect 16037 22117 16071 22151
rect 1409 22049 1443 22083
rect 6561 22049 6595 22083
rect 8033 22049 8067 22083
rect 9137 22049 9171 22083
rect 10609 22049 10643 22083
rect 12081 22049 12115 22083
rect 12725 22049 12759 22083
rect 13001 22049 13035 22083
rect 13277 22049 13311 22083
rect 15393 22049 15427 22083
rect 16430 22049 16464 22083
rect 16589 22049 16623 22083
rect 17325 22049 17359 22083
rect 1685 21981 1719 22015
rect 2329 21981 2363 22015
rect 2605 21981 2639 22015
rect 3249 21957 3283 21991
rect 5365 21981 5399 22015
rect 5457 21981 5491 22015
rect 6835 21981 6869 22015
rect 7941 21981 7975 22015
rect 8125 21981 8159 22015
rect 9379 21981 9413 22015
rect 10851 21981 10885 22015
rect 12265 21981 12299 22015
rect 13118 21981 13152 22015
rect 15577 21981 15611 22015
rect 16313 21981 16347 22015
rect 17599 21981 17633 22015
rect 18889 21981 18923 22015
rect 19441 21981 19475 22015
rect 20913 21981 20947 22015
rect 21281 21981 21315 22015
rect 2973 21913 3007 21947
rect 5825 21913 5859 21947
rect 19708 21913 19742 21947
rect 2513 21845 2547 21879
rect 3065 21845 3099 21879
rect 5089 21845 5123 21879
rect 6193 21845 6227 21879
rect 7573 21845 7607 21879
rect 11621 21845 11655 21879
rect 13921 21845 13955 21879
rect 17233 21845 17267 21879
rect 18337 21845 18371 21879
rect 18981 21845 19015 21879
rect 20821 21845 20855 21879
rect 21097 21845 21131 21879
rect 3893 21641 3927 21675
rect 5825 21641 5859 21675
rect 10241 21641 10275 21675
rect 10425 21641 10459 21675
rect 12817 21641 12851 21675
rect 9137 21573 9171 21607
rect 9873 21573 9907 21607
rect 11713 21573 11747 21607
rect 12449 21573 12483 21607
rect 1775 21505 1809 21539
rect 2881 21505 2915 21539
rect 3155 21505 3189 21539
rect 4535 21515 4569 21549
rect 7815 21505 7849 21539
rect 9413 21505 9447 21539
rect 9505 21505 9539 21539
rect 11989 21505 12023 21539
rect 12081 21505 12115 21539
rect 16681 21505 16715 21539
rect 17601 21505 17635 21539
rect 19867 21515 19901 21549
rect 21005 21505 21039 21539
rect 21557 21505 21591 21539
rect 1501 21437 1535 21471
rect 4261 21437 4295 21471
rect 7573 21437 7607 21471
rect 16865 21437 16899 21471
rect 17718 21437 17752 21471
rect 17877 21437 17911 21471
rect 19625 21437 19659 21471
rect 21281 21437 21315 21471
rect 5273 21369 5307 21403
rect 8585 21369 8619 21403
rect 17325 21369 17359 21403
rect 20637 21369 20671 21403
rect 2513 21301 2547 21335
rect 10793 21301 10827 21335
rect 13001 21301 13035 21335
rect 18521 21301 18555 21335
rect 21097 21301 21131 21335
rect 21189 21301 21223 21335
rect 21373 21301 21407 21335
rect 3985 21097 4019 21131
rect 5733 21097 5767 21131
rect 9965 21097 9999 21131
rect 12265 21097 12299 21131
rect 17693 21097 17727 21131
rect 20177 21097 20211 21131
rect 20729 21097 20763 21131
rect 5089 21029 5123 21063
rect 1409 20961 1443 20995
rect 1685 20961 1719 20995
rect 14105 20961 14139 20995
rect 16681 20961 16715 20995
rect 2329 20893 2363 20927
rect 2603 20893 2637 20927
rect 3801 20893 3835 20927
rect 4077 20893 4111 20927
rect 4351 20893 4385 20927
rect 6561 20893 6595 20927
rect 6929 20893 6963 20927
rect 8953 20893 8987 20927
rect 9227 20893 9261 20927
rect 11253 20893 11287 20927
rect 11527 20893 11561 20927
rect 14347 20893 14381 20927
rect 16037 20893 16071 20927
rect 16129 20893 16163 20927
rect 16313 20893 16347 20927
rect 16955 20893 16989 20927
rect 20085 20893 20119 20927
rect 6469 20825 6503 20859
rect 15669 20825 15703 20859
rect 20453 20825 20487 20859
rect 21005 20825 21039 20859
rect 21373 20825 21407 20859
rect 3341 20757 3375 20791
rect 6193 20757 6227 20791
rect 7297 20757 7331 20791
rect 7481 20757 7515 20791
rect 15117 20757 15151 20791
rect 15853 20757 15887 20791
rect 16313 20757 16347 20791
rect 2329 20553 2363 20587
rect 3985 20553 4019 20587
rect 5089 20553 5123 20587
rect 17785 20553 17819 20587
rect 19257 20553 19291 20587
rect 2605 20485 2639 20519
rect 3433 20485 3467 20519
rect 4261 20485 4295 20519
rect 4721 20485 4755 20519
rect 5549 20485 5583 20519
rect 5733 20485 5767 20519
rect 7573 20485 7607 20519
rect 7849 20485 7883 20519
rect 8309 20485 8343 20519
rect 8677 20485 8711 20519
rect 14933 20485 14967 20519
rect 1409 20417 1443 20451
rect 2053 20417 2087 20451
rect 2697 20417 2731 20451
rect 3065 20417 3099 20451
rect 4353 20417 4387 20451
rect 7941 20417 7975 20451
rect 10057 20417 10091 20451
rect 10331 20417 10365 20451
rect 11787 20447 11821 20481
rect 13277 20417 13311 20451
rect 15025 20417 15059 20451
rect 15299 20417 15333 20451
rect 17015 20417 17049 20451
rect 19441 20417 19475 20451
rect 19791 20447 19825 20481
rect 21189 20417 21223 20451
rect 21281 20417 21315 20451
rect 11529 20349 11563 20383
rect 13093 20349 13127 20383
rect 14013 20349 14047 20383
rect 14151 20349 14185 20383
rect 14289 20349 14323 20383
rect 16773 20349 16807 20383
rect 19533 20349 19567 20383
rect 1593 20281 1627 20315
rect 13737 20281 13771 20315
rect 3617 20213 3651 20247
rect 5273 20213 5307 20247
rect 6653 20213 6687 20247
rect 8861 20213 8895 20247
rect 11069 20213 11103 20247
rect 12541 20213 12575 20247
rect 16037 20213 16071 20247
rect 20545 20213 20579 20247
rect 21005 20213 21039 20247
rect 21465 20213 21499 20247
rect 1593 20009 1627 20043
rect 3341 20009 3375 20043
rect 11253 20009 11287 20043
rect 15945 20009 15979 20043
rect 20637 20009 20671 20043
rect 2053 19941 2087 19975
rect 3985 19941 4019 19975
rect 5549 19941 5583 19975
rect 13645 19941 13679 19975
rect 14749 19941 14783 19975
rect 17509 19941 17543 19975
rect 2329 19873 2363 19907
rect 4537 19873 4571 19907
rect 12633 19873 12667 19907
rect 14105 19873 14139 19907
rect 15025 19873 15059 19907
rect 15142 19873 15176 19907
rect 15301 19873 15335 19907
rect 19257 19873 19291 19907
rect 1501 19805 1535 19839
rect 2587 19775 2621 19809
rect 3801 19805 3835 19839
rect 4779 19805 4813 19839
rect 6377 19805 6411 19839
rect 10241 19805 10275 19839
rect 10333 19805 10367 19839
rect 11529 19805 11563 19839
rect 12891 19775 12925 19809
rect 14289 19805 14323 19839
rect 18797 19805 18831 19839
rect 19073 19805 19107 19839
rect 19513 19805 19547 19839
rect 20913 19805 20947 19839
rect 21097 19805 21131 19839
rect 21281 19805 21315 19839
rect 1869 19737 1903 19771
rect 6055 19737 6089 19771
rect 6469 19737 6503 19771
rect 6837 19737 6871 19771
rect 7205 19737 7239 19771
rect 10701 19737 10735 19771
rect 11713 19737 11747 19771
rect 16497 19737 16531 19771
rect 16589 19737 16623 19771
rect 16957 19737 16991 19771
rect 17325 19737 17359 19771
rect 21005 19737 21039 19771
rect 7389 19669 7423 19703
rect 9965 19669 9999 19703
rect 11069 19669 11103 19703
rect 16221 19669 16255 19703
rect 18613 19669 18647 19703
rect 18889 19669 18923 19703
rect 21465 19669 21499 19703
rect 2513 19465 2547 19499
rect 3065 19465 3099 19499
rect 5917 19465 5951 19499
rect 8493 19465 8527 19499
rect 17693 19465 17727 19499
rect 16313 19397 16347 19431
rect 19318 19397 19352 19431
rect 1501 19329 1535 19363
rect 1775 19329 1809 19363
rect 2881 19329 2915 19363
rect 3525 19329 3559 19363
rect 3767 19329 3801 19363
rect 4905 19329 4939 19363
rect 5179 19329 5213 19363
rect 7481 19329 7515 19363
rect 7755 19329 7789 19363
rect 10299 19339 10333 19373
rect 12633 19329 12667 19363
rect 13507 19329 13541 19363
rect 14381 19329 14415 19363
rect 14655 19329 14689 19363
rect 15945 19329 15979 19363
rect 16129 19329 16163 19363
rect 16681 19329 16715 19363
rect 16955 19329 16989 19363
rect 18797 19329 18831 19363
rect 20545 19329 20579 19363
rect 21189 19329 21223 19363
rect 10057 19261 10091 19295
rect 12449 19261 12483 19295
rect 13369 19261 13403 19295
rect 13645 19261 13679 19295
rect 19073 19261 19107 19295
rect 20821 19261 20855 19295
rect 13093 19193 13127 19227
rect 20637 19193 20671 19227
rect 4537 19125 4571 19159
rect 7389 19125 7423 19159
rect 11069 19125 11103 19159
rect 14289 19125 14323 19159
rect 15393 19125 15427 19159
rect 16221 19125 16255 19159
rect 18889 19125 18923 19159
rect 20453 19125 20487 19159
rect 20729 19125 20763 19159
rect 21465 19125 21499 19159
rect 5733 18921 5767 18955
rect 7113 18921 7147 18955
rect 10425 18921 10459 18955
rect 13553 18921 13587 18955
rect 15393 18921 15427 18955
rect 16773 18921 16807 18955
rect 21097 18921 21131 18955
rect 11713 18853 11747 18887
rect 1409 18785 1443 18819
rect 1685 18785 1719 18819
rect 2329 18785 2363 18819
rect 3801 18785 3835 18819
rect 4077 18785 4111 18819
rect 4721 18785 4755 18819
rect 6101 18785 6135 18819
rect 9413 18785 9447 18819
rect 11069 18785 11103 18819
rect 11989 18785 12023 18819
rect 12106 18785 12140 18819
rect 12265 18785 12299 18819
rect 15761 18785 15795 18819
rect 17417 18785 17451 18819
rect 19257 18785 19291 18819
rect 20729 18785 20763 18819
rect 21005 18785 21039 18819
rect 21189 18785 21223 18819
rect 2571 18717 2605 18751
rect 4995 18717 5029 18751
rect 6359 18687 6393 18721
rect 7481 18717 7515 18751
rect 7755 18717 7789 18751
rect 9137 18717 9171 18751
rect 9687 18717 9721 18751
rect 11253 18717 11287 18751
rect 12909 18717 12943 18751
rect 15301 18717 15335 18751
rect 16035 18717 16069 18751
rect 17141 18717 17175 18751
rect 19499 18717 19533 18751
rect 20637 18717 20671 18751
rect 20913 18717 20947 18751
rect 21281 18717 21315 18751
rect 3341 18581 3375 18615
rect 8493 18581 8527 18615
rect 20269 18581 20303 18615
rect 21465 18581 21499 18615
rect 5641 18377 5675 18411
rect 8401 18377 8435 18411
rect 9505 18377 9539 18411
rect 9689 18377 9723 18411
rect 13093 18377 13127 18411
rect 16129 18377 16163 18411
rect 20545 18377 20579 18411
rect 2053 18309 2087 18343
rect 2237 18309 2271 18343
rect 8677 18309 8711 18343
rect 9137 18309 9171 18343
rect 18950 18309 18984 18343
rect 21189 18309 21223 18343
rect 1501 18241 1535 18275
rect 2663 18241 2697 18275
rect 3801 18241 3835 18275
rect 4997 18241 5031 18275
rect 7111 18241 7145 18275
rect 8769 18241 8803 18275
rect 10331 18241 10365 18275
rect 12323 18241 12357 18275
rect 14163 18241 14197 18275
rect 16313 18241 16347 18275
rect 16939 18271 16973 18305
rect 20361 18241 20395 18275
rect 20545 18241 20579 18275
rect 20821 18241 20855 18275
rect 2421 18173 2455 18207
rect 3985 18173 4019 18207
rect 4721 18173 4755 18207
rect 4838 18173 4872 18207
rect 6837 18173 6871 18207
rect 10057 18173 10091 18207
rect 12081 18173 12115 18207
rect 13921 18173 13955 18207
rect 16681 18173 16715 18207
rect 18705 18173 18739 18207
rect 4445 18105 4479 18139
rect 20085 18105 20119 18139
rect 20637 18105 20671 18139
rect 1593 18037 1627 18071
rect 3433 18037 3467 18071
rect 7849 18037 7883 18071
rect 11069 18037 11103 18071
rect 14933 18037 14967 18071
rect 17693 18037 17727 18071
rect 21465 18037 21499 18071
rect 9965 17833 9999 17867
rect 21005 17833 21039 17867
rect 1593 17765 1627 17799
rect 6745 17765 6779 17799
rect 8677 17765 8711 17799
rect 13645 17765 13679 17799
rect 14749 17765 14783 17799
rect 19717 17765 19751 17799
rect 1777 17697 1811 17731
rect 2421 17697 2455 17731
rect 2697 17697 2731 17731
rect 2835 17697 2869 17731
rect 5733 17697 5767 17731
rect 12633 17697 12667 17731
rect 15025 17697 15059 17731
rect 15301 17697 15335 17731
rect 20085 17697 20119 17731
rect 20453 17697 20487 17731
rect 20637 17697 20671 17731
rect 1409 17629 1443 17663
rect 1961 17629 1995 17663
rect 2973 17629 3007 17663
rect 4813 17629 4847 17663
rect 6007 17629 6041 17663
rect 7665 17629 7699 17663
rect 7757 17629 7791 17663
rect 8125 17629 8159 17663
rect 8953 17629 8987 17663
rect 9227 17629 9261 17663
rect 10701 17629 10735 17663
rect 10975 17629 11009 17663
rect 12875 17629 12909 17663
rect 14105 17629 14139 17663
rect 14289 17629 14323 17663
rect 15142 17629 15176 17663
rect 17693 17629 17727 17663
rect 17967 17629 18001 17663
rect 19441 17629 19475 17663
rect 19901 17629 19935 17663
rect 19993 17629 20027 17663
rect 20361 17629 20395 17663
rect 20913 17629 20947 17663
rect 21097 17629 21131 17663
rect 21281 17629 21315 17663
rect 7389 17561 7423 17595
rect 16497 17561 16531 17595
rect 16589 17561 16623 17595
rect 16957 17561 16991 17595
rect 3617 17493 3651 17527
rect 4629 17493 4663 17527
rect 5365 17493 5399 17527
rect 8493 17493 8527 17527
rect 11713 17493 11747 17527
rect 15945 17493 15979 17527
rect 16221 17493 16255 17527
rect 17325 17493 17359 17527
rect 17509 17493 17543 17527
rect 18705 17493 18739 17527
rect 19257 17493 19291 17527
rect 20637 17493 20671 17527
rect 21465 17493 21499 17527
rect 1685 17289 1719 17323
rect 3433 17289 3467 17323
rect 8493 17289 8527 17323
rect 15025 17289 15059 17323
rect 16221 17289 16255 17323
rect 20637 17289 20671 17323
rect 20729 17289 20763 17323
rect 1593 17221 1627 17255
rect 7205 17221 7239 17255
rect 7573 17221 7607 17255
rect 7941 17221 7975 17255
rect 8309 17221 8343 17255
rect 2663 17163 2697 17197
rect 3801 17153 3835 17187
rect 4997 17153 5031 17187
rect 5917 17153 5951 17187
rect 7481 17153 7515 17187
rect 10223 17183 10257 17217
rect 11529 17153 11563 17187
rect 12173 17153 12207 17187
rect 14841 17153 14875 17187
rect 15451 17153 15485 17187
rect 16681 17153 16715 17187
rect 17601 17153 17635 17187
rect 19165 17153 19199 17187
rect 19524 17153 19558 17187
rect 20913 17153 20947 17187
rect 21005 17153 21039 17187
rect 21189 17153 21223 17187
rect 21281 17153 21315 17187
rect 2421 17085 2455 17119
rect 3985 17085 4019 17119
rect 4445 17085 4479 17119
rect 4721 17085 4755 17119
rect 4838 17085 4872 17119
rect 9965 17085 9999 17119
rect 12357 17085 12391 17119
rect 13093 17085 13127 17119
rect 13231 17085 13265 17119
rect 13369 17085 13403 17119
rect 15209 17085 15243 17119
rect 16865 17085 16899 17119
rect 17718 17085 17752 17119
rect 17875 17085 17909 17119
rect 18797 17085 18831 17119
rect 19257 17085 19291 17119
rect 5733 17017 5767 17051
rect 12817 17017 12851 17051
rect 17325 17017 17359 17051
rect 5641 16949 5675 16983
rect 10977 16949 11011 16983
rect 11713 16949 11747 16983
rect 14013 16949 14047 16983
rect 18521 16949 18555 16983
rect 18981 16949 19015 16983
rect 21097 16949 21131 16983
rect 21465 16949 21499 16983
rect 2881 16745 2915 16779
rect 4537 16745 4571 16779
rect 6837 16745 6871 16779
rect 8493 16745 8527 16779
rect 13461 16745 13495 16779
rect 16773 16745 16807 16779
rect 17877 16745 17911 16779
rect 20361 16745 20395 16779
rect 10977 16677 11011 16711
rect 15577 16677 15611 16711
rect 1869 16609 1903 16643
rect 4997 16609 5031 16643
rect 5641 16609 5675 16643
rect 5917 16609 5951 16643
rect 6193 16609 6227 16643
rect 7481 16609 7515 16643
rect 8953 16609 8987 16643
rect 10333 16609 10367 16643
rect 11253 16609 11287 16643
rect 11529 16609 11563 16643
rect 15117 16609 15151 16643
rect 15970 16609 16004 16643
rect 16129 16609 16163 16643
rect 21005 16609 21039 16643
rect 21465 16609 21499 16643
rect 2143 16541 2177 16575
rect 3617 16541 3651 16575
rect 4445 16541 4479 16575
rect 5181 16541 5215 16575
rect 6055 16541 6089 16575
rect 7723 16541 7757 16575
rect 9227 16541 9261 16575
rect 10517 16541 10551 16575
rect 11370 16541 11404 16575
rect 12449 16541 12483 16575
rect 12723 16541 12757 16575
rect 14105 16541 14139 16575
rect 14933 16541 14967 16575
rect 15853 16541 15887 16575
rect 16865 16541 16899 16575
rect 17139 16531 17173 16565
rect 19349 16541 19383 16575
rect 19607 16511 19641 16545
rect 20729 16541 20763 16575
rect 20821 16541 20855 16575
rect 3893 16473 3927 16507
rect 7113 16473 7147 16507
rect 21189 16473 21223 16507
rect 3433 16405 3467 16439
rect 3985 16405 4019 16439
rect 9965 16405 9999 16439
rect 12173 16405 12207 16439
rect 14289 16405 14323 16439
rect 21005 16405 21039 16439
rect 1593 16201 1627 16235
rect 5917 16201 5951 16235
rect 11345 16201 11379 16235
rect 12909 16201 12943 16235
rect 15669 16201 15703 16235
rect 17693 16201 17727 16235
rect 18797 16201 18831 16235
rect 20637 16201 20671 16235
rect 21097 16201 21131 16235
rect 1501 16133 1535 16167
rect 2421 16065 2455 16099
rect 3433 16065 3467 16099
rect 4261 16065 4295 16099
rect 5163 16095 5197 16129
rect 8125 16065 8159 16099
rect 8399 16065 8433 16099
rect 9505 16065 9539 16099
rect 10563 16065 10597 16099
rect 11897 16065 11931 16099
rect 12171 16065 12205 16099
rect 13551 16065 13585 16099
rect 14931 16065 14965 16099
rect 16221 16065 16255 16099
rect 16923 16065 16957 16099
rect 18337 16065 18371 16099
rect 18981 16065 19015 16099
rect 19073 16065 19107 16099
rect 19257 16065 19291 16099
rect 19867 16065 19901 16099
rect 21005 16065 21039 16099
rect 21281 16065 21315 16099
rect 2237 15997 2271 16031
rect 3157 15997 3191 16031
rect 3295 15997 3329 16031
rect 4905 15997 4939 16031
rect 7757 15997 7791 16031
rect 9689 15997 9723 16031
rect 10149 15997 10183 16031
rect 10425 15997 10459 16031
rect 10701 15997 10735 16031
rect 13277 15997 13311 16031
rect 14657 15997 14691 16031
rect 16681 15997 16715 16031
rect 19625 15997 19659 16031
rect 2881 15929 2915 15963
rect 4077 15861 4111 15895
rect 4353 15861 4387 15895
rect 9137 15861 9171 15895
rect 14289 15861 14323 15895
rect 18429 15861 18463 15895
rect 19165 15861 19199 15895
rect 21465 15861 21499 15895
rect 2421 15657 2455 15691
rect 2881 15657 2915 15691
rect 5917 15657 5951 15691
rect 13921 15657 13955 15691
rect 17049 15657 17083 15691
rect 18889 15657 18923 15691
rect 20913 15657 20947 15691
rect 18705 15589 18739 15623
rect 4077 15521 4111 15555
rect 4721 15521 4755 15555
rect 4997 15521 5031 15555
rect 5114 15521 5148 15555
rect 12081 15521 12115 15555
rect 12725 15521 12759 15555
rect 13001 15521 13035 15555
rect 13277 15521 13311 15555
rect 14565 15521 14599 15555
rect 19073 15521 19107 15555
rect 1409 15453 1443 15487
rect 1683 15453 1717 15487
rect 3065 15453 3099 15487
rect 3985 15453 4019 15487
rect 4261 15453 4295 15487
rect 5273 15453 5307 15487
rect 6193 15453 6227 15487
rect 7021 15453 7055 15487
rect 9229 15453 9263 15487
rect 9471 15453 9505 15487
rect 12265 15453 12299 15487
rect 13139 15453 13173 15487
rect 14105 15453 14139 15487
rect 14807 15453 14841 15487
rect 17233 15453 17267 15487
rect 17325 15453 17359 15487
rect 18797 15453 18831 15487
rect 19257 15453 19291 15487
rect 19524 15453 19558 15487
rect 20821 15453 20855 15487
rect 21005 15453 21039 15487
rect 21189 15453 21223 15487
rect 3249 15385 3283 15419
rect 6653 15385 6687 15419
rect 6929 15385 6963 15419
rect 7389 15385 7423 15419
rect 7757 15385 7791 15419
rect 17570 15385 17604 15419
rect 21557 15385 21591 15419
rect 3341 15317 3375 15351
rect 3801 15317 3835 15351
rect 6009 15317 6043 15351
rect 7941 15317 7975 15351
rect 10241 15317 10275 15351
rect 14289 15317 14323 15351
rect 15577 15317 15611 15351
rect 19073 15317 19107 15351
rect 20637 15317 20671 15351
rect 4813 15113 4847 15147
rect 13093 15113 13127 15147
rect 18797 15113 18831 15147
rect 1851 15007 1885 15041
rect 4010 14977 4044 15011
rect 4169 14977 4203 15011
rect 5179 14977 5213 15011
rect 6561 14977 6595 15011
rect 8935 15007 8969 15041
rect 10057 14977 10091 15011
rect 10315 15007 10349 15041
rect 12081 14977 12115 15011
rect 12355 14977 12389 15011
rect 18059 14977 18093 15011
rect 19809 14977 19843 15011
rect 20269 14977 20303 15011
rect 20821 14977 20855 15011
rect 20913 14977 20947 15011
rect 21097 14977 21131 15011
rect 21281 14977 21315 15011
rect 1593 14909 1627 14943
rect 2973 14909 3007 14943
rect 3157 14909 3191 14943
rect 3893 14909 3927 14943
rect 4905 14909 4939 14943
rect 6377 14909 6411 14943
rect 7297 14909 7331 14943
rect 7435 14909 7469 14943
rect 7573 14909 7607 14943
rect 8677 14909 8711 14943
rect 13737 14909 13771 14943
rect 13921 14909 13955 14943
rect 14657 14909 14691 14943
rect 14795 14909 14829 14943
rect 14933 14909 14967 14943
rect 17785 14909 17819 14943
rect 2605 14841 2639 14875
rect 3597 14841 3631 14875
rect 7021 14841 7055 14875
rect 14381 14841 14415 14875
rect 19625 14841 19659 14875
rect 20637 14841 20671 14875
rect 5917 14773 5951 14807
rect 8217 14773 8251 14807
rect 9689 14773 9723 14807
rect 11069 14773 11103 14807
rect 15577 14773 15611 14807
rect 20361 14773 20395 14807
rect 21005 14773 21039 14807
rect 21465 14773 21499 14807
rect 1777 14569 1811 14603
rect 3341 14569 3375 14603
rect 5273 14569 5307 14603
rect 6653 14569 6687 14603
rect 8033 14569 8067 14603
rect 13645 14569 13679 14603
rect 15117 14569 15151 14603
rect 10517 14501 10551 14535
rect 15669 14501 15703 14535
rect 20545 14501 20579 14535
rect 10057 14433 10091 14467
rect 10910 14433 10944 14467
rect 12449 14433 12483 14467
rect 12725 14433 12759 14467
rect 12863 14433 12897 14467
rect 19533 14433 19567 14467
rect 21189 14433 21223 14467
rect 1685 14365 1719 14399
rect 2329 14365 2363 14399
rect 2603 14365 2637 14399
rect 4261 14365 4295 14399
rect 4519 14335 4553 14369
rect 5641 14365 5675 14399
rect 5915 14365 5949 14399
rect 7021 14365 7055 14399
rect 7263 14365 7297 14399
rect 9873 14365 9907 14399
rect 10793 14365 10827 14399
rect 11069 14365 11103 14399
rect 11805 14365 11839 14399
rect 11989 14365 12023 14399
rect 13001 14365 13035 14399
rect 14105 14365 14139 14399
rect 14347 14365 14381 14399
rect 15485 14365 15519 14399
rect 15761 14365 15795 14399
rect 19775 14365 19809 14399
rect 20913 14365 20947 14399
rect 21005 14365 21039 14399
rect 21281 14365 21315 14399
rect 11713 14229 11747 14263
rect 15945 14229 15979 14263
rect 21189 14229 21223 14263
rect 21465 14229 21499 14263
rect 1869 14025 1903 14059
rect 4261 14025 4295 14059
rect 5917 14025 5951 14059
rect 8033 14025 8067 14059
rect 11253 14025 11287 14059
rect 12909 14025 12943 14059
rect 15117 14025 15151 14059
rect 20821 14025 20855 14059
rect 6745 13957 6779 13991
rect 7021 13957 7055 13991
rect 15393 13957 15427 13991
rect 15485 13957 15519 13991
rect 16221 13957 16255 13991
rect 19073 13957 19107 13991
rect 1593 13889 1627 13923
rect 1777 13889 1811 13923
rect 3249 13889 3283 13923
rect 3523 13889 3557 13923
rect 5179 13889 5213 13923
rect 7113 13889 7147 13923
rect 7481 13889 7515 13923
rect 7863 13889 7897 13923
rect 9919 13889 9953 13923
rect 10057 13889 10091 13923
rect 10701 13889 10735 13923
rect 10793 13889 10827 13923
rect 11069 13889 11103 13923
rect 11897 13889 11931 13923
rect 12155 13919 12189 13953
rect 15853 13889 15887 13923
rect 16681 13889 16715 13923
rect 16955 13889 16989 13923
rect 18981 13889 19015 13923
rect 19441 13889 19475 13923
rect 19708 13889 19742 13923
rect 21189 13889 21223 13923
rect 4905 13821 4939 13855
rect 8861 13821 8895 13855
rect 9045 13821 9079 13855
rect 9781 13821 9815 13855
rect 1409 13753 1443 13787
rect 9505 13753 9539 13787
rect 16405 13753 16439 13787
rect 17693 13753 17727 13787
rect 2881 13685 2915 13719
rect 10977 13685 11011 13719
rect 21465 13685 21499 13719
rect 1777 13481 1811 13515
rect 3249 13481 3283 13515
rect 5825 13481 5859 13515
rect 7113 13481 7147 13515
rect 8493 13481 8527 13515
rect 12725 13481 12759 13515
rect 15945 13481 15979 13515
rect 17141 13481 17175 13515
rect 19257 13481 19291 13515
rect 21189 13481 21223 13515
rect 14749 13413 14783 13447
rect 2237 13345 2271 13379
rect 4445 13345 4479 13379
rect 4721 13345 4755 13379
rect 4859 13345 4893 13379
rect 5007 13345 5041 13379
rect 6101 13345 6135 13379
rect 7481 13345 7515 13379
rect 9781 13345 9815 13379
rect 10425 13345 10459 13379
rect 10701 13345 10735 13379
rect 10839 13345 10873 13379
rect 11713 13345 11747 13379
rect 14105 13345 14139 13379
rect 14289 13345 14323 13379
rect 15142 13345 15176 13379
rect 16129 13345 16163 13379
rect 1685 13277 1719 13311
rect 2511 13277 2545 13311
rect 3801 13277 3835 13311
rect 3985 13277 4019 13311
rect 6009 13277 6043 13311
rect 6375 13277 6409 13311
rect 7755 13277 7789 13311
rect 9137 13277 9171 13311
rect 9965 13277 9999 13311
rect 10977 13277 11011 13311
rect 11955 13277 11989 13311
rect 15025 13277 15059 13311
rect 15301 13277 15335 13311
rect 16387 13247 16421 13281
rect 17693 13277 17727 13311
rect 17960 13277 17994 13311
rect 19441 13277 19475 13311
rect 19625 13277 19659 13311
rect 19899 13277 19933 13311
rect 21557 13277 21591 13311
rect 5641 13141 5675 13175
rect 8953 13141 8987 13175
rect 11621 13141 11655 13175
rect 19073 13141 19107 13175
rect 20637 13141 20671 13175
rect 21373 13141 21407 13175
rect 14473 12937 14507 12971
rect 15853 12937 15887 12971
rect 1685 12869 1719 12903
rect 4169 12869 4203 12903
rect 6653 12869 6687 12903
rect 6929 12869 6963 12903
rect 7389 12869 7423 12903
rect 7757 12869 7791 12903
rect 20821 12869 20855 12903
rect 21557 12869 21591 12903
rect 2513 12801 2547 12835
rect 3249 12801 3283 12835
rect 3525 12801 3559 12835
rect 4963 12801 4997 12835
rect 7021 12801 7055 12835
rect 8951 12801 8985 12835
rect 10331 12801 10365 12835
rect 12081 12801 12115 12835
rect 12355 12801 12389 12835
rect 13735 12801 13769 12835
rect 14841 12801 14875 12835
rect 15115 12801 15149 12835
rect 17785 12801 17819 12835
rect 18337 12801 18371 12835
rect 18611 12801 18645 12835
rect 19717 12801 19751 12835
rect 19809 12801 19843 12835
rect 20269 12801 20303 12835
rect 20453 12801 20487 12835
rect 21281 12801 21315 12835
rect 2329 12733 2363 12767
rect 3387 12733 3421 12767
rect 4721 12733 4755 12767
rect 8677 12733 8711 12767
rect 10057 12733 10091 12767
rect 13461 12733 13495 12767
rect 17969 12733 18003 12767
rect 19993 12733 20027 12767
rect 21557 12733 21591 12767
rect 2973 12665 3007 12699
rect 5733 12665 5767 12699
rect 7941 12665 7975 12699
rect 9689 12665 9723 12699
rect 11069 12665 11103 12699
rect 19349 12665 19383 12699
rect 20545 12665 20579 12699
rect 21373 12665 21407 12699
rect 1777 12597 1811 12631
rect 13093 12597 13127 12631
rect 19901 12597 19935 12631
rect 20085 12597 20119 12631
rect 21097 12597 21131 12631
rect 1593 12393 1627 12427
rect 3341 12393 3375 12427
rect 4353 12393 4387 12427
rect 5733 12393 5767 12427
rect 7113 12393 7147 12427
rect 19533 12393 19567 12427
rect 20361 12393 20395 12427
rect 21465 12393 21499 12427
rect 8493 12325 8527 12359
rect 13645 12325 13679 12359
rect 16037 12325 16071 12359
rect 2329 12257 2363 12291
rect 4721 12257 4755 12291
rect 7481 12257 7515 12291
rect 10057 12257 10091 12291
rect 10517 12257 10551 12291
rect 10793 12257 10827 12291
rect 11069 12257 11103 12291
rect 12633 12257 12667 12291
rect 15025 12257 15059 12291
rect 16865 12257 16899 12291
rect 2237 12189 2271 12223
rect 2603 12189 2637 12223
rect 3985 12189 4019 12223
rect 4995 12189 5029 12223
rect 6101 12189 6135 12223
rect 6375 12189 6409 12223
rect 7755 12189 7789 12223
rect 9873 12189 9907 12223
rect 10931 12189 10965 12223
rect 12907 12189 12941 12223
rect 15283 12159 15317 12193
rect 17107 12189 17141 12223
rect 18245 12189 18279 12223
rect 18429 12189 18463 12223
rect 18705 12189 18739 12223
rect 19441 12189 19475 12223
rect 19625 12189 19659 12223
rect 19901 12189 19935 12223
rect 19993 12189 20027 12223
rect 20177 12189 20211 12223
rect 20269 12189 20303 12223
rect 20453 12189 20487 12223
rect 20545 12189 20579 12223
rect 20913 12189 20947 12223
rect 21281 12189 21315 12223
rect 1501 12121 1535 12155
rect 4261 12121 4295 12155
rect 2053 12053 2087 12087
rect 3801 12053 3835 12087
rect 11713 12053 11747 12087
rect 17877 12053 17911 12087
rect 18337 12053 18371 12087
rect 18521 12053 18555 12087
rect 19717 12053 19751 12087
rect 20177 12053 20211 12087
rect 20729 12053 20763 12087
rect 21097 12053 21131 12087
rect 1409 11849 1443 11883
rect 2697 11849 2731 11883
rect 5733 11849 5767 11883
rect 6929 11849 6963 11883
rect 14289 11849 14323 11883
rect 21373 11849 21407 11883
rect 15025 11781 15059 11815
rect 15393 11781 15427 11815
rect 16129 11781 16163 11815
rect 1593 11713 1627 11747
rect 1685 11713 1719 11747
rect 1959 11713 1993 11747
rect 3341 11713 3375 11747
rect 3615 11713 3649 11747
rect 4721 11713 4755 11747
rect 4995 11713 5029 11747
rect 6451 11713 6485 11747
rect 7113 11713 7147 11747
rect 7389 11713 7423 11747
rect 8585 11713 8619 11747
rect 10057 11713 10091 11747
rect 10315 11713 10349 11747
rect 13369 11713 13403 11747
rect 13507 11713 13541 11747
rect 13645 11713 13679 11747
rect 15301 11713 15335 11747
rect 15761 11713 15795 11747
rect 16957 11713 16991 11747
rect 17233 11713 17267 11747
rect 17500 11713 17534 11747
rect 19071 11723 19105 11757
rect 20545 11713 20579 11747
rect 21005 11713 21039 11747
rect 21557 11713 21591 11747
rect 7573 11645 7607 11679
rect 8309 11645 8343 11679
rect 8447 11645 8481 11679
rect 12449 11645 12483 11679
rect 12633 11645 12667 11679
rect 18797 11645 18831 11679
rect 20269 11645 20303 11679
rect 8033 11577 8067 11611
rect 13093 11577 13127 11611
rect 19809 11577 19843 11611
rect 21005 11577 21039 11611
rect 4353 11509 4387 11543
rect 6561 11509 6595 11543
rect 9229 11509 9263 11543
rect 11069 11509 11103 11543
rect 16313 11509 16347 11543
rect 17049 11509 17083 11543
rect 18613 11509 18647 11543
rect 3341 11305 3375 11339
rect 6745 11305 6779 11339
rect 7205 11305 7239 11339
rect 8953 11305 8987 11339
rect 13001 11305 13035 11339
rect 15117 11305 15151 11339
rect 16589 11305 16623 11339
rect 18705 11305 18739 11339
rect 19809 11305 19843 11339
rect 1869 11237 1903 11271
rect 8493 11237 8527 11271
rect 9873 11237 9907 11271
rect 11805 11237 11839 11271
rect 19441 11237 19475 11271
rect 2329 11169 2363 11203
rect 4905 11169 4939 11203
rect 5549 11169 5583 11203
rect 5825 11169 5859 11203
rect 5963 11169 5997 11203
rect 7481 11169 7515 11203
rect 10149 11169 10183 11203
rect 10287 11169 10321 11203
rect 11345 11169 11379 11203
rect 12081 11169 12115 11203
rect 14105 11169 14139 11203
rect 15577 11169 15611 11203
rect 17601 11169 17635 11203
rect 19993 11169 20027 11203
rect 1685 11101 1719 11135
rect 2587 11071 2621 11105
rect 4629 11101 4663 11135
rect 5089 11101 5123 11135
rect 6101 11101 6135 11135
rect 6929 11101 6963 11135
rect 7755 11101 7789 11135
rect 9137 11101 9171 11135
rect 9229 11101 9263 11135
rect 9413 11101 9447 11135
rect 10425 11101 10459 11135
rect 11161 11101 11195 11135
rect 12219 11101 12253 11135
rect 12357 11101 12391 11135
rect 14379 11101 14413 11135
rect 15819 11101 15853 11135
rect 17877 11101 17911 11135
rect 18337 11101 18371 11135
rect 18889 11101 18923 11135
rect 19625 11101 19659 11135
rect 19717 11101 19751 11135
rect 4261 11033 4295 11067
rect 11069 11033 11103 11067
rect 18613 11033 18647 11067
rect 20238 11033 20272 11067
rect 21373 10965 21407 10999
rect 6193 10761 6227 10795
rect 8309 10761 8343 10795
rect 9689 10761 9723 10795
rect 11069 10761 11103 10795
rect 20545 10761 20579 10795
rect 21465 10761 21499 10795
rect 1685 10693 1719 10727
rect 21189 10693 21223 10727
rect 2329 10625 2363 10659
rect 3525 10625 3559 10659
rect 4537 10625 4571 10659
rect 5390 10625 5424 10659
rect 5549 10625 5583 10659
rect 6653 10625 6687 10659
rect 7539 10625 7573 10659
rect 8951 10625 8985 10659
rect 10057 10625 10091 10659
rect 10331 10625 10365 10659
rect 12633 10625 12667 10659
rect 13553 10625 13587 10659
rect 13670 10625 13704 10659
rect 14565 10625 14599 10659
rect 14839 10625 14873 10659
rect 17567 10625 17601 10659
rect 19441 10625 19475 10659
rect 19775 10625 19809 10659
rect 2513 10557 2547 10591
rect 3249 10557 3283 10591
rect 3387 10557 3421 10591
rect 4353 10557 4387 10591
rect 5273 10557 5307 10591
rect 7297 10557 7331 10591
rect 8677 10557 8711 10591
rect 12817 10557 12851 10591
rect 13277 10557 13311 10591
rect 13829 10557 13863 10591
rect 17325 10557 17359 10591
rect 19533 10557 19567 10591
rect 2973 10489 3007 10523
rect 4997 10489 5031 10523
rect 1777 10421 1811 10455
rect 4169 10421 4203 10455
rect 6469 10421 6503 10455
rect 6929 10421 6963 10455
rect 14473 10421 14507 10455
rect 15577 10421 15611 10455
rect 18337 10421 18371 10455
rect 19257 10421 19291 10455
rect 1685 10217 1719 10251
rect 2145 10217 2179 10251
rect 3341 10217 3375 10251
rect 3985 10217 4019 10251
rect 4537 10217 4571 10251
rect 6101 10217 6135 10251
rect 10425 10217 10459 10251
rect 20913 10217 20947 10251
rect 8585 10149 8619 10183
rect 18153 10149 18187 10183
rect 2329 10081 2363 10115
rect 5089 10081 5123 10115
rect 6653 10081 6687 10115
rect 6837 10081 6871 10115
rect 7297 10081 7331 10115
rect 7573 10081 7607 10115
rect 7690 10081 7724 10115
rect 11897 10081 11931 10115
rect 12357 10081 12391 10115
rect 12633 10081 12667 10115
rect 12771 10081 12805 10115
rect 13553 10081 13587 10115
rect 1869 10013 1903 10047
rect 2603 10013 2637 10047
rect 5363 10013 5397 10047
rect 7849 10013 7883 10047
rect 8769 10013 8803 10047
rect 9413 10013 9447 10047
rect 9687 10013 9721 10047
rect 11713 10013 11747 10047
rect 12909 10013 12943 10047
rect 14933 10013 14967 10047
rect 16037 10013 16071 10047
rect 16311 10013 16345 10047
rect 17969 10013 18003 10047
rect 18153 10013 18187 10047
rect 18613 10013 18647 10047
rect 18797 10013 18831 10047
rect 19073 10013 19107 10047
rect 19257 10013 19291 10047
rect 19515 9983 19549 10017
rect 20729 10013 20763 10047
rect 3893 9945 3927 9979
rect 4445 9945 4479 9979
rect 14841 9945 14875 9979
rect 15301 9945 15335 9979
rect 18521 9945 18555 9979
rect 18705 9945 18739 9979
rect 21189 9945 21223 9979
rect 21557 9945 21591 9979
rect 8493 9877 8527 9911
rect 14565 9877 14599 9911
rect 15669 9877 15703 9911
rect 15853 9877 15887 9911
rect 17049 9877 17083 9911
rect 18889 9877 18923 9911
rect 20269 9877 20303 9911
rect 10609 9673 10643 9707
rect 19165 9673 19199 9707
rect 20545 9673 20579 9707
rect 1501 9605 1535 9639
rect 1869 9605 1903 9639
rect 13921 9605 13955 9639
rect 14841 9605 14875 9639
rect 15117 9605 15151 9639
rect 15945 9605 15979 9639
rect 2237 9537 2271 9571
rect 2605 9537 2639 9571
rect 3479 9537 3513 9571
rect 4261 9537 4295 9571
rect 5273 9537 5307 9571
rect 5411 9537 5445 9571
rect 6469 9537 6503 9571
rect 7113 9537 7147 9571
rect 7663 9537 7697 9571
rect 8953 9537 8987 9571
rect 9965 9537 9999 9571
rect 10885 9537 10919 9571
rect 12081 9537 12115 9571
rect 13277 9537 13311 9571
rect 15209 9537 15243 9571
rect 15577 9537 15611 9571
rect 17693 9537 17727 9571
rect 18052 9537 18086 9571
rect 19441 9537 19475 9571
rect 19533 9537 19567 9571
rect 19807 9537 19841 9571
rect 20913 9537 20947 9571
rect 21097 9537 21131 9571
rect 21465 9537 21499 9571
rect 2421 9469 2455 9503
rect 3341 9469 3375 9503
rect 3617 9469 3651 9503
rect 4353 9469 4387 9503
rect 4537 9469 4571 9503
rect 5549 9469 5583 9503
rect 7389 9469 7423 9503
rect 8769 9469 8803 9503
rect 9689 9469 9723 9503
rect 9827 9469 9861 9503
rect 12265 9469 12299 9503
rect 13001 9469 13035 9503
rect 13139 9469 13173 9503
rect 17785 9469 17819 9503
rect 3065 9401 3099 9435
rect 4997 9401 5031 9435
rect 6193 9401 6227 9435
rect 6929 9401 6963 9435
rect 8401 9401 8435 9435
rect 9413 9401 9447 9435
rect 12725 9401 12759 9435
rect 16129 9401 16163 9435
rect 21097 9401 21131 9435
rect 2053 9333 2087 9367
rect 6561 9333 6595 9367
rect 10701 9333 10735 9367
rect 17509 9333 17543 9367
rect 19257 9333 19291 9367
rect 1777 9129 1811 9163
rect 4813 9129 4847 9163
rect 8033 9129 8067 9163
rect 10057 9129 10091 9163
rect 11621 9129 11655 9163
rect 13001 9129 13035 9163
rect 15117 9129 15151 9163
rect 16497 9129 16531 9163
rect 18337 9129 18371 9163
rect 19441 9129 19475 9163
rect 21465 9129 21499 9163
rect 5181 9061 5215 9095
rect 18797 9061 18831 9095
rect 21005 9061 21039 9095
rect 2145 8993 2179 9027
rect 3801 8993 3835 9027
rect 5641 8993 5675 9027
rect 7021 8993 7055 9027
rect 9045 8993 9079 9027
rect 10609 8993 10643 9027
rect 11989 8993 12023 9027
rect 14105 8993 14139 9027
rect 15485 8993 15519 9027
rect 2387 8925 2421 8959
rect 4075 8925 4109 8959
rect 5365 8925 5399 8959
rect 5915 8925 5949 8959
rect 7295 8925 7329 8959
rect 8585 8925 8619 8959
rect 9319 8925 9353 8959
rect 10851 8915 10885 8949
rect 12263 8925 12297 8959
rect 14347 8925 14381 8959
rect 15759 8925 15793 8959
rect 16865 8925 16899 8959
rect 17123 8895 17157 8929
rect 18245 8925 18279 8959
rect 18521 8925 18555 8959
rect 18705 8925 18739 8959
rect 18981 8925 19015 8959
rect 19349 8915 19383 8949
rect 19533 8925 19567 8959
rect 19625 8925 19659 8959
rect 19899 8925 19933 8959
rect 21189 8925 21223 8959
rect 21281 8925 21315 8959
rect 1501 8857 1535 8891
rect 3157 8789 3191 8823
rect 6653 8789 6687 8823
rect 8401 8789 8435 8823
rect 17877 8789 17911 8823
rect 18613 8789 18647 8823
rect 20637 8789 20671 8823
rect 1777 8585 1811 8619
rect 4445 8585 4479 8619
rect 7481 8585 7515 8619
rect 11253 8585 11287 8619
rect 12541 8585 12575 8619
rect 13921 8585 13955 8619
rect 15301 8585 15335 8619
rect 18337 8585 18371 8619
rect 21373 8585 21407 8619
rect 1501 8449 1535 8483
rect 2513 8449 2547 8483
rect 3387 8449 3421 8483
rect 3525 8449 3559 8483
rect 4353 8449 4387 8483
rect 5055 8449 5089 8483
rect 6711 8449 6745 8483
rect 8033 8449 8067 8483
rect 8307 8449 8341 8483
rect 9413 8449 9447 8483
rect 10333 8449 10367 8483
rect 11529 8449 11563 8483
rect 11803 8449 11837 8483
rect 13183 8449 13217 8483
rect 14289 8449 14323 8483
rect 14531 8459 14565 8493
rect 16865 8449 16899 8483
rect 17224 8449 17258 8483
rect 18855 8449 18889 8483
rect 20235 8449 20269 8483
rect 21557 8449 21591 8483
rect 2329 8381 2363 8415
rect 3249 8381 3283 8415
rect 4813 8381 4847 8415
rect 6469 8381 6503 8415
rect 9597 8381 9631 8415
rect 10471 8381 10505 8415
rect 10609 8381 10643 8415
rect 12909 8381 12943 8415
rect 16957 8381 16991 8415
rect 18613 8381 18647 8415
rect 19993 8381 20027 8415
rect 2973 8313 3007 8347
rect 5825 8313 5859 8347
rect 9045 8313 9079 8347
rect 10057 8313 10091 8347
rect 19625 8313 19659 8347
rect 21005 8313 21039 8347
rect 4169 8245 4203 8279
rect 16681 8245 16715 8279
rect 3341 8041 3375 8075
rect 3893 8041 3927 8075
rect 5181 8041 5215 8075
rect 10609 8041 10643 8075
rect 21465 8041 21499 8075
rect 6837 7973 6871 8007
rect 8401 7973 8435 8007
rect 11805 7973 11839 8007
rect 15853 7973 15887 8007
rect 18797 7973 18831 8007
rect 2329 7905 2363 7939
rect 4169 7905 4203 7939
rect 6193 7905 6227 7939
rect 9597 7905 9631 7939
rect 11161 7905 11195 7939
rect 12081 7905 12115 7939
rect 12357 7905 12391 7939
rect 16313 7905 16347 7939
rect 19441 7905 19475 7939
rect 2603 7837 2637 7871
rect 4077 7837 4111 7871
rect 4411 7837 4445 7871
rect 6377 7837 6411 7871
rect 7113 7837 7147 7871
rect 7251 7837 7285 7871
rect 7389 7837 7423 7871
rect 8309 7837 8343 7871
rect 8585 7837 8619 7871
rect 9137 7837 9171 7871
rect 9871 7837 9905 7871
rect 11345 7837 11379 7871
rect 12198 7837 12232 7871
rect 13737 7837 13771 7871
rect 14105 7837 14139 7871
rect 14347 7837 14381 7871
rect 15669 7837 15703 7871
rect 15853 7837 15887 7871
rect 16555 7837 16589 7871
rect 17693 7837 17727 7871
rect 18153 7837 18187 7871
rect 18521 7837 18555 7871
rect 18889 7837 18923 7871
rect 21097 7837 21131 7871
rect 21373 7837 21407 7871
rect 1501 7769 1535 7803
rect 2145 7769 2179 7803
rect 5733 7769 5767 7803
rect 16221 7769 16255 7803
rect 19686 7769 19720 7803
rect 1777 7701 1811 7735
rect 5825 7701 5859 7735
rect 8033 7701 8067 7735
rect 8125 7701 8159 7735
rect 8953 7701 8987 7735
rect 13001 7701 13035 7735
rect 13921 7701 13955 7735
rect 15117 7701 15151 7735
rect 17325 7701 17359 7735
rect 17785 7701 17819 7735
rect 20821 7701 20855 7735
rect 20913 7701 20947 7735
rect 1869 7497 1903 7531
rect 3893 7497 3927 7531
rect 4445 7497 4479 7531
rect 5825 7497 5859 7531
rect 9413 7497 9447 7531
rect 12541 7497 12575 7531
rect 16129 7497 16163 7531
rect 17969 7497 18003 7531
rect 1593 7429 1627 7463
rect 7021 7429 7055 7463
rect 14841 7429 14875 7463
rect 14933 7429 14967 7463
rect 15117 7429 15151 7463
rect 2053 7361 2087 7395
rect 3249 7361 3283 7395
rect 4169 7361 4203 7395
rect 4353 7361 4387 7395
rect 5087 7361 5121 7395
rect 6469 7361 6503 7395
rect 8769 7361 8803 7395
rect 10425 7361 10459 7395
rect 10542 7361 10576 7395
rect 11529 7361 11563 7395
rect 11803 7361 11837 7395
rect 14565 7361 14599 7395
rect 14749 7361 14783 7395
rect 15025 7361 15059 7395
rect 15209 7361 15243 7395
rect 16027 7361 16061 7395
rect 16221 7361 16255 7395
rect 16497 7361 16531 7395
rect 16865 7361 16899 7395
rect 17233 7361 17267 7395
rect 17601 7361 17635 7395
rect 17877 7361 17911 7395
rect 18337 7361 18371 7395
rect 18887 7361 18921 7395
rect 19993 7361 20027 7395
rect 20249 7361 20283 7395
rect 2237 7293 2271 7327
rect 2973 7293 3007 7327
rect 3111 7293 3145 7327
rect 4813 7293 4847 7327
rect 7573 7293 7607 7327
rect 7757 7293 7791 7327
rect 8493 7293 8527 7327
rect 8631 7293 8665 7327
rect 9505 7293 9539 7327
rect 9689 7293 9723 7327
rect 10701 7293 10735 7327
rect 18613 7293 18647 7327
rect 2697 7225 2731 7259
rect 3985 7225 4019 7259
rect 8217 7225 8251 7259
rect 10149 7225 10183 7259
rect 16313 7225 16347 7259
rect 17509 7225 17543 7259
rect 18153 7225 18187 7259
rect 6561 7157 6595 7191
rect 7113 7157 7147 7191
rect 11345 7157 11379 7191
rect 19625 7157 19659 7191
rect 21373 7157 21407 7191
rect 7113 6953 7147 6987
rect 8493 6953 8527 6987
rect 10609 6953 10643 6987
rect 11989 6953 12023 6987
rect 13829 6953 13863 6987
rect 15485 6953 15519 6987
rect 17969 6953 18003 6987
rect 18705 6953 18739 6987
rect 4077 6885 4111 6919
rect 6009 6885 6043 6919
rect 18889 6885 18923 6919
rect 20545 6885 20579 6919
rect 4813 6817 4847 6851
rect 5089 6817 5123 6851
rect 5227 6817 5261 6851
rect 7481 6817 7515 6851
rect 9597 6817 9631 6851
rect 10977 6817 11011 6851
rect 19533 6817 19567 6851
rect 21005 6817 21039 6851
rect 2329 6749 2363 6783
rect 2603 6749 2637 6783
rect 4169 6749 4203 6783
rect 4353 6749 4387 6783
rect 5365 6749 5399 6783
rect 6101 6749 6135 6783
rect 6375 6749 6409 6783
rect 7755 6749 7789 6783
rect 9871 6749 9905 6783
rect 11251 6749 11285 6783
rect 13737 6749 13771 6783
rect 14105 6749 14139 6783
rect 14347 6749 14381 6783
rect 15669 6749 15703 6783
rect 16589 6749 16623 6783
rect 18245 6749 18279 6783
rect 18337 6749 18371 6783
rect 18613 6749 18647 6783
rect 19073 6749 19107 6783
rect 19441 6749 19475 6783
rect 19717 6749 19751 6783
rect 20085 6749 20119 6783
rect 20637 6749 20671 6783
rect 20913 6749 20947 6783
rect 21097 6749 21131 6783
rect 21373 6749 21407 6783
rect 1501 6681 1535 6715
rect 3893 6681 3927 6715
rect 16834 6681 16868 6715
rect 1777 6613 1811 6647
rect 3341 6613 3375 6647
rect 15117 6613 15151 6647
rect 18061 6613 18095 6647
rect 18521 6613 18555 6647
rect 21189 6613 21223 6647
rect 2513 6409 2547 6443
rect 3433 6409 3467 6443
rect 3985 6409 4019 6443
rect 5365 6409 5399 6443
rect 10333 6409 10367 6443
rect 14013 6409 14047 6443
rect 15669 6409 15703 6443
rect 18153 6409 18187 6443
rect 21281 6409 21315 6443
rect 21373 6409 21407 6443
rect 5825 6341 5859 6375
rect 6561 6341 6595 6375
rect 7665 6341 7699 6375
rect 17785 6341 17819 6375
rect 20168 6341 20202 6375
rect 1501 6273 1535 6307
rect 1759 6303 1793 6337
rect 3157 6273 3191 6307
rect 3617 6273 3651 6307
rect 3893 6273 3927 6307
rect 4353 6273 4387 6307
rect 4627 6273 4661 6307
rect 6837 6273 6871 6307
rect 6929 6273 6963 6307
rect 7297 6273 7331 6307
rect 9321 6273 9355 6307
rect 9579 6303 9613 6337
rect 10885 6273 10919 6307
rect 11161 6273 11195 6307
rect 11621 6273 11655 6307
rect 14197 6273 14231 6307
rect 14556 6273 14590 6307
rect 15761 6273 15795 6307
rect 15945 6273 15979 6307
rect 17049 6273 17083 6307
rect 17509 6273 17543 6307
rect 17969 6273 18003 6307
rect 18153 6273 18187 6307
rect 18429 6273 18463 6307
rect 18795 6273 18829 6307
rect 19901 6273 19935 6307
rect 21557 6273 21591 6307
rect 14289 6205 14323 6239
rect 16865 6205 16899 6239
rect 18521 6205 18555 6239
rect 7849 6137 7883 6171
rect 5917 6069 5951 6103
rect 10701 6069 10735 6103
rect 10977 6069 11011 6103
rect 11805 6069 11839 6103
rect 15853 6069 15887 6103
rect 18245 6069 18279 6103
rect 19533 6069 19567 6103
rect 1501 5865 1535 5899
rect 6193 5865 6227 5899
rect 7573 5865 7607 5899
rect 15393 5865 15427 5899
rect 15577 5865 15611 5899
rect 15945 5865 15979 5899
rect 17141 5865 17175 5899
rect 21373 5865 21407 5899
rect 4721 5797 4755 5831
rect 14473 5797 14507 5831
rect 18337 5797 18371 5831
rect 19073 5797 19107 5831
rect 1777 5729 1811 5763
rect 2421 5729 2455 5763
rect 2697 5729 2731 5763
rect 2835 5729 2869 5763
rect 4077 5729 4111 5763
rect 5135 5729 5169 5763
rect 6561 5729 6595 5763
rect 13829 5729 13863 5763
rect 14657 5729 14691 5763
rect 16129 5729 16163 5763
rect 17601 5729 17635 5763
rect 19257 5729 19291 5763
rect 1685 5661 1719 5695
rect 1961 5661 1995 5695
rect 2973 5661 3007 5695
rect 3985 5661 4019 5695
rect 4261 5661 4295 5695
rect 4997 5661 5031 5695
rect 5273 5661 5307 5695
rect 5917 5661 5951 5695
rect 6803 5661 6837 5695
rect 8125 5661 8159 5695
rect 10609 5661 10643 5695
rect 13737 5661 13771 5695
rect 14473 5661 14507 5695
rect 14841 5661 14875 5695
rect 14933 5661 14967 5695
rect 15117 5661 15151 5695
rect 15761 5661 15795 5695
rect 15853 5661 15887 5695
rect 16371 5661 16405 5695
rect 17877 5661 17911 5695
rect 18337 5661 18371 5695
rect 18889 5661 18923 5695
rect 19499 5661 19533 5695
rect 20637 5661 20671 5695
rect 20821 5661 20855 5695
rect 21097 5661 21131 5695
rect 21557 5661 21591 5695
rect 6101 5593 6135 5627
rect 15485 5593 15519 5627
rect 3617 5525 3651 5559
rect 3801 5525 3835 5559
rect 7941 5525 7975 5559
rect 10425 5525 10459 5559
rect 20269 5525 20303 5559
rect 20821 5525 20855 5559
rect 20913 5525 20947 5559
rect 1777 5321 1811 5355
rect 3157 5321 3191 5355
rect 4537 5321 4571 5355
rect 13921 5321 13955 5355
rect 15669 5321 15703 5355
rect 16405 5321 16439 5355
rect 19165 5321 19199 5355
rect 1501 5253 1535 5287
rect 21465 5253 21499 5287
rect 2419 5185 2453 5219
rect 3525 5185 3559 5219
rect 3799 5185 3833 5219
rect 5179 5185 5213 5219
rect 13183 5185 13217 5219
rect 14289 5185 14323 5219
rect 14556 5185 14590 5219
rect 15945 5185 15979 5219
rect 16037 5185 16071 5219
rect 16313 5185 16347 5219
rect 16497 5185 16531 5219
rect 16937 5185 16971 5219
rect 18411 5215 18445 5249
rect 19807 5185 19841 5219
rect 20913 5185 20947 5219
rect 21097 5185 21131 5219
rect 21373 5185 21407 5219
rect 2145 5117 2179 5151
rect 4905 5117 4939 5151
rect 12909 5117 12943 5151
rect 16129 5117 16163 5151
rect 16681 5117 16715 5151
rect 18153 5117 18187 5151
rect 19533 5117 19567 5151
rect 5917 5049 5951 5083
rect 15761 4981 15795 5015
rect 18061 4981 18095 5015
rect 20545 4981 20579 5015
rect 2145 4777 2179 4811
rect 3341 4777 3375 4811
rect 4905 4777 4939 4811
rect 6285 4777 6319 4811
rect 15669 4777 15703 4811
rect 16405 4777 16439 4811
rect 16957 4777 16991 4811
rect 15577 4709 15611 4743
rect 16221 4709 16255 4743
rect 16589 4709 16623 4743
rect 19257 4709 19291 4743
rect 2329 4641 2363 4675
rect 3893 4641 3927 4675
rect 17141 4641 17175 4675
rect 19993 4641 20027 4675
rect 1593 4573 1627 4607
rect 1869 4573 1903 4607
rect 2603 4573 2637 4607
rect 4167 4573 4201 4607
rect 5273 4573 5307 4607
rect 5547 4573 5581 4607
rect 14197 4573 14231 4607
rect 14453 4573 14487 4607
rect 15853 4573 15887 4607
rect 16037 4573 16071 4607
rect 16313 4573 16347 4607
rect 16497 4573 16531 4607
rect 16773 4573 16807 4607
rect 16865 4573 16899 4607
rect 17049 4573 17083 4607
rect 18797 4573 18831 4607
rect 18889 4573 18923 4607
rect 19073 4573 19107 4607
rect 19441 4573 19475 4607
rect 19533 4573 19567 4607
rect 20249 4573 20283 4607
rect 17408 4505 17442 4539
rect 18981 4505 19015 4539
rect 1409 4437 1443 4471
rect 18521 4437 18555 4471
rect 18613 4437 18647 4471
rect 19625 4437 19659 4471
rect 21373 4437 21407 4471
rect 2605 4233 2639 4267
rect 14473 4233 14507 4267
rect 14933 4233 14967 4267
rect 15301 4233 15335 4267
rect 19165 4233 19199 4267
rect 21097 4233 21131 4267
rect 19892 4165 19926 4199
rect 1867 4097 1901 4131
rect 2973 4097 3007 4131
rect 3247 4097 3281 4131
rect 4595 4097 4629 4131
rect 5917 4097 5951 4131
rect 14381 4097 14415 4131
rect 14657 4097 14691 4131
rect 15117 4097 15151 4131
rect 15209 4097 15243 4131
rect 15485 4097 15519 4131
rect 15577 4097 15611 4131
rect 15945 4097 15979 4131
rect 16221 4097 16255 4131
rect 16497 4097 16531 4131
rect 17049 4097 17083 4131
rect 17325 4097 17359 4131
rect 17877 4097 17911 4131
rect 18429 4097 18463 4131
rect 18705 4097 18739 4131
rect 18889 4097 18923 4131
rect 18981 4097 19015 4131
rect 19441 4097 19475 4131
rect 21281 4097 21315 4131
rect 21557 4097 21591 4131
rect 1593 4029 1627 4063
rect 4353 4029 4387 4063
rect 17693 4029 17727 4063
rect 18797 4029 18831 4063
rect 19625 4029 19659 4063
rect 14197 3961 14231 3995
rect 16037 3961 16071 3995
rect 17141 3961 17175 3995
rect 18337 3961 18371 3995
rect 19257 3961 19291 3995
rect 3985 3893 4019 3927
rect 5365 3893 5399 3927
rect 5733 3893 5767 3927
rect 15761 3893 15795 3927
rect 16313 3893 16347 3927
rect 16865 3893 16899 3927
rect 21005 3893 21039 3927
rect 21373 3893 21407 3927
rect 2605 3689 2639 3723
rect 3341 3689 3375 3723
rect 5549 3689 5583 3723
rect 5733 3689 5767 3723
rect 8953 3689 8987 3723
rect 14657 3689 14691 3723
rect 17693 3689 17727 3723
rect 18429 3689 18463 3723
rect 20637 3689 20671 3723
rect 4813 3621 4847 3655
rect 13369 3621 13403 3655
rect 14289 3621 14323 3655
rect 14381 3621 14415 3655
rect 16773 3621 16807 3655
rect 18889 3621 18923 3655
rect 21373 3621 21407 3655
rect 1593 3553 1627 3587
rect 3801 3553 3835 3587
rect 21005 3553 21039 3587
rect 1835 3485 1869 3519
rect 4059 3455 4093 3489
rect 5273 3485 5307 3519
rect 5917 3485 5951 3519
rect 7665 3485 7699 3519
rect 8033 3485 8067 3519
rect 8493 3485 8527 3519
rect 8769 3485 8803 3519
rect 9137 3485 9171 3519
rect 9413 3485 9447 3519
rect 9689 3485 9723 3519
rect 10057 3485 10091 3519
rect 13093 3485 13127 3519
rect 13553 3485 13587 3519
rect 13921 3485 13955 3519
rect 14105 3485 14139 3519
rect 14565 3485 14599 3519
rect 14841 3485 14875 3519
rect 15117 3485 15151 3519
rect 15393 3485 15427 3519
rect 15669 3485 15703 3519
rect 16681 3485 16715 3519
rect 16957 3485 16991 3519
rect 17233 3485 17267 3519
rect 17509 3485 17543 3519
rect 17601 3485 17635 3519
rect 18061 3485 18095 3519
rect 18337 3485 18371 3519
rect 18613 3485 18647 3519
rect 18705 3485 18739 3519
rect 19257 3485 19291 3519
rect 20821 3485 20855 3519
rect 3249 3417 3283 3451
rect 16037 3417 16071 3451
rect 19502 3417 19536 3451
rect 21189 3417 21223 3451
rect 7481 3349 7515 3383
rect 7849 3349 7883 3383
rect 8309 3349 8343 3383
rect 8585 3349 8619 3383
rect 9229 3349 9263 3383
rect 9873 3349 9907 3383
rect 12909 3349 12943 3383
rect 13737 3349 13771 3383
rect 14933 3349 14967 3383
rect 15209 3349 15243 3383
rect 15485 3349 15519 3383
rect 16129 3349 16163 3383
rect 16497 3349 16531 3383
rect 17049 3349 17083 3383
rect 17325 3349 17359 3383
rect 17877 3349 17911 3383
rect 18153 3349 18187 3383
rect 2697 3145 2731 3179
rect 4997 3145 5031 3179
rect 5273 3145 5307 3179
rect 6561 3145 6595 3179
rect 7113 3145 7147 3179
rect 11529 3145 11563 3179
rect 13277 3145 13311 3179
rect 13737 3145 13771 3179
rect 14105 3145 14139 3179
rect 14657 3145 14691 3179
rect 16129 3145 16163 3179
rect 18061 3145 18095 3179
rect 18521 3145 18555 3179
rect 20085 3145 20119 3179
rect 20453 3145 20487 3179
rect 20821 3145 20855 3179
rect 4537 3077 4571 3111
rect 15669 3077 15703 3111
rect 17325 3077 17359 3111
rect 19993 3077 20027 3111
rect 1685 3009 1719 3043
rect 1943 3039 1977 3073
rect 3065 3009 3099 3043
rect 3323 3039 3357 3073
rect 5181 3009 5215 3043
rect 5457 3009 5491 3043
rect 6745 3009 6779 3043
rect 7021 3009 7055 3043
rect 7297 3009 7331 3043
rect 7573 3009 7607 3043
rect 7849 3009 7883 3043
rect 8125 3009 8159 3043
rect 8401 3009 8435 3043
rect 8677 3009 8711 3043
rect 8953 3009 8987 3043
rect 9229 3009 9263 3043
rect 9505 3009 9539 3043
rect 9597 3009 9631 3043
rect 10241 3009 10275 3043
rect 10701 3009 10735 3043
rect 11069 3009 11103 3043
rect 11713 3009 11747 3043
rect 12541 3009 12575 3043
rect 12817 3009 12851 3043
rect 13553 3009 13587 3043
rect 14013 3009 14047 3043
rect 14289 3009 14323 3043
rect 14565 3009 14599 3043
rect 14841 3009 14875 3043
rect 15117 3009 15151 3043
rect 15393 3009 15427 3043
rect 16313 3009 16347 3043
rect 16773 3009 16807 3043
rect 17969 3009 18003 3043
rect 18245 3009 18279 3043
rect 18429 3009 18463 3043
rect 18889 3009 18923 3043
rect 19165 3009 19199 3043
rect 19533 3009 19567 3043
rect 20361 3009 20395 3043
rect 20729 3009 20763 3043
rect 21097 3009 21131 3043
rect 21557 3009 21591 3043
rect 9321 2873 9355 2907
rect 9781 2873 9815 2907
rect 16957 2873 16991 2907
rect 19533 2873 19567 2907
rect 21281 2873 21315 2907
rect 4077 2805 4111 2839
rect 4629 2805 4663 2839
rect 6837 2805 6871 2839
rect 7389 2805 7423 2839
rect 7665 2805 7699 2839
rect 7941 2805 7975 2839
rect 8217 2805 8251 2839
rect 8493 2805 8527 2839
rect 8769 2805 8803 2839
rect 9045 2805 9079 2839
rect 10057 2805 10091 2839
rect 10517 2805 10551 2839
rect 11253 2805 11287 2839
rect 12357 2805 12391 2839
rect 12633 2805 12667 2839
rect 13829 2805 13863 2839
rect 14381 2805 14415 2839
rect 14933 2805 14967 2839
rect 15209 2805 15243 2839
rect 15761 2805 15795 2839
rect 17417 2805 17451 2839
rect 17785 2805 17819 2839
rect 21373 2805 21407 2839
rect 2329 2601 2363 2635
rect 3341 2601 3375 2635
rect 4169 2601 4203 2635
rect 4537 2601 4571 2635
rect 5181 2601 5215 2635
rect 5457 2601 5491 2635
rect 7573 2601 7607 2635
rect 7941 2601 7975 2635
rect 8677 2601 8711 2635
rect 10793 2601 10827 2635
rect 12541 2601 12575 2635
rect 12909 2601 12943 2635
rect 14473 2601 14507 2635
rect 15577 2601 15611 2635
rect 16681 2601 16715 2635
rect 18981 2601 19015 2635
rect 9321 2533 9355 2567
rect 2881 2465 2915 2499
rect 8401 2465 8435 2499
rect 11253 2465 11287 2499
rect 17601 2465 17635 2499
rect 20085 2465 20119 2499
rect 21189 2465 21223 2499
rect 1685 2397 1719 2431
rect 2053 2397 2087 2431
rect 2605 2397 2639 2431
rect 3893 2397 3927 2431
rect 4353 2397 4387 2431
rect 4905 2397 4939 2431
rect 4997 2397 5031 2431
rect 5641 2397 5675 2431
rect 6929 2397 6963 2431
rect 7481 2397 7515 2431
rect 7757 2397 7791 2431
rect 8217 2397 8251 2431
rect 8493 2397 8527 2431
rect 9689 2397 9723 2431
rect 10149 2397 10183 2431
rect 10425 2397 10459 2431
rect 10701 2397 10735 2431
rect 10977 2397 11011 2431
rect 11621 2397 11655 2431
rect 11897 2397 11931 2431
rect 12265 2397 12299 2431
rect 13369 2397 13403 2431
rect 13829 2397 13863 2431
rect 14657 2397 14691 2431
rect 14841 2397 14875 2431
rect 16019 2397 16053 2431
rect 16589 2397 16623 2431
rect 17233 2397 17267 2431
rect 18521 2397 18555 2431
rect 18889 2397 18923 2431
rect 19257 2397 19291 2431
rect 20361 2397 20395 2431
rect 3249 2329 3283 2363
rect 6101 2329 6135 2363
rect 6285 2329 6319 2363
rect 6469 2329 6503 2363
rect 6653 2329 6687 2363
rect 14289 2329 14323 2363
rect 15485 2329 15519 2363
rect 4721 2261 4755 2295
rect 7021 2261 7055 2295
rect 9965 2261 9999 2295
rect 10241 2261 10275 2295
rect 10517 2261 10551 2295
rect 11437 2261 11471 2295
rect 11713 2261 11747 2295
rect 12081 2261 12115 2295
rect 13645 2261 13679 2295
rect 15025 2261 15059 2295
rect 16129 2261 16163 2295
rect 18337 2261 18371 2295
rect 1593 2057 1627 2091
rect 2881 2057 2915 2091
rect 3433 2057 3467 2091
rect 4353 2057 4387 2091
rect 4721 2057 4755 2091
rect 6837 2057 6871 2091
rect 8677 2057 8711 2091
rect 13001 2057 13035 2091
rect 20913 2057 20947 2091
rect 21281 2057 21315 2091
rect 1501 1989 1535 2023
rect 2053 1989 2087 2023
rect 2421 1989 2455 2023
rect 7113 1989 7147 2023
rect 7481 1989 7515 2023
rect 7849 1989 7883 2023
rect 8217 1989 8251 2023
rect 9321 1989 9355 2023
rect 10425 1989 10459 2023
rect 10977 1989 11011 2023
rect 11621 1989 11655 2023
rect 13829 1989 13863 2023
rect 14381 1989 14415 2023
rect 15485 1989 15519 2023
rect 16037 1989 16071 2023
rect 20453 1989 20487 2023
rect 20821 1989 20855 2023
rect 2605 1921 2639 1955
rect 3249 1921 3283 1955
rect 3709 1921 3743 1955
rect 4169 1921 4203 1955
rect 4629 1921 4663 1955
rect 4905 1921 4939 1955
rect 5549 1921 5583 1955
rect 6653 1921 6687 1955
rect 8493 1921 8527 1955
rect 8861 1921 8895 1955
rect 9873 1921 9907 1955
rect 12173 1921 12207 1955
rect 12817 1921 12851 1955
rect 13277 1921 13311 1955
rect 14933 1921 14967 1955
rect 16681 1921 16715 1955
rect 17785 1921 17819 1955
rect 19625 1921 19659 1955
rect 21189 1921 21223 1955
rect 5273 1853 5307 1887
rect 7665 1853 7699 1887
rect 17049 1853 17083 1887
rect 19533 1853 19567 1887
rect 3985 1785 4019 1819
rect 5089 1785 5123 1819
rect 9045 1785 9079 1819
rect 7205 1717 7239 1751
rect 7941 1717 7975 1751
rect 8309 1717 8343 1751
rect 9597 1717 9631 1751
rect 10149 1717 10183 1751
rect 10517 1717 10551 1751
rect 11069 1717 11103 1751
rect 11713 1717 11747 1751
rect 12265 1717 12299 1751
rect 13369 1717 13403 1751
rect 13921 1717 13955 1751
rect 14473 1717 14507 1751
rect 15025 1717 15059 1751
rect 15577 1717 15611 1751
rect 16129 1717 16163 1751
rect 1593 1513 1627 1547
rect 5365 1513 5399 1547
rect 6101 1513 6135 1547
rect 6653 1513 6687 1547
rect 8033 1513 8067 1547
rect 12449 1513 12483 1547
rect 14289 1513 14323 1547
rect 14841 1513 14875 1547
rect 15209 1513 15243 1547
rect 16865 1513 16899 1547
rect 18797 1513 18831 1547
rect 9689 1445 9723 1479
rect 4353 1377 4387 1411
rect 8677 1377 8711 1411
rect 10241 1377 10275 1411
rect 11069 1377 11103 1411
rect 15853 1377 15887 1411
rect 2881 1309 2915 1343
rect 4445 1309 4479 1343
rect 5089 1309 5123 1343
rect 5181 1309 5215 1343
rect 5825 1309 5859 1343
rect 7113 1309 7147 1343
rect 7389 1309 7423 1343
rect 8217 1309 8251 1343
rect 8953 1309 8987 1343
rect 9413 1309 9447 1343
rect 9965 1309 9999 1343
rect 10793 1309 10827 1343
rect 11529 1309 11563 1343
rect 11897 1309 11931 1343
rect 12817 1309 12851 1343
rect 13185 1309 13219 1343
rect 13553 1309 13587 1343
rect 14197 1309 14231 1343
rect 14749 1309 14783 1343
rect 15393 1309 15427 1343
rect 15669 1309 15703 1343
rect 16773 1309 16807 1343
rect 19349 1309 19383 1343
rect 20361 1309 20395 1343
rect 21189 1309 21223 1343
rect 1501 1241 1535 1275
rect 2329 1241 2363 1275
rect 2697 1241 2731 1275
rect 3065 1241 3099 1275
rect 3249 1241 3283 1275
rect 3433 1241 3467 1275
rect 4169 1241 4203 1275
rect 4905 1241 4939 1275
rect 5641 1241 5675 1275
rect 6009 1241 6043 1275
rect 6561 1241 6595 1275
rect 8401 1241 8435 1275
rect 12357 1241 12391 1275
rect 17325 1241 17359 1275
rect 20085 1241 20119 1275
rect 2421 1173 2455 1207
rect 3525 1173 3559 1207
rect 4629 1173 4663 1207
rect 9137 1173 9171 1207
rect 11713 1173 11747 1207
rect 12081 1173 12115 1207
rect 13001 1173 13035 1207
rect 13369 1173 13403 1207
rect 13737 1173 13771 1207
<< metal1 >>
rect 13354 43868 13360 43920
rect 13412 43908 13418 43920
rect 15194 43908 15200 43920
rect 13412 43880 15200 43908
rect 13412 43868 13418 43880
rect 15194 43868 15200 43880
rect 15252 43868 15258 43920
rect 16942 43868 16948 43920
rect 17000 43908 17006 43920
rect 17402 43908 17408 43920
rect 17000 43880 17408 43908
rect 17000 43868 17006 43880
rect 17402 43868 17408 43880
rect 17460 43868 17466 43920
rect 5074 43800 5080 43852
rect 5132 43840 5138 43852
rect 6270 43840 6276 43852
rect 5132 43812 6276 43840
rect 5132 43800 5138 43812
rect 6270 43800 6276 43812
rect 6328 43800 6334 43852
rect 16758 43800 16764 43852
rect 16816 43840 16822 43852
rect 17770 43840 17776 43852
rect 16816 43812 17776 43840
rect 16816 43800 16822 43812
rect 17770 43800 17776 43812
rect 17828 43800 17834 43852
rect 1394 43732 1400 43784
rect 1452 43772 1458 43784
rect 1452 43744 2774 43772
rect 1452 43732 1458 43744
rect 2746 43636 2774 43744
rect 12158 43732 12164 43784
rect 12216 43772 12222 43784
rect 12342 43772 12348 43784
rect 12216 43744 12348 43772
rect 12216 43732 12222 43744
rect 12342 43732 12348 43744
rect 12400 43732 12406 43784
rect 12434 43636 12440 43648
rect 2746 43608 12440 43636
rect 12434 43596 12440 43608
rect 12492 43596 12498 43648
rect 18966 43596 18972 43648
rect 19024 43636 19030 43648
rect 20806 43636 20812 43648
rect 19024 43608 20812 43636
rect 19024 43596 19030 43608
rect 20806 43596 20812 43608
rect 20864 43596 20870 43648
rect 1104 43546 22056 43568
rect 1104 43494 6148 43546
rect 6200 43494 6212 43546
rect 6264 43494 6276 43546
rect 6328 43494 6340 43546
rect 6392 43494 6404 43546
rect 6456 43494 11346 43546
rect 11398 43494 11410 43546
rect 11462 43494 11474 43546
rect 11526 43494 11538 43546
rect 11590 43494 11602 43546
rect 11654 43494 16544 43546
rect 16596 43494 16608 43546
rect 16660 43494 16672 43546
rect 16724 43494 16736 43546
rect 16788 43494 16800 43546
rect 16852 43494 21742 43546
rect 21794 43494 21806 43546
rect 21858 43494 21870 43546
rect 21922 43494 21934 43546
rect 21986 43494 21998 43546
rect 22050 43494 22056 43546
rect 1104 43472 22056 43494
rect 2222 43392 2228 43444
rect 2280 43392 2286 43444
rect 3142 43392 3148 43444
rect 3200 43392 3206 43444
rect 3326 43392 3332 43444
rect 3384 43392 3390 43444
rect 3973 43435 4031 43441
rect 3973 43401 3985 43435
rect 4019 43432 4031 43435
rect 5166 43432 5172 43444
rect 4019 43404 5172 43432
rect 4019 43401 4031 43404
rect 3973 43395 4031 43401
rect 5166 43392 5172 43404
rect 5224 43392 5230 43444
rect 5258 43392 5264 43444
rect 5316 43392 5322 43444
rect 5442 43392 5448 43444
rect 5500 43392 5506 43444
rect 5810 43392 5816 43444
rect 5868 43392 5874 43444
rect 6825 43435 6883 43441
rect 6825 43401 6837 43435
rect 6871 43432 6883 43435
rect 7374 43432 7380 43444
rect 6871 43404 7380 43432
rect 6871 43401 6883 43404
rect 6825 43395 6883 43401
rect 7374 43392 7380 43404
rect 7432 43392 7438 43444
rect 8297 43435 8355 43441
rect 8297 43401 8309 43435
rect 8343 43432 8355 43435
rect 8570 43432 8576 43444
rect 8343 43404 8576 43432
rect 8343 43401 8355 43404
rect 8297 43395 8355 43401
rect 8570 43392 8576 43404
rect 8628 43392 8634 43444
rect 8665 43435 8723 43441
rect 8665 43401 8677 43435
rect 8711 43432 8723 43435
rect 9030 43432 9036 43444
rect 8711 43404 9036 43432
rect 8711 43401 8723 43404
rect 8665 43395 8723 43401
rect 9030 43392 9036 43404
rect 9088 43392 9094 43444
rect 9125 43435 9183 43441
rect 9125 43401 9137 43435
rect 9171 43432 9183 43435
rect 9398 43432 9404 43444
rect 9171 43404 9404 43432
rect 9171 43401 9183 43404
rect 9125 43395 9183 43401
rect 9398 43392 9404 43404
rect 9456 43392 9462 43444
rect 10042 43392 10048 43444
rect 10100 43432 10106 43444
rect 12161 43435 12219 43441
rect 12161 43432 12173 43435
rect 10100 43404 12173 43432
rect 10100 43392 10106 43404
rect 12161 43401 12173 43404
rect 12207 43401 12219 43435
rect 12161 43395 12219 43401
rect 12434 43392 12440 43444
rect 12492 43392 12498 43444
rect 13722 43392 13728 43444
rect 13780 43432 13786 43444
rect 13780 43404 13860 43432
rect 13780 43392 13786 43404
rect 2869 43367 2927 43373
rect 2869 43333 2881 43367
rect 2915 43364 2927 43367
rect 3344 43364 3372 43392
rect 2915 43336 3372 43364
rect 4985 43367 5043 43373
rect 2915 43333 2927 43336
rect 2869 43327 2927 43333
rect 4985 43333 4997 43367
rect 5031 43364 5043 43367
rect 5460 43364 5488 43392
rect 5031 43336 5488 43364
rect 7837 43367 7895 43373
rect 5031 43333 5043 43336
rect 4985 43327 5043 43333
rect 7837 43333 7849 43367
rect 7883 43364 7895 43367
rect 8386 43364 8392 43376
rect 7883 43336 8392 43364
rect 7883 43333 7895 43336
rect 7837 43327 7895 43333
rect 8386 43324 8392 43336
rect 8444 43324 8450 43376
rect 9766 43324 9772 43376
rect 9824 43324 9830 43376
rect 10318 43324 10324 43376
rect 10376 43324 10382 43376
rect 10870 43324 10876 43376
rect 10928 43324 10934 43376
rect 12342 43324 12348 43376
rect 12400 43324 12406 43376
rect 12894 43324 12900 43376
rect 12952 43324 12958 43376
rect 13078 43324 13084 43376
rect 13136 43364 13142 43376
rect 13832 43364 13860 43404
rect 13906 43392 13912 43444
rect 13964 43392 13970 43444
rect 14274 43392 14280 43444
rect 14332 43432 14338 43444
rect 14332 43404 16436 43432
rect 14332 43392 14338 43404
rect 13136 43336 13768 43364
rect 13832 43336 14504 43364
rect 13136 43324 13142 43336
rect 1949 43299 2007 43305
rect 1949 43265 1961 43299
rect 1995 43265 2007 43299
rect 1949 43259 2007 43265
rect 1964 43228 1992 43259
rect 2038 43256 2044 43308
rect 2096 43256 2102 43308
rect 2498 43256 2504 43308
rect 2556 43256 2562 43308
rect 3050 43256 3056 43308
rect 3108 43256 3114 43308
rect 3789 43299 3847 43305
rect 3789 43265 3801 43299
rect 3835 43296 3847 43299
rect 3970 43296 3976 43308
rect 3835 43268 3976 43296
rect 3835 43265 3847 43268
rect 3789 43259 3847 43265
rect 3970 43256 3976 43268
rect 4028 43256 4034 43308
rect 4157 43299 4215 43305
rect 4157 43265 4169 43299
rect 4203 43296 4215 43299
rect 4338 43296 4344 43308
rect 4203 43268 4344 43296
rect 4203 43265 4215 43268
rect 4157 43259 4215 43265
rect 4338 43256 4344 43268
rect 4396 43256 4402 43308
rect 4617 43299 4675 43305
rect 4617 43265 4629 43299
rect 4663 43265 4675 43299
rect 4617 43259 4675 43265
rect 2590 43228 2596 43240
rect 1964 43200 2596 43228
rect 2590 43188 2596 43200
rect 2648 43188 2654 43240
rect 1765 43163 1823 43169
rect 1765 43129 1777 43163
rect 1811 43160 1823 43163
rect 2958 43160 2964 43172
rect 1811 43132 2964 43160
rect 1811 43129 1823 43132
rect 1765 43123 1823 43129
rect 2958 43120 2964 43132
rect 3016 43120 3022 43172
rect 4154 43120 4160 43172
rect 4212 43160 4218 43172
rect 4632 43160 4660 43259
rect 4706 43256 4712 43308
rect 4764 43296 4770 43308
rect 5169 43299 5227 43305
rect 5169 43296 5181 43299
rect 4764 43268 5181 43296
rect 4764 43256 4770 43268
rect 5169 43265 5181 43268
rect 5215 43265 5227 43299
rect 5169 43259 5227 43265
rect 5534 43256 5540 43308
rect 5592 43296 5598 43308
rect 5721 43299 5779 43305
rect 5721 43296 5733 43299
rect 5592 43268 5733 43296
rect 5592 43256 5598 43268
rect 5721 43265 5733 43268
rect 5767 43265 5779 43299
rect 5721 43259 5779 43265
rect 6549 43299 6607 43305
rect 6549 43265 6561 43299
rect 6595 43265 6607 43299
rect 6549 43259 6607 43265
rect 7009 43299 7067 43305
rect 7009 43265 7021 43299
rect 7055 43296 7067 43299
rect 7374 43296 7380 43308
rect 7055 43268 7380 43296
rect 7055 43265 7067 43268
rect 7009 43259 7067 43265
rect 5074 43188 5080 43240
rect 5132 43188 5138 43240
rect 4212 43132 4660 43160
rect 4212 43120 4218 43132
rect 4341 43095 4399 43101
rect 4341 43061 4353 43095
rect 4387 43092 4399 43095
rect 5092 43092 5120 43188
rect 6564 43160 6592 43259
rect 7374 43256 7380 43268
rect 7432 43256 7438 43308
rect 7469 43299 7527 43305
rect 7469 43265 7481 43299
rect 7515 43296 7527 43299
rect 7650 43296 7656 43308
rect 7515 43268 7656 43296
rect 7515 43265 7527 43268
rect 7469 43259 7527 43265
rect 7650 43256 7656 43268
rect 7708 43256 7714 43308
rect 8021 43299 8079 43305
rect 8021 43265 8033 43299
rect 8067 43265 8079 43299
rect 8021 43259 8079 43265
rect 8481 43299 8539 43305
rect 8481 43265 8493 43299
rect 8527 43265 8539 43299
rect 8481 43259 8539 43265
rect 7466 43160 7472 43172
rect 6564 43132 7472 43160
rect 7466 43120 7472 43132
rect 7524 43120 7530 43172
rect 8036 43160 8064 43259
rect 8496 43228 8524 43259
rect 8938 43256 8944 43308
rect 8996 43256 9002 43308
rect 9309 43299 9367 43305
rect 9309 43265 9321 43299
rect 9355 43296 9367 43299
rect 9674 43296 9680 43308
rect 9355 43268 9680 43296
rect 9355 43265 9367 43268
rect 9309 43259 9367 43265
rect 9674 43256 9680 43268
rect 9732 43256 9738 43308
rect 11333 43299 11391 43305
rect 11333 43265 11345 43299
rect 11379 43296 11391 43299
rect 11606 43296 11612 43308
rect 11379 43268 11612 43296
rect 11379 43265 11391 43268
rect 11333 43259 11391 43265
rect 11606 43256 11612 43268
rect 11664 43256 11670 43308
rect 11701 43299 11759 43305
rect 11701 43265 11713 43299
rect 11747 43296 11759 43299
rect 11882 43296 11888 43308
rect 11747 43268 11888 43296
rect 11747 43265 11759 43268
rect 11701 43259 11759 43265
rect 11882 43256 11888 43268
rect 11940 43256 11946 43308
rect 11977 43299 12035 43305
rect 11977 43265 11989 43299
rect 12023 43296 12035 43299
rect 12066 43296 12072 43308
rect 12023 43268 12072 43296
rect 12023 43265 12035 43268
rect 11977 43259 12035 43265
rect 12066 43256 12072 43268
rect 12124 43256 12130 43308
rect 13354 43256 13360 43308
rect 13412 43296 13418 43308
rect 13740 43305 13768 43336
rect 14476 43305 14504 43336
rect 13633 43299 13691 43305
rect 13633 43296 13645 43299
rect 13412 43268 13645 43296
rect 13412 43256 13418 43268
rect 13633 43265 13645 43268
rect 13679 43265 13691 43299
rect 13633 43259 13691 43265
rect 13725 43299 13783 43305
rect 13725 43265 13737 43299
rect 13771 43265 13783 43299
rect 13725 43259 13783 43265
rect 14093 43299 14151 43305
rect 14093 43265 14105 43299
rect 14139 43265 14151 43299
rect 14093 43259 14151 43265
rect 14461 43299 14519 43305
rect 14461 43265 14473 43299
rect 14507 43265 14519 43299
rect 14461 43259 14519 43265
rect 10594 43228 10600 43240
rect 8496 43200 10600 43228
rect 10594 43188 10600 43200
rect 10652 43188 10658 43240
rect 13262 43188 13268 43240
rect 13320 43228 13326 43240
rect 14108 43228 14136 43259
rect 14734 43256 14740 43308
rect 14792 43296 14798 43308
rect 15013 43299 15071 43305
rect 15013 43296 15025 43299
rect 14792 43268 15025 43296
rect 14792 43256 14798 43268
rect 15013 43265 15025 43268
rect 15059 43265 15071 43299
rect 15013 43259 15071 43265
rect 15286 43256 15292 43308
rect 15344 43256 15350 43308
rect 15562 43256 15568 43308
rect 15620 43256 15626 43308
rect 15654 43256 15660 43308
rect 15712 43296 15718 43308
rect 15841 43299 15899 43305
rect 15841 43296 15853 43299
rect 15712 43268 15853 43296
rect 15712 43256 15718 43268
rect 15841 43265 15853 43268
rect 15887 43265 15899 43299
rect 15841 43259 15899 43265
rect 16114 43256 16120 43308
rect 16172 43256 16178 43308
rect 16408 43305 16436 43404
rect 16574 43392 16580 43444
rect 16632 43432 16638 43444
rect 16853 43435 16911 43441
rect 16853 43432 16865 43435
rect 16632 43404 16865 43432
rect 16632 43392 16638 43404
rect 16853 43401 16865 43404
rect 16899 43401 16911 43435
rect 16853 43395 16911 43401
rect 16942 43392 16948 43444
rect 17000 43432 17006 43444
rect 17405 43435 17463 43441
rect 17405 43432 17417 43435
rect 17000 43404 17417 43432
rect 17000 43392 17006 43404
rect 17405 43401 17417 43404
rect 17451 43401 17463 43435
rect 17405 43395 17463 43401
rect 17770 43392 17776 43444
rect 17828 43392 17834 43444
rect 18141 43435 18199 43441
rect 18141 43401 18153 43435
rect 18187 43401 18199 43435
rect 18141 43395 18199 43401
rect 17310 43324 17316 43376
rect 17368 43364 17374 43376
rect 18156 43364 18184 43395
rect 18414 43392 18420 43444
rect 18472 43432 18478 43444
rect 19429 43435 19487 43441
rect 19429 43432 19441 43435
rect 18472 43404 19441 43432
rect 18472 43392 18478 43404
rect 19429 43401 19441 43404
rect 19475 43401 19487 43435
rect 19429 43395 19487 43401
rect 20714 43364 20720 43376
rect 17368 43336 18184 43364
rect 19352 43336 20720 43364
rect 17368 43324 17374 43336
rect 16393 43299 16451 43305
rect 16393 43265 16405 43299
rect 16439 43265 16451 43299
rect 16393 43259 16451 43265
rect 16761 43299 16819 43305
rect 16761 43265 16773 43299
rect 16807 43265 16819 43299
rect 16761 43259 16819 43265
rect 17221 43299 17279 43305
rect 17221 43265 17233 43299
rect 17267 43265 17279 43299
rect 17221 43259 17279 43265
rect 17589 43299 17647 43305
rect 17589 43265 17601 43299
rect 17635 43296 17647 43299
rect 17770 43296 17776 43308
rect 17635 43268 17776 43296
rect 17635 43265 17647 43268
rect 17589 43259 17647 43265
rect 13320 43200 14136 43228
rect 13320 43188 13326 43200
rect 14274 43188 14280 43240
rect 14332 43228 14338 43240
rect 14642 43228 14648 43240
rect 14332 43200 14648 43228
rect 14332 43188 14338 43200
rect 14642 43188 14648 43200
rect 14700 43188 14706 43240
rect 16298 43188 16304 43240
rect 16356 43228 16362 43240
rect 16776 43228 16804 43259
rect 16356 43200 16804 43228
rect 17236 43228 17264 43259
rect 17770 43256 17776 43268
rect 17828 43256 17834 43308
rect 18049 43299 18107 43305
rect 18049 43265 18061 43299
rect 18095 43296 18107 43299
rect 18414 43296 18420 43308
rect 18095 43268 18420 43296
rect 18095 43265 18107 43268
rect 18049 43259 18107 43265
rect 18414 43256 18420 43268
rect 18472 43256 18478 43308
rect 18598 43256 18604 43308
rect 18656 43256 18662 43308
rect 19352 43305 19380 43336
rect 20714 43324 20720 43336
rect 20772 43324 20778 43376
rect 20806 43324 20812 43376
rect 20864 43324 20870 43376
rect 19337 43299 19395 43305
rect 19337 43265 19349 43299
rect 19383 43265 19395 43299
rect 19337 43259 19395 43265
rect 19889 43299 19947 43305
rect 19889 43265 19901 43299
rect 19935 43265 19947 43299
rect 19889 43259 19947 43265
rect 20441 43299 20499 43305
rect 20441 43265 20453 43299
rect 20487 43265 20499 43299
rect 20441 43259 20499 43265
rect 17310 43228 17316 43240
rect 17236 43200 17316 43228
rect 16356 43188 16362 43200
rect 17310 43188 17316 43200
rect 17368 43188 17374 43240
rect 18506 43188 18512 43240
rect 18564 43228 18570 43240
rect 19904 43228 19932 43259
rect 18564 43200 19932 43228
rect 20456 43228 20484 43259
rect 20990 43256 20996 43308
rect 21048 43256 21054 43308
rect 21634 43228 21640 43240
rect 20456 43200 21640 43228
rect 18564 43188 18570 43200
rect 21634 43188 21640 43200
rect 21692 43188 21698 43240
rect 8478 43160 8484 43172
rect 8036 43132 8484 43160
rect 8478 43120 8484 43132
rect 8536 43120 8542 43172
rect 8570 43120 8576 43172
rect 8628 43160 8634 43172
rect 8628 43132 9904 43160
rect 8628 43120 8634 43132
rect 4387 43064 5120 43092
rect 7193 43095 7251 43101
rect 4387 43061 4399 43064
rect 4341 43055 4399 43061
rect 7193 43061 7205 43095
rect 7239 43092 7251 43095
rect 8110 43092 8116 43104
rect 7239 43064 8116 43092
rect 7239 43061 7251 43064
rect 7193 43055 7251 43061
rect 8110 43052 8116 43064
rect 8168 43052 8174 43104
rect 8202 43052 8208 43104
rect 8260 43092 8266 43104
rect 9876 43101 9904 43132
rect 10226 43120 10232 43172
rect 10284 43160 10290 43172
rect 11057 43163 11115 43169
rect 11057 43160 11069 43163
rect 10284 43132 11069 43160
rect 10284 43120 10290 43132
rect 11057 43129 11069 43132
rect 11103 43129 11115 43163
rect 11057 43123 11115 43129
rect 13078 43120 13084 43172
rect 13136 43120 13142 43172
rect 13446 43120 13452 43172
rect 13504 43120 13510 43172
rect 13538 43120 13544 43172
rect 13596 43160 13602 43172
rect 16209 43163 16267 43169
rect 16209 43160 16221 43163
rect 13596 43132 16221 43160
rect 13596 43120 13602 43132
rect 16209 43129 16221 43132
rect 16255 43129 16267 43163
rect 16209 43123 16267 43129
rect 17678 43120 17684 43172
rect 17736 43160 17742 43172
rect 17736 43132 18736 43160
rect 17736 43120 17742 43132
rect 9493 43095 9551 43101
rect 9493 43092 9505 43095
rect 8260 43064 9505 43092
rect 8260 43052 8266 43064
rect 9493 43061 9505 43064
rect 9539 43061 9551 43095
rect 9493 43055 9551 43061
rect 9861 43095 9919 43101
rect 9861 43061 9873 43095
rect 9907 43061 9919 43095
rect 9861 43055 9919 43061
rect 10413 43095 10471 43101
rect 10413 43061 10425 43095
rect 10459 43092 10471 43095
rect 10778 43092 10784 43104
rect 10459 43064 10784 43092
rect 10459 43061 10471 43064
rect 10413 43055 10471 43061
rect 10778 43052 10784 43064
rect 10836 43052 10842 43104
rect 11146 43052 11152 43104
rect 11204 43052 11210 43104
rect 11698 43052 11704 43104
rect 11756 43092 11762 43104
rect 11885 43095 11943 43101
rect 11885 43092 11897 43095
rect 11756 43064 11897 43092
rect 11756 43052 11762 43064
rect 11885 43061 11897 43064
rect 11931 43061 11943 43095
rect 11885 43055 11943 43061
rect 13354 43052 13360 43104
rect 13412 43092 13418 43104
rect 14277 43095 14335 43101
rect 14277 43092 14289 43095
rect 13412 43064 14289 43092
rect 13412 43052 13418 43064
rect 14277 43061 14289 43064
rect 14323 43061 14335 43095
rect 14277 43055 14335 43061
rect 14642 43052 14648 43104
rect 14700 43052 14706 43104
rect 14826 43052 14832 43104
rect 14884 43052 14890 43104
rect 15105 43095 15163 43101
rect 15105 43061 15117 43095
rect 15151 43092 15163 43095
rect 15286 43092 15292 43104
rect 15151 43064 15292 43092
rect 15151 43061 15163 43064
rect 15105 43055 15163 43061
rect 15286 43052 15292 43064
rect 15344 43052 15350 43104
rect 15378 43052 15384 43104
rect 15436 43052 15442 43104
rect 15654 43052 15660 43104
rect 15712 43052 15718 43104
rect 15930 43052 15936 43104
rect 15988 43052 15994 43104
rect 18708 43101 18736 43132
rect 19426 43120 19432 43172
rect 19484 43160 19490 43172
rect 19484 43132 21128 43160
rect 19484 43120 19490 43132
rect 18693 43095 18751 43101
rect 18693 43061 18705 43095
rect 18739 43061 18751 43095
rect 18693 43055 18751 43061
rect 18782 43052 18788 43104
rect 18840 43092 18846 43104
rect 21100 43101 21128 43132
rect 19981 43095 20039 43101
rect 19981 43092 19993 43095
rect 18840 43064 19993 43092
rect 18840 43052 18846 43064
rect 19981 43061 19993 43064
rect 20027 43061 20039 43095
rect 19981 43055 20039 43061
rect 21085 43095 21143 43101
rect 21085 43061 21097 43095
rect 21131 43061 21143 43095
rect 21085 43055 21143 43061
rect 1104 43002 21896 43024
rect 1104 42950 3549 43002
rect 3601 42950 3613 43002
rect 3665 42950 3677 43002
rect 3729 42950 3741 43002
rect 3793 42950 3805 43002
rect 3857 42950 8747 43002
rect 8799 42950 8811 43002
rect 8863 42950 8875 43002
rect 8927 42950 8939 43002
rect 8991 42950 9003 43002
rect 9055 42950 13945 43002
rect 13997 42950 14009 43002
rect 14061 42950 14073 43002
rect 14125 42950 14137 43002
rect 14189 42950 14201 43002
rect 14253 42950 19143 43002
rect 19195 42950 19207 43002
rect 19259 42950 19271 43002
rect 19323 42950 19335 43002
rect 19387 42950 19399 43002
rect 19451 42950 21896 43002
rect 1104 42928 21896 42950
rect 5353 42891 5411 42897
rect 5353 42857 5365 42891
rect 5399 42888 5411 42891
rect 5994 42888 6000 42900
rect 5399 42860 6000 42888
rect 5399 42857 5411 42860
rect 5353 42851 5411 42857
rect 5994 42848 6000 42860
rect 6052 42848 6058 42900
rect 6104 42860 7052 42888
rect 2961 42823 3019 42829
rect 2961 42789 2973 42823
rect 3007 42789 3019 42823
rect 2961 42783 3019 42789
rect 2866 42752 2872 42764
rect 2516 42724 2872 42752
rect 1946 42644 1952 42696
rect 2004 42644 2010 42696
rect 2516 42693 2544 42724
rect 2866 42712 2872 42724
rect 2924 42712 2930 42764
rect 2976 42752 3004 42783
rect 4430 42780 4436 42832
rect 4488 42820 4494 42832
rect 6104 42820 6132 42860
rect 4488 42792 6132 42820
rect 7024 42820 7052 42860
rect 7650 42848 7656 42900
rect 7708 42888 7714 42900
rect 9674 42888 9680 42900
rect 7708 42860 9680 42888
rect 7708 42848 7714 42860
rect 9674 42848 9680 42860
rect 9732 42848 9738 42900
rect 11517 42891 11575 42897
rect 11517 42888 11529 42891
rect 11256 42860 11529 42888
rect 8570 42820 8576 42832
rect 7024 42792 8576 42820
rect 4488 42780 4494 42792
rect 8570 42780 8576 42792
rect 8628 42780 8634 42832
rect 9140 42792 9812 42820
rect 3142 42752 3148 42764
rect 2976 42724 3148 42752
rect 3142 42712 3148 42724
rect 3200 42712 3206 42764
rect 3418 42712 3424 42764
rect 3476 42752 3482 42764
rect 3513 42755 3571 42761
rect 3513 42752 3525 42755
rect 3476 42724 3525 42752
rect 3476 42712 3482 42724
rect 3513 42721 3525 42724
rect 3559 42721 3571 42755
rect 3513 42715 3571 42721
rect 4249 42755 4307 42761
rect 4249 42721 4261 42755
rect 4295 42752 4307 42755
rect 4614 42752 4620 42764
rect 4295 42724 4620 42752
rect 4295 42721 4307 42724
rect 4249 42715 4307 42721
rect 4614 42712 4620 42724
rect 4672 42712 4678 42764
rect 4801 42755 4859 42761
rect 4801 42721 4813 42755
rect 4847 42752 4859 42755
rect 4982 42752 4988 42764
rect 4847 42724 4988 42752
rect 4847 42721 4859 42724
rect 4801 42715 4859 42721
rect 4982 42712 4988 42724
rect 5040 42712 5046 42764
rect 6457 42755 6515 42761
rect 6457 42721 6469 42755
rect 6503 42752 6515 42755
rect 6822 42752 6828 42764
rect 6503 42724 6828 42752
rect 6503 42721 6515 42724
rect 6457 42715 6515 42721
rect 6822 42712 6828 42724
rect 6880 42712 6886 42764
rect 7006 42712 7012 42764
rect 7064 42712 7070 42764
rect 7558 42712 7564 42764
rect 7616 42712 7622 42764
rect 8113 42755 8171 42761
rect 8113 42721 8125 42755
rect 8159 42752 8171 42755
rect 8202 42752 8208 42764
rect 8159 42724 8208 42752
rect 8159 42721 8171 42724
rect 8113 42715 8171 42721
rect 8202 42712 8208 42724
rect 8260 42712 8266 42764
rect 8662 42712 8668 42764
rect 8720 42712 8726 42764
rect 8754 42712 8760 42764
rect 8812 42752 8818 42764
rect 9140 42752 9168 42792
rect 8812 42724 9168 42752
rect 8812 42712 8818 42724
rect 9214 42712 9220 42764
rect 9272 42752 9278 42764
rect 9677 42755 9735 42761
rect 9677 42752 9689 42755
rect 9272 42724 9689 42752
rect 9272 42712 9278 42724
rect 9677 42721 9689 42724
rect 9723 42721 9735 42755
rect 9784 42752 9812 42792
rect 11256 42752 11284 42860
rect 11517 42857 11529 42860
rect 11563 42857 11575 42891
rect 11517 42851 11575 42857
rect 12158 42848 12164 42900
rect 12216 42888 12222 42900
rect 14642 42888 14648 42900
rect 12216 42860 14648 42888
rect 12216 42848 12222 42860
rect 14642 42848 14648 42860
rect 14700 42848 14706 42900
rect 15654 42848 15660 42900
rect 15712 42848 15718 42900
rect 16022 42848 16028 42900
rect 16080 42888 16086 42900
rect 16390 42888 16396 42900
rect 16080 42860 16396 42888
rect 16080 42848 16086 42860
rect 16390 42848 16396 42860
rect 16448 42848 16454 42900
rect 17218 42848 17224 42900
rect 17276 42848 17282 42900
rect 17494 42848 17500 42900
rect 17552 42888 17558 42900
rect 17773 42891 17831 42897
rect 17773 42888 17785 42891
rect 17552 42860 17785 42888
rect 17552 42848 17558 42860
rect 17773 42857 17785 42860
rect 17819 42857 17831 42891
rect 18782 42888 18788 42900
rect 17773 42851 17831 42857
rect 17880 42860 18788 42888
rect 11330 42780 11336 42832
rect 11388 42780 11394 42832
rect 15672 42820 15700 42848
rect 15120 42792 15700 42820
rect 9784 42724 11284 42752
rect 11348 42752 11376 42780
rect 11348 42724 12204 42752
rect 9677 42715 9735 42721
rect 2501 42687 2559 42693
rect 2056 42656 2360 42684
rect 382 42576 388 42628
rect 440 42616 446 42628
rect 1394 42616 1400 42628
rect 440 42588 1400 42616
rect 440 42576 446 42588
rect 1394 42576 1400 42588
rect 1452 42576 1458 42628
rect 2056 42616 2084 42656
rect 1780 42588 2084 42616
rect 1780 42557 1808 42588
rect 2130 42576 2136 42628
rect 2188 42576 2194 42628
rect 1765 42551 1823 42557
rect 1765 42517 1777 42551
rect 1811 42517 1823 42551
rect 2332 42548 2360 42656
rect 2501 42653 2513 42687
rect 2547 42653 2559 42687
rect 2501 42647 2559 42653
rect 2958 42644 2964 42696
rect 3016 42684 3022 42696
rect 3237 42687 3295 42693
rect 3237 42684 3249 42687
rect 3016 42656 3249 42684
rect 3016 42644 3022 42656
rect 3237 42653 3249 42656
rect 3283 42653 3295 42687
rect 3237 42647 3295 42653
rect 5997 42687 6055 42693
rect 5997 42653 6009 42687
rect 6043 42684 6055 42687
rect 6546 42684 6552 42696
rect 6043 42656 6552 42684
rect 6043 42653 6055 42656
rect 5997 42647 6055 42653
rect 6546 42644 6552 42656
rect 6604 42644 6610 42696
rect 9122 42644 9128 42696
rect 9180 42644 9186 42696
rect 9582 42644 9588 42696
rect 9640 42684 9646 42696
rect 9861 42687 9919 42693
rect 9861 42684 9873 42687
rect 9640 42656 9873 42684
rect 9640 42644 9646 42656
rect 9861 42653 9873 42656
rect 9907 42653 9919 42687
rect 9861 42647 9919 42653
rect 10410 42644 10416 42696
rect 10468 42684 10474 42696
rect 10505 42687 10563 42693
rect 10505 42684 10517 42687
rect 10468 42656 10517 42684
rect 10468 42644 10474 42656
rect 10505 42653 10517 42656
rect 10551 42653 10563 42687
rect 10505 42647 10563 42653
rect 10686 42644 10692 42696
rect 10744 42684 10750 42696
rect 10781 42687 10839 42693
rect 10781 42684 10793 42687
rect 10744 42656 10793 42684
rect 10744 42644 10750 42656
rect 10781 42653 10793 42656
rect 10827 42653 10839 42687
rect 10781 42647 10839 42653
rect 10962 42644 10968 42696
rect 11020 42684 11026 42696
rect 11057 42687 11115 42693
rect 11057 42684 11069 42687
rect 11020 42656 11069 42684
rect 11020 42644 11026 42656
rect 11057 42653 11069 42656
rect 11103 42653 11115 42687
rect 11057 42647 11115 42653
rect 11146 42644 11152 42696
rect 11204 42684 11210 42696
rect 11333 42687 11391 42693
rect 11333 42684 11345 42687
rect 11204 42656 11345 42684
rect 11204 42644 11210 42656
rect 11333 42653 11345 42656
rect 11379 42653 11391 42687
rect 11333 42647 11391 42653
rect 11422 42644 11428 42696
rect 11480 42684 11486 42696
rect 11701 42687 11759 42693
rect 11701 42684 11713 42687
rect 11480 42656 11713 42684
rect 11480 42644 11486 42656
rect 11701 42653 11713 42656
rect 11747 42653 11759 42687
rect 11701 42647 11759 42653
rect 11882 42644 11888 42696
rect 11940 42644 11946 42696
rect 12176 42693 12204 42724
rect 12250 42712 12256 42764
rect 12308 42752 12314 42764
rect 15120 42752 15148 42792
rect 15746 42780 15752 42832
rect 15804 42820 15810 42832
rect 17880 42820 17908 42860
rect 18782 42848 18788 42860
rect 18840 42848 18846 42900
rect 19702 42848 19708 42900
rect 19760 42888 19766 42900
rect 20533 42891 20591 42897
rect 20533 42888 20545 42891
rect 19760 42860 20545 42888
rect 19760 42848 19766 42860
rect 20533 42857 20545 42860
rect 20579 42857 20591 42891
rect 20533 42851 20591 42857
rect 15804 42792 17908 42820
rect 15804 42780 15810 42792
rect 18230 42780 18236 42832
rect 18288 42820 18294 42832
rect 18288 42792 19334 42820
rect 18288 42780 18294 42792
rect 12308 42724 13768 42752
rect 12308 42712 12314 42724
rect 12161 42687 12219 42693
rect 12161 42653 12173 42687
rect 12207 42653 12219 42687
rect 12161 42647 12219 42653
rect 12618 42644 12624 42696
rect 12676 42644 12682 42696
rect 13081 42687 13139 42693
rect 13081 42653 13093 42687
rect 13127 42653 13139 42687
rect 13081 42647 13139 42653
rect 2682 42576 2688 42628
rect 2740 42576 2746 42628
rect 2774 42576 2780 42628
rect 2832 42616 2838 42628
rect 3973 42619 4031 42625
rect 3973 42616 3985 42619
rect 2832 42588 3985 42616
rect 2832 42576 2838 42588
rect 3973 42585 3985 42588
rect 4019 42585 4031 42619
rect 3973 42579 4031 42585
rect 4525 42619 4583 42625
rect 4525 42585 4537 42619
rect 4571 42616 4583 42619
rect 4890 42616 4896 42628
rect 4571 42588 4896 42616
rect 4571 42585 4583 42588
rect 4525 42579 4583 42585
rect 4890 42576 4896 42588
rect 4948 42576 4954 42628
rect 5074 42576 5080 42628
rect 5132 42576 5138 42628
rect 5629 42619 5687 42625
rect 5629 42585 5641 42619
rect 5675 42616 5687 42619
rect 5810 42616 5816 42628
rect 5675 42588 5816 42616
rect 5675 42585 5687 42588
rect 5629 42579 5687 42585
rect 5810 42576 5816 42588
rect 5868 42576 5874 42628
rect 5902 42576 5908 42628
rect 5960 42616 5966 42628
rect 6181 42619 6239 42625
rect 6181 42616 6193 42619
rect 5960 42588 6193 42616
rect 5960 42576 5966 42588
rect 6181 42585 6193 42588
rect 6227 42585 6239 42619
rect 6181 42579 6239 42585
rect 6730 42576 6736 42628
rect 6788 42576 6794 42628
rect 7285 42619 7343 42625
rect 7285 42585 7297 42619
rect 7331 42585 7343 42619
rect 7285 42579 7343 42585
rect 3050 42548 3056 42560
rect 2332 42520 3056 42548
rect 1765 42511 1823 42517
rect 3050 42508 3056 42520
rect 3108 42508 3114 42560
rect 5994 42508 6000 42560
rect 6052 42548 6058 42560
rect 7300 42548 7328 42579
rect 7834 42576 7840 42628
rect 7892 42576 7898 42628
rect 8386 42576 8392 42628
rect 8444 42576 8450 42628
rect 8754 42616 8760 42628
rect 8496 42588 8760 42616
rect 6052 42520 7328 42548
rect 6052 42508 6058 42520
rect 8018 42508 8024 42560
rect 8076 42548 8082 42560
rect 8496 42548 8524 42588
rect 8754 42576 8760 42588
rect 8812 42576 8818 42628
rect 9306 42576 9312 42628
rect 9364 42616 9370 42628
rect 9401 42619 9459 42625
rect 9401 42616 9413 42619
rect 9364 42588 9413 42616
rect 9364 42576 9370 42588
rect 9401 42585 9413 42588
rect 9447 42585 9459 42619
rect 9401 42579 9459 42585
rect 9490 42576 9496 42628
rect 9548 42616 9554 42628
rect 13096 42616 13124 42647
rect 13170 42644 13176 42696
rect 13228 42644 13234 42696
rect 13538 42644 13544 42696
rect 13596 42644 13602 42696
rect 13630 42644 13636 42696
rect 13688 42644 13694 42696
rect 13556 42616 13584 42644
rect 9548 42588 10364 42616
rect 9548 42576 9554 42588
rect 8076 42520 8524 42548
rect 8076 42508 8082 42520
rect 8662 42508 8668 42560
rect 8720 42548 8726 42560
rect 8941 42551 8999 42557
rect 8941 42548 8953 42551
rect 8720 42520 8953 42548
rect 8720 42508 8726 42520
rect 8941 42517 8953 42520
rect 8987 42517 8999 42551
rect 8941 42511 8999 42517
rect 9214 42508 9220 42560
rect 9272 42548 9278 42560
rect 9858 42548 9864 42560
rect 9272 42520 9864 42548
rect 9272 42508 9278 42520
rect 9858 42508 9864 42520
rect 9916 42508 9922 42560
rect 10042 42508 10048 42560
rect 10100 42508 10106 42560
rect 10336 42557 10364 42588
rect 11256 42588 12848 42616
rect 13096 42588 13584 42616
rect 11256 42560 11284 42588
rect 10321 42551 10379 42557
rect 10321 42517 10333 42551
rect 10367 42517 10379 42551
rect 10321 42511 10379 42517
rect 10502 42508 10508 42560
rect 10560 42548 10566 42560
rect 10597 42551 10655 42557
rect 10597 42548 10609 42551
rect 10560 42520 10609 42548
rect 10560 42508 10566 42520
rect 10597 42517 10609 42520
rect 10643 42517 10655 42551
rect 10597 42511 10655 42517
rect 10686 42508 10692 42560
rect 10744 42548 10750 42560
rect 10873 42551 10931 42557
rect 10873 42548 10885 42551
rect 10744 42520 10885 42548
rect 10744 42508 10750 42520
rect 10873 42517 10885 42520
rect 10919 42517 10931 42551
rect 10873 42511 10931 42517
rect 11146 42508 11152 42560
rect 11204 42508 11210 42560
rect 11238 42508 11244 42560
rect 11296 42508 11302 42560
rect 12066 42508 12072 42560
rect 12124 42508 12130 42560
rect 12342 42508 12348 42560
rect 12400 42508 12406 42560
rect 12820 42557 12848 42588
rect 12805 42551 12863 42557
rect 12805 42517 12817 42551
rect 12851 42517 12863 42551
rect 12805 42511 12863 42517
rect 12894 42508 12900 42560
rect 12952 42508 12958 42560
rect 12986 42508 12992 42560
rect 13044 42548 13050 42560
rect 13740 42557 13768 42724
rect 14660 42724 15148 42752
rect 13814 42644 13820 42696
rect 13872 42684 13878 42696
rect 14660 42693 14688 42724
rect 15470 42712 15476 42764
rect 15528 42752 15534 42764
rect 17126 42752 17132 42764
rect 15528 42724 17132 42752
rect 15528 42712 15534 42724
rect 17126 42712 17132 42724
rect 17184 42712 17190 42764
rect 18046 42712 18052 42764
rect 18104 42752 18110 42764
rect 18509 42755 18567 42761
rect 18509 42752 18521 42755
rect 18104 42724 18521 42752
rect 18104 42712 18110 42724
rect 18509 42721 18521 42724
rect 18555 42721 18567 42755
rect 19306 42752 19334 42792
rect 19613 42755 19671 42761
rect 19613 42752 19625 42755
rect 19306 42724 19625 42752
rect 18509 42715 18567 42721
rect 19613 42721 19625 42724
rect 19659 42721 19671 42755
rect 19613 42715 19671 42721
rect 19978 42712 19984 42764
rect 20036 42752 20042 42764
rect 21269 42755 21327 42761
rect 21269 42752 21281 42755
rect 20036 42724 21281 42752
rect 20036 42712 20042 42724
rect 21269 42721 21281 42724
rect 21315 42721 21327 42755
rect 21269 42715 21327 42721
rect 14185 42687 14243 42693
rect 14185 42684 14197 42687
rect 13872 42656 14197 42684
rect 13872 42644 13878 42656
rect 14185 42653 14197 42656
rect 14231 42653 14243 42687
rect 14185 42647 14243 42653
rect 14645 42687 14703 42693
rect 14645 42653 14657 42687
rect 14691 42653 14703 42687
rect 14645 42647 14703 42653
rect 14921 42687 14979 42693
rect 14921 42653 14933 42687
rect 14967 42653 14979 42687
rect 14921 42647 14979 42653
rect 14090 42576 14096 42628
rect 14148 42616 14154 42628
rect 14936 42616 14964 42647
rect 18322 42644 18328 42696
rect 18380 42684 18386 42696
rect 18877 42687 18935 42693
rect 18877 42684 18889 42687
rect 18380 42656 18889 42684
rect 18380 42644 18386 42656
rect 18877 42653 18889 42656
rect 18923 42653 18935 42687
rect 18877 42647 18935 42653
rect 19058 42644 19064 42696
rect 19116 42684 19122 42696
rect 19116 42656 20024 42684
rect 19116 42644 19122 42656
rect 14148 42588 14964 42616
rect 14148 42576 14154 42588
rect 15102 42576 15108 42628
rect 15160 42576 15166 42628
rect 15470 42576 15476 42628
rect 15528 42616 15534 42628
rect 16853 42619 16911 42625
rect 15528 42588 16528 42616
rect 15528 42576 15534 42588
rect 13357 42551 13415 42557
rect 13357 42548 13369 42551
rect 13044 42520 13369 42548
rect 13044 42508 13050 42520
rect 13357 42517 13369 42520
rect 13403 42517 13415 42551
rect 13357 42511 13415 42517
rect 13725 42551 13783 42557
rect 13725 42517 13737 42551
rect 13771 42517 13783 42551
rect 13725 42511 13783 42517
rect 13814 42508 13820 42560
rect 13872 42548 13878 42560
rect 14277 42551 14335 42557
rect 14277 42548 14289 42551
rect 13872 42520 14289 42548
rect 13872 42508 13878 42520
rect 14277 42517 14289 42520
rect 14323 42517 14335 42551
rect 14277 42511 14335 42517
rect 14458 42508 14464 42560
rect 14516 42508 14522 42560
rect 14734 42508 14740 42560
rect 14792 42508 14798 42560
rect 16500 42548 16528 42588
rect 16853 42585 16865 42619
rect 16899 42616 16911 42619
rect 17034 42616 17040 42628
rect 16899 42588 17040 42616
rect 16899 42585 16911 42588
rect 16853 42579 16911 42585
rect 17034 42576 17040 42588
rect 17092 42576 17098 42628
rect 17129 42619 17187 42625
rect 17129 42585 17141 42619
rect 17175 42616 17187 42619
rect 17494 42616 17500 42628
rect 17175 42588 17500 42616
rect 17175 42585 17187 42588
rect 17129 42579 17187 42585
rect 17494 42576 17500 42588
rect 17552 42576 17558 42628
rect 17586 42576 17592 42628
rect 17644 42616 17650 42628
rect 17681 42619 17739 42625
rect 17681 42616 17693 42619
rect 17644 42588 17693 42616
rect 17644 42576 17650 42588
rect 17681 42585 17693 42588
rect 17727 42585 17739 42619
rect 17681 42579 17739 42585
rect 18046 42576 18052 42628
rect 18104 42616 18110 42628
rect 18233 42619 18291 42625
rect 18233 42616 18245 42619
rect 18104 42588 18245 42616
rect 18104 42576 18110 42588
rect 18233 42585 18245 42588
rect 18279 42585 18291 42619
rect 18233 42579 18291 42585
rect 19334 42576 19340 42628
rect 19392 42576 19398 42628
rect 19610 42576 19616 42628
rect 19668 42616 19674 42628
rect 19889 42619 19947 42625
rect 19889 42616 19901 42619
rect 19668 42588 19901 42616
rect 19668 42576 19674 42588
rect 19889 42585 19901 42588
rect 19935 42585 19947 42619
rect 19889 42579 19947 42585
rect 19996 42557 20024 42656
rect 20438 42576 20444 42628
rect 20496 42576 20502 42628
rect 20993 42619 21051 42625
rect 20993 42585 21005 42619
rect 21039 42616 21051 42619
rect 21358 42616 21364 42628
rect 21039 42588 21364 42616
rect 21039 42585 21051 42588
rect 20993 42579 21051 42585
rect 21358 42576 21364 42588
rect 21416 42576 21422 42628
rect 18693 42551 18751 42557
rect 18693 42548 18705 42551
rect 16500 42520 18705 42548
rect 18693 42517 18705 42520
rect 18739 42517 18751 42551
rect 18693 42511 18751 42517
rect 19981 42551 20039 42557
rect 19981 42517 19993 42551
rect 20027 42517 20039 42551
rect 19981 42511 20039 42517
rect 1104 42458 22056 42480
rect 1104 42406 6148 42458
rect 6200 42406 6212 42458
rect 6264 42406 6276 42458
rect 6328 42406 6340 42458
rect 6392 42406 6404 42458
rect 6456 42406 11346 42458
rect 11398 42406 11410 42458
rect 11462 42406 11474 42458
rect 11526 42406 11538 42458
rect 11590 42406 11602 42458
rect 11654 42406 16544 42458
rect 16596 42406 16608 42458
rect 16660 42406 16672 42458
rect 16724 42406 16736 42458
rect 16788 42406 16800 42458
rect 16852 42406 21742 42458
rect 21794 42406 21806 42458
rect 21858 42406 21870 42458
rect 21922 42406 21934 42458
rect 21986 42406 21998 42458
rect 22050 42406 22056 42458
rect 1104 42384 22056 42406
rect 2038 42304 2044 42356
rect 2096 42344 2102 42356
rect 2501 42347 2559 42353
rect 2501 42344 2513 42347
rect 2096 42316 2513 42344
rect 2096 42304 2102 42316
rect 2501 42313 2513 42316
rect 2547 42313 2559 42347
rect 2501 42307 2559 42313
rect 2774 42304 2780 42356
rect 2832 42304 2838 42356
rect 3053 42347 3111 42353
rect 3053 42313 3065 42347
rect 3099 42313 3111 42347
rect 3053 42307 3111 42313
rect 3513 42347 3571 42353
rect 3513 42313 3525 42347
rect 3559 42344 3571 42347
rect 4062 42344 4068 42356
rect 3559 42316 4068 42344
rect 3559 42313 3571 42316
rect 3513 42307 3571 42313
rect 3068 42276 3096 42307
rect 4062 42304 4068 42316
rect 4120 42304 4126 42356
rect 4157 42347 4215 42353
rect 4157 42313 4169 42347
rect 4203 42344 4215 42347
rect 4246 42344 4252 42356
rect 4203 42316 4252 42344
rect 4203 42313 4215 42316
rect 4157 42307 4215 42313
rect 4246 42304 4252 42316
rect 4304 42304 4310 42356
rect 4522 42304 4528 42356
rect 4580 42304 4586 42356
rect 4798 42304 4804 42356
rect 4856 42344 4862 42356
rect 5077 42347 5135 42353
rect 5077 42344 5089 42347
rect 4856 42316 5089 42344
rect 4856 42304 4862 42316
rect 5077 42313 5089 42316
rect 5123 42313 5135 42347
rect 5077 42307 5135 42313
rect 5626 42304 5632 42356
rect 5684 42304 5690 42356
rect 5994 42304 6000 42356
rect 6052 42304 6058 42356
rect 6549 42347 6607 42353
rect 6549 42313 6561 42347
rect 6595 42344 6607 42347
rect 6638 42344 6644 42356
rect 6595 42316 6644 42344
rect 6595 42313 6607 42316
rect 6549 42307 6607 42313
rect 6638 42304 6644 42316
rect 6696 42304 6702 42356
rect 7190 42304 7196 42356
rect 7248 42344 7254 42356
rect 7469 42347 7527 42353
rect 7469 42344 7481 42347
rect 7248 42316 7481 42344
rect 7248 42304 7254 42316
rect 7469 42313 7481 42316
rect 7515 42313 7527 42347
rect 10321 42347 10379 42353
rect 10321 42344 10333 42347
rect 7469 42307 7527 42313
rect 9232 42316 10333 42344
rect 9232 42276 9260 42316
rect 10321 42313 10333 42316
rect 10367 42313 10379 42347
rect 10321 42307 10379 42313
rect 10594 42304 10600 42356
rect 10652 42304 10658 42356
rect 12894 42304 12900 42356
rect 12952 42304 12958 42356
rect 14458 42344 14464 42356
rect 13556 42316 14464 42344
rect 3068 42248 4936 42276
rect 1854 42168 1860 42220
rect 1912 42208 1918 42220
rect 2685 42211 2743 42217
rect 2685 42208 2697 42211
rect 1912 42180 2697 42208
rect 1912 42168 1918 42180
rect 2685 42177 2697 42180
rect 2731 42177 2743 42211
rect 2685 42171 2743 42177
rect 2961 42211 3019 42217
rect 2961 42177 2973 42211
rect 3007 42177 3019 42211
rect 2961 42171 3019 42177
rect 658 42100 664 42152
rect 716 42140 722 42152
rect 2976 42140 3004 42171
rect 3234 42168 3240 42220
rect 3292 42168 3298 42220
rect 3326 42168 3332 42220
rect 3384 42168 3390 42220
rect 3878 42168 3884 42220
rect 3936 42168 3942 42220
rect 4908 42217 4936 42248
rect 5644 42248 9260 42276
rect 4433 42211 4491 42217
rect 4433 42177 4445 42211
rect 4479 42177 4491 42211
rect 4433 42171 4491 42177
rect 4893 42211 4951 42217
rect 4893 42177 4905 42211
rect 4939 42177 4951 42211
rect 4893 42171 4951 42177
rect 716 42112 3004 42140
rect 4448 42140 4476 42171
rect 5258 42168 5264 42220
rect 5316 42208 5322 42220
rect 5537 42211 5595 42217
rect 5537 42208 5549 42211
rect 5316 42180 5549 42208
rect 5316 42168 5322 42180
rect 5537 42177 5549 42180
rect 5583 42177 5595 42211
rect 5537 42171 5595 42177
rect 5644 42140 5672 42248
rect 9858 42236 9864 42288
rect 9916 42276 9922 42288
rect 9916 42248 10088 42276
rect 9916 42236 9922 42248
rect 6178 42168 6184 42220
rect 6236 42168 6242 42220
rect 6365 42211 6423 42217
rect 6365 42177 6377 42211
rect 6411 42177 6423 42211
rect 6365 42171 6423 42177
rect 6917 42211 6975 42217
rect 6917 42177 6929 42211
rect 6963 42208 6975 42211
rect 7282 42208 7288 42220
rect 6963 42180 7288 42208
rect 6963 42177 6975 42180
rect 6917 42171 6975 42177
rect 4448 42112 5672 42140
rect 716 42100 722 42112
rect 5718 42100 5724 42152
rect 5776 42140 5782 42152
rect 6380 42140 6408 42171
rect 7282 42168 7288 42180
rect 7340 42168 7346 42220
rect 7377 42211 7435 42217
rect 7377 42177 7389 42211
rect 7423 42177 7435 42211
rect 7377 42171 7435 42177
rect 8297 42211 8355 42217
rect 8297 42177 8309 42211
rect 8343 42208 8355 42211
rect 9125 42211 9183 42217
rect 9125 42208 9137 42211
rect 8343 42180 9137 42208
rect 8343 42177 8355 42180
rect 8297 42171 8355 42177
rect 9125 42177 9137 42180
rect 9171 42208 9183 42211
rect 9171 42192 9260 42208
rect 9171 42180 9352 42192
rect 9171 42177 9183 42180
rect 9125 42171 9183 42177
rect 7392 42140 7420 42171
rect 9232 42164 9352 42180
rect 9398 42168 9404 42220
rect 9456 42168 9462 42220
rect 9677 42211 9735 42217
rect 9677 42177 9689 42211
rect 9723 42208 9735 42211
rect 10060 42208 10088 42248
rect 10686 42236 10692 42288
rect 10744 42276 10750 42288
rect 11238 42276 11244 42288
rect 10744 42248 11244 42276
rect 10744 42236 10750 42248
rect 11238 42236 11244 42248
rect 11296 42236 11302 42288
rect 10505 42211 10563 42217
rect 10505 42208 10517 42211
rect 9723 42180 9996 42208
rect 10060 42180 10517 42208
rect 9723 42177 9735 42180
rect 9677 42171 9735 42177
rect 5776 42112 6408 42140
rect 6472 42112 7420 42140
rect 5776 42100 5782 42112
rect 5994 42032 6000 42084
rect 6052 42072 6058 42084
rect 6472 42072 6500 42112
rect 7742 42100 7748 42152
rect 7800 42100 7806 42152
rect 9324 42140 9352 42164
rect 9324 42112 9904 42140
rect 6052 42044 6500 42072
rect 7101 42075 7159 42081
rect 6052 42032 6058 42044
rect 7101 42041 7113 42075
rect 7147 42072 7159 42075
rect 7760 42072 7788 42100
rect 7147 42044 7788 42072
rect 7147 42041 7159 42044
rect 7101 42035 7159 42041
rect 8938 42032 8944 42084
rect 8996 42032 9002 42084
rect 9030 42032 9036 42084
rect 9088 42072 9094 42084
rect 9088 42044 9168 42072
rect 9088 42032 9094 42044
rect 1026 41964 1032 42016
rect 1084 42004 1090 42016
rect 7742 42004 7748 42016
rect 1084 41976 7748 42004
rect 1084 41964 1090 41976
rect 7742 41964 7748 41976
rect 7800 41964 7806 42016
rect 8570 41964 8576 42016
rect 8628 41964 8634 42016
rect 9140 42004 9168 42044
rect 9876 42016 9904 42112
rect 9968 42016 9996 42180
rect 10505 42177 10517 42180
rect 10551 42177 10563 42211
rect 10505 42171 10563 42177
rect 10781 42211 10839 42217
rect 10781 42177 10793 42211
rect 10827 42177 10839 42211
rect 10781 42171 10839 42177
rect 10134 42100 10140 42152
rect 10192 42140 10198 42152
rect 10796 42140 10824 42171
rect 10192 42112 10824 42140
rect 12912 42140 12940 42304
rect 13556 42217 13584 42316
rect 14458 42304 14464 42316
rect 14516 42304 14522 42356
rect 14734 42304 14740 42356
rect 14792 42304 14798 42356
rect 17310 42304 17316 42356
rect 17368 42304 17374 42356
rect 17402 42304 17408 42356
rect 17460 42344 17466 42356
rect 17957 42347 18015 42353
rect 17957 42344 17969 42347
rect 17460 42316 17969 42344
rect 17460 42304 17466 42316
rect 17957 42313 17969 42316
rect 18003 42313 18015 42347
rect 17957 42307 18015 42313
rect 18138 42304 18144 42356
rect 18196 42344 18202 42356
rect 18325 42347 18383 42353
rect 18325 42344 18337 42347
rect 18196 42316 18337 42344
rect 18196 42304 18202 42316
rect 18325 42313 18337 42316
rect 18371 42313 18383 42347
rect 18325 42307 18383 42313
rect 18969 42347 19027 42353
rect 18969 42313 18981 42347
rect 19015 42313 19027 42347
rect 18969 42307 19027 42313
rect 14185 42279 14243 42285
rect 14185 42245 14197 42279
rect 14231 42276 14243 42279
rect 14752 42276 14780 42304
rect 14231 42248 14780 42276
rect 14231 42245 14243 42248
rect 14185 42239 14243 42245
rect 14826 42236 14832 42288
rect 14884 42276 14890 42288
rect 15105 42279 15163 42285
rect 15105 42276 15117 42279
rect 14884 42248 15117 42276
rect 14884 42236 14890 42248
rect 15105 42245 15117 42248
rect 15151 42245 15163 42279
rect 15105 42239 15163 42245
rect 15194 42236 15200 42288
rect 15252 42276 15258 42288
rect 17328 42276 17356 42304
rect 18984 42276 19012 42307
rect 19150 42304 19156 42356
rect 19208 42344 19214 42356
rect 19613 42347 19671 42353
rect 19613 42344 19625 42347
rect 19208 42316 19625 42344
rect 19208 42304 19214 42316
rect 19613 42313 19625 42316
rect 19659 42313 19671 42347
rect 19613 42307 19671 42313
rect 20165 42347 20223 42353
rect 20165 42313 20177 42347
rect 20211 42344 20223 42347
rect 22186 42344 22192 42356
rect 20211 42316 22192 42344
rect 20211 42313 20223 42316
rect 20165 42307 20223 42313
rect 22186 42304 22192 42316
rect 22244 42304 22250 42356
rect 22370 42304 22376 42356
rect 22428 42304 22434 42356
rect 15252 42248 17172 42276
rect 17328 42248 19012 42276
rect 15252 42236 15258 42248
rect 13541 42211 13599 42217
rect 13541 42177 13553 42211
rect 13587 42177 13599 42211
rect 13541 42171 13599 42177
rect 13722 42168 13728 42220
rect 13780 42208 13786 42220
rect 14090 42208 14096 42220
rect 13780 42180 14096 42208
rect 13780 42168 13786 42180
rect 14090 42168 14096 42180
rect 14148 42168 14154 42220
rect 14645 42211 14703 42217
rect 14645 42177 14657 42211
rect 14691 42177 14703 42211
rect 14645 42171 14703 42177
rect 14660 42140 14688 42171
rect 15286 42168 15292 42220
rect 15344 42208 15350 42220
rect 15381 42211 15439 42217
rect 15381 42208 15393 42211
rect 15344 42180 15393 42208
rect 15344 42168 15350 42180
rect 15381 42177 15393 42180
rect 15427 42177 15439 42211
rect 15381 42171 15439 42177
rect 15749 42211 15807 42217
rect 15749 42177 15761 42211
rect 15795 42208 15807 42211
rect 15930 42208 15936 42220
rect 15795 42180 15936 42208
rect 15795 42177 15807 42180
rect 15749 42171 15807 42177
rect 15930 42168 15936 42180
rect 15988 42168 15994 42220
rect 16022 42168 16028 42220
rect 16080 42208 16086 42220
rect 16209 42211 16267 42217
rect 16209 42208 16221 42211
rect 16080 42180 16221 42208
rect 16080 42168 16086 42180
rect 16209 42177 16221 42180
rect 16255 42177 16267 42211
rect 16209 42171 16267 42177
rect 16758 42168 16764 42220
rect 16816 42168 16822 42220
rect 12912 42112 14688 42140
rect 10192 42100 10198 42112
rect 15654 42100 15660 42152
rect 15712 42140 15718 42152
rect 16298 42140 16304 42152
rect 15712 42112 16304 42140
rect 15712 42100 15718 42112
rect 16298 42100 16304 42112
rect 16356 42100 16362 42152
rect 10686 42032 10692 42084
rect 10744 42072 10750 42084
rect 11698 42072 11704 42084
rect 10744 42044 11704 42072
rect 10744 42032 10750 42044
rect 11698 42032 11704 42044
rect 11756 42032 11762 42084
rect 11974 42032 11980 42084
rect 12032 42072 12038 42084
rect 13814 42072 13820 42084
rect 12032 42044 13820 42072
rect 12032 42032 12038 42044
rect 13814 42032 13820 42044
rect 13872 42032 13878 42084
rect 14936 42044 16344 42072
rect 14936 42016 14964 42044
rect 9217 42007 9275 42013
rect 9217 42004 9229 42007
rect 9140 41976 9229 42004
rect 9217 41973 9229 41976
rect 9263 41973 9275 42007
rect 9217 41967 9275 41973
rect 9493 42007 9551 42013
rect 9493 41973 9505 42007
rect 9539 42004 9551 42007
rect 9582 42004 9588 42016
rect 9539 41976 9588 42004
rect 9539 41973 9551 41976
rect 9493 41967 9551 41973
rect 9582 41964 9588 41976
rect 9640 41964 9646 42016
rect 9858 41964 9864 42016
rect 9916 41964 9922 42016
rect 9950 41964 9956 42016
rect 10008 41964 10014 42016
rect 13538 41964 13544 42016
rect 13596 42004 13602 42016
rect 13725 42007 13783 42013
rect 13725 42004 13737 42007
rect 13596 41976 13737 42004
rect 13596 41964 13602 41976
rect 13725 41973 13737 41976
rect 13771 41973 13783 42007
rect 13725 41967 13783 41973
rect 13998 41964 14004 42016
rect 14056 42004 14062 42016
rect 14277 42007 14335 42013
rect 14277 42004 14289 42007
rect 14056 41976 14289 42004
rect 14056 41964 14062 41976
rect 14277 41973 14289 41976
rect 14323 41973 14335 42007
rect 14277 41967 14335 41973
rect 14458 41964 14464 42016
rect 14516 42004 14522 42016
rect 14829 42007 14887 42013
rect 14829 42004 14841 42007
rect 14516 41976 14841 42004
rect 14516 41964 14522 41976
rect 14829 41973 14841 41976
rect 14875 41973 14887 42007
rect 14829 41967 14887 41973
rect 14918 41964 14924 42016
rect 14976 41964 14982 42016
rect 15194 41964 15200 42016
rect 15252 41964 15258 42016
rect 15565 42007 15623 42013
rect 15565 41973 15577 42007
rect 15611 42004 15623 42007
rect 15746 42004 15752 42016
rect 15611 41976 15752 42004
rect 15611 41973 15623 41976
rect 15565 41967 15623 41973
rect 15746 41964 15752 41976
rect 15804 41964 15810 42016
rect 15930 41964 15936 42016
rect 15988 41964 15994 42016
rect 16316 42013 16344 42044
rect 16301 42007 16359 42013
rect 16301 41973 16313 42007
rect 16347 41973 16359 42007
rect 16301 41967 16359 41973
rect 16850 41964 16856 42016
rect 16908 41964 16914 42016
rect 16942 41964 16948 42016
rect 17000 42004 17006 42016
rect 17037 42007 17095 42013
rect 17037 42004 17049 42007
rect 17000 41976 17049 42004
rect 17000 41964 17006 41976
rect 17037 41973 17049 41976
rect 17083 41973 17095 42007
rect 17144 42004 17172 42248
rect 19058 42236 19064 42288
rect 19116 42276 19122 42288
rect 19116 42248 19656 42276
rect 19116 42236 19122 42248
rect 17221 42211 17279 42217
rect 17221 42177 17233 42211
rect 17267 42177 17279 42211
rect 17221 42171 17279 42177
rect 17236 42072 17264 42171
rect 17494 42168 17500 42220
rect 17552 42168 17558 42220
rect 17770 42168 17776 42220
rect 17828 42168 17834 42220
rect 18233 42211 18291 42217
rect 18233 42177 18245 42211
rect 18279 42208 18291 42211
rect 18598 42208 18604 42220
rect 18279 42180 18604 42208
rect 18279 42177 18291 42180
rect 18233 42171 18291 42177
rect 18598 42168 18604 42180
rect 18656 42168 18662 42220
rect 18874 42168 18880 42220
rect 18932 42168 18938 42220
rect 18966 42168 18972 42220
rect 19024 42208 19030 42220
rect 19153 42211 19211 42217
rect 19153 42208 19165 42211
rect 19024 42180 19165 42208
rect 19024 42168 19030 42180
rect 19153 42177 19165 42180
rect 19199 42177 19211 42211
rect 19153 42171 19211 42177
rect 19518 42168 19524 42220
rect 19576 42168 19582 42220
rect 17402 42100 17408 42152
rect 17460 42140 17466 42152
rect 18322 42140 18328 42152
rect 17460 42112 18328 42140
rect 17460 42100 17466 42112
rect 18322 42100 18328 42112
rect 18380 42100 18386 42152
rect 19628 42140 19656 42248
rect 19702 42236 19708 42288
rect 19760 42276 19766 42288
rect 20809 42279 20867 42285
rect 20809 42276 20821 42279
rect 19760 42248 20821 42276
rect 19760 42236 19766 42248
rect 20809 42245 20821 42248
rect 20855 42245 20867 42279
rect 20809 42239 20867 42245
rect 21361 42279 21419 42285
rect 21361 42245 21373 42279
rect 21407 42276 21419 42279
rect 22388 42276 22416 42304
rect 21407 42248 22416 42276
rect 21407 42245 21419 42248
rect 21361 42239 21419 42245
rect 19978 42168 19984 42220
rect 20036 42168 20042 42220
rect 20438 42168 20444 42220
rect 20496 42168 20502 42220
rect 20898 42168 20904 42220
rect 20956 42208 20962 42220
rect 20993 42211 21051 42217
rect 20993 42208 21005 42211
rect 20956 42180 21005 42208
rect 20956 42168 20962 42180
rect 20993 42177 21005 42180
rect 21039 42177 21051 42211
rect 20993 42171 21051 42177
rect 21542 42140 21548 42152
rect 19628 42112 21548 42140
rect 21542 42100 21548 42112
rect 21600 42100 21606 42152
rect 18693 42075 18751 42081
rect 18693 42072 18705 42075
rect 17236 42044 18705 42072
rect 18693 42041 18705 42044
rect 18739 42041 18751 42075
rect 18693 42035 18751 42041
rect 18874 42032 18880 42084
rect 18932 42072 18938 42084
rect 20806 42072 20812 42084
rect 18932 42044 20812 42072
rect 18932 42032 18938 42044
rect 20806 42032 20812 42044
rect 20864 42032 20870 42084
rect 17313 42007 17371 42013
rect 17313 42004 17325 42007
rect 17144 41976 17325 42004
rect 17037 41967 17095 41973
rect 17313 41973 17325 41976
rect 17359 41973 17371 42007
rect 17313 41967 17371 41973
rect 17770 41964 17776 42016
rect 17828 42004 17834 42016
rect 19702 42004 19708 42016
rect 17828 41976 19708 42004
rect 17828 41964 17834 41976
rect 19702 41964 19708 41976
rect 19760 41964 19766 42016
rect 1104 41914 21896 41936
rect 1104 41862 3549 41914
rect 3601 41862 3613 41914
rect 3665 41862 3677 41914
rect 3729 41862 3741 41914
rect 3793 41862 3805 41914
rect 3857 41862 8747 41914
rect 8799 41862 8811 41914
rect 8863 41862 8875 41914
rect 8927 41862 8939 41914
rect 8991 41862 9003 41914
rect 9055 41862 13945 41914
rect 13997 41862 14009 41914
rect 14061 41862 14073 41914
rect 14125 41862 14137 41914
rect 14189 41862 14201 41914
rect 14253 41862 19143 41914
rect 19195 41862 19207 41914
rect 19259 41862 19271 41914
rect 19323 41862 19335 41914
rect 19387 41862 19399 41914
rect 19451 41862 21896 41914
rect 1104 41840 21896 41862
rect 2682 41760 2688 41812
rect 2740 41800 2746 41812
rect 3145 41803 3203 41809
rect 2740 41760 2774 41800
rect 3145 41769 3157 41803
rect 3191 41800 3203 41803
rect 3326 41800 3332 41812
rect 3191 41772 3332 41800
rect 3191 41769 3203 41772
rect 3145 41763 3203 41769
rect 3326 41760 3332 41772
rect 3384 41760 3390 41812
rect 3789 41803 3847 41809
rect 3789 41769 3801 41803
rect 3835 41800 3847 41803
rect 3878 41800 3884 41812
rect 3835 41772 3884 41800
rect 3835 41769 3847 41772
rect 3789 41763 3847 41769
rect 3878 41760 3884 41772
rect 3936 41760 3942 41812
rect 3970 41760 3976 41812
rect 4028 41800 4034 41812
rect 4341 41803 4399 41809
rect 4341 41800 4353 41803
rect 4028 41772 4353 41800
rect 4028 41760 4034 41772
rect 4341 41769 4353 41772
rect 4387 41769 4399 41803
rect 4341 41763 4399 41769
rect 4617 41803 4675 41809
rect 4617 41769 4629 41803
rect 4663 41800 4675 41803
rect 4706 41800 4712 41812
rect 4663 41772 4712 41800
rect 4663 41769 4675 41772
rect 4617 41763 4675 41769
rect 4706 41760 4712 41772
rect 4764 41760 4770 41812
rect 4893 41803 4951 41809
rect 4893 41769 4905 41803
rect 4939 41800 4951 41803
rect 5258 41800 5264 41812
rect 4939 41772 5264 41800
rect 4939 41769 4951 41772
rect 4893 41763 4951 41769
rect 5258 41760 5264 41772
rect 5316 41760 5322 41812
rect 5445 41803 5503 41809
rect 5445 41769 5457 41803
rect 5491 41800 5503 41803
rect 5491 41772 5672 41800
rect 5491 41769 5503 41772
rect 5445 41763 5503 41769
rect 2746 41732 2774 41760
rect 3421 41735 3479 41741
rect 3421 41732 3433 41735
rect 2746 41704 3433 41732
rect 3421 41701 3433 41704
rect 3467 41701 3479 41735
rect 3421 41695 3479 41701
rect 4062 41692 4068 41744
rect 4120 41692 4126 41744
rect 5169 41735 5227 41741
rect 5169 41701 5181 41735
rect 5215 41732 5227 41735
rect 5534 41732 5540 41744
rect 5215 41704 5540 41732
rect 5215 41701 5227 41704
rect 5169 41695 5227 41701
rect 5534 41692 5540 41704
rect 5592 41692 5598 41744
rect 5644 41732 5672 41772
rect 5718 41760 5724 41812
rect 5776 41760 5782 41812
rect 5902 41760 5908 41812
rect 5960 41760 5966 41812
rect 5997 41803 6055 41809
rect 5997 41769 6009 41803
rect 6043 41800 6055 41803
rect 6178 41800 6184 41812
rect 6043 41772 6184 41800
rect 6043 41769 6055 41772
rect 5997 41763 6055 41769
rect 6178 41760 6184 41772
rect 6236 41760 6242 41812
rect 6454 41760 6460 41812
rect 6512 41800 6518 41812
rect 6512 41772 7052 41800
rect 6512 41760 6518 41772
rect 5920 41732 5948 41760
rect 5644 41704 5948 41732
rect 6825 41735 6883 41741
rect 6825 41701 6837 41735
rect 6871 41701 6883 41735
rect 6825 41695 6883 41701
rect 6840 41664 6868 41695
rect 5644 41636 6868 41664
rect 750 41556 756 41608
rect 808 41596 814 41608
rect 1397 41599 1455 41605
rect 1397 41596 1409 41599
rect 808 41568 1409 41596
rect 808 41556 814 41568
rect 1397 41565 1409 41568
rect 1443 41565 1455 41599
rect 1397 41559 1455 41565
rect 1949 41599 2007 41605
rect 1949 41565 1961 41599
rect 1995 41596 2007 41599
rect 2958 41596 2964 41608
rect 1995 41568 2964 41596
rect 1995 41565 2007 41568
rect 1949 41559 2007 41565
rect 2958 41556 2964 41568
rect 3016 41556 3022 41608
rect 3329 41599 3387 41605
rect 3329 41565 3341 41599
rect 3375 41565 3387 41599
rect 3329 41559 3387 41565
rect 1486 41488 1492 41540
rect 1544 41528 1550 41540
rect 1673 41531 1731 41537
rect 1673 41528 1685 41531
rect 1544 41500 1685 41528
rect 1544 41488 1550 41500
rect 1673 41497 1685 41500
rect 1719 41497 1731 41531
rect 1673 41491 1731 41497
rect 2222 41488 2228 41540
rect 2280 41488 2286 41540
rect 3344 41528 3372 41559
rect 3602 41556 3608 41608
rect 3660 41556 3666 41608
rect 3970 41556 3976 41608
rect 4028 41556 4034 41608
rect 4246 41556 4252 41608
rect 4304 41556 4310 41608
rect 4522 41556 4528 41608
rect 4580 41556 4586 41608
rect 4798 41556 4804 41608
rect 4856 41556 4862 41608
rect 5077 41599 5135 41605
rect 5077 41565 5089 41599
rect 5123 41596 5135 41599
rect 5166 41596 5172 41608
rect 5123 41568 5172 41596
rect 5123 41565 5135 41568
rect 5077 41559 5135 41565
rect 5166 41556 5172 41568
rect 5224 41556 5230 41608
rect 5350 41556 5356 41608
rect 5408 41556 5414 41608
rect 5644 41605 5672 41636
rect 5629 41599 5687 41605
rect 5629 41565 5641 41599
rect 5675 41565 5687 41599
rect 5629 41559 5687 41565
rect 5902 41556 5908 41608
rect 5960 41556 5966 41608
rect 7024 41605 7052 41772
rect 7116 41772 7328 41800
rect 6181 41599 6239 41605
rect 6181 41565 6193 41599
rect 6227 41565 6239 41599
rect 6181 41559 6239 41565
rect 7009 41599 7067 41605
rect 7009 41565 7021 41599
rect 7055 41565 7067 41599
rect 7009 41559 7067 41565
rect 4154 41528 4160 41540
rect 3344 41500 4160 41528
rect 4154 41488 4160 41500
rect 4212 41488 4218 41540
rect 5258 41488 5264 41540
rect 5316 41528 5322 41540
rect 6196 41528 6224 41559
rect 5316 41500 6224 41528
rect 5316 41488 5322 41500
rect 4982 41420 4988 41472
rect 5040 41460 5046 41472
rect 7116 41460 7144 41772
rect 7193 41735 7251 41741
rect 7193 41701 7205 41735
rect 7239 41701 7251 41735
rect 7300 41732 7328 41772
rect 7374 41760 7380 41812
rect 7432 41800 7438 41812
rect 7745 41803 7803 41809
rect 7745 41800 7757 41803
rect 7432 41772 7757 41800
rect 7432 41760 7438 41772
rect 7745 41769 7757 41772
rect 7791 41769 7803 41803
rect 7745 41763 7803 41769
rect 7834 41760 7840 41812
rect 7892 41800 7898 41812
rect 8573 41803 8631 41809
rect 8573 41800 8585 41803
rect 7892 41772 8585 41800
rect 7892 41760 7898 41772
rect 8573 41769 8585 41772
rect 8619 41769 8631 41803
rect 12250 41800 12256 41812
rect 8573 41763 8631 41769
rect 8772 41772 12256 41800
rect 8772 41732 8800 41772
rect 12250 41760 12256 41772
rect 12308 41760 12314 41812
rect 13722 41760 13728 41812
rect 13780 41800 13786 41812
rect 14185 41803 14243 41809
rect 14185 41800 14197 41803
rect 13780 41772 14197 41800
rect 13780 41760 13786 41772
rect 14185 41769 14197 41772
rect 14231 41769 14243 41803
rect 15378 41800 15384 41812
rect 14185 41763 14243 41769
rect 15212 41772 15384 41800
rect 7300 41704 8800 41732
rect 8941 41735 8999 41741
rect 7193 41695 7251 41701
rect 8941 41701 8953 41735
rect 8987 41701 8999 41735
rect 8941 41695 8999 41701
rect 7208 41664 7236 41695
rect 7208 41636 7696 41664
rect 7374 41556 7380 41608
rect 7432 41556 7438 41608
rect 7668 41605 7696 41636
rect 7742 41624 7748 41676
rect 7800 41664 7806 41676
rect 8956 41664 8984 41695
rect 9122 41692 9128 41744
rect 9180 41732 9186 41744
rect 9180 41704 9996 41732
rect 9180 41692 9186 41704
rect 9306 41664 9312 41676
rect 7800 41636 8892 41664
rect 8956 41636 9312 41664
rect 7800 41624 7806 41636
rect 7653 41599 7711 41605
rect 7653 41565 7665 41599
rect 7699 41565 7711 41599
rect 7653 41559 7711 41565
rect 7929 41599 7987 41605
rect 7929 41565 7941 41599
rect 7975 41596 7987 41599
rect 7975 41568 8616 41596
rect 7975 41565 7987 41568
rect 7929 41559 7987 41565
rect 8113 41531 8171 41537
rect 8113 41528 8125 41531
rect 7484 41500 8125 41528
rect 7484 41469 7512 41500
rect 8113 41497 8125 41500
rect 8159 41497 8171 41531
rect 8113 41491 8171 41497
rect 8478 41488 8484 41540
rect 8536 41488 8542 41540
rect 8588 41528 8616 41568
rect 8662 41556 8668 41608
rect 8720 41596 8726 41608
rect 8757 41599 8815 41605
rect 8757 41596 8769 41599
rect 8720 41568 8769 41596
rect 8720 41556 8726 41568
rect 8757 41565 8769 41568
rect 8803 41565 8815 41599
rect 8864 41596 8892 41636
rect 9306 41624 9312 41636
rect 9364 41624 9370 41676
rect 9582 41624 9588 41676
rect 9640 41664 9646 41676
rect 9640 41636 9812 41664
rect 9640 41624 9646 41636
rect 9125 41599 9183 41605
rect 9125 41596 9137 41599
rect 8864 41568 9137 41596
rect 8757 41559 8815 41565
rect 9125 41565 9137 41568
rect 9171 41565 9183 41599
rect 9125 41559 9183 41565
rect 9398 41556 9404 41608
rect 9456 41605 9462 41608
rect 9456 41596 9467 41605
rect 9456 41568 9501 41596
rect 9456 41559 9467 41568
rect 9456 41556 9462 41559
rect 9674 41556 9680 41608
rect 9732 41556 9738 41608
rect 8588 41500 9536 41528
rect 5040 41432 7144 41460
rect 7469 41463 7527 41469
rect 5040 41420 5046 41432
rect 7469 41429 7481 41463
rect 7515 41429 7527 41463
rect 7469 41423 7527 41429
rect 7926 41420 7932 41472
rect 7984 41460 7990 41472
rect 8389 41463 8447 41469
rect 8389 41460 8401 41463
rect 7984 41432 8401 41460
rect 7984 41420 7990 41432
rect 8389 41429 8401 41432
rect 8435 41429 8447 41463
rect 8496 41460 8524 41488
rect 9508 41469 9536 41500
rect 9784 41469 9812 41636
rect 9968 41605 9996 41704
rect 13906 41624 13912 41676
rect 13964 41664 13970 41676
rect 15105 41667 15163 41673
rect 15105 41664 15117 41667
rect 13964 41636 15117 41664
rect 13964 41624 13970 41636
rect 15105 41633 15117 41636
rect 15151 41633 15163 41667
rect 15105 41627 15163 41633
rect 9953 41599 10011 41605
rect 9953 41565 9965 41599
rect 9999 41565 10011 41599
rect 9953 41559 10011 41565
rect 14366 41556 14372 41608
rect 14424 41556 14430 41608
rect 14553 41599 14611 41605
rect 14553 41565 14565 41599
rect 14599 41596 14611 41599
rect 15212 41596 15240 41772
rect 15378 41760 15384 41772
rect 15436 41760 15442 41812
rect 15933 41803 15991 41809
rect 15933 41769 15945 41803
rect 15979 41800 15991 41803
rect 16022 41800 16028 41812
rect 15979 41772 16028 41800
rect 15979 41769 15991 41772
rect 15933 41763 15991 41769
rect 16022 41760 16028 41772
rect 16080 41760 16086 41812
rect 16209 41803 16267 41809
rect 16209 41769 16221 41803
rect 16255 41800 16267 41803
rect 16758 41800 16764 41812
rect 16255 41772 16764 41800
rect 16255 41769 16267 41772
rect 16209 41763 16267 41769
rect 16758 41760 16764 41772
rect 16816 41760 16822 41812
rect 16942 41760 16948 41812
rect 17000 41760 17006 41812
rect 17052 41772 18368 41800
rect 16960 41732 16988 41760
rect 17052 41741 17080 41772
rect 15304 41704 16988 41732
rect 17037 41735 17095 41741
rect 15304 41605 15332 41704
rect 17037 41701 17049 41735
rect 17083 41701 17095 41735
rect 17037 41695 17095 41701
rect 17126 41692 17132 41744
rect 17184 41732 17190 41744
rect 17184 41704 17540 41732
rect 17184 41692 17190 41704
rect 15378 41624 15384 41676
rect 15436 41624 15442 41676
rect 15470 41624 15476 41676
rect 15528 41664 15534 41676
rect 17310 41664 17316 41676
rect 15528 41636 15792 41664
rect 15528 41624 15534 41636
rect 14599 41568 15240 41596
rect 15289 41599 15347 41605
rect 14599 41565 14611 41568
rect 14553 41559 14611 41565
rect 15289 41565 15301 41599
rect 15335 41565 15347 41599
rect 15396 41596 15424 41624
rect 15657 41599 15715 41605
rect 15657 41596 15669 41599
rect 15396 41568 15669 41596
rect 15289 41559 15347 41565
rect 15657 41565 15669 41568
rect 15703 41565 15715 41599
rect 15657 41559 15715 41565
rect 14921 41531 14979 41537
rect 14921 41497 14933 41531
rect 14967 41528 14979 41531
rect 15764 41528 15792 41636
rect 16592 41636 17316 41664
rect 16125 41595 16183 41601
rect 16125 41561 16137 41595
rect 16171 41592 16183 41595
rect 16298 41592 16304 41608
rect 16171 41564 16304 41592
rect 16171 41561 16183 41564
rect 16125 41555 16183 41561
rect 16298 41556 16304 41564
rect 16356 41556 16362 41608
rect 16393 41599 16451 41605
rect 16393 41565 16405 41599
rect 16439 41596 16451 41599
rect 16592 41596 16620 41636
rect 17310 41624 17316 41636
rect 17368 41624 17374 41676
rect 17402 41624 17408 41676
rect 17460 41624 17466 41676
rect 17512 41664 17540 41704
rect 17586 41692 17592 41744
rect 17644 41692 17650 41744
rect 17862 41692 17868 41744
rect 17920 41692 17926 41744
rect 18340 41732 18368 41772
rect 18414 41760 18420 41812
rect 18472 41800 18478 41812
rect 18693 41803 18751 41809
rect 18693 41800 18705 41803
rect 18472 41772 18705 41800
rect 18472 41760 18478 41772
rect 18693 41769 18705 41772
rect 18739 41769 18751 41803
rect 18693 41763 18751 41769
rect 19260 41772 20484 41800
rect 18874 41732 18880 41744
rect 18340 41704 18880 41732
rect 18874 41692 18880 41704
rect 18932 41692 18938 41744
rect 17512 41636 17908 41664
rect 16439 41568 16620 41596
rect 16439 41565 16451 41568
rect 16393 41559 16451 41565
rect 16666 41556 16672 41608
rect 16724 41556 16730 41608
rect 16942 41556 16948 41608
rect 17000 41556 17006 41608
rect 17218 41556 17224 41608
rect 17276 41556 17282 41608
rect 17420 41596 17448 41624
rect 17880 41612 17908 41636
rect 18414 41624 18420 41676
rect 18472 41624 18478 41676
rect 19260 41664 19288 41772
rect 19334 41692 19340 41744
rect 19392 41732 19398 41744
rect 20073 41735 20131 41741
rect 20073 41732 20085 41735
rect 19392 41704 20085 41732
rect 19392 41692 19398 41704
rect 20073 41701 20085 41704
rect 20119 41701 20131 41735
rect 20456 41732 20484 41772
rect 20530 41760 20536 41812
rect 20588 41760 20594 41812
rect 20901 41803 20959 41809
rect 20901 41769 20913 41803
rect 20947 41800 20959 41803
rect 21910 41800 21916 41812
rect 20947 41772 21916 41800
rect 20947 41769 20959 41772
rect 20901 41763 20959 41769
rect 21910 41760 21916 41772
rect 21968 41760 21974 41812
rect 21450 41732 21456 41744
rect 20456 41704 21456 41732
rect 20073 41695 20131 41701
rect 21450 41692 21456 41704
rect 21508 41692 21514 41744
rect 22646 41664 22652 41676
rect 18616 41636 19288 41664
rect 19444 41636 22652 41664
rect 18049 41615 18107 41621
rect 18049 41612 18061 41615
rect 17328 41568 17448 41596
rect 17497 41599 17555 41605
rect 14967 41500 15792 41528
rect 16500 41500 17080 41528
rect 14967 41497 14979 41500
rect 14921 41491 14979 41497
rect 9217 41463 9275 41469
rect 9217 41460 9229 41463
rect 8496 41432 9229 41460
rect 8389 41423 8447 41429
rect 9217 41429 9229 41432
rect 9263 41429 9275 41463
rect 9217 41423 9275 41429
rect 9493 41463 9551 41469
rect 9493 41429 9505 41463
rect 9539 41429 9551 41463
rect 9493 41423 9551 41429
rect 9769 41463 9827 41469
rect 9769 41429 9781 41463
rect 9815 41429 9827 41463
rect 9769 41423 9827 41429
rect 9858 41420 9864 41472
rect 9916 41460 9922 41472
rect 12526 41460 12532 41472
rect 9916 41432 12532 41460
rect 9916 41420 9922 41432
rect 12526 41420 12532 41432
rect 12584 41420 12590 41472
rect 14182 41420 14188 41472
rect 14240 41460 14246 41472
rect 14645 41463 14703 41469
rect 14645 41460 14657 41463
rect 14240 41432 14657 41460
rect 14240 41420 14246 41432
rect 14645 41429 14657 41432
rect 14691 41429 14703 41463
rect 14645 41423 14703 41429
rect 14826 41420 14832 41472
rect 14884 41460 14890 41472
rect 15194 41460 15200 41472
rect 14884 41432 15200 41460
rect 14884 41420 14890 41432
rect 15194 41420 15200 41432
rect 15252 41420 15258 41472
rect 15378 41420 15384 41472
rect 15436 41420 15442 41472
rect 15470 41420 15476 41472
rect 15528 41460 15534 41472
rect 16500 41469 16528 41500
rect 17052 41472 17080 41500
rect 15749 41463 15807 41469
rect 15749 41460 15761 41463
rect 15528 41432 15761 41460
rect 15528 41420 15534 41432
rect 15749 41429 15761 41432
rect 15795 41429 15807 41463
rect 15749 41423 15807 41429
rect 16485 41463 16543 41469
rect 16485 41429 16497 41463
rect 16531 41429 16543 41463
rect 16485 41423 16543 41429
rect 16761 41463 16819 41469
rect 16761 41429 16773 41463
rect 16807 41460 16819 41463
rect 16850 41460 16856 41472
rect 16807 41432 16856 41460
rect 16807 41429 16819 41432
rect 16761 41423 16819 41429
rect 16850 41420 16856 41432
rect 16908 41420 16914 41472
rect 17034 41420 17040 41472
rect 17092 41420 17098 41472
rect 17328 41469 17356 41568
rect 17497 41565 17509 41599
rect 17543 41565 17555 41599
rect 17497 41559 17555 41565
rect 17402 41488 17408 41540
rect 17460 41528 17466 41540
rect 17512 41528 17540 41559
rect 17770 41556 17776 41608
rect 17828 41556 17834 41608
rect 17880 41584 18061 41612
rect 18049 41581 18061 41584
rect 18095 41581 18107 41615
rect 18049 41575 18107 41581
rect 18322 41556 18328 41608
rect 18380 41556 18386 41608
rect 17460 41500 17540 41528
rect 18432 41528 18460 41624
rect 18616 41605 18644 41636
rect 19444 41605 19472 41636
rect 22646 41624 22652 41636
rect 22704 41624 22710 41676
rect 18601 41599 18659 41605
rect 18601 41565 18613 41599
rect 18647 41565 18659 41599
rect 18601 41559 18659 41565
rect 18877 41599 18935 41605
rect 18877 41565 18889 41599
rect 18923 41565 18935 41599
rect 18877 41559 18935 41565
rect 19429 41599 19487 41605
rect 19429 41565 19441 41599
rect 19475 41565 19487 41599
rect 19429 41559 19487 41565
rect 18892 41528 18920 41559
rect 19794 41556 19800 41608
rect 19852 41556 19858 41608
rect 20257 41599 20315 41605
rect 20257 41565 20269 41599
rect 20303 41565 20315 41599
rect 20257 41559 20315 41565
rect 19812 41528 19840 41556
rect 18432 41500 18920 41528
rect 19352 41500 19840 41528
rect 17460 41488 17466 41500
rect 17313 41463 17371 41469
rect 17313 41429 17325 41463
rect 17359 41429 17371 41463
rect 17313 41423 17371 41429
rect 18141 41463 18199 41469
rect 18141 41429 18153 41463
rect 18187 41460 18199 41463
rect 18230 41460 18236 41472
rect 18187 41432 18236 41460
rect 18187 41429 18199 41432
rect 18141 41423 18199 41429
rect 18230 41420 18236 41432
rect 18288 41420 18294 41472
rect 18414 41420 18420 41472
rect 18472 41420 18478 41472
rect 19245 41463 19303 41469
rect 19245 41429 19257 41463
rect 19291 41460 19303 41463
rect 19352 41460 19380 41500
rect 19291 41432 19380 41460
rect 19797 41463 19855 41469
rect 19291 41429 19303 41432
rect 19245 41423 19303 41429
rect 19797 41429 19809 41463
rect 19843 41460 19855 41463
rect 20272 41460 20300 41559
rect 20346 41556 20352 41608
rect 20404 41556 20410 41608
rect 20717 41599 20775 41605
rect 20717 41565 20729 41599
rect 20763 41596 20775 41599
rect 21082 41596 21088 41608
rect 20763 41568 21088 41596
rect 20763 41565 20775 41568
rect 20717 41559 20775 41565
rect 21082 41556 21088 41568
rect 21140 41556 21146 41608
rect 21174 41488 21180 41540
rect 21232 41488 21238 41540
rect 21545 41531 21603 41537
rect 21545 41497 21557 41531
rect 21591 41528 21603 41531
rect 22278 41528 22284 41540
rect 21591 41500 22284 41528
rect 21591 41497 21603 41500
rect 21545 41491 21603 41497
rect 22278 41488 22284 41500
rect 22336 41488 22342 41540
rect 22554 41460 22560 41472
rect 19843 41432 22560 41460
rect 19843 41429 19855 41432
rect 19797 41423 19855 41429
rect 22554 41420 22560 41432
rect 22612 41420 22618 41472
rect 1104 41370 22056 41392
rect 1104 41318 6148 41370
rect 6200 41318 6212 41370
rect 6264 41318 6276 41370
rect 6328 41318 6340 41370
rect 6392 41318 6404 41370
rect 6456 41318 11346 41370
rect 11398 41318 11410 41370
rect 11462 41318 11474 41370
rect 11526 41318 11538 41370
rect 11590 41318 11602 41370
rect 11654 41318 16544 41370
rect 16596 41318 16608 41370
rect 16660 41318 16672 41370
rect 16724 41318 16736 41370
rect 16788 41318 16800 41370
rect 16852 41318 21742 41370
rect 21794 41318 21806 41370
rect 21858 41318 21870 41370
rect 21922 41318 21934 41370
rect 21986 41318 21998 41370
rect 22050 41318 22056 41370
rect 1104 41296 22056 41318
rect 2498 41216 2504 41268
rect 2556 41256 2562 41268
rect 3973 41259 4031 41265
rect 3973 41256 3985 41259
rect 2556 41228 3985 41256
rect 2556 41216 2562 41228
rect 3973 41225 3985 41228
rect 4019 41225 4031 41259
rect 3973 41219 4031 41225
rect 4890 41216 4896 41268
rect 4948 41256 4954 41268
rect 5169 41259 5227 41265
rect 5169 41256 5181 41259
rect 4948 41228 5181 41256
rect 4948 41216 4954 41228
rect 5169 41225 5181 41228
rect 5215 41225 5227 41259
rect 5169 41219 5227 41225
rect 5445 41259 5503 41265
rect 5445 41225 5457 41259
rect 5491 41225 5503 41259
rect 5445 41219 5503 41225
rect 5721 41259 5779 41265
rect 5721 41225 5733 41259
rect 5767 41225 5779 41259
rect 5721 41219 5779 41225
rect 2225 41191 2283 41197
rect 2225 41157 2237 41191
rect 2271 41188 2283 41191
rect 4706 41188 4712 41200
rect 2271 41160 4712 41188
rect 2271 41157 2283 41160
rect 2225 41151 2283 41157
rect 4706 41148 4712 41160
rect 4764 41148 4770 41200
rect 5074 41148 5080 41200
rect 5132 41188 5138 41200
rect 5460 41188 5488 41219
rect 5132 41160 5488 41188
rect 5736 41188 5764 41219
rect 5994 41216 6000 41268
rect 6052 41216 6058 41268
rect 6730 41256 6736 41268
rect 6104 41228 6736 41256
rect 6104 41188 6132 41228
rect 6730 41216 6736 41228
rect 6788 41216 6794 41268
rect 8113 41259 8171 41265
rect 8113 41256 8125 41259
rect 6840 41228 8125 41256
rect 6840 41188 6868 41228
rect 8113 41225 8125 41228
rect 8159 41225 8171 41259
rect 8113 41219 8171 41225
rect 8386 41216 8392 41268
rect 8444 41216 8450 41268
rect 14642 41216 14648 41268
rect 14700 41216 14706 41268
rect 14921 41259 14979 41265
rect 14921 41225 14933 41259
rect 14967 41256 14979 41259
rect 15010 41256 15016 41268
rect 14967 41228 15016 41256
rect 14967 41225 14979 41228
rect 14921 41219 14979 41225
rect 15010 41216 15016 41228
rect 15068 41216 15074 41268
rect 15197 41259 15255 41265
rect 15197 41225 15209 41259
rect 15243 41256 15255 41259
rect 15562 41256 15568 41268
rect 15243 41228 15568 41256
rect 15243 41225 15255 41228
rect 15197 41219 15255 41225
rect 15562 41216 15568 41228
rect 15620 41216 15626 41268
rect 15933 41259 15991 41265
rect 15933 41225 15945 41259
rect 15979 41256 15991 41259
rect 17310 41256 17316 41268
rect 15979 41228 17316 41256
rect 15979 41225 15991 41228
rect 15933 41219 15991 41225
rect 17310 41216 17316 41228
rect 17368 41216 17374 41268
rect 17405 41259 17463 41265
rect 17405 41225 17417 41259
rect 17451 41225 17463 41259
rect 17405 41219 17463 41225
rect 5736 41160 6132 41188
rect 6196 41160 6868 41188
rect 5132 41148 5138 41160
rect 1210 41080 1216 41132
rect 1268 41120 1274 41132
rect 1397 41123 1455 41129
rect 1397 41120 1409 41123
rect 1268 41092 1409 41120
rect 1268 41080 1274 41092
rect 1397 41089 1409 41092
rect 1443 41089 1455 41123
rect 1397 41083 1455 41089
rect 1949 41123 2007 41129
rect 1949 41089 1961 41123
rect 1995 41089 2007 41123
rect 1949 41083 2007 41089
rect 2501 41123 2559 41129
rect 2501 41089 2513 41123
rect 2547 41120 2559 41123
rect 2774 41120 2780 41132
rect 2547 41092 2780 41120
rect 2547 41089 2559 41092
rect 2501 41083 2559 41089
rect 1578 41012 1584 41064
rect 1636 41012 1642 41064
rect 1964 40984 1992 41083
rect 2774 41080 2780 41092
rect 2832 41080 2838 41132
rect 4154 41080 4160 41132
rect 4212 41080 4218 41132
rect 4893 41123 4951 41129
rect 4893 41089 4905 41123
rect 4939 41120 4951 41123
rect 5258 41120 5264 41132
rect 4939 41092 5264 41120
rect 4939 41089 4951 41092
rect 4893 41083 4951 41089
rect 5258 41080 5264 41092
rect 5316 41120 5322 41132
rect 5353 41123 5411 41129
rect 5353 41120 5365 41123
rect 5316 41092 5365 41120
rect 5316 41080 5322 41092
rect 5353 41089 5365 41092
rect 5399 41089 5411 41123
rect 5353 41083 5411 41089
rect 5629 41123 5687 41129
rect 5629 41089 5641 41123
rect 5675 41089 5687 41123
rect 5629 41083 5687 41089
rect 2685 41055 2743 41061
rect 2685 41021 2697 41055
rect 2731 41052 2743 41055
rect 4062 41052 4068 41064
rect 2731 41024 4068 41052
rect 2731 41021 2743 41024
rect 2685 41015 2743 41021
rect 4062 41012 4068 41024
rect 4120 41012 4126 41064
rect 5644 41052 5672 41083
rect 5718 41080 5724 41132
rect 5776 41120 5782 41132
rect 6196 41129 6224 41160
rect 7650 41148 7656 41200
rect 7708 41188 7714 41200
rect 7708 41160 11192 41188
rect 7708 41148 7714 41160
rect 11164 41132 11192 41160
rect 14274 41148 14280 41200
rect 14332 41188 14338 41200
rect 14332 41160 15148 41188
rect 14332 41148 14338 41160
rect 5905 41123 5963 41129
rect 5905 41120 5917 41123
rect 5776 41092 5917 41120
rect 5776 41080 5782 41092
rect 5905 41089 5917 41092
rect 5951 41089 5963 41123
rect 5905 41083 5963 41089
rect 6181 41123 6239 41129
rect 6181 41089 6193 41123
rect 6227 41089 6239 41123
rect 6181 41083 6239 41089
rect 6546 41080 6552 41132
rect 6604 41080 6610 41132
rect 6917 41123 6975 41129
rect 6917 41089 6929 41123
rect 6963 41120 6975 41123
rect 7193 41123 7251 41129
rect 7193 41120 7205 41123
rect 6963 41092 7205 41120
rect 6963 41089 6975 41092
rect 6917 41083 6975 41089
rect 7193 41089 7205 41092
rect 7239 41120 7251 41123
rect 7282 41120 7288 41132
rect 7239 41092 7288 41120
rect 7239 41089 7251 41092
rect 7193 41083 7251 41089
rect 7282 41080 7288 41092
rect 7340 41080 7346 41132
rect 7469 41123 7527 41129
rect 7469 41089 7481 41123
rect 7515 41089 7527 41123
rect 8297 41123 8355 41129
rect 8297 41120 8309 41123
rect 7469 41083 7527 41089
rect 7760 41092 8309 41120
rect 7484 41052 7512 41083
rect 7760 41064 7788 41092
rect 8297 41089 8309 41092
rect 8343 41089 8355 41123
rect 8297 41083 8355 41089
rect 8570 41080 8576 41132
rect 8628 41080 8634 41132
rect 11146 41080 11152 41132
rect 11204 41080 11210 41132
rect 14550 41080 14556 41132
rect 14608 41120 14614 41132
rect 15120 41129 15148 41160
rect 15470 41148 15476 41200
rect 15528 41188 15534 41200
rect 15528 41160 16252 41188
rect 15528 41148 15534 41160
rect 14829 41123 14887 41129
rect 14829 41120 14841 41123
rect 14608 41092 14841 41120
rect 14608 41080 14614 41092
rect 14829 41089 14841 41092
rect 14875 41089 14887 41123
rect 14829 41083 14887 41089
rect 15105 41123 15163 41129
rect 15105 41089 15117 41123
rect 15151 41089 15163 41123
rect 15105 41083 15163 41089
rect 15194 41080 15200 41132
rect 15252 41120 15258 41132
rect 15381 41123 15439 41129
rect 15381 41120 15393 41123
rect 15252 41092 15393 41120
rect 15252 41080 15258 41092
rect 15381 41089 15393 41092
rect 15427 41089 15439 41123
rect 15381 41083 15439 41089
rect 15657 41123 15715 41129
rect 15657 41089 15669 41123
rect 15703 41089 15715 41123
rect 15657 41083 15715 41089
rect 5644 41024 6960 41052
rect 2866 40984 2872 40996
rect 1964 40956 2872 40984
rect 2866 40944 2872 40956
rect 2924 40944 2930 40996
rect 5902 40944 5908 40996
rect 5960 40984 5966 40996
rect 6365 40987 6423 40993
rect 6365 40984 6377 40987
rect 5960 40956 6377 40984
rect 5960 40944 5966 40956
rect 6365 40953 6377 40956
rect 6411 40953 6423 40987
rect 6365 40947 6423 40953
rect 6932 40916 6960 41024
rect 7024 41024 7512 41052
rect 7024 40993 7052 41024
rect 7742 41012 7748 41064
rect 7800 41012 7806 41064
rect 14734 41012 14740 41064
rect 14792 41052 14798 41064
rect 15672 41052 15700 41083
rect 15838 41080 15844 41132
rect 15896 41120 15902 41132
rect 16117 41123 16175 41129
rect 16117 41120 16129 41123
rect 15896 41092 16129 41120
rect 15896 41080 15902 41092
rect 16117 41089 16129 41092
rect 16163 41089 16175 41123
rect 16224 41120 16252 41160
rect 16390 41148 16396 41200
rect 16448 41188 16454 41200
rect 16448 41160 17172 41188
rect 16448 41148 16454 41160
rect 16485 41123 16543 41129
rect 16485 41120 16497 41123
rect 16224 41092 16497 41120
rect 16117 41083 16175 41089
rect 16485 41089 16497 41092
rect 16531 41089 16543 41123
rect 16485 41083 16543 41089
rect 16850 41080 16856 41132
rect 16908 41080 16914 41132
rect 17144 41129 17172 41160
rect 17129 41123 17187 41129
rect 17129 41089 17141 41123
rect 17175 41089 17187 41123
rect 17129 41083 17187 41089
rect 17221 41123 17279 41129
rect 17221 41089 17233 41123
rect 17267 41120 17279 41123
rect 17310 41120 17316 41132
rect 17267 41092 17316 41120
rect 17267 41089 17279 41092
rect 17221 41083 17279 41089
rect 17310 41080 17316 41092
rect 17368 41080 17374 41132
rect 14792 41024 15700 41052
rect 14792 41012 14798 41024
rect 16574 41012 16580 41064
rect 16632 41052 16638 41064
rect 17420 41052 17448 41219
rect 17586 41216 17592 41268
rect 17644 41216 17650 41268
rect 17681 41259 17739 41265
rect 17681 41225 17693 41259
rect 17727 41256 17739 41259
rect 17862 41256 17868 41268
rect 17727 41228 17868 41256
rect 17727 41225 17739 41228
rect 17681 41219 17739 41225
rect 17862 41216 17868 41228
rect 17920 41216 17926 41268
rect 17954 41216 17960 41268
rect 18012 41256 18018 41268
rect 18233 41259 18291 41265
rect 18233 41256 18245 41259
rect 18012 41228 18245 41256
rect 18012 41216 18018 41228
rect 18233 41225 18245 41228
rect 18279 41225 18291 41259
rect 18233 41219 18291 41225
rect 18690 41216 18696 41268
rect 18748 41216 18754 41268
rect 18782 41216 18788 41268
rect 18840 41256 18846 41268
rect 19058 41256 19064 41268
rect 18840 41228 19064 41256
rect 18840 41216 18846 41228
rect 19058 41216 19064 41228
rect 19116 41216 19122 41268
rect 19429 41259 19487 41265
rect 19429 41256 19441 41259
rect 19306 41228 19441 41256
rect 17604 41188 17632 41216
rect 17604 41160 18000 41188
rect 17972 41144 18000 41160
rect 18141 41147 18199 41153
rect 18141 41144 18153 41147
rect 17586 41080 17592 41132
rect 17644 41120 17650 41132
rect 17865 41123 17923 41129
rect 17865 41120 17877 41123
rect 17644 41092 17877 41120
rect 17644 41080 17650 41092
rect 17865 41089 17877 41092
rect 17911 41089 17923 41123
rect 17972 41116 18153 41144
rect 18141 41113 18153 41116
rect 18187 41113 18199 41147
rect 18141 41107 18199 41113
rect 17865 41083 17923 41089
rect 18230 41080 18236 41132
rect 18288 41120 18294 41132
rect 18417 41123 18475 41129
rect 18417 41120 18429 41123
rect 18288 41092 18429 41120
rect 18288 41080 18294 41092
rect 18417 41089 18429 41092
rect 18463 41089 18475 41123
rect 18417 41083 18475 41089
rect 16632 41024 17448 41052
rect 16632 41012 16638 41024
rect 17494 41012 17500 41064
rect 17552 41012 17558 41064
rect 17678 41012 17684 41064
rect 17736 41012 17742 41064
rect 18708 41052 18736 41216
rect 19306 41188 19334 41228
rect 19429 41225 19441 41228
rect 19475 41225 19487 41259
rect 19429 41219 19487 41225
rect 19702 41216 19708 41268
rect 19760 41256 19766 41268
rect 20257 41259 20315 41265
rect 20257 41256 20269 41259
rect 19760 41228 20269 41256
rect 19760 41216 19766 41228
rect 20257 41225 20269 41228
rect 20303 41225 20315 41259
rect 20257 41219 20315 41225
rect 20809 41259 20867 41265
rect 20809 41225 20821 41259
rect 20855 41256 20867 41259
rect 21542 41256 21548 41268
rect 20855 41228 21548 41256
rect 20855 41225 20867 41228
rect 20809 41219 20867 41225
rect 21542 41216 21548 41228
rect 21600 41216 21606 41268
rect 18800 41160 19334 41188
rect 18800 41129 18828 41160
rect 18785 41123 18843 41129
rect 18785 41089 18797 41123
rect 18831 41089 18843 41123
rect 18785 41083 18843 41089
rect 19058 41080 19064 41132
rect 19116 41080 19122 41132
rect 19337 41107 19395 41113
rect 19337 41073 19349 41107
rect 19383 41104 19395 41107
rect 19383 41076 19472 41104
rect 19518 41080 19524 41132
rect 19576 41120 19582 41132
rect 19613 41123 19671 41129
rect 19613 41120 19625 41123
rect 19576 41092 19625 41120
rect 19576 41080 19582 41092
rect 19613 41089 19625 41092
rect 19659 41089 19671 41123
rect 19613 41083 19671 41089
rect 19886 41080 19892 41132
rect 19944 41080 19950 41132
rect 20162 41080 20168 41132
rect 20220 41080 20226 41132
rect 20438 41080 20444 41132
rect 20496 41080 20502 41132
rect 20717 41123 20775 41129
rect 20717 41089 20729 41123
rect 20763 41089 20775 41123
rect 20717 41083 20775 41089
rect 19383 41073 19395 41076
rect 19337 41067 19395 41073
rect 17880 41024 18736 41052
rect 7009 40987 7067 40993
rect 7009 40953 7021 40987
rect 7055 40953 7067 40987
rect 7009 40947 7067 40953
rect 7285 40987 7343 40993
rect 7285 40953 7297 40987
rect 7331 40984 7343 40987
rect 7374 40984 7380 40996
rect 7331 40956 7380 40984
rect 7331 40953 7343 40956
rect 7285 40947 7343 40953
rect 7374 40944 7380 40956
rect 7432 40944 7438 40996
rect 11054 40984 11060 40996
rect 7668 40956 11060 40984
rect 7668 40916 7696 40956
rect 11054 40944 11060 40956
rect 11112 40944 11118 40996
rect 15473 40987 15531 40993
rect 15473 40953 15485 40987
rect 15519 40984 15531 40987
rect 16114 40984 16120 40996
rect 15519 40956 16120 40984
rect 15519 40953 15531 40956
rect 15473 40947 15531 40953
rect 16114 40944 16120 40956
rect 16172 40944 16178 40996
rect 16669 40987 16727 40993
rect 16669 40953 16681 40987
rect 16715 40984 16727 40987
rect 17218 40984 17224 40996
rect 16715 40956 17224 40984
rect 16715 40953 16727 40956
rect 16669 40947 16727 40953
rect 17218 40944 17224 40956
rect 17276 40944 17282 40996
rect 17512 40984 17540 41012
rect 17328 40956 17540 40984
rect 6932 40888 7696 40916
rect 7742 40876 7748 40928
rect 7800 40876 7806 40928
rect 16301 40919 16359 40925
rect 16301 40885 16313 40919
rect 16347 40916 16359 40919
rect 16758 40916 16764 40928
rect 16347 40888 16764 40916
rect 16347 40885 16359 40888
rect 16301 40879 16359 40885
rect 16758 40876 16764 40888
rect 16816 40876 16822 40928
rect 16945 40919 17003 40925
rect 16945 40885 16957 40919
rect 16991 40916 17003 40919
rect 17328 40916 17356 40956
rect 16991 40888 17356 40916
rect 17696 40916 17724 41012
rect 17880 40996 17908 41024
rect 17862 40944 17868 40996
rect 17920 40944 17926 40996
rect 18690 40944 18696 40996
rect 18748 40984 18754 40996
rect 19153 40987 19211 40993
rect 18748 40956 19012 40984
rect 18748 40944 18754 40956
rect 17957 40919 18015 40925
rect 17957 40916 17969 40919
rect 17696 40888 17969 40916
rect 16991 40885 17003 40888
rect 16945 40879 17003 40885
rect 17957 40885 17969 40888
rect 18003 40885 18015 40919
rect 17957 40879 18015 40885
rect 18601 40919 18659 40925
rect 18601 40885 18613 40919
rect 18647 40916 18659 40919
rect 18782 40916 18788 40928
rect 18647 40888 18788 40916
rect 18647 40885 18659 40888
rect 18601 40879 18659 40885
rect 18782 40876 18788 40888
rect 18840 40876 18846 40928
rect 18874 40876 18880 40928
rect 18932 40876 18938 40928
rect 18984 40916 19012 40956
rect 19153 40953 19165 40987
rect 19199 40984 19211 40987
rect 19334 40984 19340 40996
rect 19199 40956 19340 40984
rect 19199 40953 19211 40956
rect 19153 40947 19211 40953
rect 19334 40944 19340 40956
rect 19392 40944 19398 40996
rect 19444 40984 19472 41076
rect 19978 41012 19984 41064
rect 20036 41052 20042 41064
rect 20732 41052 20760 41083
rect 20806 41080 20812 41132
rect 20864 41120 20870 41132
rect 20993 41123 21051 41129
rect 20993 41120 21005 41123
rect 20864 41092 21005 41120
rect 20864 41080 20870 41092
rect 20993 41089 21005 41092
rect 21039 41089 21051 41123
rect 20993 41083 21051 41089
rect 21266 41080 21272 41132
rect 21324 41080 21330 41132
rect 21634 41052 21640 41064
rect 20036 41024 20668 41052
rect 20732 41024 21640 41052
rect 20036 41012 20042 41024
rect 20533 40987 20591 40993
rect 20533 40984 20545 40987
rect 19444 40956 20545 40984
rect 20533 40953 20545 40956
rect 20579 40953 20591 40987
rect 20640 40984 20668 41024
rect 21634 41012 21640 41024
rect 21692 41012 21698 41064
rect 20898 40984 20904 40996
rect 20640 40956 20904 40984
rect 20533 40947 20591 40953
rect 20898 40944 20904 40956
rect 20956 40944 20962 40996
rect 20990 40944 20996 40996
rect 21048 40944 21054 40996
rect 19705 40919 19763 40925
rect 19705 40916 19717 40919
rect 18984 40888 19717 40916
rect 19705 40885 19717 40888
rect 19751 40885 19763 40919
rect 19705 40879 19763 40885
rect 19981 40919 20039 40925
rect 19981 40885 19993 40919
rect 20027 40916 20039 40919
rect 21008 40916 21036 40944
rect 20027 40888 21036 40916
rect 21453 40919 21511 40925
rect 20027 40885 20039 40888
rect 19981 40879 20039 40885
rect 21453 40885 21465 40919
rect 21499 40916 21511 40919
rect 22186 40916 22192 40928
rect 21499 40888 22192 40916
rect 21499 40885 21511 40888
rect 21453 40879 21511 40885
rect 22186 40876 22192 40888
rect 22244 40876 22250 40928
rect 1104 40826 21896 40848
rect 1104 40774 3549 40826
rect 3601 40774 3613 40826
rect 3665 40774 3677 40826
rect 3729 40774 3741 40826
rect 3793 40774 3805 40826
rect 3857 40774 8747 40826
rect 8799 40774 8811 40826
rect 8863 40774 8875 40826
rect 8927 40774 8939 40826
rect 8991 40774 9003 40826
rect 9055 40774 13945 40826
rect 13997 40774 14009 40826
rect 14061 40774 14073 40826
rect 14125 40774 14137 40826
rect 14189 40774 14201 40826
rect 14253 40774 19143 40826
rect 19195 40774 19207 40826
rect 19259 40774 19271 40826
rect 19323 40774 19335 40826
rect 19387 40774 19399 40826
rect 19451 40774 21896 40826
rect 1104 40752 21896 40774
rect 5442 40672 5448 40724
rect 5500 40672 5506 40724
rect 7101 40715 7159 40721
rect 7101 40681 7113 40715
rect 7147 40712 7159 40715
rect 8570 40712 8576 40724
rect 7147 40684 8576 40712
rect 7147 40681 7159 40684
rect 7101 40675 7159 40681
rect 8570 40672 8576 40684
rect 8628 40672 8634 40724
rect 16206 40672 16212 40724
rect 16264 40712 16270 40724
rect 19061 40715 19119 40721
rect 19061 40712 19073 40715
rect 16264 40684 19073 40712
rect 16264 40672 16270 40684
rect 19061 40681 19073 40684
rect 19107 40681 19119 40715
rect 19705 40715 19763 40721
rect 19705 40712 19717 40715
rect 19061 40675 19119 40681
rect 19536 40684 19717 40712
rect 1946 40604 1952 40656
rect 2004 40644 2010 40656
rect 4338 40644 4344 40656
rect 2004 40616 4344 40644
rect 2004 40604 2010 40616
rect 4338 40604 4344 40616
rect 4396 40604 4402 40656
rect 7466 40604 7472 40656
rect 7524 40644 7530 40656
rect 7742 40644 7748 40656
rect 7524 40616 7748 40644
rect 7524 40604 7530 40616
rect 7742 40604 7748 40616
rect 7800 40604 7806 40656
rect 17126 40604 17132 40656
rect 17184 40604 17190 40656
rect 17494 40604 17500 40656
rect 17552 40604 17558 40656
rect 17773 40647 17831 40653
rect 17773 40613 17785 40647
rect 17819 40644 17831 40647
rect 17862 40644 17868 40656
rect 17819 40616 17868 40644
rect 17819 40613 17831 40616
rect 17773 40607 17831 40613
rect 17862 40604 17868 40616
rect 17920 40604 17926 40656
rect 18325 40647 18383 40653
rect 18325 40613 18337 40647
rect 18371 40644 18383 40647
rect 19426 40644 19432 40656
rect 18371 40616 19432 40644
rect 18371 40613 18383 40616
rect 18325 40607 18383 40613
rect 19426 40604 19432 40616
rect 19484 40604 19490 40656
rect 7374 40536 7380 40588
rect 7432 40576 7438 40588
rect 8202 40576 8208 40588
rect 7432 40548 8208 40576
rect 7432 40536 7438 40548
rect 8202 40536 8208 40548
rect 8260 40536 8266 40588
rect 17144 40576 17172 40604
rect 19536 40576 19564 40684
rect 19705 40681 19717 40684
rect 19751 40681 19763 40715
rect 19705 40675 19763 40681
rect 20438 40672 20444 40724
rect 20496 40712 20502 40724
rect 20714 40712 20720 40724
rect 20496 40684 20720 40712
rect 20496 40672 20502 40684
rect 20714 40672 20720 40684
rect 20772 40672 20778 40724
rect 20809 40715 20867 40721
rect 20809 40681 20821 40715
rect 20855 40712 20867 40715
rect 21266 40712 21272 40724
rect 20855 40684 21272 40712
rect 20855 40681 20867 40684
rect 20809 40675 20867 40681
rect 21266 40672 21272 40684
rect 21324 40672 21330 40724
rect 19794 40604 19800 40656
rect 19852 40644 19858 40656
rect 19981 40647 20039 40653
rect 19852 40616 19932 40644
rect 19852 40604 19858 40616
rect 17144 40548 18920 40576
rect 290 40468 296 40520
rect 348 40508 354 40520
rect 1397 40511 1455 40517
rect 1397 40508 1409 40511
rect 348 40480 1409 40508
rect 348 40468 354 40480
rect 1397 40477 1409 40480
rect 1443 40477 1455 40511
rect 1397 40471 1455 40477
rect 1946 40468 1952 40520
rect 2004 40468 2010 40520
rect 2038 40468 2044 40520
rect 2096 40508 2102 40520
rect 2501 40511 2559 40517
rect 2501 40508 2513 40511
rect 2096 40480 2513 40508
rect 2096 40468 2102 40480
rect 2501 40477 2513 40480
rect 2547 40477 2559 40511
rect 2501 40471 2559 40477
rect 5626 40468 5632 40520
rect 5684 40468 5690 40520
rect 6825 40511 6883 40517
rect 6825 40477 6837 40511
rect 6871 40508 6883 40511
rect 7285 40511 7343 40517
rect 7285 40508 7297 40511
rect 6871 40480 7297 40508
rect 6871 40477 6883 40480
rect 6825 40471 6883 40477
rect 7285 40477 7297 40480
rect 7331 40508 7343 40511
rect 17405 40511 17463 40517
rect 7331 40480 8248 40508
rect 7331 40477 7343 40480
rect 7285 40471 7343 40477
rect 1670 40400 1676 40452
rect 1728 40400 1734 40452
rect 2222 40400 2228 40452
rect 2280 40400 2286 40452
rect 2777 40443 2835 40449
rect 2777 40409 2789 40443
rect 2823 40440 2835 40443
rect 6546 40440 6552 40452
rect 2823 40412 6552 40440
rect 2823 40409 2835 40412
rect 2777 40403 2835 40409
rect 6546 40400 6552 40412
rect 6604 40400 6610 40452
rect 8220 40384 8248 40480
rect 17405 40477 17417 40511
rect 17451 40477 17463 40511
rect 17405 40471 17463 40477
rect 17420 40440 17448 40471
rect 17678 40468 17684 40520
rect 17736 40468 17742 40520
rect 17954 40468 17960 40520
rect 18012 40468 18018 40520
rect 18230 40468 18236 40520
rect 18288 40468 18294 40520
rect 18322 40468 18328 40520
rect 18380 40508 18386 40520
rect 18509 40511 18567 40517
rect 18509 40508 18521 40511
rect 18380 40480 18521 40508
rect 18380 40468 18386 40480
rect 18509 40477 18521 40480
rect 18555 40477 18567 40511
rect 18509 40471 18567 40477
rect 18782 40468 18788 40520
rect 18840 40468 18846 40520
rect 18892 40517 18920 40548
rect 19306 40548 19564 40576
rect 19904 40576 19932 40616
rect 19981 40613 19993 40647
rect 20027 40644 20039 40647
rect 21174 40644 21180 40656
rect 20027 40616 21180 40644
rect 20027 40613 20039 40616
rect 19981 40607 20039 40613
rect 21174 40604 21180 40616
rect 21232 40604 21238 40656
rect 19904 40548 20484 40576
rect 18877 40511 18935 40517
rect 18877 40477 18889 40511
rect 18923 40477 18935 40511
rect 19306 40508 19334 40548
rect 18877 40471 18935 40477
rect 18984 40480 19334 40508
rect 18984 40440 19012 40480
rect 19610 40468 19616 40520
rect 19668 40468 19674 40520
rect 19889 40511 19947 40517
rect 19889 40477 19901 40511
rect 19935 40504 19947 40511
rect 20070 40504 20076 40520
rect 19935 40477 20076 40504
rect 19889 40476 20076 40477
rect 19889 40471 19947 40476
rect 20070 40468 20076 40476
rect 20128 40468 20134 40520
rect 20456 40517 20484 40548
rect 20165 40511 20223 40517
rect 20165 40477 20177 40511
rect 20211 40477 20223 40511
rect 20165 40471 20223 40477
rect 20441 40511 20499 40517
rect 20441 40477 20453 40511
rect 20487 40477 20499 40511
rect 20441 40471 20499 40477
rect 17420 40412 19012 40440
rect 19150 40400 19156 40452
rect 19208 40440 19214 40452
rect 20180 40440 20208 40471
rect 20714 40468 20720 40520
rect 20772 40468 20778 40520
rect 20806 40468 20812 40520
rect 20864 40508 20870 40520
rect 20993 40511 21051 40517
rect 20993 40508 21005 40511
rect 20864 40480 21005 40508
rect 20864 40468 20870 40480
rect 20993 40477 21005 40480
rect 21039 40477 21051 40511
rect 20993 40471 21051 40477
rect 21266 40468 21272 40520
rect 21324 40468 21330 40520
rect 19208 40412 20208 40440
rect 19208 40400 19214 40412
rect 8202 40332 8208 40384
rect 8260 40332 8266 40384
rect 17218 40332 17224 40384
rect 17276 40332 17282 40384
rect 18049 40375 18107 40381
rect 18049 40341 18061 40375
rect 18095 40372 18107 40375
rect 18506 40372 18512 40384
rect 18095 40344 18512 40372
rect 18095 40341 18107 40344
rect 18049 40335 18107 40341
rect 18506 40332 18512 40344
rect 18564 40332 18570 40384
rect 18598 40332 18604 40384
rect 18656 40332 18662 40384
rect 19426 40332 19432 40384
rect 19484 40332 19490 40384
rect 20254 40332 20260 40384
rect 20312 40332 20318 40384
rect 20530 40332 20536 40384
rect 20588 40332 20594 40384
rect 21453 40375 21511 40381
rect 21453 40341 21465 40375
rect 21499 40372 21511 40375
rect 22186 40372 22192 40384
rect 21499 40344 22192 40372
rect 21499 40341 21511 40344
rect 21453 40335 21511 40341
rect 22186 40332 22192 40344
rect 22244 40332 22250 40384
rect 1104 40282 22056 40304
rect 1104 40230 6148 40282
rect 6200 40230 6212 40282
rect 6264 40230 6276 40282
rect 6328 40230 6340 40282
rect 6392 40230 6404 40282
rect 6456 40230 11346 40282
rect 11398 40230 11410 40282
rect 11462 40230 11474 40282
rect 11526 40230 11538 40282
rect 11590 40230 11602 40282
rect 11654 40230 16544 40282
rect 16596 40230 16608 40282
rect 16660 40230 16672 40282
rect 16724 40230 16736 40282
rect 16788 40230 16800 40282
rect 16852 40230 21742 40282
rect 21794 40230 21806 40282
rect 21858 40230 21870 40282
rect 21922 40230 21934 40282
rect 21986 40230 21998 40282
rect 22050 40230 22056 40282
rect 1104 40208 22056 40230
rect 2130 40128 2136 40180
rect 2188 40168 2194 40180
rect 9214 40168 9220 40180
rect 2188 40140 9220 40168
rect 2188 40128 2194 40140
rect 9214 40128 9220 40140
rect 9272 40128 9278 40180
rect 15654 40128 15660 40180
rect 15712 40168 15718 40180
rect 16117 40171 16175 40177
rect 16117 40168 16129 40171
rect 15712 40140 16129 40168
rect 15712 40128 15718 40140
rect 16117 40137 16129 40140
rect 16163 40137 16175 40171
rect 16117 40131 16175 40137
rect 17497 40171 17555 40177
rect 17497 40137 17509 40171
rect 17543 40168 17555 40171
rect 17586 40168 17592 40180
rect 17543 40140 17592 40168
rect 17543 40137 17555 40140
rect 17497 40131 17555 40137
rect 17586 40128 17592 40140
rect 17644 40128 17650 40180
rect 17678 40128 17684 40180
rect 17736 40128 17742 40180
rect 17770 40128 17776 40180
rect 17828 40128 17834 40180
rect 18046 40128 18052 40180
rect 18104 40128 18110 40180
rect 18325 40171 18383 40177
rect 18325 40137 18337 40171
rect 18371 40168 18383 40171
rect 18414 40168 18420 40180
rect 18371 40140 18420 40168
rect 18371 40137 18383 40140
rect 18325 40131 18383 40137
rect 18414 40128 18420 40140
rect 18472 40128 18478 40180
rect 18601 40171 18659 40177
rect 18601 40137 18613 40171
rect 18647 40168 18659 40171
rect 18782 40168 18788 40180
rect 18647 40140 18788 40168
rect 18647 40137 18659 40140
rect 18601 40131 18659 40137
rect 18782 40128 18788 40140
rect 18840 40128 18846 40180
rect 18874 40128 18880 40180
rect 18932 40128 18938 40180
rect 18966 40128 18972 40180
rect 19024 40128 19030 40180
rect 19150 40128 19156 40180
rect 19208 40128 19214 40180
rect 19429 40171 19487 40177
rect 19429 40137 19441 40171
rect 19475 40137 19487 40171
rect 19429 40131 19487 40137
rect 2041 40103 2099 40109
rect 2041 40069 2053 40103
rect 2087 40100 2099 40103
rect 3142 40100 3148 40112
rect 2087 40072 3148 40100
rect 2087 40069 2099 40072
rect 2041 40063 2099 40069
rect 3142 40060 3148 40072
rect 3200 40060 3206 40112
rect 17696 40100 17724 40128
rect 18138 40100 18144 40112
rect 17696 40072 17908 40100
rect 1762 39992 1768 40044
rect 1820 39992 1826 40044
rect 2317 40035 2375 40041
rect 2317 40001 2329 40035
rect 2363 40032 2375 40035
rect 2682 40032 2688 40044
rect 2363 40004 2688 40032
rect 2363 40001 2375 40004
rect 2317 39995 2375 40001
rect 2682 39992 2688 40004
rect 2740 39992 2746 40044
rect 3053 40035 3111 40041
rect 3053 40001 3065 40035
rect 3099 40001 3111 40035
rect 3053 39995 3111 40001
rect 2590 39924 2596 39976
rect 2648 39924 2654 39976
rect 1118 39856 1124 39908
rect 1176 39896 1182 39908
rect 3068 39896 3096 39995
rect 16298 39992 16304 40044
rect 16356 39992 16362 40044
rect 17678 39992 17684 40044
rect 17736 39992 17742 40044
rect 3329 39967 3387 39973
rect 3329 39933 3341 39967
rect 3375 39964 3387 39967
rect 3418 39964 3424 39976
rect 3375 39936 3424 39964
rect 3375 39933 3387 39936
rect 3329 39927 3387 39933
rect 3418 39924 3424 39936
rect 3476 39924 3482 39976
rect 1176 39868 3096 39896
rect 1176 39856 1182 39868
rect 4706 39856 4712 39908
rect 4764 39896 4770 39908
rect 5534 39896 5540 39908
rect 4764 39868 5540 39896
rect 4764 39856 4770 39868
rect 5534 39856 5540 39868
rect 5592 39896 5598 39908
rect 5592 39868 12434 39896
rect 5592 39856 5598 39868
rect 4062 39788 4068 39840
rect 4120 39828 4126 39840
rect 6822 39828 6828 39840
rect 4120 39800 6828 39828
rect 4120 39788 4126 39800
rect 6822 39788 6828 39800
rect 6880 39788 6886 39840
rect 12406 39828 12434 39868
rect 13538 39856 13544 39908
rect 13596 39896 13602 39908
rect 15930 39896 15936 39908
rect 13596 39868 15936 39896
rect 13596 39856 13602 39868
rect 15930 39856 15936 39868
rect 15988 39856 15994 39908
rect 17880 39896 17908 40072
rect 17972 40072 18144 40100
rect 17972 40041 18000 40072
rect 18138 40060 18144 40072
rect 18196 40060 18202 40112
rect 18892 40100 18920 40128
rect 18248 40072 18920 40100
rect 18984 40100 19012 40128
rect 19444 40100 19472 40131
rect 20254 40128 20260 40180
rect 20312 40128 20318 40180
rect 20346 40128 20352 40180
rect 20404 40168 20410 40180
rect 20533 40171 20591 40177
rect 20533 40168 20545 40171
rect 20404 40140 20545 40168
rect 20404 40128 20410 40140
rect 20533 40137 20545 40140
rect 20579 40137 20591 40171
rect 20533 40131 20591 40137
rect 20809 40171 20867 40177
rect 20809 40137 20821 40171
rect 20855 40168 20867 40171
rect 20855 40140 21220 40168
rect 20855 40137 20867 40140
rect 20809 40131 20867 40137
rect 20272 40100 20300 40128
rect 20898 40100 20904 40112
rect 18984 40072 19472 40100
rect 19904 40072 20116 40100
rect 20272 40072 20484 40100
rect 18248 40041 18276 40072
rect 17957 40035 18015 40041
rect 17957 40001 17969 40035
rect 18003 40001 18015 40035
rect 17957 39995 18015 40001
rect 18233 40035 18291 40041
rect 18233 40001 18245 40035
rect 18279 40001 18291 40035
rect 18233 39995 18291 40001
rect 18509 40035 18567 40041
rect 18509 40001 18521 40035
rect 18555 40032 18567 40035
rect 18690 40032 18696 40044
rect 18555 40004 18696 40032
rect 18555 40001 18567 40004
rect 18509 39995 18567 40001
rect 18690 39992 18696 40004
rect 18748 39992 18754 40044
rect 18782 39992 18788 40044
rect 18840 39992 18846 40044
rect 18966 39992 18972 40044
rect 19024 40032 19030 40044
rect 19061 40035 19119 40041
rect 19061 40032 19073 40035
rect 19024 40004 19073 40032
rect 19024 39992 19030 40004
rect 19061 40001 19073 40004
rect 19107 40001 19119 40035
rect 19061 39995 19119 40001
rect 19337 40035 19395 40041
rect 19337 40001 19349 40035
rect 19383 40001 19395 40035
rect 19337 39995 19395 40001
rect 19613 40035 19671 40041
rect 19613 40001 19625 40035
rect 19659 40032 19671 40035
rect 19702 40032 19708 40044
rect 19659 40004 19708 40032
rect 19659 40001 19671 40004
rect 19613 39995 19671 40001
rect 18046 39924 18052 39976
rect 18104 39964 18110 39976
rect 19352 39964 19380 39995
rect 19702 39992 19708 40004
rect 19760 39992 19766 40044
rect 18104 39936 19380 39964
rect 18104 39924 18110 39936
rect 19426 39924 19432 39976
rect 19484 39964 19490 39976
rect 19904 39964 19932 40072
rect 19981 40035 20039 40041
rect 19981 40001 19993 40035
rect 20027 40001 20039 40035
rect 19981 39995 20039 40001
rect 19484 39936 19932 39964
rect 19484 39924 19490 39936
rect 18877 39899 18935 39905
rect 17880 39868 18460 39896
rect 16206 39828 16212 39840
rect 12406 39800 16212 39828
rect 16206 39788 16212 39800
rect 16264 39788 16270 39840
rect 18432 39828 18460 39868
rect 18877 39865 18889 39899
rect 18923 39896 18935 39899
rect 19886 39896 19892 39908
rect 18923 39868 19892 39896
rect 18923 39865 18935 39868
rect 18877 39859 18935 39865
rect 19886 39856 19892 39868
rect 19944 39856 19950 39908
rect 19797 39831 19855 39837
rect 19797 39828 19809 39831
rect 18432 39800 19809 39828
rect 19797 39797 19809 39800
rect 19843 39797 19855 39831
rect 19996 39828 20024 39995
rect 20088 39964 20116 40072
rect 20456 40041 20484 40072
rect 20732 40072 20904 40100
rect 20732 40041 20760 40072
rect 20898 40060 20904 40072
rect 20956 40060 20962 40112
rect 21192 40109 21220 40140
rect 21177 40103 21235 40109
rect 21177 40069 21189 40103
rect 21223 40069 21235 40103
rect 21177 40063 21235 40069
rect 20441 40035 20499 40041
rect 20441 40001 20453 40035
rect 20487 40001 20499 40035
rect 20441 39995 20499 40001
rect 20717 40035 20775 40041
rect 20717 40001 20729 40035
rect 20763 40001 20775 40035
rect 20717 39995 20775 40001
rect 20993 40035 21051 40041
rect 20993 40001 21005 40035
rect 21039 40032 21051 40035
rect 21082 40032 21088 40044
rect 21039 40004 21088 40032
rect 21039 40001 21051 40004
rect 20993 39995 21051 40001
rect 21082 39992 21088 40004
rect 21140 39992 21146 40044
rect 21358 39964 21364 39976
rect 20088 39936 21364 39964
rect 21358 39924 21364 39936
rect 21416 39924 21422 39976
rect 20257 39899 20315 39905
rect 20257 39865 20269 39899
rect 20303 39896 20315 39899
rect 20990 39896 20996 39908
rect 20303 39868 20996 39896
rect 20303 39865 20315 39868
rect 20257 39859 20315 39865
rect 20990 39856 20996 39868
rect 21048 39856 21054 39908
rect 22462 39896 22468 39908
rect 21376 39868 22468 39896
rect 21376 39828 21404 39868
rect 22462 39856 22468 39868
rect 22520 39856 22526 39908
rect 19996 39800 21404 39828
rect 19797 39791 19855 39797
rect 21450 39788 21456 39840
rect 21508 39788 21514 39840
rect 1104 39738 21896 39760
rect 1104 39686 3549 39738
rect 3601 39686 3613 39738
rect 3665 39686 3677 39738
rect 3729 39686 3741 39738
rect 3793 39686 3805 39738
rect 3857 39686 8747 39738
rect 8799 39686 8811 39738
rect 8863 39686 8875 39738
rect 8927 39686 8939 39738
rect 8991 39686 9003 39738
rect 9055 39686 13945 39738
rect 13997 39686 14009 39738
rect 14061 39686 14073 39738
rect 14125 39686 14137 39738
rect 14189 39686 14201 39738
rect 14253 39686 19143 39738
rect 19195 39686 19207 39738
rect 19259 39686 19271 39738
rect 19323 39686 19335 39738
rect 19387 39686 19399 39738
rect 19451 39686 21896 39738
rect 1104 39664 21896 39686
rect 5810 39584 5816 39636
rect 5868 39624 5874 39636
rect 6181 39627 6239 39633
rect 6181 39624 6193 39627
rect 5868 39596 6193 39624
rect 5868 39584 5874 39596
rect 6181 39593 6193 39596
rect 6227 39593 6239 39627
rect 10134 39624 10140 39636
rect 6181 39587 6239 39593
rect 8128 39596 10140 39624
rect 8128 39568 8156 39596
rect 10134 39584 10140 39596
rect 10192 39584 10198 39636
rect 15933 39627 15991 39633
rect 15933 39593 15945 39627
rect 15979 39624 15991 39627
rect 16298 39624 16304 39636
rect 15979 39596 16304 39624
rect 15979 39593 15991 39596
rect 15933 39587 15991 39593
rect 16298 39584 16304 39596
rect 16356 39584 16362 39636
rect 17405 39627 17463 39633
rect 17405 39593 17417 39627
rect 17451 39624 17463 39627
rect 17678 39624 17684 39636
rect 17451 39596 17684 39624
rect 17451 39593 17463 39596
rect 17405 39587 17463 39593
rect 17678 39584 17684 39596
rect 17736 39584 17742 39636
rect 18046 39584 18052 39636
rect 18104 39584 18110 39636
rect 18877 39627 18935 39633
rect 18877 39593 18889 39627
rect 18923 39624 18935 39627
rect 19610 39624 19616 39636
rect 18923 39596 19616 39624
rect 18923 39593 18935 39596
rect 18877 39587 18935 39593
rect 19610 39584 19616 39596
rect 19668 39584 19674 39636
rect 19797 39627 19855 39633
rect 19797 39593 19809 39627
rect 19843 39624 19855 39627
rect 20714 39624 20720 39636
rect 19843 39596 20720 39624
rect 19843 39593 19855 39596
rect 19797 39587 19855 39593
rect 20714 39584 20720 39596
rect 20772 39584 20778 39636
rect 21266 39584 21272 39636
rect 21324 39584 21330 39636
rect 8110 39516 8116 39568
rect 8168 39516 8174 39568
rect 18966 39556 18972 39568
rect 12406 39528 18972 39556
rect 3050 39488 3056 39500
rect 2884 39460 3056 39488
rect 1489 39423 1547 39429
rect 1489 39389 1501 39423
rect 1535 39420 1547 39423
rect 1670 39420 1676 39432
rect 1535 39392 1676 39420
rect 1535 39389 1547 39392
rect 1489 39383 1547 39389
rect 1670 39380 1676 39392
rect 1728 39380 1734 39432
rect 1763 39423 1821 39429
rect 1763 39389 1775 39423
rect 1809 39420 1821 39423
rect 1854 39420 1860 39432
rect 1809 39392 1860 39420
rect 1809 39389 1821 39392
rect 1763 39383 1821 39389
rect 1854 39380 1860 39392
rect 1912 39380 1918 39432
rect 2884 39429 2912 39460
rect 3050 39448 3056 39460
rect 3108 39448 3114 39500
rect 3694 39448 3700 39500
rect 3752 39488 3758 39500
rect 4065 39491 4123 39497
rect 4065 39488 4077 39491
rect 3752 39460 4077 39488
rect 3752 39448 3758 39460
rect 4065 39457 4077 39460
rect 4111 39488 4123 39491
rect 12406 39488 12434 39528
rect 18966 39516 18972 39528
rect 19024 39516 19030 39568
rect 19334 39516 19340 39568
rect 19392 39556 19398 39568
rect 19521 39559 19579 39565
rect 19521 39556 19533 39559
rect 19392 39528 19533 39556
rect 19392 39516 19398 39528
rect 19521 39525 19533 39528
rect 19567 39525 19579 39559
rect 19521 39519 19579 39525
rect 20073 39559 20131 39565
rect 20073 39525 20085 39559
rect 20119 39556 20131 39559
rect 21284 39556 21312 39584
rect 20119 39528 21312 39556
rect 20119 39525 20131 39528
rect 20073 39519 20131 39525
rect 19610 39488 19616 39500
rect 4111 39460 12434 39488
rect 18616 39460 19616 39488
rect 4111 39457 4123 39460
rect 4065 39451 4123 39457
rect 2869 39423 2927 39429
rect 2869 39389 2881 39423
rect 2915 39389 2927 39423
rect 3789 39423 3847 39429
rect 3789 39420 3801 39423
rect 2869 39383 2927 39389
rect 3068 39392 3801 39420
rect 1302 39312 1308 39364
rect 1360 39352 1366 39364
rect 3068 39352 3096 39392
rect 3789 39389 3801 39392
rect 3835 39389 3847 39423
rect 3789 39383 3847 39389
rect 5718 39380 5724 39432
rect 5776 39420 5782 39432
rect 6365 39423 6423 39429
rect 6365 39420 6377 39423
rect 5776 39392 6377 39420
rect 5776 39380 5782 39392
rect 6365 39389 6377 39392
rect 6411 39389 6423 39423
rect 6365 39383 6423 39389
rect 16114 39380 16120 39432
rect 16172 39380 16178 39432
rect 17494 39380 17500 39432
rect 17552 39420 17558 39432
rect 17589 39423 17647 39429
rect 17589 39420 17601 39423
rect 17552 39392 17601 39420
rect 17552 39380 17558 39392
rect 17589 39389 17601 39392
rect 17635 39389 17647 39423
rect 17589 39383 17647 39389
rect 17678 39380 17684 39432
rect 17736 39420 17742 39432
rect 17865 39423 17923 39429
rect 17865 39420 17877 39423
rect 17736 39392 17877 39420
rect 17736 39380 17742 39392
rect 17865 39389 17877 39392
rect 17911 39389 17923 39423
rect 17865 39383 17923 39389
rect 18233 39423 18291 39429
rect 18233 39389 18245 39423
rect 18279 39389 18291 39423
rect 18233 39383 18291 39389
rect 1360 39324 3096 39352
rect 3145 39355 3203 39361
rect 1360 39312 1366 39324
rect 3145 39321 3157 39355
rect 3191 39352 3203 39355
rect 3970 39352 3976 39364
rect 3191 39324 3976 39352
rect 3191 39321 3203 39324
rect 3145 39315 3203 39321
rect 3970 39312 3976 39324
rect 4028 39312 4034 39364
rect 18248 39352 18276 39383
rect 17052 39324 18276 39352
rect 17052 39296 17080 39324
rect 2498 39244 2504 39296
rect 2556 39244 2562 39296
rect 4154 39244 4160 39296
rect 4212 39284 4218 39296
rect 8386 39284 8392 39296
rect 4212 39256 8392 39284
rect 4212 39244 4218 39256
rect 8386 39244 8392 39256
rect 8444 39244 8450 39296
rect 17034 39244 17040 39296
rect 17092 39244 17098 39296
rect 17681 39287 17739 39293
rect 17681 39253 17693 39287
rect 17727 39284 17739 39287
rect 18616 39284 18644 39460
rect 19610 39448 19616 39460
rect 19668 39448 19674 39500
rect 18874 39380 18880 39432
rect 18932 39420 18938 39432
rect 19061 39423 19119 39429
rect 19061 39420 19073 39423
rect 18932 39392 19073 39420
rect 18932 39380 18938 39392
rect 19061 39389 19073 39392
rect 19107 39389 19119 39423
rect 19061 39383 19119 39389
rect 19429 39423 19487 39429
rect 19429 39389 19441 39423
rect 19475 39420 19487 39423
rect 19518 39420 19524 39432
rect 19475 39392 19524 39420
rect 19475 39389 19487 39392
rect 19429 39383 19487 39389
rect 19518 39380 19524 39392
rect 19576 39380 19582 39432
rect 19702 39380 19708 39432
rect 19760 39380 19766 39432
rect 19794 39380 19800 39432
rect 19852 39420 19858 39432
rect 19981 39423 20039 39429
rect 19981 39420 19993 39423
rect 19852 39392 19993 39420
rect 19852 39380 19858 39392
rect 19981 39389 19993 39392
rect 20027 39389 20039 39423
rect 20257 39423 20315 39429
rect 20257 39420 20269 39423
rect 19981 39383 20039 39389
rect 20088 39392 20269 39420
rect 18782 39312 18788 39364
rect 18840 39352 18846 39364
rect 20088 39352 20116 39392
rect 20257 39389 20269 39392
rect 20303 39389 20315 39423
rect 20257 39383 20315 39389
rect 20346 39380 20352 39432
rect 20404 39420 20410 39432
rect 20533 39423 20591 39429
rect 20533 39420 20545 39423
rect 20404 39392 20545 39420
rect 20404 39380 20410 39392
rect 20533 39389 20545 39392
rect 20579 39389 20591 39423
rect 20806 39420 20812 39432
rect 20533 39383 20591 39389
rect 20640 39392 20812 39420
rect 20438 39352 20444 39364
rect 18840 39324 20116 39352
rect 20180 39324 20444 39352
rect 18840 39312 18846 39324
rect 17727 39256 18644 39284
rect 19245 39287 19303 39293
rect 17727 39253 17739 39256
rect 17681 39247 17739 39253
rect 19245 39253 19257 39287
rect 19291 39284 19303 39287
rect 20180 39284 20208 39324
rect 20438 39312 20444 39324
rect 20496 39312 20502 39364
rect 19291 39256 20208 39284
rect 20349 39287 20407 39293
rect 19291 39253 19303 39256
rect 19245 39247 19303 39253
rect 20349 39253 20361 39287
rect 20395 39284 20407 39287
rect 20640 39284 20668 39392
rect 20806 39380 20812 39392
rect 20864 39380 20870 39432
rect 20990 39380 20996 39432
rect 21048 39380 21054 39432
rect 21269 39423 21327 39429
rect 21269 39389 21281 39423
rect 21315 39389 21327 39423
rect 21269 39383 21327 39389
rect 20714 39312 20720 39364
rect 20772 39352 20778 39364
rect 21284 39352 21312 39383
rect 20772 39324 21312 39352
rect 20772 39312 20778 39324
rect 20395 39256 20668 39284
rect 20395 39253 20407 39256
rect 20349 39247 20407 39253
rect 20806 39244 20812 39296
rect 20864 39244 20870 39296
rect 21453 39287 21511 39293
rect 21453 39253 21465 39287
rect 21499 39284 21511 39287
rect 22186 39284 22192 39296
rect 21499 39256 22192 39284
rect 21499 39253 21511 39256
rect 21453 39247 21511 39253
rect 22186 39244 22192 39256
rect 22244 39244 22250 39296
rect 1104 39194 22056 39216
rect 1104 39142 6148 39194
rect 6200 39142 6212 39194
rect 6264 39142 6276 39194
rect 6328 39142 6340 39194
rect 6392 39142 6404 39194
rect 6456 39142 11346 39194
rect 11398 39142 11410 39194
rect 11462 39142 11474 39194
rect 11526 39142 11538 39194
rect 11590 39142 11602 39194
rect 11654 39142 16544 39194
rect 16596 39142 16608 39194
rect 16660 39142 16672 39194
rect 16724 39142 16736 39194
rect 16788 39142 16800 39194
rect 16852 39142 21742 39194
rect 21794 39142 21806 39194
rect 21858 39142 21870 39194
rect 21922 39142 21934 39194
rect 21986 39142 21998 39194
rect 22050 39142 22056 39194
rect 1104 39120 22056 39142
rect 1578 39040 1584 39092
rect 1636 39040 1642 39092
rect 5074 39080 5080 39092
rect 1688 39052 5080 39080
rect 1397 38947 1455 38953
rect 1397 38913 1409 38947
rect 1443 38913 1455 38947
rect 1397 38907 1455 38913
rect 1412 38740 1440 38907
rect 1596 38808 1624 39040
rect 1688 39021 1716 39052
rect 5074 39040 5080 39052
rect 5132 39040 5138 39092
rect 5994 39040 6000 39092
rect 6052 39040 6058 39092
rect 15657 39083 15715 39089
rect 15657 39049 15669 39083
rect 15703 39080 15715 39083
rect 16114 39080 16120 39092
rect 15703 39052 16120 39080
rect 15703 39049 15715 39052
rect 15657 39043 15715 39049
rect 16114 39040 16120 39052
rect 16172 39040 16178 39092
rect 18782 39040 18788 39092
rect 18840 39040 18846 39092
rect 19705 39083 19763 39089
rect 19705 39049 19717 39083
rect 19751 39049 19763 39083
rect 19705 39043 19763 39049
rect 20073 39083 20131 39089
rect 20073 39049 20085 39083
rect 20119 39080 20131 39083
rect 20162 39080 20168 39092
rect 20119 39052 20168 39080
rect 20119 39049 20131 39052
rect 20073 39043 20131 39049
rect 1673 39015 1731 39021
rect 1673 38981 1685 39015
rect 1719 38981 1731 39015
rect 1673 38975 1731 38981
rect 1854 38972 1860 39024
rect 1912 39012 1918 39024
rect 2958 39012 2964 39024
rect 1912 38984 2964 39012
rect 1912 38972 1918 38984
rect 2958 38972 2964 38984
rect 3016 38972 3022 39024
rect 3142 38972 3148 39024
rect 3200 39012 3206 39024
rect 3326 39012 3332 39024
rect 3200 38984 3332 39012
rect 3200 38972 3206 38984
rect 3326 38972 3332 38984
rect 3384 39012 3390 39024
rect 3384 38984 3832 39012
rect 3384 38972 3390 38984
rect 2223 38947 2281 38953
rect 2223 38913 2235 38947
rect 2269 38944 2281 38947
rect 2590 38944 2596 38956
rect 2269 38916 2596 38944
rect 2269 38913 2281 38916
rect 2223 38907 2281 38913
rect 2590 38904 2596 38916
rect 2648 38944 2654 38956
rect 3694 38944 3700 38956
rect 2648 38916 3700 38944
rect 2648 38904 2654 38916
rect 3694 38904 3700 38916
rect 3752 38904 3758 38956
rect 3804 38944 3832 38984
rect 8294 38972 8300 39024
rect 8352 39012 8358 39024
rect 19720 39012 19748 39043
rect 20162 39040 20168 39052
rect 20220 39040 20226 39092
rect 20346 39040 20352 39092
rect 20404 39040 20410 39092
rect 20533 39083 20591 39089
rect 20533 39049 20545 39083
rect 20579 39080 20591 39083
rect 20714 39080 20720 39092
rect 20579 39052 20720 39080
rect 20579 39049 20591 39052
rect 20533 39043 20591 39049
rect 20714 39040 20720 39052
rect 20772 39040 20778 39092
rect 20806 39040 20812 39092
rect 20864 39080 20870 39092
rect 20864 39052 21220 39080
rect 20864 39040 20870 39052
rect 20364 39012 20392 39040
rect 21192 39021 21220 39052
rect 8352 38984 19104 39012
rect 19720 38984 20392 39012
rect 21177 39015 21235 39021
rect 8352 38972 8358 38984
rect 4047 38947 4105 38953
rect 4047 38944 4059 38947
rect 3804 38916 4059 38944
rect 4047 38913 4059 38916
rect 4093 38913 4105 38947
rect 4047 38907 4105 38913
rect 5994 38904 6000 38956
rect 6052 38944 6058 38956
rect 6181 38947 6239 38953
rect 6181 38944 6193 38947
rect 6052 38916 6193 38944
rect 6052 38904 6058 38916
rect 6181 38913 6193 38916
rect 6227 38913 6239 38947
rect 6181 38907 6239 38913
rect 6365 38947 6423 38953
rect 6365 38913 6377 38947
rect 6411 38913 6423 38947
rect 6365 38907 6423 38913
rect 1670 38836 1676 38888
rect 1728 38876 1734 38888
rect 1949 38879 2007 38885
rect 1949 38876 1961 38879
rect 1728 38848 1961 38876
rect 1728 38836 1734 38848
rect 1949 38845 1961 38848
rect 1995 38845 2007 38879
rect 1949 38839 2007 38845
rect 1596 38780 1716 38808
rect 1688 38752 1716 38780
rect 1486 38740 1492 38752
rect 1412 38712 1492 38740
rect 1486 38700 1492 38712
rect 1544 38700 1550 38752
rect 1670 38700 1676 38752
rect 1728 38700 1734 38752
rect 1964 38740 1992 38839
rect 2958 38836 2964 38888
rect 3016 38876 3022 38888
rect 3418 38876 3424 38888
rect 3016 38848 3424 38876
rect 3016 38836 3022 38848
rect 3418 38836 3424 38848
rect 3476 38836 3482 38888
rect 3789 38879 3847 38885
rect 3789 38845 3801 38879
rect 3835 38845 3847 38879
rect 3789 38839 3847 38845
rect 3804 38808 3832 38839
rect 3804 38780 3924 38808
rect 3896 38752 3924 38780
rect 5258 38768 5264 38820
rect 5316 38808 5322 38820
rect 6380 38808 6408 38907
rect 6546 38904 6552 38956
rect 6604 38944 6610 38956
rect 6639 38947 6697 38953
rect 6639 38944 6651 38947
rect 6604 38916 6651 38944
rect 6604 38904 6610 38916
rect 6639 38913 6651 38916
rect 6685 38944 6697 38947
rect 6730 38944 6736 38956
rect 6685 38916 6736 38944
rect 6685 38913 6697 38916
rect 6639 38907 6697 38913
rect 6730 38904 6736 38916
rect 6788 38944 6794 38956
rect 6788 38916 12434 38944
rect 6788 38904 6794 38916
rect 12406 38876 12434 38916
rect 15838 38904 15844 38956
rect 15896 38904 15902 38956
rect 17034 38944 17040 38956
rect 16132 38916 17040 38944
rect 16132 38876 16160 38916
rect 17034 38904 17040 38916
rect 17092 38904 17098 38956
rect 18966 38904 18972 38956
rect 19024 38904 19030 38956
rect 19076 38944 19104 38984
rect 21177 38981 21189 39015
rect 21223 38981 21235 39015
rect 21177 38975 21235 38981
rect 19794 38944 19800 38956
rect 19076 38916 19800 38944
rect 19794 38904 19800 38916
rect 19852 38904 19858 38956
rect 19889 38947 19947 38953
rect 19889 38913 19901 38947
rect 19935 38913 19947 38947
rect 19889 38907 19947 38913
rect 12406 38848 16160 38876
rect 16206 38836 16212 38888
rect 16264 38876 16270 38888
rect 19904 38876 19932 38907
rect 20254 38904 20260 38956
rect 20312 38904 20318 38956
rect 20714 38904 20720 38956
rect 20772 38904 20778 38956
rect 20898 38904 20904 38956
rect 20956 38944 20962 38956
rect 20993 38947 21051 38953
rect 20993 38944 21005 38947
rect 20956 38916 21005 38944
rect 20956 38904 20962 38916
rect 20993 38913 21005 38916
rect 21039 38913 21051 38947
rect 20993 38907 21051 38913
rect 16264 38848 19932 38876
rect 16264 38836 16270 38848
rect 5316 38780 6408 38808
rect 5316 38768 5322 38780
rect 2314 38740 2320 38752
rect 1964 38712 2320 38740
rect 2314 38700 2320 38712
rect 2372 38700 2378 38752
rect 2961 38743 3019 38749
rect 2961 38709 2973 38743
rect 3007 38740 3019 38743
rect 3142 38740 3148 38752
rect 3007 38712 3148 38740
rect 3007 38709 3019 38712
rect 2961 38703 3019 38709
rect 3142 38700 3148 38712
rect 3200 38700 3206 38752
rect 3878 38700 3884 38752
rect 3936 38700 3942 38752
rect 4522 38700 4528 38752
rect 4580 38740 4586 38752
rect 4801 38743 4859 38749
rect 4801 38740 4813 38743
rect 4580 38712 4813 38740
rect 4580 38700 4586 38712
rect 4801 38709 4813 38712
rect 4847 38709 4859 38743
rect 4801 38703 4859 38709
rect 5166 38700 5172 38752
rect 5224 38740 5230 38752
rect 5902 38740 5908 38752
rect 5224 38712 5908 38740
rect 5224 38700 5230 38712
rect 5902 38700 5908 38712
rect 5960 38700 5966 38752
rect 6380 38740 6408 38780
rect 11882 38768 11888 38820
rect 11940 38808 11946 38820
rect 12250 38808 12256 38820
rect 11940 38780 12256 38808
rect 11940 38768 11946 38780
rect 12250 38768 12256 38780
rect 12308 38768 12314 38820
rect 6638 38740 6644 38752
rect 6380 38712 6644 38740
rect 6638 38700 6644 38712
rect 6696 38700 6702 38752
rect 7374 38700 7380 38752
rect 7432 38700 7438 38752
rect 7558 38700 7564 38752
rect 7616 38740 7622 38752
rect 12618 38740 12624 38752
rect 7616 38712 12624 38740
rect 7616 38700 7622 38712
rect 12618 38700 12624 38712
rect 12676 38700 12682 38752
rect 15746 38700 15752 38752
rect 15804 38740 15810 38752
rect 16206 38740 16212 38752
rect 15804 38712 16212 38740
rect 15804 38700 15810 38712
rect 16206 38700 16212 38712
rect 16264 38700 16270 38752
rect 20809 38743 20867 38749
rect 20809 38709 20821 38743
rect 20855 38740 20867 38743
rect 21174 38740 21180 38752
rect 20855 38712 21180 38740
rect 20855 38709 20867 38712
rect 20809 38703 20867 38709
rect 21174 38700 21180 38712
rect 21232 38700 21238 38752
rect 21450 38700 21456 38752
rect 21508 38700 21514 38752
rect 1104 38650 21896 38672
rect 1104 38598 3549 38650
rect 3601 38598 3613 38650
rect 3665 38598 3677 38650
rect 3729 38598 3741 38650
rect 3793 38598 3805 38650
rect 3857 38598 8747 38650
rect 8799 38598 8811 38650
rect 8863 38598 8875 38650
rect 8927 38598 8939 38650
rect 8991 38598 9003 38650
rect 9055 38598 13945 38650
rect 13997 38598 14009 38650
rect 14061 38598 14073 38650
rect 14125 38598 14137 38650
rect 14189 38598 14201 38650
rect 14253 38598 19143 38650
rect 19195 38598 19207 38650
rect 19259 38598 19271 38650
rect 19323 38598 19335 38650
rect 19387 38598 19399 38650
rect 19451 38598 21896 38650
rect 1104 38576 21896 38598
rect 1688 38508 2774 38536
rect 1118 38360 1124 38412
rect 1176 38400 1182 38412
rect 1688 38409 1716 38508
rect 1673 38403 1731 38409
rect 1673 38400 1685 38403
rect 1176 38372 1685 38400
rect 1176 38360 1182 38372
rect 1673 38369 1685 38372
rect 1719 38369 1731 38403
rect 2746 38400 2774 38508
rect 6822 38496 6828 38548
rect 6880 38536 6886 38548
rect 9674 38536 9680 38548
rect 6880 38508 9680 38536
rect 6880 38496 6886 38508
rect 9674 38496 9680 38508
rect 9732 38536 9738 38548
rect 13170 38536 13176 38548
rect 9732 38508 13176 38536
rect 9732 38496 9738 38508
rect 13170 38496 13176 38508
rect 13228 38496 13234 38548
rect 16022 38496 16028 38548
rect 16080 38536 16086 38548
rect 16117 38539 16175 38545
rect 16117 38536 16129 38539
rect 16080 38508 16129 38536
rect 16080 38496 16086 38508
rect 16117 38505 16129 38508
rect 16163 38505 16175 38539
rect 16117 38499 16175 38505
rect 17313 38539 17371 38545
rect 17313 38505 17325 38539
rect 17359 38536 17371 38539
rect 17678 38536 17684 38548
rect 17359 38508 17684 38536
rect 17359 38505 17371 38508
rect 17313 38499 17371 38505
rect 17678 38496 17684 38508
rect 17736 38496 17742 38548
rect 17865 38539 17923 38545
rect 17865 38505 17877 38539
rect 17911 38536 17923 38539
rect 18966 38536 18972 38548
rect 17911 38508 18972 38536
rect 17911 38505 17923 38508
rect 17865 38499 17923 38505
rect 18966 38496 18972 38508
rect 19024 38496 19030 38548
rect 19705 38539 19763 38545
rect 19705 38505 19717 38539
rect 19751 38536 19763 38539
rect 20714 38536 20720 38548
rect 19751 38508 20720 38536
rect 19751 38505 19763 38508
rect 19705 38499 19763 38505
rect 20714 38496 20720 38508
rect 20772 38496 20778 38548
rect 20990 38496 20996 38548
rect 21048 38496 21054 38548
rect 19978 38428 19984 38480
rect 20036 38428 20042 38480
rect 20257 38471 20315 38477
rect 20257 38437 20269 38471
rect 20303 38468 20315 38471
rect 21008 38468 21036 38496
rect 20303 38440 21036 38468
rect 20303 38437 20315 38440
rect 20257 38431 20315 38437
rect 3878 38400 3884 38412
rect 2746 38372 3884 38400
rect 1673 38363 1731 38369
rect 3878 38360 3884 38372
rect 3936 38360 3942 38412
rect 5258 38360 5264 38412
rect 5316 38400 5322 38412
rect 5353 38403 5411 38409
rect 5353 38400 5365 38403
rect 5316 38372 5365 38400
rect 5316 38360 5322 38372
rect 5353 38369 5365 38372
rect 5399 38369 5411 38403
rect 5353 38363 5411 38369
rect 7558 38360 7564 38412
rect 7616 38400 7622 38412
rect 12710 38400 12716 38412
rect 7616 38372 12716 38400
rect 7616 38360 7622 38372
rect 12710 38360 12716 38372
rect 12768 38360 12774 38412
rect 14550 38360 14556 38412
rect 14608 38400 14614 38412
rect 16022 38400 16028 38412
rect 14608 38372 16028 38400
rect 14608 38360 14614 38372
rect 16022 38360 16028 38372
rect 16080 38400 16086 38412
rect 16080 38372 17540 38400
rect 16080 38360 16086 38372
rect 1854 38292 1860 38344
rect 1912 38332 1918 38344
rect 1947 38335 2005 38341
rect 1947 38332 1959 38335
rect 1912 38304 1959 38332
rect 1912 38292 1918 38304
rect 1947 38301 1959 38304
rect 1993 38301 2005 38335
rect 3145 38335 3203 38341
rect 3145 38332 3157 38335
rect 1947 38295 2005 38301
rect 2746 38304 3157 38332
rect 1302 38224 1308 38276
rect 1360 38264 1366 38276
rect 2746 38264 2774 38304
rect 3145 38301 3157 38304
rect 3191 38301 3203 38335
rect 3145 38295 3203 38301
rect 4062 38292 4068 38344
rect 4120 38332 4126 38344
rect 4155 38335 4213 38341
rect 4155 38332 4167 38335
rect 4120 38304 4167 38332
rect 4120 38292 4126 38304
rect 4155 38301 4167 38304
rect 4201 38332 4213 38335
rect 4890 38332 4896 38344
rect 4201 38304 4896 38332
rect 4201 38301 4213 38304
rect 4155 38295 4213 38301
rect 4890 38292 4896 38304
rect 4948 38292 4954 38344
rect 5534 38332 5540 38344
rect 5460 38304 5540 38332
rect 1360 38236 2774 38264
rect 1360 38224 1366 38236
rect 3418 38224 3424 38276
rect 3476 38224 3482 38276
rect 5460 38264 5488 38304
rect 5534 38292 5540 38304
rect 5592 38341 5598 38344
rect 5592 38335 5653 38341
rect 5592 38301 5607 38335
rect 5641 38301 5653 38335
rect 5592 38295 5653 38301
rect 5592 38292 5598 38295
rect 6638 38292 6644 38344
rect 6696 38332 6702 38344
rect 6733 38335 6791 38341
rect 6733 38332 6745 38335
rect 6696 38304 6745 38332
rect 6696 38292 6702 38304
rect 6733 38301 6745 38304
rect 6779 38301 6791 38335
rect 6733 38295 6791 38301
rect 5276 38236 5488 38264
rect 6748 38264 6776 38295
rect 6914 38292 6920 38344
rect 6972 38332 6978 38344
rect 7007 38335 7065 38341
rect 7007 38332 7019 38335
rect 6972 38304 7019 38332
rect 6972 38292 6978 38304
rect 7007 38301 7019 38304
rect 7053 38332 7065 38335
rect 9122 38332 9128 38344
rect 7053 38304 9128 38332
rect 7053 38301 7065 38304
rect 7007 38295 7065 38301
rect 9122 38292 9128 38304
rect 9180 38292 9186 38344
rect 13538 38292 13544 38344
rect 13596 38332 13602 38344
rect 17512 38341 17540 38372
rect 16301 38335 16359 38341
rect 16301 38332 16313 38335
rect 13596 38304 16313 38332
rect 13596 38292 13602 38304
rect 16301 38301 16313 38304
rect 16347 38301 16359 38335
rect 16301 38295 16359 38301
rect 17497 38335 17555 38341
rect 17497 38301 17509 38335
rect 17543 38301 17555 38335
rect 17497 38295 17555 38301
rect 18049 38335 18107 38341
rect 18049 38301 18061 38335
rect 18095 38301 18107 38335
rect 18049 38295 18107 38301
rect 6748 38236 7236 38264
rect 5276 38208 5304 38236
rect 7208 38208 7236 38236
rect 7834 38224 7840 38276
rect 7892 38264 7898 38276
rect 11698 38264 11704 38276
rect 7892 38236 11704 38264
rect 7892 38224 7898 38236
rect 11698 38224 11704 38236
rect 11756 38224 11762 38276
rect 18064 38264 18092 38295
rect 18598 38292 18604 38344
rect 18656 38332 18662 38344
rect 19889 38335 19947 38341
rect 19889 38332 19901 38335
rect 18656 38304 19901 38332
rect 18656 38292 18662 38304
rect 19889 38301 19901 38304
rect 19935 38301 19947 38335
rect 19889 38295 19947 38301
rect 20162 38292 20168 38344
rect 20220 38292 20226 38344
rect 20438 38292 20444 38344
rect 20496 38292 20502 38344
rect 20714 38292 20720 38344
rect 20772 38292 20778 38344
rect 20806 38292 20812 38344
rect 20864 38332 20870 38344
rect 20993 38335 21051 38341
rect 20993 38332 21005 38335
rect 20864 38304 21005 38332
rect 20864 38292 20870 38304
rect 20993 38301 21005 38304
rect 21039 38301 21051 38335
rect 20993 38295 21051 38301
rect 21269 38335 21327 38341
rect 21269 38301 21281 38335
rect 21315 38301 21327 38335
rect 21269 38295 21327 38301
rect 21284 38264 21312 38295
rect 15212 38236 18092 38264
rect 20548 38236 21312 38264
rect 15212 38208 15240 38236
rect 2682 38156 2688 38208
rect 2740 38156 2746 38208
rect 4893 38199 4951 38205
rect 4893 38165 4905 38199
rect 4939 38196 4951 38199
rect 4982 38196 4988 38208
rect 4939 38168 4988 38196
rect 4939 38165 4951 38168
rect 4893 38159 4951 38165
rect 4982 38156 4988 38168
rect 5040 38156 5046 38208
rect 5258 38156 5264 38208
rect 5316 38156 5322 38208
rect 6365 38199 6423 38205
rect 6365 38165 6377 38199
rect 6411 38196 6423 38199
rect 6546 38196 6552 38208
rect 6411 38168 6552 38196
rect 6411 38165 6423 38168
rect 6365 38159 6423 38165
rect 6546 38156 6552 38168
rect 6604 38156 6610 38208
rect 7190 38156 7196 38208
rect 7248 38156 7254 38208
rect 7742 38156 7748 38208
rect 7800 38156 7806 38208
rect 8202 38156 8208 38208
rect 8260 38196 8266 38208
rect 14826 38196 14832 38208
rect 8260 38168 14832 38196
rect 8260 38156 8266 38168
rect 14826 38156 14832 38168
rect 14884 38156 14890 38208
rect 15194 38156 15200 38208
rect 15252 38156 15258 38208
rect 20548 38205 20576 38236
rect 20533 38199 20591 38205
rect 20533 38165 20545 38199
rect 20579 38165 20591 38199
rect 20533 38159 20591 38165
rect 20809 38199 20867 38205
rect 20809 38165 20821 38199
rect 20855 38196 20867 38199
rect 21082 38196 21088 38208
rect 20855 38168 21088 38196
rect 20855 38165 20867 38168
rect 20809 38159 20867 38165
rect 21082 38156 21088 38168
rect 21140 38156 21146 38208
rect 21453 38199 21511 38205
rect 21453 38165 21465 38199
rect 21499 38196 21511 38199
rect 22186 38196 22192 38208
rect 21499 38168 22192 38196
rect 21499 38165 21511 38168
rect 21453 38159 21511 38165
rect 22186 38156 22192 38168
rect 22244 38156 22250 38208
rect 1104 38106 22056 38128
rect 1104 38054 6148 38106
rect 6200 38054 6212 38106
rect 6264 38054 6276 38106
rect 6328 38054 6340 38106
rect 6392 38054 6404 38106
rect 6456 38054 11346 38106
rect 11398 38054 11410 38106
rect 11462 38054 11474 38106
rect 11526 38054 11538 38106
rect 11590 38054 11602 38106
rect 11654 38054 16544 38106
rect 16596 38054 16608 38106
rect 16660 38054 16672 38106
rect 16724 38054 16736 38106
rect 16788 38054 16800 38106
rect 16852 38054 21742 38106
rect 21794 38054 21806 38106
rect 21858 38054 21870 38106
rect 21922 38054 21934 38106
rect 21986 38054 21998 38106
rect 22050 38054 22056 38106
rect 1104 38032 22056 38054
rect 3234 37952 3240 38004
rect 3292 37992 3298 38004
rect 3789 37995 3847 38001
rect 3789 37992 3801 37995
rect 3292 37964 3801 37992
rect 3292 37952 3298 37964
rect 3789 37961 3801 37964
rect 3835 37961 3847 37995
rect 3789 37955 3847 37961
rect 5994 37952 6000 38004
rect 6052 37952 6058 38004
rect 8205 37995 8263 38001
rect 8205 37992 8217 37995
rect 6196 37964 8217 37992
rect 6196 37924 6224 37964
rect 8205 37961 8217 37964
rect 8251 37961 8263 37995
rect 10042 37992 10048 38004
rect 8205 37955 8263 37961
rect 9692 37964 10048 37992
rect 3896 37896 6224 37924
rect 3896 37868 3924 37896
rect 1397 37859 1455 37865
rect 1397 37825 1409 37859
rect 1443 37856 1455 37859
rect 1486 37856 1492 37868
rect 1443 37828 1492 37856
rect 1443 37825 1455 37828
rect 1397 37819 1455 37825
rect 1486 37816 1492 37828
rect 1544 37816 1550 37868
rect 3142 37816 3148 37868
rect 3200 37816 3206 37868
rect 3878 37816 3884 37868
rect 3936 37816 3942 37868
rect 4890 37856 4896 37868
rect 4851 37828 4896 37856
rect 4890 37816 4896 37828
rect 4948 37816 4954 37868
rect 6196 37865 6224 37896
rect 7098 37884 7104 37936
rect 7156 37884 7162 37936
rect 7377 37927 7435 37933
rect 7377 37893 7389 37927
rect 7423 37893 7435 37927
rect 7377 37887 7435 37893
rect 7469 37927 7527 37933
rect 7469 37893 7481 37927
rect 7515 37924 7527 37927
rect 7515 37896 8156 37924
rect 7515 37893 7527 37896
rect 7469 37887 7527 37893
rect 6181 37859 6239 37865
rect 6181 37825 6193 37859
rect 6227 37825 6239 37859
rect 6181 37819 6239 37825
rect 6270 37816 6276 37868
rect 6328 37856 6334 37868
rect 7282 37856 7288 37868
rect 6328 37828 7288 37856
rect 6328 37816 6334 37828
rect 7282 37816 7288 37828
rect 7340 37816 7346 37868
rect 7392 37856 7420 37887
rect 7650 37856 7656 37868
rect 7392 37828 7656 37856
rect 7650 37816 7656 37828
rect 7708 37816 7714 37868
rect 7834 37816 7840 37868
rect 7892 37816 7898 37868
rect 8128 37856 8156 37896
rect 8294 37856 8300 37868
rect 8128 37828 8300 37856
rect 8294 37816 8300 37828
rect 8352 37816 8358 37868
rect 9692 37865 9720 37964
rect 10042 37952 10048 37964
rect 10100 37992 10106 38004
rect 15838 37992 15844 38004
rect 10100 37964 15844 37992
rect 10100 37952 10106 37964
rect 15838 37952 15844 37964
rect 15896 37952 15902 38004
rect 18598 37952 18604 38004
rect 18656 37952 18662 38004
rect 19889 37995 19947 38001
rect 19889 37961 19901 37995
rect 19935 37992 19947 37995
rect 20162 37992 20168 38004
rect 19935 37964 20168 37992
rect 19935 37961 19947 37964
rect 19889 37955 19947 37961
rect 20162 37952 20168 37964
rect 20220 37952 20226 38004
rect 20533 37995 20591 38001
rect 20533 37961 20545 37995
rect 20579 37992 20591 37995
rect 20714 37992 20720 38004
rect 20579 37964 20720 37992
rect 20579 37961 20591 37964
rect 20533 37955 20591 37961
rect 20714 37952 20720 37964
rect 20772 37952 20778 38004
rect 13538 37924 13544 37936
rect 13004 37896 13544 37924
rect 9677 37859 9735 37865
rect 9677 37825 9689 37859
rect 9723 37825 9735 37859
rect 9677 37819 9735 37825
rect 9951 37859 10009 37865
rect 9951 37825 9963 37859
rect 9997 37856 10009 37859
rect 11238 37856 11244 37868
rect 9997 37828 11244 37856
rect 9997 37825 10009 37828
rect 9951 37819 10009 37825
rect 11238 37816 11244 37828
rect 11296 37816 11302 37868
rect 12250 37816 12256 37868
rect 12308 37856 12314 37868
rect 13004 37865 13032 37896
rect 13538 37884 13544 37896
rect 13596 37884 13602 37936
rect 14182 37884 14188 37936
rect 14240 37924 14246 37936
rect 14240 37896 14504 37924
rect 14240 37884 14246 37896
rect 12989 37859 13047 37865
rect 12989 37856 13001 37859
rect 12308 37828 13001 37856
rect 12308 37816 12314 37828
rect 12989 37825 13001 37828
rect 13035 37825 13047 37859
rect 12989 37819 13047 37825
rect 13170 37816 13176 37868
rect 13228 37856 13234 37868
rect 13263 37859 13321 37865
rect 13263 37856 13275 37859
rect 13228 37828 13275 37856
rect 13228 37816 13234 37828
rect 13263 37825 13275 37828
rect 13309 37856 13321 37859
rect 14476 37856 14504 37896
rect 14827 37869 14885 37875
rect 14827 37856 14839 37869
rect 13309 37828 14410 37856
rect 14476 37835 14839 37856
rect 14873 37856 14885 37869
rect 15194 37856 15200 37868
rect 14873 37835 15200 37856
rect 14476 37828 15200 37835
rect 13309 37825 13321 37828
rect 13263 37819 13321 37825
rect 1673 37791 1731 37797
rect 1673 37757 1685 37791
rect 1719 37788 1731 37791
rect 1854 37788 1860 37800
rect 1719 37760 1860 37788
rect 1719 37757 1731 37760
rect 1673 37751 1731 37757
rect 1854 37748 1860 37760
rect 1912 37748 1918 37800
rect 1949 37791 2007 37797
rect 1949 37757 1961 37791
rect 1995 37757 2007 37791
rect 1949 37751 2007 37757
rect 2133 37791 2191 37797
rect 2133 37757 2145 37791
rect 2179 37757 2191 37791
rect 2133 37751 2191 37757
rect 1964 37652 1992 37751
rect 2148 37720 2176 37751
rect 2498 37748 2504 37800
rect 2556 37788 2562 37800
rect 2593 37791 2651 37797
rect 2593 37788 2605 37791
rect 2556 37760 2605 37788
rect 2556 37748 2562 37760
rect 2593 37757 2605 37760
rect 2639 37757 2651 37791
rect 2593 37751 2651 37757
rect 2866 37748 2872 37800
rect 2924 37748 2930 37800
rect 3007 37791 3065 37797
rect 3007 37757 3019 37791
rect 3053 37788 3065 37791
rect 3053 37760 4108 37788
rect 3053 37757 3065 37760
rect 3007 37751 3065 37757
rect 2406 37720 2412 37732
rect 2148 37692 2412 37720
rect 2406 37680 2412 37692
rect 2464 37680 2470 37732
rect 4080 37720 4108 37760
rect 4154 37748 4160 37800
rect 4212 37788 4218 37800
rect 4617 37791 4675 37797
rect 4617 37788 4629 37791
rect 4212 37760 4629 37788
rect 4212 37748 4218 37760
rect 4617 37757 4629 37760
rect 4663 37757 4675 37791
rect 4617 37751 4675 37757
rect 7742 37748 7748 37800
rect 7800 37748 7806 37800
rect 4080 37692 4660 37720
rect 3142 37652 3148 37664
rect 1964 37624 3148 37652
rect 3142 37612 3148 37624
rect 3200 37612 3206 37664
rect 4522 37612 4528 37664
rect 4580 37612 4586 37664
rect 4632 37652 4660 37692
rect 5276 37692 6960 37720
rect 5276 37652 5304 37692
rect 6932 37664 6960 37692
rect 4632 37624 5304 37652
rect 5534 37612 5540 37664
rect 5592 37652 5598 37664
rect 5629 37655 5687 37661
rect 5629 37652 5641 37655
rect 5592 37624 5641 37652
rect 5592 37612 5598 37624
rect 5629 37621 5641 37624
rect 5675 37621 5687 37655
rect 5629 37615 5687 37621
rect 6638 37612 6644 37664
rect 6696 37612 6702 37664
rect 6914 37612 6920 37664
rect 6972 37612 6978 37664
rect 8389 37655 8447 37661
rect 8389 37621 8401 37655
rect 8435 37652 8447 37655
rect 8478 37652 8484 37664
rect 8435 37624 8484 37652
rect 8435 37621 8447 37624
rect 8389 37615 8447 37621
rect 8478 37612 8484 37624
rect 8536 37652 8542 37664
rect 9214 37652 9220 37664
rect 8536 37624 9220 37652
rect 8536 37612 8542 37624
rect 9214 37612 9220 37624
rect 9272 37612 9278 37664
rect 10686 37612 10692 37664
rect 10744 37612 10750 37664
rect 11146 37612 11152 37664
rect 11204 37652 11210 37664
rect 12066 37652 12072 37664
rect 11204 37624 12072 37652
rect 11204 37612 11210 37624
rect 12066 37612 12072 37624
rect 12124 37612 12130 37664
rect 14001 37655 14059 37661
rect 14001 37621 14013 37655
rect 14047 37652 14059 37655
rect 14274 37652 14280 37664
rect 14047 37624 14280 37652
rect 14047 37621 14059 37624
rect 14001 37615 14059 37621
rect 14274 37612 14280 37624
rect 14332 37612 14338 37664
rect 14382 37652 14410 37828
rect 15194 37816 15200 37828
rect 15252 37816 15258 37868
rect 18782 37816 18788 37868
rect 18840 37816 18846 37868
rect 20070 37816 20076 37868
rect 20128 37816 20134 37868
rect 20162 37816 20168 37868
rect 20220 37856 20226 37868
rect 20441 37859 20499 37865
rect 20441 37856 20453 37859
rect 20220 37828 20453 37856
rect 20220 37816 20226 37828
rect 20441 37825 20453 37828
rect 20487 37825 20499 37859
rect 20441 37819 20499 37825
rect 20714 37816 20720 37868
rect 20772 37816 20778 37868
rect 20990 37816 20996 37868
rect 21048 37816 21054 37868
rect 21174 37816 21180 37868
rect 21232 37856 21238 37868
rect 21269 37859 21327 37865
rect 21269 37856 21281 37859
rect 21232 37828 21281 37856
rect 21232 37816 21238 37828
rect 21269 37825 21281 37828
rect 21315 37825 21327 37859
rect 21269 37819 21327 37825
rect 14550 37748 14556 37800
rect 14608 37748 14614 37800
rect 19702 37748 19708 37800
rect 19760 37788 19766 37800
rect 20806 37788 20812 37800
rect 19760 37760 20812 37788
rect 19760 37748 19766 37760
rect 20806 37748 20812 37760
rect 20864 37748 20870 37800
rect 18322 37720 18328 37732
rect 15212 37692 18328 37720
rect 15212 37652 15240 37692
rect 18322 37680 18328 37692
rect 18380 37680 18386 37732
rect 20257 37723 20315 37729
rect 20257 37689 20269 37723
rect 20303 37720 20315 37723
rect 20898 37720 20904 37732
rect 20303 37692 20904 37720
rect 20303 37689 20315 37692
rect 20257 37683 20315 37689
rect 20898 37680 20904 37692
rect 20956 37680 20962 37732
rect 14382 37624 15240 37652
rect 15562 37612 15568 37664
rect 15620 37612 15626 37664
rect 20806 37612 20812 37664
rect 20864 37612 20870 37664
rect 21450 37612 21456 37664
rect 21508 37612 21514 37664
rect 1104 37562 21896 37584
rect 1104 37510 3549 37562
rect 3601 37510 3613 37562
rect 3665 37510 3677 37562
rect 3729 37510 3741 37562
rect 3793 37510 3805 37562
rect 3857 37510 8747 37562
rect 8799 37510 8811 37562
rect 8863 37510 8875 37562
rect 8927 37510 8939 37562
rect 8991 37510 9003 37562
rect 9055 37510 13945 37562
rect 13997 37510 14009 37562
rect 14061 37510 14073 37562
rect 14125 37510 14137 37562
rect 14189 37510 14201 37562
rect 14253 37510 19143 37562
rect 19195 37510 19207 37562
rect 19259 37510 19271 37562
rect 19323 37510 19335 37562
rect 19387 37510 19399 37562
rect 19451 37510 21896 37562
rect 1104 37488 21896 37510
rect 1854 37408 1860 37460
rect 1912 37448 1918 37460
rect 4246 37448 4252 37460
rect 1912 37420 4252 37448
rect 1912 37408 1918 37420
rect 4246 37408 4252 37420
rect 4304 37408 4310 37460
rect 5442 37448 5448 37460
rect 4354 37420 5448 37448
rect 2314 37340 2320 37392
rect 2372 37380 2378 37392
rect 2866 37380 2872 37392
rect 2372 37352 2872 37380
rect 2372 37340 2378 37352
rect 2866 37340 2872 37352
rect 2924 37380 2930 37392
rect 4354 37380 4382 37420
rect 5442 37408 5448 37420
rect 5500 37408 5506 37460
rect 5718 37408 5724 37460
rect 5776 37408 5782 37460
rect 11517 37451 11575 37457
rect 11517 37417 11529 37451
rect 11563 37448 11575 37451
rect 13998 37448 14004 37460
rect 11563 37420 14004 37448
rect 11563 37417 11575 37420
rect 11517 37411 11575 37417
rect 13998 37408 14004 37420
rect 14056 37408 14062 37460
rect 19702 37408 19708 37460
rect 19760 37408 19766 37460
rect 19981 37451 20039 37457
rect 19981 37417 19993 37451
rect 20027 37448 20039 37451
rect 20162 37448 20168 37460
rect 20027 37420 20168 37448
rect 20027 37417 20039 37420
rect 19981 37411 20039 37417
rect 20162 37408 20168 37420
rect 20220 37408 20226 37460
rect 20257 37451 20315 37457
rect 20257 37417 20269 37451
rect 20303 37448 20315 37451
rect 20438 37448 20444 37460
rect 20303 37420 20444 37448
rect 20303 37417 20315 37420
rect 20257 37411 20315 37417
rect 20438 37408 20444 37420
rect 20496 37408 20502 37460
rect 20533 37451 20591 37457
rect 20533 37417 20545 37451
rect 20579 37448 20591 37451
rect 20714 37448 20720 37460
rect 20579 37420 20720 37448
rect 20579 37417 20591 37420
rect 20533 37411 20591 37417
rect 20714 37408 20720 37420
rect 20772 37408 20778 37460
rect 2924 37352 4382 37380
rect 2924 37340 2930 37352
rect 4430 37340 4436 37392
rect 4488 37340 4494 37392
rect 4522 37340 4528 37392
rect 4580 37340 4586 37392
rect 15654 37340 15660 37392
rect 15712 37380 15718 37392
rect 16942 37380 16948 37392
rect 15712 37352 16948 37380
rect 15712 37340 15718 37352
rect 16942 37340 16948 37352
rect 17000 37340 17006 37392
rect 4062 37312 4068 37324
rect 2976 37284 4068 37312
rect 1489 37247 1547 37253
rect 1489 37213 1501 37247
rect 1535 37213 1547 37247
rect 1489 37207 1547 37213
rect 1763 37247 1821 37253
rect 1763 37213 1775 37247
rect 1809 37244 1821 37247
rect 2976 37244 3004 37284
rect 4062 37272 4068 37284
rect 4120 37272 4126 37324
rect 4540 37312 4568 37340
rect 4709 37315 4767 37321
rect 4709 37312 4721 37315
rect 4540 37284 4721 37312
rect 4709 37281 4721 37284
rect 4755 37281 4767 37315
rect 4709 37275 4767 37281
rect 4982 37272 4988 37324
rect 5040 37272 5046 37324
rect 5629 37315 5687 37321
rect 5629 37281 5641 37315
rect 5675 37312 5687 37315
rect 5675 37284 5856 37312
rect 5675 37281 5687 37284
rect 5629 37275 5687 37281
rect 1809 37216 3004 37244
rect 1809 37213 1821 37216
rect 1763 37207 1821 37213
rect 1504 37176 1532 37207
rect 3050 37204 3056 37256
rect 3108 37204 3114 37256
rect 3142 37204 3148 37256
rect 3200 37244 3206 37256
rect 3789 37247 3847 37253
rect 3789 37244 3801 37247
rect 3200 37216 3801 37244
rect 3200 37204 3206 37216
rect 3789 37213 3801 37216
rect 3835 37244 3847 37247
rect 3835 37216 3924 37244
rect 3835 37213 3847 37216
rect 3789 37207 3847 37213
rect 1504 37148 1900 37176
rect 1872 37120 1900 37148
rect 3234 37136 3240 37188
rect 3292 37176 3298 37188
rect 3329 37179 3387 37185
rect 3329 37176 3341 37179
rect 3292 37148 3341 37176
rect 3292 37136 3298 37148
rect 3329 37145 3341 37148
rect 3375 37145 3387 37179
rect 3329 37139 3387 37145
rect 3896 37120 3924 37216
rect 3970 37204 3976 37256
rect 4028 37204 4034 37256
rect 4890 37253 4896 37256
rect 4847 37247 4896 37253
rect 4847 37213 4859 37247
rect 4893 37213 4896 37247
rect 4847 37207 4896 37213
rect 4862 37206 4896 37207
rect 4890 37204 4896 37206
rect 4948 37204 4954 37256
rect 1854 37068 1860 37120
rect 1912 37068 1918 37120
rect 2501 37111 2559 37117
rect 2501 37077 2513 37111
rect 2547 37108 2559 37111
rect 2958 37108 2964 37120
rect 2547 37080 2964 37108
rect 2547 37077 2559 37080
rect 2501 37071 2559 37077
rect 2958 37068 2964 37080
rect 3016 37068 3022 37120
rect 3878 37068 3884 37120
rect 3936 37068 3942 37120
rect 3988 37108 4016 37204
rect 5828 37176 5856 37284
rect 6546 37272 6552 37324
rect 6604 37272 6610 37324
rect 7374 37272 7380 37324
rect 7432 37272 7438 37324
rect 9950 37312 9956 37324
rect 7484 37284 9956 37312
rect 5905 37247 5963 37253
rect 5905 37213 5917 37247
rect 5951 37244 5963 37247
rect 6362 37244 6368 37256
rect 5951 37216 6368 37244
rect 5951 37213 5963 37216
rect 5905 37207 5963 37213
rect 6362 37204 6368 37216
rect 6420 37204 6426 37256
rect 6457 37247 6515 37253
rect 6457 37213 6469 37247
rect 6503 37244 6515 37247
rect 6638 37244 6644 37256
rect 6503 37216 6644 37244
rect 6503 37213 6515 37216
rect 6457 37207 6515 37213
rect 6638 37204 6644 37216
rect 6696 37204 6702 37256
rect 7392 37244 7420 37272
rect 6840 37216 7420 37244
rect 6549 37179 6607 37185
rect 5828 37148 6500 37176
rect 4706 37108 4712 37120
rect 3988 37080 4712 37108
rect 4706 37068 4712 37080
rect 4764 37068 4770 37120
rect 5442 37068 5448 37120
rect 5500 37108 5506 37120
rect 6181 37111 6239 37117
rect 6181 37108 6193 37111
rect 5500 37080 6193 37108
rect 5500 37068 5506 37080
rect 6181 37077 6193 37080
rect 6227 37108 6239 37111
rect 6270 37108 6276 37120
rect 6227 37080 6276 37108
rect 6227 37077 6239 37080
rect 6181 37071 6239 37077
rect 6270 37068 6276 37080
rect 6328 37068 6334 37120
rect 6472 37108 6500 37148
rect 6549 37145 6561 37179
rect 6595 37176 6607 37179
rect 6840 37176 6868 37216
rect 6595 37148 6868 37176
rect 6595 37145 6607 37148
rect 6549 37139 6607 37145
rect 6914 37136 6920 37188
rect 6972 37136 6978 37188
rect 7484 37176 7512 37284
rect 9950 37272 9956 37284
rect 10008 37272 10014 37324
rect 10686 37272 10692 37324
rect 10744 37272 10750 37324
rect 12250 37272 12256 37324
rect 12308 37312 12314 37324
rect 12345 37315 12403 37321
rect 12345 37312 12357 37315
rect 12308 37284 12357 37312
rect 12308 37272 12314 37284
rect 12345 37281 12357 37284
rect 12391 37281 12403 37315
rect 12345 37275 12403 37281
rect 13078 37272 13084 37324
rect 13136 37312 13142 37324
rect 13136 37284 13676 37312
rect 13136 37272 13142 37284
rect 10505 37247 10563 37253
rect 10505 37213 10517 37247
rect 10551 37244 10563 37247
rect 10870 37244 10876 37256
rect 10551 37216 10876 37244
rect 10551 37213 10563 37216
rect 10505 37207 10563 37213
rect 10870 37204 10876 37216
rect 10928 37204 10934 37256
rect 11698 37204 11704 37256
rect 11756 37204 11762 37256
rect 12603 37217 12661 37223
rect 7024 37148 7512 37176
rect 7024 37108 7052 37148
rect 10410 37136 10416 37188
rect 10468 37176 10474 37188
rect 10597 37179 10655 37185
rect 10597 37176 10609 37179
rect 10468 37148 10609 37176
rect 10468 37136 10474 37148
rect 10597 37145 10609 37148
rect 10643 37145 10655 37179
rect 10597 37139 10655 37145
rect 10962 37136 10968 37188
rect 11020 37136 11026 37188
rect 12603 37183 12615 37217
rect 12649 37188 12661 37217
rect 12603 37177 12624 37183
rect 12618 37136 12624 37177
rect 12676 37176 12682 37188
rect 13648 37176 13676 37284
rect 15562 37272 15568 37324
rect 15620 37312 15626 37324
rect 15620 37284 16068 37312
rect 15620 37272 15626 37284
rect 14277 37247 14335 37253
rect 14277 37213 14289 37247
rect 14323 37244 14335 37247
rect 15102 37244 15108 37256
rect 14323 37216 15108 37244
rect 14323 37213 14335 37216
rect 14277 37207 14335 37213
rect 15102 37204 15108 37216
rect 15160 37204 15166 37256
rect 15746 37204 15752 37256
rect 15804 37204 15810 37256
rect 16040 37253 16068 37284
rect 16132 37284 16436 37312
rect 16025 37247 16083 37253
rect 16025 37213 16037 37247
rect 16071 37213 16083 37247
rect 16025 37207 16083 37213
rect 14550 37185 14556 37188
rect 14522 37179 14556 37185
rect 14522 37176 14534 37179
rect 12676 37148 13584 37176
rect 13648 37148 14534 37176
rect 12676 37136 12682 37148
rect 6472 37080 7052 37108
rect 7098 37068 7104 37120
rect 7156 37108 7162 37120
rect 7285 37111 7343 37117
rect 7285 37108 7297 37111
rect 7156 37080 7297 37108
rect 7156 37068 7162 37080
rect 7285 37077 7297 37080
rect 7331 37077 7343 37111
rect 7285 37071 7343 37077
rect 7469 37111 7527 37117
rect 7469 37077 7481 37111
rect 7515 37108 7527 37111
rect 7742 37108 7748 37120
rect 7515 37080 7748 37108
rect 7515 37077 7527 37080
rect 7469 37071 7527 37077
rect 7742 37068 7748 37080
rect 7800 37068 7806 37120
rect 8570 37068 8576 37120
rect 8628 37108 8634 37120
rect 8846 37108 8852 37120
rect 8628 37080 8852 37108
rect 8628 37068 8634 37080
rect 8846 37068 8852 37080
rect 8904 37068 8910 37120
rect 9766 37068 9772 37120
rect 9824 37068 9830 37120
rect 10226 37068 10232 37120
rect 10284 37068 10290 37120
rect 11330 37068 11336 37120
rect 11388 37068 11394 37120
rect 11885 37111 11943 37117
rect 11885 37077 11897 37111
rect 11931 37108 11943 37111
rect 12066 37108 12072 37120
rect 11931 37080 12072 37108
rect 11931 37077 11943 37080
rect 11885 37071 11943 37077
rect 12066 37068 12072 37080
rect 12124 37068 12130 37120
rect 13357 37111 13415 37117
rect 13357 37077 13369 37111
rect 13403 37108 13415 37111
rect 13446 37108 13452 37120
rect 13403 37080 13452 37108
rect 13403 37077 13415 37080
rect 13357 37071 13415 37077
rect 13446 37068 13452 37080
rect 13504 37068 13510 37120
rect 13556 37108 13584 37148
rect 14522 37145 14534 37148
rect 14522 37139 14556 37145
rect 14550 37136 14556 37139
rect 14608 37136 14614 37188
rect 16132 37176 16160 37284
rect 16209 37247 16267 37253
rect 16209 37213 16221 37247
rect 16255 37244 16267 37247
rect 16408 37244 16436 37284
rect 19812 37284 20024 37312
rect 16485 37247 16543 37253
rect 16485 37244 16497 37247
rect 16255 37216 16344 37244
rect 16408 37216 16497 37244
rect 16255 37213 16267 37216
rect 16209 37207 16267 37213
rect 15672 37148 16160 37176
rect 13906 37108 13912 37120
rect 13556 37080 13912 37108
rect 13906 37068 13912 37080
rect 13964 37068 13970 37120
rect 13998 37068 14004 37120
rect 14056 37108 14062 37120
rect 14366 37108 14372 37120
rect 14056 37080 14372 37108
rect 14056 37068 14062 37080
rect 14366 37068 14372 37080
rect 14424 37068 14430 37120
rect 15672 37117 15700 37148
rect 15657 37111 15715 37117
rect 15657 37077 15669 37111
rect 15703 37077 15715 37111
rect 15657 37071 15715 37077
rect 15838 37068 15844 37120
rect 15896 37068 15902 37120
rect 16114 37068 16120 37120
rect 16172 37068 16178 37120
rect 16316 37117 16344 37216
rect 16485 37213 16497 37216
rect 16531 37213 16543 37247
rect 16485 37207 16543 37213
rect 17218 37204 17224 37256
rect 17276 37204 17282 37256
rect 17862 37204 17868 37256
rect 17920 37204 17926 37256
rect 17957 37247 18015 37253
rect 17957 37213 17969 37247
rect 18003 37244 18015 37247
rect 18046 37244 18052 37256
rect 18003 37216 18052 37244
rect 18003 37213 18015 37216
rect 17957 37207 18015 37213
rect 18046 37204 18052 37216
rect 18104 37204 18110 37256
rect 18141 37247 18199 37253
rect 18141 37213 18153 37247
rect 18187 37213 18199 37247
rect 18141 37207 18199 37213
rect 18156 37176 18184 37207
rect 18230 37204 18236 37256
rect 18288 37244 18294 37256
rect 18969 37247 19027 37253
rect 18969 37244 18981 37247
rect 18288 37216 18981 37244
rect 18288 37204 18294 37216
rect 18969 37213 18981 37216
rect 19015 37213 19027 37247
rect 18969 37207 19027 37213
rect 19702 37204 19708 37256
rect 19760 37244 19766 37256
rect 19812 37244 19840 37284
rect 19760 37216 19840 37244
rect 19889 37247 19947 37253
rect 19760 37204 19766 37216
rect 19889 37213 19901 37247
rect 19935 37213 19947 37247
rect 19996 37244 20024 37284
rect 20165 37247 20223 37253
rect 20165 37244 20177 37247
rect 19996 37216 20177 37244
rect 19889 37207 19947 37213
rect 20165 37213 20177 37216
rect 20211 37213 20223 37247
rect 20165 37207 20223 37213
rect 19904 37176 19932 37207
rect 20438 37204 20444 37256
rect 20496 37204 20502 37256
rect 20530 37204 20536 37256
rect 20588 37244 20594 37256
rect 20717 37247 20775 37253
rect 20717 37244 20729 37247
rect 20588 37216 20729 37244
rect 20588 37204 20594 37216
rect 20717 37213 20729 37216
rect 20763 37213 20775 37247
rect 20717 37207 20775 37213
rect 20898 37204 20904 37256
rect 20956 37244 20962 37256
rect 20993 37247 21051 37253
rect 20993 37244 21005 37247
rect 20956 37216 21005 37244
rect 20956 37204 20962 37216
rect 20993 37213 21005 37216
rect 21039 37213 21051 37247
rect 20993 37207 21051 37213
rect 21082 37204 21088 37256
rect 21140 37244 21146 37256
rect 21177 37247 21235 37253
rect 21177 37244 21189 37247
rect 21140 37216 21189 37244
rect 21140 37204 21146 37216
rect 21177 37213 21189 37216
rect 21223 37213 21235 37247
rect 21177 37207 21235 37213
rect 17696 37148 18184 37176
rect 18800 37148 19932 37176
rect 21545 37179 21603 37185
rect 16301 37111 16359 37117
rect 16301 37077 16313 37111
rect 16347 37077 16359 37111
rect 16301 37071 16359 37077
rect 17310 37068 17316 37120
rect 17368 37068 17374 37120
rect 17696 37117 17724 37148
rect 17681 37111 17739 37117
rect 17681 37077 17693 37111
rect 17727 37077 17739 37111
rect 17681 37071 17739 37077
rect 18138 37068 18144 37120
rect 18196 37068 18202 37120
rect 18800 37117 18828 37148
rect 21545 37145 21557 37179
rect 21591 37176 21603 37179
rect 22278 37176 22284 37188
rect 21591 37148 22284 37176
rect 21591 37145 21603 37148
rect 21545 37139 21603 37145
rect 22278 37136 22284 37148
rect 22336 37136 22342 37188
rect 18785 37111 18843 37117
rect 18785 37077 18797 37111
rect 18831 37077 18843 37111
rect 18785 37071 18843 37077
rect 20809 37111 20867 37117
rect 20809 37077 20821 37111
rect 20855 37108 20867 37111
rect 21082 37108 21088 37120
rect 20855 37080 21088 37108
rect 20855 37077 20867 37080
rect 20809 37071 20867 37077
rect 21082 37068 21088 37080
rect 21140 37068 21146 37120
rect 1104 37018 22056 37040
rect 1104 36966 6148 37018
rect 6200 36966 6212 37018
rect 6264 36966 6276 37018
rect 6328 36966 6340 37018
rect 6392 36966 6404 37018
rect 6456 36966 11346 37018
rect 11398 36966 11410 37018
rect 11462 36966 11474 37018
rect 11526 36966 11538 37018
rect 11590 36966 11602 37018
rect 11654 36966 16544 37018
rect 16596 36966 16608 37018
rect 16660 36966 16672 37018
rect 16724 36966 16736 37018
rect 16788 36966 16800 37018
rect 16852 36966 21742 37018
rect 21794 36966 21806 37018
rect 21858 36966 21870 37018
rect 21922 36966 21934 37018
rect 21986 36966 21998 37018
rect 22050 36966 22056 37018
rect 1104 36944 22056 36966
rect 3786 36904 3792 36916
rect 584 36876 3792 36904
rect 584 36780 612 36876
rect 3786 36864 3792 36876
rect 3844 36864 3850 36916
rect 5626 36864 5632 36916
rect 5684 36904 5690 36916
rect 5997 36907 6055 36913
rect 5997 36904 6009 36907
rect 5684 36876 6009 36904
rect 5684 36864 5690 36876
rect 5997 36873 6009 36876
rect 6043 36873 6055 36907
rect 5997 36867 6055 36873
rect 8294 36864 8300 36916
rect 8352 36864 8358 36916
rect 9950 36904 9956 36916
rect 8680 36876 9956 36904
rect 1688 36808 6960 36836
rect 1688 36780 1716 36808
rect 566 36728 572 36780
rect 624 36728 630 36780
rect 1670 36728 1676 36780
rect 1728 36728 1734 36780
rect 2498 36728 2504 36780
rect 2556 36768 2562 36780
rect 2927 36771 2985 36777
rect 2927 36768 2939 36771
rect 2556 36740 2939 36768
rect 2556 36728 2562 36740
rect 2927 36737 2939 36740
rect 2973 36768 2985 36771
rect 3326 36768 3332 36780
rect 2973 36740 3332 36768
rect 2973 36737 2985 36740
rect 2927 36731 2985 36737
rect 3326 36728 3332 36740
rect 3384 36728 3390 36780
rect 4338 36768 4344 36780
rect 4299 36740 4344 36768
rect 4338 36728 4344 36740
rect 4396 36728 4402 36780
rect 4890 36728 4896 36780
rect 4948 36768 4954 36780
rect 5442 36768 5448 36780
rect 4948 36740 5448 36768
rect 4948 36728 4954 36740
rect 5442 36728 5448 36740
rect 5500 36728 5506 36780
rect 5721 36771 5779 36777
rect 5721 36737 5733 36771
rect 5767 36768 5779 36771
rect 5994 36768 6000 36780
rect 5767 36740 6000 36768
rect 5767 36737 5779 36740
rect 5721 36731 5779 36737
rect 5994 36728 6000 36740
rect 6052 36768 6058 36780
rect 6181 36771 6239 36777
rect 6181 36768 6193 36771
rect 6052 36740 6193 36768
rect 6052 36728 6058 36740
rect 6181 36737 6193 36740
rect 6227 36737 6239 36771
rect 6181 36731 6239 36737
rect 6362 36728 6368 36780
rect 6420 36728 6426 36780
rect 6932 36772 6960 36808
rect 7558 36777 7564 36780
rect 6932 36768 7052 36772
rect 7527 36771 7564 36777
rect 7527 36768 7539 36771
rect 6932 36744 7539 36768
rect 7024 36740 7539 36744
rect 7527 36737 7539 36740
rect 7527 36731 7564 36737
rect 7558 36728 7564 36731
rect 7616 36728 7622 36780
rect 7650 36728 7656 36780
rect 7708 36768 7714 36780
rect 8680 36777 8708 36876
rect 9950 36864 9956 36876
rect 10008 36864 10014 36916
rect 10226 36864 10232 36916
rect 10284 36904 10290 36916
rect 10284 36876 10362 36904
rect 10284 36864 10290 36876
rect 9122 36796 9128 36848
rect 9180 36836 9186 36848
rect 10334 36836 10362 36876
rect 10410 36864 10416 36916
rect 10468 36904 10474 36916
rect 11057 36907 11115 36913
rect 11057 36904 11069 36907
rect 10468 36876 11069 36904
rect 10468 36864 10474 36876
rect 11057 36873 11069 36876
rect 11103 36873 11115 36907
rect 11057 36867 11115 36873
rect 14550 36864 14556 36916
rect 14608 36864 14614 36916
rect 14829 36907 14887 36913
rect 14829 36873 14841 36907
rect 14875 36904 14887 36907
rect 15746 36904 15752 36916
rect 14875 36876 15752 36904
rect 14875 36873 14887 36876
rect 14829 36867 14887 36873
rect 15746 36864 15752 36876
rect 15804 36864 15810 36916
rect 15838 36864 15844 36916
rect 15896 36864 15902 36916
rect 16114 36864 16120 36916
rect 16172 36864 16178 36916
rect 16209 36907 16267 36913
rect 16209 36873 16221 36907
rect 16255 36904 16267 36907
rect 16390 36904 16396 36916
rect 16255 36876 16396 36904
rect 16255 36873 16267 36876
rect 16209 36867 16267 36873
rect 16390 36864 16396 36876
rect 16448 36864 16454 36916
rect 16574 36864 16580 36916
rect 16632 36904 16638 36916
rect 17218 36904 17224 36916
rect 16632 36876 17224 36904
rect 16632 36864 16638 36876
rect 17218 36864 17224 36876
rect 17276 36864 17282 36916
rect 17310 36864 17316 36916
rect 17368 36864 17374 36916
rect 17862 36864 17868 36916
rect 17920 36904 17926 36916
rect 18049 36907 18107 36913
rect 18049 36904 18061 36907
rect 17920 36876 18061 36904
rect 17920 36864 17926 36876
rect 18049 36873 18061 36876
rect 18095 36873 18107 36907
rect 18049 36867 18107 36873
rect 18138 36864 18144 36916
rect 18196 36864 18202 36916
rect 19889 36907 19947 36913
rect 19889 36873 19901 36907
rect 19935 36873 19947 36907
rect 19889 36867 19947 36873
rect 11609 36839 11667 36845
rect 11609 36836 11621 36839
rect 9180 36808 9996 36836
rect 10334 36808 11621 36836
rect 9180 36796 9186 36808
rect 8665 36771 8723 36777
rect 8665 36768 8677 36771
rect 7708 36740 8677 36768
rect 7708 36728 7714 36740
rect 8665 36737 8677 36740
rect 8711 36737 8723 36771
rect 8665 36731 8723 36737
rect 8846 36728 8852 36780
rect 8904 36768 8910 36780
rect 8939 36771 8997 36777
rect 8939 36768 8951 36771
rect 8904 36740 8951 36768
rect 8904 36728 8910 36740
rect 8939 36737 8951 36740
rect 8985 36768 8997 36771
rect 9398 36768 9404 36780
rect 8985 36740 9404 36768
rect 8985 36737 8997 36740
rect 8939 36731 8997 36737
rect 9398 36728 9404 36740
rect 9456 36728 9462 36780
rect 1854 36660 1860 36712
rect 1912 36700 1918 36712
rect 2406 36700 2412 36712
rect 1912 36672 2412 36700
rect 1912 36660 1918 36672
rect 2406 36660 2412 36672
rect 2464 36700 2470 36712
rect 2685 36703 2743 36709
rect 2685 36700 2697 36703
rect 2464 36672 2697 36700
rect 2464 36660 2470 36672
rect 2685 36669 2697 36672
rect 2731 36669 2743 36703
rect 2685 36663 2743 36669
rect 3418 36660 3424 36712
rect 3476 36660 3482 36712
rect 4062 36660 4068 36712
rect 4120 36660 4126 36712
rect 6549 36703 6607 36709
rect 6549 36700 6561 36703
rect 4908 36672 6561 36700
rect 3436 36632 3464 36660
rect 3436 36604 4200 36632
rect 2406 36524 2412 36576
rect 2464 36564 2470 36576
rect 3697 36567 3755 36573
rect 3697 36564 3709 36567
rect 2464 36536 3709 36564
rect 2464 36524 2470 36536
rect 3697 36533 3709 36536
rect 3743 36533 3755 36567
rect 4172 36564 4200 36604
rect 4908 36564 4936 36672
rect 6549 36669 6561 36672
rect 6595 36700 6607 36703
rect 6822 36700 6828 36712
rect 6595 36672 6828 36700
rect 6595 36669 6607 36672
rect 6549 36663 6607 36669
rect 6822 36660 6828 36672
rect 6880 36660 6886 36712
rect 7190 36660 7196 36712
rect 7248 36700 7254 36712
rect 7285 36703 7343 36709
rect 7285 36700 7297 36703
rect 7248 36672 7297 36700
rect 7248 36660 7254 36672
rect 7285 36669 7297 36672
rect 7331 36669 7343 36703
rect 7285 36663 7343 36669
rect 5442 36592 5448 36644
rect 5500 36632 5506 36644
rect 6914 36632 6920 36644
rect 5500 36604 6920 36632
rect 5500 36592 5506 36604
rect 6914 36592 6920 36604
rect 6972 36592 6978 36644
rect 9508 36604 9904 36632
rect 4172 36536 4936 36564
rect 3697 36527 3755 36533
rect 4982 36524 4988 36576
rect 5040 36564 5046 36576
rect 5077 36567 5135 36573
rect 5077 36564 5089 36567
rect 5040 36536 5089 36564
rect 5040 36524 5046 36536
rect 5077 36533 5089 36536
rect 5123 36533 5135 36567
rect 5077 36527 5135 36533
rect 5718 36524 5724 36576
rect 5776 36564 5782 36576
rect 9508 36564 9536 36604
rect 9876 36576 9904 36604
rect 5776 36536 9536 36564
rect 5776 36524 5782 36536
rect 9582 36524 9588 36576
rect 9640 36564 9646 36576
rect 9677 36567 9735 36573
rect 9677 36564 9689 36567
rect 9640 36536 9689 36564
rect 9640 36524 9646 36536
rect 9677 36533 9689 36536
rect 9723 36533 9735 36567
rect 9677 36527 9735 36533
rect 9858 36524 9864 36576
rect 9916 36524 9922 36576
rect 9968 36564 9996 36808
rect 11609 36805 11621 36808
rect 11655 36836 11667 36839
rect 12986 36836 12992 36848
rect 11655 36808 12992 36836
rect 11655 36805 11667 36808
rect 11609 36799 11667 36805
rect 12986 36796 12992 36808
rect 13044 36796 13050 36848
rect 14568 36836 14596 36864
rect 14568 36808 15056 36836
rect 10042 36728 10048 36780
rect 10100 36728 10106 36780
rect 10226 36728 10232 36780
rect 10284 36768 10290 36780
rect 10319 36771 10377 36777
rect 10319 36768 10331 36771
rect 10284 36740 10331 36768
rect 10284 36728 10290 36740
rect 10319 36737 10331 36740
rect 10365 36768 10377 36771
rect 11698 36768 11704 36780
rect 10365 36740 11704 36768
rect 10365 36737 10377 36740
rect 10319 36731 10377 36737
rect 11698 36728 11704 36740
rect 11756 36728 11762 36780
rect 13998 36777 14004 36780
rect 13955 36771 14004 36777
rect 13955 36737 13967 36771
rect 14001 36737 14004 36771
rect 13955 36731 14004 36737
rect 13998 36728 14004 36731
rect 14056 36728 14062 36780
rect 15028 36777 15056 36808
rect 15013 36771 15071 36777
rect 15013 36737 15025 36771
rect 15059 36737 15071 36771
rect 15013 36731 15071 36737
rect 15102 36728 15108 36780
rect 15160 36768 15166 36780
rect 15657 36771 15715 36777
rect 15160 36740 15608 36768
rect 15160 36728 15166 36740
rect 12897 36703 12955 36709
rect 12897 36669 12909 36703
rect 12943 36669 12955 36703
rect 12897 36663 12955 36669
rect 13081 36703 13139 36709
rect 13081 36669 13093 36703
rect 13127 36700 13139 36703
rect 13170 36700 13176 36712
rect 13127 36672 13176 36700
rect 13127 36669 13139 36672
rect 13081 36663 13139 36669
rect 11790 36592 11796 36644
rect 11848 36592 11854 36644
rect 12912 36632 12940 36663
rect 13170 36660 13176 36672
rect 13228 36660 13234 36712
rect 13446 36660 13452 36712
rect 13504 36700 13510 36712
rect 13541 36703 13599 36709
rect 13541 36700 13553 36703
rect 13504 36672 13553 36700
rect 13504 36660 13510 36672
rect 13541 36669 13553 36672
rect 13587 36669 13599 36703
rect 13541 36663 13599 36669
rect 13630 36660 13636 36712
rect 13688 36660 13694 36712
rect 13814 36660 13820 36712
rect 13872 36660 13878 36712
rect 14093 36703 14151 36709
rect 14093 36669 14105 36703
rect 14139 36700 14151 36703
rect 14274 36700 14280 36712
rect 14139 36672 14280 36700
rect 14139 36669 14151 36672
rect 14093 36663 14151 36669
rect 14274 36660 14280 36672
rect 14332 36660 14338 36712
rect 15473 36703 15531 36709
rect 15473 36669 15485 36703
rect 15519 36669 15531 36703
rect 15580 36700 15608 36740
rect 15657 36737 15669 36771
rect 15703 36768 15715 36771
rect 15856 36768 15884 36864
rect 16025 36839 16083 36845
rect 16025 36805 16037 36839
rect 16071 36836 16083 36839
rect 16132 36836 16160 36864
rect 16071 36808 16160 36836
rect 16071 36805 16083 36808
rect 16025 36799 16083 36805
rect 15703 36740 15884 36768
rect 15933 36771 15991 36777
rect 15703 36737 15715 36740
rect 15657 36731 15715 36737
rect 15933 36737 15945 36771
rect 15979 36768 15991 36771
rect 16298 36768 16304 36780
rect 15979 36740 16304 36768
rect 15979 36737 15991 36740
rect 15933 36731 15991 36737
rect 16298 36728 16304 36740
rect 16356 36728 16362 36780
rect 16390 36728 16396 36780
rect 16448 36728 16454 36780
rect 16482 36728 16488 36780
rect 16540 36768 16546 36780
rect 16925 36771 16983 36777
rect 16925 36768 16937 36771
rect 16540 36740 16937 36768
rect 16540 36728 16546 36740
rect 16925 36737 16937 36740
rect 16971 36737 16983 36771
rect 17328 36768 17356 36864
rect 18156 36836 18184 36864
rect 18693 36839 18751 36845
rect 18693 36836 18705 36839
rect 18156 36808 18705 36836
rect 18693 36805 18705 36808
rect 18739 36805 18751 36839
rect 19904 36836 19932 36867
rect 20806 36864 20812 36916
rect 20864 36864 20870 36916
rect 20901 36907 20959 36913
rect 20901 36873 20913 36907
rect 20947 36904 20959 36907
rect 20990 36904 20996 36916
rect 20947 36876 20996 36904
rect 20947 36873 20959 36876
rect 20901 36867 20959 36873
rect 20990 36864 20996 36876
rect 21048 36864 21054 36916
rect 20824 36836 20852 36864
rect 19904 36808 20760 36836
rect 20824 36808 21312 36836
rect 18693 36799 18751 36805
rect 18325 36771 18383 36777
rect 18325 36768 18337 36771
rect 17328 36740 18337 36768
rect 16925 36731 16983 36737
rect 18325 36737 18337 36740
rect 18371 36737 18383 36771
rect 18325 36731 18383 36737
rect 19610 36728 19616 36780
rect 19668 36768 19674 36780
rect 20073 36771 20131 36777
rect 20073 36768 20085 36771
rect 19668 36740 20085 36768
rect 19668 36728 19674 36740
rect 20073 36737 20085 36740
rect 20119 36737 20131 36771
rect 20073 36731 20131 36737
rect 20346 36728 20352 36780
rect 20404 36728 20410 36780
rect 20533 36772 20591 36777
rect 20533 36771 20668 36772
rect 20533 36737 20545 36771
rect 20579 36744 20668 36771
rect 20579 36737 20591 36744
rect 20533 36731 20591 36737
rect 16669 36703 16727 36709
rect 16669 36700 16681 36703
rect 15580 36672 16681 36700
rect 15473 36663 15531 36669
rect 16669 36669 16681 36672
rect 16715 36669 16727 36703
rect 16669 36663 16727 36669
rect 18141 36703 18199 36709
rect 18141 36669 18153 36703
rect 18187 36669 18199 36703
rect 18141 36663 18199 36669
rect 13648 36632 13676 36660
rect 12912 36604 13676 36632
rect 15488 36632 15516 36663
rect 15562 36632 15568 36644
rect 15488 36604 15568 36632
rect 15562 36592 15568 36604
rect 15620 36592 15626 36644
rect 14550 36564 14556 36576
rect 9968 36536 14556 36564
rect 14550 36524 14556 36536
rect 14608 36524 14614 36576
rect 14737 36567 14795 36573
rect 14737 36533 14749 36567
rect 14783 36564 14795 36567
rect 16482 36564 16488 36576
rect 14783 36536 16488 36564
rect 14783 36533 14795 36536
rect 14737 36527 14795 36533
rect 16482 36524 16488 36536
rect 16540 36524 16546 36576
rect 16684 36564 16712 36663
rect 18156 36576 18184 36663
rect 18506 36660 18512 36712
rect 18564 36700 18570 36712
rect 20438 36700 20444 36712
rect 18564 36672 20444 36700
rect 18564 36660 18570 36672
rect 20438 36660 20444 36672
rect 20496 36660 20502 36712
rect 18601 36635 18659 36641
rect 18601 36601 18613 36635
rect 18647 36632 18659 36635
rect 19794 36632 19800 36644
rect 18647 36604 19800 36632
rect 18647 36601 18659 36604
rect 18601 36595 18659 36601
rect 19794 36592 19800 36604
rect 19852 36592 19858 36644
rect 20640 36641 20668 36744
rect 20732 36700 20760 36808
rect 20806 36728 20812 36780
rect 20864 36728 20870 36780
rect 21284 36777 21312 36808
rect 21085 36771 21143 36777
rect 21085 36737 21097 36771
rect 21131 36737 21143 36771
rect 21085 36731 21143 36737
rect 21269 36771 21327 36777
rect 21269 36737 21281 36771
rect 21315 36737 21327 36771
rect 21269 36731 21327 36737
rect 21100 36700 21128 36731
rect 20732 36672 21128 36700
rect 20625 36635 20683 36641
rect 20625 36601 20637 36635
rect 20671 36601 20683 36635
rect 20625 36595 20683 36601
rect 17954 36564 17960 36576
rect 16684 36536 17960 36564
rect 17954 36524 17960 36536
rect 18012 36524 18018 36576
rect 18138 36524 18144 36576
rect 18196 36524 18202 36576
rect 19702 36524 19708 36576
rect 19760 36564 19766 36576
rect 19978 36564 19984 36576
rect 19760 36536 19984 36564
rect 19760 36524 19766 36536
rect 19978 36524 19984 36536
rect 20036 36524 20042 36576
rect 20441 36567 20499 36573
rect 20441 36533 20453 36567
rect 20487 36564 20499 36567
rect 20898 36564 20904 36576
rect 20487 36536 20904 36564
rect 20487 36533 20499 36536
rect 20441 36527 20499 36533
rect 20898 36524 20904 36536
rect 20956 36524 20962 36576
rect 21450 36524 21456 36576
rect 21508 36524 21514 36576
rect 1104 36474 21896 36496
rect 1104 36422 3549 36474
rect 3601 36422 3613 36474
rect 3665 36422 3677 36474
rect 3729 36422 3741 36474
rect 3793 36422 3805 36474
rect 3857 36422 8747 36474
rect 8799 36422 8811 36474
rect 8863 36422 8875 36474
rect 8927 36422 8939 36474
rect 8991 36422 9003 36474
rect 9055 36422 13945 36474
rect 13997 36422 14009 36474
rect 14061 36422 14073 36474
rect 14125 36422 14137 36474
rect 14189 36422 14201 36474
rect 14253 36422 19143 36474
rect 19195 36422 19207 36474
rect 19259 36422 19271 36474
rect 19323 36422 19335 36474
rect 19387 36422 19399 36474
rect 19451 36422 21896 36474
rect 1104 36400 21896 36422
rect 1210 36320 1216 36372
rect 1268 36360 1274 36372
rect 1578 36360 1584 36372
rect 1268 36332 1584 36360
rect 1268 36320 1274 36332
rect 1578 36320 1584 36332
rect 1636 36320 1642 36372
rect 3973 36363 4031 36369
rect 3973 36329 3985 36363
rect 4019 36360 4031 36363
rect 4798 36360 4804 36372
rect 4019 36332 4804 36360
rect 4019 36329 4031 36332
rect 3973 36323 4031 36329
rect 4798 36320 4804 36332
rect 4856 36320 4862 36372
rect 5626 36320 5632 36372
rect 5684 36320 5690 36372
rect 5810 36320 5816 36372
rect 5868 36320 5874 36372
rect 7101 36363 7159 36369
rect 7101 36329 7113 36363
rect 7147 36329 7159 36363
rect 7101 36323 7159 36329
rect 7208 36332 9674 36360
rect 5644 36292 5672 36320
rect 4080 36264 5672 36292
rect 2225 36227 2283 36233
rect 2225 36224 2237 36227
rect 1136 36196 2237 36224
rect 1136 36168 1164 36196
rect 2225 36193 2237 36196
rect 2271 36193 2283 36227
rect 2225 36187 2283 36193
rect 1118 36116 1124 36168
rect 1176 36116 1182 36168
rect 1394 36116 1400 36168
rect 1452 36116 1458 36168
rect 2499 36159 2557 36165
rect 2499 36125 2511 36159
rect 2545 36156 2557 36159
rect 2590 36156 2596 36168
rect 2545 36128 2596 36156
rect 2545 36125 2557 36128
rect 2499 36119 2557 36125
rect 2590 36116 2596 36128
rect 2648 36156 2654 36168
rect 4080 36156 4108 36264
rect 5442 36224 5448 36236
rect 4172 36196 5448 36224
rect 4172 36165 4200 36196
rect 5442 36184 5448 36196
rect 5500 36184 5506 36236
rect 5828 36210 5856 36320
rect 6914 36184 6920 36236
rect 6972 36224 6978 36236
rect 7116 36224 7144 36323
rect 7208 36236 7236 36332
rect 6972 36196 7144 36224
rect 6972 36184 6978 36196
rect 7190 36184 7196 36236
rect 7248 36184 7254 36236
rect 8956 36233 8984 36332
rect 9646 36292 9674 36332
rect 9766 36320 9772 36372
rect 9824 36360 9830 36372
rect 10962 36360 10968 36372
rect 9824 36332 10968 36360
rect 9824 36320 9830 36332
rect 10962 36320 10968 36332
rect 11020 36320 11026 36372
rect 13814 36320 13820 36372
rect 13872 36360 13878 36372
rect 14277 36363 14335 36369
rect 14277 36360 14289 36363
rect 13872 36332 14289 36360
rect 13872 36320 13878 36332
rect 14277 36329 14289 36332
rect 14323 36329 14335 36363
rect 14277 36323 14335 36329
rect 14734 36320 14740 36372
rect 14792 36360 14798 36372
rect 15010 36360 15016 36372
rect 14792 36332 15016 36360
rect 14792 36320 14798 36332
rect 15010 36320 15016 36332
rect 15068 36320 15074 36372
rect 15933 36363 15991 36369
rect 15933 36329 15945 36363
rect 15979 36360 15991 36363
rect 16390 36360 16396 36372
rect 15979 36332 16396 36360
rect 15979 36329 15991 36332
rect 15933 36323 15991 36329
rect 16390 36320 16396 36332
rect 16448 36320 16454 36372
rect 16574 36320 16580 36372
rect 16632 36320 16638 36372
rect 17865 36363 17923 36369
rect 16684 36332 17538 36360
rect 10042 36292 10048 36304
rect 9646 36264 10048 36292
rect 10042 36252 10048 36264
rect 10100 36252 10106 36304
rect 12250 36252 12256 36304
rect 12308 36252 12314 36304
rect 14550 36252 14556 36304
rect 14608 36292 14614 36304
rect 16684 36292 16712 36332
rect 14608 36264 16712 36292
rect 17510 36292 17538 36332
rect 17865 36329 17877 36363
rect 17911 36360 17923 36363
rect 18138 36360 18144 36372
rect 17911 36332 18144 36360
rect 17911 36329 17923 36332
rect 17865 36323 17923 36329
rect 18138 36320 18144 36332
rect 18196 36320 18202 36372
rect 19521 36363 19579 36369
rect 19521 36329 19533 36363
rect 19567 36360 19579 36363
rect 21174 36360 21180 36372
rect 19567 36332 21180 36360
rect 19567 36329 19579 36332
rect 19521 36323 19579 36329
rect 21174 36320 21180 36332
rect 21232 36320 21238 36372
rect 19702 36292 19708 36304
rect 17510 36264 19708 36292
rect 14608 36252 14614 36264
rect 19702 36252 19708 36264
rect 19760 36252 19766 36304
rect 19797 36295 19855 36301
rect 19797 36261 19809 36295
rect 19843 36261 19855 36295
rect 19797 36255 19855 36261
rect 8941 36227 8999 36233
rect 8941 36193 8953 36227
rect 8987 36193 8999 36227
rect 8941 36187 8999 36193
rect 9646 36196 11192 36224
rect 2648 36128 4108 36156
rect 4157 36159 4215 36165
rect 2648 36116 2654 36128
rect 4157 36125 4169 36159
rect 4203 36125 4215 36159
rect 4157 36119 4215 36125
rect 5092 36128 6040 36156
rect 1673 36091 1731 36097
rect 1673 36057 1685 36091
rect 1719 36088 1731 36091
rect 4062 36088 4068 36100
rect 1719 36060 4068 36088
rect 1719 36057 1731 36060
rect 1673 36051 1731 36057
rect 4062 36048 4068 36060
rect 4120 36048 4126 36100
rect 1578 35980 1584 36032
rect 1636 36020 1642 36032
rect 2222 36020 2228 36032
rect 1636 35992 2228 36020
rect 1636 35980 1642 35992
rect 2222 35980 2228 35992
rect 2280 35980 2286 36032
rect 2590 35980 2596 36032
rect 2648 36020 2654 36032
rect 3237 36023 3295 36029
rect 3237 36020 3249 36023
rect 2648 35992 3249 36020
rect 2648 35980 2654 35992
rect 3237 35989 3249 35992
rect 3283 35989 3295 36023
rect 3237 35983 3295 35989
rect 3326 35980 3332 36032
rect 3384 36020 3390 36032
rect 5092 36020 5120 36128
rect 6012 36088 6040 36128
rect 6086 36116 6092 36168
rect 6144 36116 6150 36168
rect 6181 36159 6239 36165
rect 6181 36125 6193 36159
rect 6227 36156 6239 36159
rect 7282 36156 7288 36168
rect 6227 36128 7288 36156
rect 6227 36125 6239 36128
rect 6181 36119 6239 36125
rect 7282 36116 7288 36128
rect 7340 36116 7346 36168
rect 7469 36159 7527 36165
rect 7469 36125 7481 36159
rect 7515 36156 7527 36159
rect 7650 36156 7656 36168
rect 7515 36128 7656 36156
rect 7515 36125 7527 36128
rect 7469 36119 7527 36125
rect 6549 36091 6607 36097
rect 6549 36088 6561 36091
rect 6012 36060 6561 36088
rect 6549 36057 6561 36060
rect 6595 36057 6607 36091
rect 7484 36088 7512 36119
rect 7650 36116 7656 36128
rect 7708 36116 7714 36168
rect 7742 36116 7748 36168
rect 7800 36156 7806 36168
rect 9183 36159 9241 36165
rect 9183 36156 9195 36159
rect 7800 36128 7843 36156
rect 8036 36128 9195 36156
rect 7800 36116 7806 36128
rect 8036 36100 8064 36128
rect 9183 36125 9195 36128
rect 9229 36156 9241 36159
rect 9646 36156 9674 36196
rect 9229 36128 9674 36156
rect 10505 36159 10563 36165
rect 9229 36125 9241 36128
rect 9183 36119 9241 36125
rect 10505 36125 10517 36159
rect 10551 36156 10563 36159
rect 10594 36156 10600 36168
rect 10551 36128 10600 36156
rect 10551 36125 10563 36128
rect 10505 36119 10563 36125
rect 10594 36116 10600 36128
rect 10652 36116 10658 36168
rect 6549 36051 6607 36057
rect 6840 36060 7512 36088
rect 5261 36023 5319 36029
rect 5261 36020 5273 36023
rect 3384 35992 5273 36020
rect 3384 35980 3390 35992
rect 5261 35989 5273 35992
rect 5307 35989 5319 36023
rect 5261 35983 5319 35989
rect 5718 35980 5724 36032
rect 5776 36020 5782 36032
rect 5813 36023 5871 36029
rect 5813 36020 5825 36023
rect 5776 35992 5825 36020
rect 5776 35980 5782 35992
rect 5813 35989 5825 35992
rect 5859 35989 5871 36023
rect 5813 35983 5871 35989
rect 6178 35980 6184 36032
rect 6236 36020 6242 36032
rect 6840 36020 6868 36060
rect 8018 36048 8024 36100
rect 8076 36048 8082 36100
rect 8294 36048 8300 36100
rect 8352 36088 8358 36100
rect 8352 36060 10088 36088
rect 8352 36048 8358 36060
rect 6236 35992 6868 36020
rect 6236 35980 6242 35992
rect 6914 35980 6920 36032
rect 6972 36020 6978 36032
rect 7834 36020 7840 36032
rect 6972 35992 7840 36020
rect 6972 35980 6978 35992
rect 7834 35980 7840 35992
rect 7892 35980 7898 36032
rect 8481 36023 8539 36029
rect 8481 35989 8493 36023
rect 8527 36020 8539 36023
rect 8754 36020 8760 36032
rect 8527 35992 8760 36020
rect 8527 35989 8539 35992
rect 8481 35983 8539 35989
rect 8754 35980 8760 35992
rect 8812 35980 8818 36032
rect 9122 35980 9128 36032
rect 9180 36020 9186 36032
rect 9306 36020 9312 36032
rect 9180 35992 9312 36020
rect 9180 35980 9186 35992
rect 9306 35980 9312 35992
rect 9364 35980 9370 36032
rect 9766 35980 9772 36032
rect 9824 36020 9830 36032
rect 9953 36023 10011 36029
rect 9953 36020 9965 36023
rect 9824 35992 9965 36020
rect 9824 35980 9830 35992
rect 9953 35989 9965 35992
rect 9999 35989 10011 36023
rect 10060 36020 10088 36060
rect 10597 36023 10655 36029
rect 10597 36020 10609 36023
rect 10060 35992 10609 36020
rect 9953 35983 10011 35989
rect 10597 35989 10609 35992
rect 10643 35989 10655 36023
rect 11164 36020 11192 36196
rect 12084 36196 13952 36224
rect 11241 36159 11299 36165
rect 11241 36125 11253 36159
rect 11287 36125 11299 36159
rect 11241 36119 11299 36125
rect 11256 36088 11284 36119
rect 11422 36116 11428 36168
rect 11480 36156 11486 36168
rect 11515 36159 11573 36165
rect 11515 36156 11527 36159
rect 11480 36128 11527 36156
rect 11480 36116 11486 36128
rect 11515 36125 11527 36128
rect 11561 36156 11573 36159
rect 12084 36156 12112 36196
rect 11561 36128 12112 36156
rect 11561 36125 11573 36128
rect 11515 36119 11573 36125
rect 12158 36116 12164 36168
rect 12216 36116 12222 36168
rect 12176 36088 12204 36116
rect 11256 36060 12204 36088
rect 13814 36020 13820 36032
rect 11164 35992 13820 36020
rect 10597 35983 10655 35989
rect 13814 35980 13820 35992
rect 13872 35980 13878 36032
rect 13924 36020 13952 36196
rect 16022 36184 16028 36236
rect 16080 36224 16086 36236
rect 16206 36224 16212 36236
rect 16080 36196 16212 36224
rect 16080 36184 16086 36196
rect 16206 36184 16212 36196
rect 16264 36224 16270 36236
rect 16853 36227 16911 36233
rect 16853 36224 16865 36227
rect 16264 36196 16865 36224
rect 16264 36184 16270 36196
rect 16853 36193 16865 36196
rect 16899 36193 16911 36227
rect 16853 36187 16911 36193
rect 18046 36184 18052 36236
rect 18104 36224 18110 36236
rect 19334 36224 19340 36236
rect 18104 36196 19340 36224
rect 18104 36184 18110 36196
rect 19334 36184 19340 36196
rect 19392 36184 19398 36236
rect 19812 36224 19840 36255
rect 19886 36252 19892 36304
rect 19944 36292 19950 36304
rect 20990 36292 20996 36304
rect 19944 36264 20996 36292
rect 19944 36252 19950 36264
rect 20990 36252 20996 36264
rect 21048 36252 21054 36304
rect 19812 36196 20300 36224
rect 16117 36159 16175 36165
rect 16117 36156 16129 36159
rect 14752 36128 16129 36156
rect 14752 36100 14780 36128
rect 16117 36125 16129 36128
rect 16163 36125 16175 36159
rect 16117 36119 16175 36125
rect 16482 36116 16488 36168
rect 16540 36156 16546 36168
rect 16761 36159 16819 36165
rect 16761 36156 16773 36159
rect 16540 36128 16773 36156
rect 16540 36116 16546 36128
rect 16761 36125 16773 36128
rect 16807 36125 16819 36159
rect 16761 36119 16819 36125
rect 17127 36159 17185 36165
rect 17127 36125 17139 36159
rect 17173 36156 17185 36159
rect 18322 36156 18328 36168
rect 17173 36128 18328 36156
rect 17173 36125 17185 36128
rect 17127 36119 17185 36125
rect 18322 36116 18328 36128
rect 18380 36116 18386 36168
rect 18966 36116 18972 36168
rect 19024 36156 19030 36168
rect 19429 36159 19487 36165
rect 19429 36156 19441 36159
rect 19024 36128 19441 36156
rect 19024 36116 19030 36128
rect 19429 36125 19441 36128
rect 19475 36125 19487 36159
rect 19429 36119 19487 36125
rect 19702 36116 19708 36168
rect 19760 36116 19766 36168
rect 20272 36165 20300 36196
rect 20249 36159 20307 36165
rect 19981 36135 20039 36141
rect 19705 36115 19763 36116
rect 19981 36101 19993 36135
rect 20027 36101 20039 36135
rect 20249 36125 20261 36159
rect 20295 36125 20307 36159
rect 20249 36119 20307 36125
rect 20438 36116 20444 36168
rect 20496 36156 20502 36168
rect 20625 36159 20683 36165
rect 20625 36156 20637 36159
rect 20496 36128 20637 36156
rect 20496 36116 20502 36128
rect 20625 36125 20637 36128
rect 20671 36125 20683 36159
rect 20625 36119 20683 36125
rect 20993 36159 21051 36165
rect 20993 36125 21005 36159
rect 21039 36156 21051 36159
rect 21358 36156 21364 36168
rect 21039 36128 21364 36156
rect 21039 36125 21051 36128
rect 20993 36119 21051 36125
rect 21358 36116 21364 36128
rect 21416 36116 21422 36168
rect 14734 36048 14740 36100
rect 14792 36048 14798 36100
rect 18414 36048 18420 36100
rect 18472 36088 18478 36100
rect 19981 36095 20039 36101
rect 18472 36060 19656 36088
rect 18472 36048 18478 36060
rect 15838 36020 15844 36032
rect 13924 35992 15844 36020
rect 15838 35980 15844 35992
rect 15896 36020 15902 36032
rect 18506 36020 18512 36032
rect 15896 35992 18512 36020
rect 15896 35980 15902 35992
rect 18506 35980 18512 35992
rect 18564 35980 18570 36032
rect 19058 35980 19064 36032
rect 19116 36020 19122 36032
rect 19245 36023 19303 36029
rect 19245 36020 19257 36023
rect 19116 35992 19257 36020
rect 19116 35980 19122 35992
rect 19245 35989 19257 35992
rect 19291 35989 19303 36023
rect 19628 36020 19656 36060
rect 19996 36020 20024 36095
rect 21177 36091 21235 36097
rect 21177 36088 21189 36091
rect 20364 36060 21189 36088
rect 19628 35992 20024 36020
rect 20073 36023 20131 36029
rect 19245 35983 19303 35989
rect 20073 35989 20085 36023
rect 20119 36020 20131 36023
rect 20364 36020 20392 36060
rect 21177 36057 21189 36060
rect 21223 36057 21235 36091
rect 21177 36051 21235 36057
rect 21545 36091 21603 36097
rect 21545 36057 21557 36091
rect 21591 36088 21603 36091
rect 22278 36088 22284 36100
rect 21591 36060 22284 36088
rect 21591 36057 21603 36060
rect 21545 36051 21603 36057
rect 22278 36048 22284 36060
rect 22336 36048 22342 36100
rect 20119 35992 20392 36020
rect 20119 35989 20131 35992
rect 20073 35983 20131 35989
rect 20438 35980 20444 36032
rect 20496 35980 20502 36032
rect 20806 35980 20812 36032
rect 20864 35980 20870 36032
rect 1104 35930 22056 35952
rect 1104 35878 6148 35930
rect 6200 35878 6212 35930
rect 6264 35878 6276 35930
rect 6328 35878 6340 35930
rect 6392 35878 6404 35930
rect 6456 35878 11346 35930
rect 11398 35878 11410 35930
rect 11462 35878 11474 35930
rect 11526 35878 11538 35930
rect 11590 35878 11602 35930
rect 11654 35878 16544 35930
rect 16596 35878 16608 35930
rect 16660 35878 16672 35930
rect 16724 35878 16736 35930
rect 16788 35878 16800 35930
rect 16852 35878 21742 35930
rect 21794 35878 21806 35930
rect 21858 35878 21870 35930
rect 21922 35878 21934 35930
rect 21986 35878 21998 35930
rect 22050 35878 22056 35930
rect 1104 35856 22056 35878
rect 2866 35816 2872 35828
rect 1964 35788 2872 35816
rect 1964 35689 1992 35788
rect 2866 35776 2872 35788
rect 2924 35776 2930 35828
rect 4614 35776 4620 35828
rect 4672 35816 4678 35828
rect 4672 35788 5396 35816
rect 4672 35776 4678 35788
rect 3510 35708 3516 35760
rect 3568 35748 3574 35760
rect 5368 35748 5396 35788
rect 5810 35776 5816 35828
rect 5868 35816 5874 35828
rect 5905 35819 5963 35825
rect 5905 35816 5917 35819
rect 5868 35788 5917 35816
rect 5868 35776 5874 35788
rect 5905 35785 5917 35788
rect 5951 35785 5963 35819
rect 13078 35816 13084 35828
rect 5905 35779 5963 35785
rect 7760 35788 13084 35816
rect 7558 35748 7564 35760
rect 3568 35720 5304 35748
rect 5368 35720 7564 35748
rect 3568 35708 3574 35720
rect 1673 35683 1731 35689
rect 1673 35649 1685 35683
rect 1719 35680 1731 35683
rect 1949 35683 2007 35689
rect 1719 35652 1900 35680
rect 1719 35649 1731 35652
rect 1673 35643 1731 35649
rect 1762 35572 1768 35624
rect 1820 35572 1826 35624
rect 1872 35612 1900 35652
rect 1949 35649 1961 35683
rect 1995 35649 2007 35683
rect 1949 35643 2007 35649
rect 2958 35640 2964 35692
rect 3016 35640 3022 35692
rect 3789 35683 3847 35689
rect 3789 35649 3801 35683
rect 3835 35649 3847 35683
rect 3789 35643 3847 35649
rect 2130 35612 2136 35624
rect 1872 35584 2136 35612
rect 2130 35572 2136 35584
rect 2188 35572 2194 35624
rect 2406 35572 2412 35624
rect 2464 35572 2470 35624
rect 2685 35615 2743 35621
rect 2685 35612 2697 35615
rect 2516 35584 2697 35612
rect 2222 35504 2228 35556
rect 2280 35544 2286 35556
rect 2516 35544 2544 35584
rect 2685 35581 2697 35584
rect 2731 35581 2743 35615
rect 2685 35575 2743 35581
rect 2774 35572 2780 35624
rect 2832 35621 2838 35624
rect 2832 35615 2860 35621
rect 2848 35581 2860 35615
rect 2832 35575 2860 35581
rect 2832 35572 2838 35575
rect 3142 35572 3148 35624
rect 3200 35612 3206 35624
rect 3804 35612 3832 35643
rect 4246 35640 4252 35692
rect 4304 35640 4310 35692
rect 4338 35640 4344 35692
rect 4396 35680 4402 35692
rect 5135 35683 5193 35689
rect 5135 35680 5147 35683
rect 4396 35652 5147 35680
rect 4396 35640 4402 35652
rect 5135 35649 5147 35652
rect 5181 35649 5193 35683
rect 5276 35680 5304 35720
rect 7558 35708 7564 35720
rect 7616 35708 7622 35760
rect 7760 35692 7788 35788
rect 13078 35776 13084 35788
rect 13136 35776 13142 35828
rect 14550 35776 14556 35828
rect 14608 35816 14614 35828
rect 14608 35788 19104 35816
rect 14608 35776 14614 35788
rect 8570 35708 8576 35760
rect 8628 35708 8634 35760
rect 18966 35757 18972 35760
rect 18938 35751 18972 35757
rect 18938 35748 18950 35751
rect 13372 35720 17908 35748
rect 12051 35713 12109 35719
rect 12051 35710 12063 35713
rect 6365 35683 6423 35689
rect 6365 35680 6377 35683
rect 5276 35652 6377 35680
rect 5135 35643 5193 35649
rect 6365 35649 6377 35652
rect 6411 35649 6423 35683
rect 6365 35643 6423 35649
rect 6641 35683 6699 35689
rect 6641 35649 6653 35683
rect 6687 35680 6699 35683
rect 7283 35683 7341 35689
rect 7283 35680 7295 35683
rect 6687 35652 7295 35680
rect 6687 35649 6699 35652
rect 6641 35643 6699 35649
rect 7283 35649 7295 35652
rect 7329 35680 7341 35683
rect 7742 35680 7748 35692
rect 7329 35652 7748 35680
rect 7329 35649 7341 35652
rect 7283 35643 7341 35649
rect 7742 35640 7748 35652
rect 7800 35640 7806 35692
rect 8389 35683 8447 35689
rect 8389 35649 8401 35683
rect 8435 35680 8447 35683
rect 8588 35680 8616 35708
rect 8435 35652 8616 35680
rect 8435 35649 8447 35652
rect 8389 35643 8447 35649
rect 9306 35640 9312 35692
rect 9364 35640 9370 35692
rect 11698 35640 11704 35692
rect 11756 35680 11762 35692
rect 12050 35680 12063 35710
rect 11756 35679 12063 35680
rect 12097 35680 12109 35713
rect 13372 35680 13400 35720
rect 12097 35679 13400 35680
rect 11756 35652 13400 35679
rect 11756 35640 11762 35652
rect 13446 35640 13452 35692
rect 13504 35680 13510 35692
rect 13504 35652 14872 35680
rect 13504 35640 13510 35652
rect 4354 35612 4382 35640
rect 3200 35584 3832 35612
rect 4080 35584 4382 35612
rect 3200 35572 3206 35584
rect 2280 35516 2544 35544
rect 2280 35504 2286 35516
rect 1302 35436 1308 35488
rect 1360 35476 1366 35488
rect 3605 35479 3663 35485
rect 3605 35476 3617 35479
rect 1360 35448 3617 35476
rect 1360 35436 1366 35448
rect 3605 35445 3617 35448
rect 3651 35445 3663 35479
rect 3605 35439 3663 35445
rect 3970 35436 3976 35488
rect 4028 35476 4034 35488
rect 4080 35485 4108 35584
rect 4522 35572 4528 35624
rect 4580 35572 4586 35624
rect 4890 35572 4896 35624
rect 4948 35572 4954 35624
rect 6822 35612 6828 35624
rect 5736 35584 6828 35612
rect 5736 35556 5764 35584
rect 6822 35572 6828 35584
rect 6880 35572 6886 35624
rect 7009 35615 7067 35621
rect 7009 35581 7021 35615
rect 7055 35581 7067 35615
rect 7009 35575 7067 35581
rect 5718 35504 5724 35556
rect 5776 35504 5782 35556
rect 6638 35504 6644 35556
rect 6696 35544 6702 35556
rect 7024 35544 7052 35575
rect 8570 35572 8576 35624
rect 8628 35572 8634 35624
rect 8754 35572 8760 35624
rect 8812 35612 8818 35624
rect 9033 35615 9091 35621
rect 9033 35612 9045 35615
rect 8812 35584 9045 35612
rect 8812 35572 8818 35584
rect 9033 35581 9045 35584
rect 9079 35581 9091 35615
rect 9033 35575 9091 35581
rect 9423 35572 9429 35624
rect 9481 35572 9487 35624
rect 9582 35572 9588 35624
rect 9640 35572 9646 35624
rect 10962 35572 10968 35624
rect 11020 35612 11026 35624
rect 11146 35612 11152 35624
rect 11020 35584 11152 35612
rect 11020 35572 11026 35584
rect 11146 35572 11152 35584
rect 11204 35572 11210 35624
rect 11793 35615 11851 35621
rect 11793 35581 11805 35615
rect 11839 35581 11851 35615
rect 14844 35612 14872 35652
rect 15194 35640 15200 35692
rect 15252 35680 15258 35692
rect 15473 35683 15531 35689
rect 15473 35680 15485 35683
rect 15252 35652 15485 35680
rect 15252 35640 15258 35652
rect 15473 35649 15485 35652
rect 15519 35649 15531 35683
rect 15473 35643 15531 35649
rect 16022 35640 16028 35692
rect 16080 35680 16086 35692
rect 16853 35683 16911 35689
rect 16853 35680 16865 35683
rect 16080 35652 16865 35680
rect 16080 35640 16086 35652
rect 16853 35649 16865 35652
rect 16899 35649 16911 35683
rect 17221 35683 17279 35689
rect 16853 35643 16911 35649
rect 16960 35652 17172 35680
rect 16960 35612 16988 35652
rect 14844 35584 16988 35612
rect 11793 35575 11851 35581
rect 6696 35516 7052 35544
rect 7668 35516 8156 35544
rect 6696 35504 6702 35516
rect 4065 35479 4123 35485
rect 4065 35476 4077 35479
rect 4028 35448 4077 35476
rect 4028 35436 4034 35448
rect 4065 35445 4077 35448
rect 4111 35445 4123 35479
rect 4065 35439 4123 35445
rect 4890 35436 4896 35488
rect 4948 35476 4954 35488
rect 7668 35476 7696 35516
rect 4948 35448 7696 35476
rect 4948 35436 4954 35448
rect 8018 35436 8024 35488
rect 8076 35436 8082 35488
rect 8128 35476 8156 35516
rect 10229 35479 10287 35485
rect 10229 35476 10241 35479
rect 8128 35448 10241 35476
rect 10229 35445 10241 35448
rect 10275 35445 10287 35479
rect 11808 35476 11836 35575
rect 17034 35572 17040 35624
rect 17092 35572 17098 35624
rect 17144 35612 17172 35652
rect 17221 35649 17233 35683
rect 17267 35680 17279 35683
rect 17267 35652 17816 35680
rect 17267 35649 17279 35652
rect 17221 35643 17279 35649
rect 17144 35584 17724 35612
rect 12526 35504 12532 35556
rect 12584 35544 12590 35556
rect 13357 35547 13415 35553
rect 13357 35544 13369 35547
rect 12584 35516 13369 35544
rect 12584 35504 12590 35516
rect 13357 35513 13369 35516
rect 13403 35513 13415 35547
rect 13357 35507 13415 35513
rect 14274 35504 14280 35556
rect 14332 35544 14338 35556
rect 17494 35544 17500 35556
rect 14332 35516 17500 35544
rect 14332 35504 14338 35516
rect 17494 35504 17500 35516
rect 17552 35504 17558 35556
rect 12158 35476 12164 35488
rect 11808 35448 12164 35476
rect 10229 35439 10287 35445
rect 12158 35436 12164 35448
rect 12216 35436 12222 35488
rect 12802 35436 12808 35488
rect 12860 35436 12866 35488
rect 15286 35436 15292 35488
rect 15344 35436 15350 35488
rect 17129 35479 17187 35485
rect 17129 35445 17141 35479
rect 17175 35476 17187 35479
rect 17586 35476 17592 35488
rect 17175 35448 17592 35476
rect 17175 35445 17187 35448
rect 17129 35439 17187 35445
rect 17586 35436 17592 35448
rect 17644 35436 17650 35488
rect 17696 35476 17724 35584
rect 17788 35556 17816 35652
rect 17770 35504 17776 35556
rect 17828 35504 17834 35556
rect 17880 35544 17908 35720
rect 18248 35720 18950 35748
rect 18248 35692 18276 35720
rect 18938 35717 18950 35720
rect 18938 35711 18972 35717
rect 18966 35708 18972 35711
rect 19024 35708 19030 35760
rect 19076 35748 19104 35788
rect 19702 35776 19708 35828
rect 19760 35816 19766 35828
rect 20165 35819 20223 35825
rect 20165 35816 20177 35819
rect 19760 35788 20177 35816
rect 19760 35776 19766 35788
rect 20165 35785 20177 35788
rect 20211 35785 20223 35819
rect 20165 35779 20223 35785
rect 20533 35819 20591 35825
rect 20533 35785 20545 35819
rect 20579 35816 20591 35819
rect 21266 35816 21272 35828
rect 20579 35788 21272 35816
rect 20579 35785 20591 35788
rect 20533 35779 20591 35785
rect 21266 35776 21272 35788
rect 21324 35776 21330 35828
rect 19076 35720 22968 35748
rect 17954 35640 17960 35692
rect 18012 35640 18018 35692
rect 18230 35640 18236 35692
rect 18288 35640 18294 35692
rect 18322 35640 18328 35692
rect 18380 35680 18386 35692
rect 18506 35680 18512 35692
rect 18380 35652 18512 35680
rect 18380 35640 18386 35652
rect 18506 35640 18512 35652
rect 18564 35680 18570 35692
rect 18601 35683 18659 35689
rect 18601 35680 18613 35683
rect 18564 35652 18613 35680
rect 18564 35640 18570 35652
rect 18601 35649 18613 35652
rect 18647 35649 18659 35683
rect 18601 35643 18659 35649
rect 19518 35640 19524 35692
rect 19576 35680 19582 35692
rect 20349 35683 20407 35689
rect 20349 35680 20361 35683
rect 19576 35652 20361 35680
rect 19576 35640 19582 35652
rect 20349 35649 20361 35652
rect 20395 35649 20407 35683
rect 20349 35643 20407 35649
rect 20438 35640 20444 35692
rect 20496 35680 20502 35692
rect 20717 35683 20775 35689
rect 20717 35680 20729 35683
rect 20496 35652 20729 35680
rect 20496 35640 20502 35652
rect 20717 35649 20729 35652
rect 20763 35649 20775 35683
rect 20717 35643 20775 35649
rect 20990 35640 20996 35692
rect 21048 35640 21054 35692
rect 21082 35640 21088 35692
rect 21140 35680 21146 35692
rect 21269 35683 21327 35689
rect 21269 35680 21281 35683
rect 21140 35652 21281 35680
rect 21140 35640 21146 35652
rect 21269 35649 21281 35652
rect 21315 35649 21327 35683
rect 21269 35643 21327 35649
rect 17972 35612 18000 35640
rect 22940 35624 22968 35720
rect 18693 35615 18751 35621
rect 18693 35612 18705 35615
rect 17972 35584 18705 35612
rect 18693 35581 18705 35584
rect 18739 35581 18751 35615
rect 22830 35612 22836 35624
rect 18693 35575 18751 35581
rect 19720 35584 22836 35612
rect 17954 35544 17960 35556
rect 17880 35516 17960 35544
rect 17954 35504 17960 35516
rect 18012 35504 18018 35556
rect 18414 35504 18420 35556
rect 18472 35504 18478 35556
rect 19720 35476 19748 35584
rect 22830 35572 22836 35584
rect 22888 35572 22894 35624
rect 22922 35572 22928 35624
rect 22980 35572 22986 35624
rect 20073 35547 20131 35553
rect 20073 35513 20085 35547
rect 20119 35544 20131 35547
rect 20714 35544 20720 35556
rect 20119 35516 20720 35544
rect 20119 35513 20131 35516
rect 20073 35507 20131 35513
rect 20714 35504 20720 35516
rect 20772 35504 20778 35556
rect 17696 35448 19748 35476
rect 20809 35479 20867 35485
rect 20809 35445 20821 35479
rect 20855 35476 20867 35479
rect 20990 35476 20996 35488
rect 20855 35448 20996 35476
rect 20855 35445 20867 35448
rect 20809 35439 20867 35445
rect 20990 35436 20996 35448
rect 21048 35436 21054 35488
rect 21450 35436 21456 35488
rect 21508 35436 21514 35488
rect 1104 35386 21896 35408
rect 1104 35334 3549 35386
rect 3601 35334 3613 35386
rect 3665 35334 3677 35386
rect 3729 35334 3741 35386
rect 3793 35334 3805 35386
rect 3857 35334 8747 35386
rect 8799 35334 8811 35386
rect 8863 35334 8875 35386
rect 8927 35334 8939 35386
rect 8991 35334 9003 35386
rect 9055 35334 13945 35386
rect 13997 35334 14009 35386
rect 14061 35334 14073 35386
rect 14125 35334 14137 35386
rect 14189 35334 14201 35386
rect 14253 35334 19143 35386
rect 19195 35334 19207 35386
rect 19259 35334 19271 35386
rect 19323 35334 19335 35386
rect 19387 35334 19399 35386
rect 19451 35334 21896 35386
rect 1104 35312 21896 35334
rect 3510 35232 3516 35284
rect 3568 35272 3574 35284
rect 4154 35272 4160 35284
rect 3568 35244 4160 35272
rect 3568 35232 3574 35244
rect 4154 35232 4160 35244
rect 4212 35272 4218 35284
rect 4212 35244 4384 35272
rect 4212 35232 4218 35244
rect 4356 35216 4384 35244
rect 4798 35232 4804 35284
rect 4856 35272 4862 35284
rect 5350 35272 5356 35284
rect 4856 35244 5356 35272
rect 4856 35232 4862 35244
rect 5350 35232 5356 35244
rect 5408 35232 5414 35284
rect 5810 35232 5816 35284
rect 5868 35272 5874 35284
rect 6638 35272 6644 35284
rect 5868 35244 6644 35272
rect 5868 35232 5874 35244
rect 1762 35164 1768 35216
rect 1820 35204 1826 35216
rect 1820 35176 1882 35204
rect 1820 35164 1826 35176
rect 1397 35071 1455 35077
rect 1397 35037 1409 35071
rect 1443 35068 1455 35071
rect 1762 35068 1768 35080
rect 1443 35040 1768 35068
rect 1443 35037 1455 35040
rect 1397 35031 1455 35037
rect 1762 35028 1768 35040
rect 1820 35028 1826 35080
rect 1670 34960 1676 35012
rect 1728 34960 1734 35012
rect 1854 35000 1882 35176
rect 4338 35164 4344 35216
rect 4396 35204 4402 35216
rect 4396 35176 4936 35204
rect 4396 35164 4402 35176
rect 2682 35096 2688 35148
rect 2740 35096 2746 35148
rect 4522 35096 4528 35148
rect 4580 35136 4586 35148
rect 4908 35145 4936 35176
rect 6288 35145 6316 35244
rect 6638 35232 6644 35244
rect 6696 35272 6702 35284
rect 7190 35272 7196 35284
rect 6696 35244 7196 35272
rect 6696 35232 6702 35244
rect 7190 35232 7196 35244
rect 7248 35232 7254 35284
rect 7282 35232 7288 35284
rect 7340 35232 7346 35284
rect 11790 35232 11796 35284
rect 11848 35272 11854 35284
rect 14550 35272 14556 35284
rect 11848 35244 14556 35272
rect 11848 35232 11854 35244
rect 14550 35232 14556 35244
rect 14608 35232 14614 35284
rect 15102 35272 15108 35284
rect 14844 35244 15108 35272
rect 7006 35164 7012 35216
rect 7064 35204 7070 35216
rect 8294 35204 8300 35216
rect 7064 35176 8300 35204
rect 7064 35164 7070 35176
rect 8294 35164 8300 35176
rect 8352 35164 8358 35216
rect 12250 35164 12256 35216
rect 12308 35164 12314 35216
rect 4893 35139 4951 35145
rect 4580 35108 4844 35136
rect 4580 35096 4586 35108
rect 2130 35028 2136 35080
rect 2188 35068 2194 35080
rect 2501 35071 2559 35077
rect 2501 35068 2513 35071
rect 2188 35040 2513 35068
rect 2188 35028 2194 35040
rect 2501 35037 2513 35040
rect 2547 35037 2559 35071
rect 2501 35031 2559 35037
rect 2590 35028 2596 35080
rect 2648 35028 2654 35080
rect 4249 35071 4307 35077
rect 4249 35037 4261 35071
rect 4295 35068 4307 35071
rect 4816 35068 4844 35108
rect 4893 35105 4905 35139
rect 4939 35105 4951 35139
rect 4893 35099 4951 35105
rect 6273 35139 6331 35145
rect 6273 35105 6285 35139
rect 6319 35105 6331 35139
rect 6273 35099 6331 35105
rect 8018 35096 8024 35148
rect 8076 35136 8082 35148
rect 8076 35108 8970 35136
rect 8076 35096 8082 35108
rect 12526 35096 12532 35148
rect 12584 35096 12590 35148
rect 12802 35096 12808 35148
rect 12860 35096 12866 35148
rect 14844 35145 14872 35244
rect 15102 35232 15108 35244
rect 15160 35232 15166 35284
rect 17034 35232 17040 35284
rect 17092 35272 17098 35284
rect 17313 35275 17371 35281
rect 17313 35272 17325 35275
rect 17092 35244 17325 35272
rect 17092 35232 17098 35244
rect 17313 35241 17325 35244
rect 17359 35241 17371 35275
rect 17313 35235 17371 35241
rect 14829 35139 14887 35145
rect 14829 35105 14841 35139
rect 14875 35105 14887 35139
rect 14829 35099 14887 35105
rect 16206 35096 16212 35148
rect 16264 35136 16270 35148
rect 16301 35139 16359 35145
rect 16301 35136 16313 35139
rect 16264 35108 16313 35136
rect 16264 35096 16270 35108
rect 16301 35105 16313 35108
rect 16347 35105 16359 35139
rect 16301 35099 16359 35105
rect 5135 35071 5193 35077
rect 5135 35068 5147 35071
rect 4295 35040 4777 35068
rect 4816 35040 5147 35068
rect 4295 35037 4307 35040
rect 4249 35031 4307 35037
rect 2961 35003 3019 35009
rect 2961 35000 2973 35003
rect 1854 34972 2973 35000
rect 2961 34969 2973 34972
rect 3007 35000 3019 35003
rect 3602 35000 3608 35012
rect 3007 34972 3608 35000
rect 3007 34969 3019 34972
rect 2961 34963 3019 34969
rect 3602 34960 3608 34972
rect 3660 34960 3666 35012
rect 3878 34960 3884 35012
rect 3936 34960 3942 35012
rect 4062 34960 4068 35012
rect 4120 35000 4126 35012
rect 4433 35003 4491 35009
rect 4433 35000 4445 35003
rect 4120 34972 4445 35000
rect 4120 34960 4126 34972
rect 4433 34969 4445 34972
rect 4479 34969 4491 35003
rect 4433 34963 4491 34969
rect 1302 34892 1308 34944
rect 1360 34932 1366 34944
rect 1854 34932 1860 34944
rect 1360 34904 1860 34932
rect 1360 34892 1366 34904
rect 1854 34892 1860 34904
rect 1912 34892 1918 34944
rect 2225 34935 2283 34941
rect 2225 34901 2237 34935
rect 2271 34932 2283 34935
rect 2314 34932 2320 34944
rect 2271 34904 2320 34932
rect 2271 34901 2283 34904
rect 2225 34895 2283 34901
rect 2314 34892 2320 34904
rect 2372 34892 2378 34944
rect 2866 34892 2872 34944
rect 2924 34932 2930 34944
rect 3050 34932 3056 34944
rect 2924 34904 3056 34932
rect 2924 34892 2930 34904
rect 3050 34892 3056 34904
rect 3108 34932 3114 34944
rect 3329 34935 3387 34941
rect 3329 34932 3341 34935
rect 3108 34904 3341 34932
rect 3108 34892 3114 34904
rect 3329 34901 3341 34904
rect 3375 34901 3387 34935
rect 3329 34895 3387 34901
rect 3510 34892 3516 34944
rect 3568 34892 3574 34944
rect 4522 34892 4528 34944
rect 4580 34892 4586 34944
rect 4749 34932 4777 35040
rect 5135 35037 5147 35040
rect 5181 35068 5193 35071
rect 6531 35071 6589 35077
rect 6531 35068 6543 35071
rect 5181 35040 6543 35068
rect 5181 35037 5193 35040
rect 5135 35031 5193 35037
rect 6531 35037 6543 35040
rect 6577 35068 6589 35071
rect 7282 35068 7288 35080
rect 6577 35040 7288 35068
rect 6577 35037 6589 35040
rect 6531 35031 6589 35037
rect 7282 35028 7288 35040
rect 7340 35028 7346 35080
rect 8662 35028 8668 35080
rect 8720 35068 8726 35080
rect 9401 35071 9459 35077
rect 9401 35068 9413 35071
rect 8720 35040 9413 35068
rect 8720 35028 8726 35040
rect 9401 35037 9413 35040
rect 9447 35037 9459 35071
rect 9401 35031 9459 35037
rect 9490 35028 9496 35080
rect 9548 35028 9554 35080
rect 10594 35068 10600 35080
rect 9784 35040 10600 35068
rect 6638 35000 6644 35012
rect 5736 34972 6644 35000
rect 5736 34932 5764 34972
rect 6638 34960 6644 34972
rect 6696 34960 6702 35012
rect 9125 35003 9183 35009
rect 9125 34969 9137 35003
rect 9171 35000 9183 35003
rect 9784 35000 9812 35040
rect 10594 35028 10600 35040
rect 10652 35068 10658 35080
rect 11057 35071 11115 35077
rect 11057 35068 11069 35071
rect 10652 35040 11069 35068
rect 10652 35028 10658 35040
rect 11057 35037 11069 35040
rect 11103 35037 11115 35071
rect 11057 35031 11115 35037
rect 11606 35028 11612 35080
rect 11664 35068 11670 35080
rect 11664 35040 11744 35068
rect 11664 35028 11670 35040
rect 9171 34972 9812 35000
rect 9171 34969 9183 34972
rect 9125 34963 9183 34969
rect 9858 34960 9864 35012
rect 9916 34960 9922 35012
rect 10226 34960 10232 35012
rect 10284 35000 10290 35012
rect 10781 35003 10839 35009
rect 10781 35000 10793 35003
rect 10284 34972 10793 35000
rect 10284 34960 10290 34972
rect 10781 34969 10793 34972
rect 10827 35000 10839 35003
rect 10870 35000 10876 35012
rect 10827 34972 10876 35000
rect 10827 34969 10839 34972
rect 10781 34963 10839 34969
rect 10870 34960 10876 34972
rect 10928 34960 10934 35012
rect 11238 34960 11244 35012
rect 11296 34960 11302 35012
rect 4749 34904 5764 34932
rect 5810 34892 5816 34944
rect 5868 34932 5874 34944
rect 5905 34935 5963 34941
rect 5905 34932 5917 34935
rect 5868 34904 5917 34932
rect 5868 34892 5874 34904
rect 5905 34901 5917 34904
rect 5951 34901 5963 34935
rect 5905 34895 5963 34901
rect 5994 34892 6000 34944
rect 6052 34932 6058 34944
rect 8018 34932 8024 34944
rect 6052 34904 8024 34932
rect 6052 34892 6058 34904
rect 8018 34892 8024 34904
rect 8076 34892 8082 34944
rect 9214 34892 9220 34944
rect 9272 34932 9278 34944
rect 9490 34932 9496 34944
rect 9272 34904 9496 34932
rect 9272 34892 9278 34904
rect 9490 34892 9496 34904
rect 9548 34892 9554 34944
rect 9950 34892 9956 34944
rect 10008 34932 10014 34944
rect 10413 34935 10471 34941
rect 10413 34932 10425 34935
rect 10008 34904 10425 34932
rect 10008 34892 10014 34904
rect 10413 34901 10425 34904
rect 10459 34932 10471 34935
rect 10502 34932 10508 34944
rect 10459 34904 10508 34932
rect 10459 34901 10471 34904
rect 10413 34895 10471 34901
rect 10502 34892 10508 34904
rect 10560 34892 10566 34944
rect 11716 34932 11744 35040
rect 11790 35028 11796 35080
rect 11848 35028 11854 35080
rect 12618 35028 12624 35080
rect 12676 35077 12682 35080
rect 12676 35071 12704 35077
rect 12692 35037 12704 35071
rect 12676 35031 12704 35037
rect 12676 35028 12682 35031
rect 13449 35003 13507 35009
rect 13449 34969 13461 35003
rect 13495 35000 13507 35003
rect 15074 35003 15132 35009
rect 15074 35000 15086 35003
rect 13495 34972 15086 35000
rect 13495 34969 13507 34972
rect 13449 34963 13507 34969
rect 15074 34969 15086 34972
rect 15120 35000 15132 35003
rect 15194 35000 15200 35012
rect 15120 34972 15200 35000
rect 15120 34969 15132 34972
rect 15074 34963 15132 34969
rect 15194 34960 15200 34972
rect 15252 34960 15258 35012
rect 12250 34932 12256 34944
rect 11716 34904 12256 34932
rect 12250 34892 12256 34904
rect 12308 34892 12314 34944
rect 16206 34892 16212 34944
rect 16264 34892 16270 34944
rect 16316 34932 16344 35099
rect 16575 35071 16633 35077
rect 16575 35037 16587 35071
rect 16621 35068 16633 35071
rect 16942 35068 16948 35080
rect 16621 35040 16948 35068
rect 16621 35037 16633 35040
rect 16575 35031 16633 35037
rect 16942 35028 16948 35040
rect 17000 35028 17006 35080
rect 17328 35068 17356 35235
rect 17494 35232 17500 35284
rect 17552 35232 17558 35284
rect 17770 35232 17776 35284
rect 17828 35232 17834 35284
rect 19702 35272 19708 35284
rect 19306 35244 19708 35272
rect 17512 35204 17540 35232
rect 19306 35204 19334 35244
rect 19702 35232 19708 35244
rect 19760 35232 19766 35284
rect 20257 35275 20315 35281
rect 20257 35241 20269 35275
rect 20303 35272 20315 35275
rect 20346 35272 20352 35284
rect 20303 35244 20352 35272
rect 20303 35241 20315 35244
rect 20257 35235 20315 35241
rect 20346 35232 20352 35244
rect 20404 35232 20410 35284
rect 21174 35232 21180 35284
rect 21232 35232 21238 35284
rect 17512 35176 19334 35204
rect 19245 35139 19303 35145
rect 19245 35136 19257 35139
rect 17972 35108 19257 35136
rect 17681 35071 17739 35077
rect 17681 35068 17693 35071
rect 17328 35040 17693 35068
rect 17681 35037 17693 35040
rect 17727 35037 17739 35071
rect 17681 35031 17739 35037
rect 17865 35071 17923 35077
rect 17865 35037 17877 35071
rect 17911 35037 17923 35071
rect 17865 35031 17923 35037
rect 16390 34960 16396 35012
rect 16448 35000 16454 35012
rect 17880 35000 17908 35031
rect 16448 34972 17908 35000
rect 16448 34960 16454 34972
rect 17034 34932 17040 34944
rect 16316 34904 17040 34932
rect 17034 34892 17040 34904
rect 17092 34932 17098 34944
rect 17972 34932 18000 35108
rect 19245 35105 19257 35108
rect 19291 35105 19303 35139
rect 20364 35136 20392 35232
rect 20625 35139 20683 35145
rect 20625 35136 20637 35139
rect 20364 35108 20637 35136
rect 19245 35099 19303 35105
rect 20625 35105 20637 35108
rect 20671 35105 20683 35139
rect 21192 35136 21220 35232
rect 21192 35108 21312 35136
rect 20625 35099 20683 35105
rect 18877 35071 18935 35077
rect 18877 35037 18889 35071
rect 18923 35068 18935 35071
rect 19058 35068 19064 35080
rect 18923 35040 19064 35068
rect 18923 35037 18935 35040
rect 18877 35031 18935 35037
rect 19058 35028 19064 35040
rect 19116 35028 19122 35080
rect 19487 35071 19545 35077
rect 19487 35037 19499 35071
rect 19533 35068 19545 35071
rect 20530 35068 20536 35080
rect 19533 35040 20536 35068
rect 19533 35037 19545 35040
rect 19487 35031 19545 35037
rect 20530 35028 20536 35040
rect 20588 35028 20594 35080
rect 20809 35071 20867 35077
rect 20809 35037 20821 35071
rect 20855 35037 20867 35071
rect 20809 35031 20867 35037
rect 18969 35003 19027 35009
rect 18969 34969 18981 35003
rect 19015 35000 19027 35003
rect 19015 34972 19748 35000
rect 19015 34969 19027 34972
rect 18969 34963 19027 34969
rect 17092 34904 18000 34932
rect 17092 34892 17098 34904
rect 18322 34892 18328 34944
rect 18380 34932 18386 34944
rect 19610 34932 19616 34944
rect 18380 34904 19616 34932
rect 18380 34892 18386 34904
rect 19610 34892 19616 34904
rect 19668 34892 19674 34944
rect 19720 34932 19748 34972
rect 20824 34932 20852 35031
rect 20898 35028 20904 35080
rect 20956 35068 20962 35080
rect 21284 35077 21312 35108
rect 21177 35071 21235 35077
rect 21177 35068 21189 35071
rect 20956 35040 21189 35068
rect 20956 35028 20962 35040
rect 21177 35037 21189 35040
rect 21223 35037 21235 35071
rect 21177 35031 21235 35037
rect 21269 35071 21327 35077
rect 21269 35037 21281 35071
rect 21315 35037 21327 35071
rect 21269 35031 21327 35037
rect 21085 35003 21143 35009
rect 21085 34969 21097 35003
rect 21131 35000 21143 35003
rect 22002 35000 22008 35012
rect 21131 34972 22008 35000
rect 21131 34969 21143 34972
rect 21085 34963 21143 34969
rect 22002 34960 22008 34972
rect 22060 34960 22066 35012
rect 19720 34904 20852 34932
rect 21453 34935 21511 34941
rect 21453 34901 21465 34935
rect 21499 34932 21511 34935
rect 22186 34932 22192 34944
rect 21499 34904 22192 34932
rect 21499 34901 21511 34904
rect 21453 34895 21511 34901
rect 22186 34892 22192 34904
rect 22244 34892 22250 34944
rect 1104 34842 22056 34864
rect 1104 34790 6148 34842
rect 6200 34790 6212 34842
rect 6264 34790 6276 34842
rect 6328 34790 6340 34842
rect 6392 34790 6404 34842
rect 6456 34790 11346 34842
rect 11398 34790 11410 34842
rect 11462 34790 11474 34842
rect 11526 34790 11538 34842
rect 11590 34790 11602 34842
rect 11654 34790 16544 34842
rect 16596 34790 16608 34842
rect 16660 34790 16672 34842
rect 16724 34790 16736 34842
rect 16788 34790 16800 34842
rect 16852 34790 21742 34842
rect 21794 34790 21806 34842
rect 21858 34790 21870 34842
rect 21922 34790 21934 34842
rect 21986 34790 21998 34842
rect 22050 34790 22056 34842
rect 1104 34768 22056 34790
rect 2130 34688 2136 34740
rect 2188 34728 2194 34740
rect 4890 34728 4896 34740
rect 2188 34700 4896 34728
rect 2188 34688 2194 34700
rect 4890 34688 4896 34700
rect 4948 34688 4954 34740
rect 5994 34688 6000 34740
rect 6052 34728 6058 34740
rect 6365 34731 6423 34737
rect 6365 34728 6377 34731
rect 6052 34700 6377 34728
rect 6052 34688 6058 34700
rect 6365 34697 6377 34700
rect 6411 34697 6423 34731
rect 6365 34691 6423 34697
rect 6454 34688 6460 34740
rect 6512 34728 6518 34740
rect 6822 34728 6828 34740
rect 6512 34700 6828 34728
rect 6512 34688 6518 34700
rect 6822 34688 6828 34700
rect 6880 34688 6886 34740
rect 7098 34688 7104 34740
rect 7156 34688 7162 34740
rect 9217 34731 9275 34737
rect 9217 34697 9229 34731
rect 9263 34728 9275 34731
rect 10410 34728 10416 34740
rect 9263 34700 10416 34728
rect 9263 34697 9275 34700
rect 9217 34691 9275 34697
rect 10410 34688 10416 34700
rect 10468 34728 10474 34740
rect 10468 34700 10824 34728
rect 10468 34688 10474 34700
rect 2314 34620 2320 34672
rect 2372 34660 2378 34672
rect 4522 34660 4528 34672
rect 2372 34632 4528 34660
rect 2372 34620 2378 34632
rect 4522 34620 4528 34632
rect 4580 34620 4586 34672
rect 4798 34620 4804 34672
rect 4856 34620 4862 34672
rect 5074 34620 5080 34672
rect 5132 34620 5138 34672
rect 5169 34663 5227 34669
rect 5169 34629 5181 34663
rect 5215 34660 5227 34663
rect 5810 34660 5816 34672
rect 5215 34632 5816 34660
rect 5215 34629 5227 34632
rect 5169 34623 5227 34629
rect 5810 34620 5816 34632
rect 5868 34620 5874 34672
rect 5905 34663 5963 34669
rect 5905 34629 5917 34663
rect 5951 34660 5963 34663
rect 6086 34660 6092 34672
rect 5951 34632 6092 34660
rect 5951 34629 5963 34632
rect 5905 34623 5963 34629
rect 6086 34620 6092 34632
rect 6144 34660 6150 34672
rect 7116 34660 7144 34688
rect 6144 34632 7144 34660
rect 6144 34620 6150 34632
rect 9398 34620 9404 34672
rect 9456 34660 9462 34672
rect 9493 34663 9551 34669
rect 9493 34660 9505 34663
rect 9456 34632 9505 34660
rect 9456 34620 9462 34632
rect 9493 34629 9505 34632
rect 9539 34629 9551 34663
rect 9493 34623 9551 34629
rect 9674 34620 9680 34672
rect 9732 34660 9738 34672
rect 10796 34669 10824 34700
rect 10870 34688 10876 34740
rect 10928 34688 10934 34740
rect 13004 34700 13400 34728
rect 10321 34663 10379 34669
rect 10321 34660 10333 34663
rect 9732 34632 10333 34660
rect 9732 34620 9738 34632
rect 10321 34629 10333 34632
rect 10367 34629 10379 34663
rect 10321 34623 10379 34629
rect 10781 34663 10839 34669
rect 10781 34629 10793 34663
rect 10827 34629 10839 34663
rect 10781 34623 10839 34629
rect 11330 34620 11336 34672
rect 11388 34660 11394 34672
rect 13004 34660 13032 34700
rect 11388 34632 13032 34660
rect 11388 34620 11394 34632
rect 1857 34595 1915 34601
rect 1857 34561 1869 34595
rect 1903 34592 1915 34595
rect 2038 34592 2044 34604
rect 1903 34564 2044 34592
rect 1903 34561 1915 34564
rect 1857 34555 1915 34561
rect 2038 34552 2044 34564
rect 2096 34552 2102 34604
rect 2131 34595 2189 34601
rect 2131 34561 2143 34595
rect 2177 34592 2189 34595
rect 2590 34592 2596 34604
rect 2177 34564 2596 34592
rect 2177 34561 2189 34564
rect 2131 34555 2189 34561
rect 2590 34552 2596 34564
rect 2648 34592 2654 34604
rect 3511 34595 3569 34601
rect 3511 34592 3523 34595
rect 2648 34564 3523 34592
rect 2648 34552 2654 34564
rect 3511 34561 3523 34564
rect 3557 34592 3569 34595
rect 4890 34592 4896 34604
rect 3557 34564 4896 34592
rect 3557 34561 3569 34564
rect 3511 34555 3569 34561
rect 4890 34552 4896 34564
rect 4948 34552 4954 34604
rect 5537 34595 5595 34601
rect 5537 34561 5549 34595
rect 5583 34592 5595 34595
rect 5994 34592 6000 34604
rect 5583 34564 6000 34592
rect 5583 34561 5595 34564
rect 5537 34555 5595 34561
rect 5994 34552 6000 34564
rect 6052 34552 6058 34604
rect 6549 34595 6607 34601
rect 6549 34561 6561 34595
rect 6595 34592 6607 34595
rect 6595 34564 6868 34592
rect 6595 34561 6607 34564
rect 6549 34555 6607 34561
rect 2958 34484 2964 34536
rect 3016 34524 3022 34536
rect 3237 34527 3295 34533
rect 3237 34524 3249 34527
rect 3016 34496 3249 34524
rect 3016 34484 3022 34496
rect 3237 34493 3249 34496
rect 3283 34493 3295 34527
rect 3237 34487 3295 34493
rect 4982 34484 4988 34536
rect 5040 34484 5046 34536
rect 5902 34484 5908 34536
rect 5960 34484 5966 34536
rect 5920 34456 5948 34484
rect 6840 34468 6868 34564
rect 7190 34552 7196 34604
rect 7248 34592 7254 34604
rect 7653 34595 7711 34601
rect 7653 34592 7665 34595
rect 7248 34564 7665 34592
rect 7248 34552 7254 34564
rect 7653 34561 7665 34564
rect 7699 34561 7711 34595
rect 7926 34592 7932 34604
rect 7887 34564 7932 34592
rect 7653 34555 7711 34561
rect 6089 34459 6147 34465
rect 6089 34456 6101 34459
rect 2746 34428 3004 34456
rect 382 34348 388 34400
rect 440 34388 446 34400
rect 2746 34388 2774 34428
rect 440 34360 2774 34388
rect 440 34348 446 34360
rect 2866 34348 2872 34400
rect 2924 34348 2930 34400
rect 2976 34388 3004 34428
rect 4172 34428 4660 34456
rect 5920 34428 6101 34456
rect 4172 34388 4200 34428
rect 4632 34400 4660 34428
rect 6089 34425 6101 34428
rect 6135 34425 6147 34459
rect 6089 34419 6147 34425
rect 6822 34416 6828 34468
rect 6880 34416 6886 34468
rect 2976 34360 4200 34388
rect 4246 34348 4252 34400
rect 4304 34348 4310 34400
rect 4614 34348 4620 34400
rect 4672 34348 4678 34400
rect 7668 34388 7696 34555
rect 7926 34552 7932 34564
rect 7984 34552 7990 34604
rect 9582 34552 9588 34604
rect 9640 34552 9646 34604
rect 9950 34552 9956 34604
rect 10008 34552 10014 34604
rect 10042 34552 10048 34604
rect 10100 34592 10106 34604
rect 10686 34592 10692 34604
rect 10100 34564 10692 34592
rect 10100 34552 10106 34564
rect 10686 34552 10692 34564
rect 10744 34592 10750 34604
rect 11348 34592 11376 34620
rect 10744 34564 11376 34592
rect 10744 34552 10750 34564
rect 12618 34552 12624 34604
rect 12676 34552 12682 34604
rect 13004 34601 13032 34632
rect 13078 34620 13084 34672
rect 13136 34620 13142 34672
rect 12989 34595 13047 34601
rect 12989 34561 13001 34595
rect 13035 34561 13047 34595
rect 13096 34592 13124 34620
rect 13231 34595 13289 34601
rect 13231 34592 13243 34595
rect 13096 34564 13243 34592
rect 12989 34555 13047 34561
rect 13231 34561 13243 34564
rect 13277 34561 13289 34595
rect 13372 34592 13400 34700
rect 15286 34688 15292 34740
rect 15344 34688 15350 34740
rect 16022 34688 16028 34740
rect 16080 34688 16086 34740
rect 16206 34688 16212 34740
rect 16264 34688 16270 34740
rect 16301 34731 16359 34737
rect 16301 34697 16313 34731
rect 16347 34728 16359 34731
rect 16390 34728 16396 34740
rect 16347 34700 16396 34728
rect 16347 34697 16359 34700
rect 16301 34691 16359 34697
rect 16390 34688 16396 34700
rect 16448 34688 16454 34740
rect 16761 34731 16819 34737
rect 16761 34697 16773 34731
rect 16807 34728 16819 34731
rect 18046 34728 18052 34740
rect 16807 34700 18052 34728
rect 16807 34697 16819 34700
rect 16761 34691 16819 34697
rect 18046 34688 18052 34700
rect 18104 34688 18110 34740
rect 18782 34688 18788 34740
rect 18840 34688 18846 34740
rect 18877 34731 18935 34737
rect 18877 34697 18889 34731
rect 18923 34728 18935 34731
rect 19518 34728 19524 34740
rect 18923 34700 19524 34728
rect 18923 34697 18935 34700
rect 18877 34691 18935 34697
rect 19518 34688 19524 34700
rect 19576 34688 19582 34740
rect 19705 34731 19763 34737
rect 19705 34697 19717 34731
rect 19751 34728 19763 34731
rect 19886 34728 19892 34740
rect 19751 34700 19892 34728
rect 19751 34697 19763 34700
rect 19705 34691 19763 34697
rect 19886 34688 19892 34700
rect 19944 34688 19950 34740
rect 19981 34731 20039 34737
rect 19981 34697 19993 34731
rect 20027 34697 20039 34731
rect 19981 34691 20039 34697
rect 13814 34620 13820 34672
rect 13872 34660 13878 34672
rect 13872 34632 14596 34660
rect 13872 34620 13878 34632
rect 14568 34622 14596 34632
rect 14627 34625 14685 34631
rect 14627 34622 14639 34625
rect 14274 34592 14280 34604
rect 13372 34564 14280 34592
rect 13231 34555 13289 34561
rect 14274 34552 14280 34564
rect 14332 34592 14338 34604
rect 14369 34595 14427 34601
rect 14369 34592 14381 34595
rect 14332 34564 14381 34592
rect 14332 34552 14338 34564
rect 14369 34561 14381 34564
rect 14415 34561 14427 34595
rect 14568 34594 14639 34622
rect 14627 34591 14639 34594
rect 14673 34591 14685 34625
rect 14627 34585 14685 34591
rect 15304 34592 15332 34688
rect 15933 34595 15991 34601
rect 15933 34592 15945 34595
rect 15304 34564 15945 34592
rect 14369 34555 14427 34561
rect 15933 34561 15945 34564
rect 15979 34561 15991 34595
rect 16224 34592 16252 34688
rect 17479 34625 17537 34631
rect 16485 34595 16543 34601
rect 16485 34592 16497 34595
rect 16224 34564 16497 34592
rect 15933 34555 15991 34561
rect 16485 34561 16497 34564
rect 16531 34561 16543 34595
rect 16485 34555 16543 34561
rect 16942 34552 16948 34604
rect 17000 34552 17006 34604
rect 17034 34552 17040 34604
rect 17092 34592 17098 34604
rect 17221 34595 17279 34601
rect 17221 34592 17233 34595
rect 17092 34564 17233 34592
rect 17092 34552 17098 34564
rect 17221 34561 17233 34564
rect 17267 34561 17279 34595
rect 17479 34591 17491 34625
rect 17525 34622 17537 34625
rect 17525 34592 17540 34622
rect 17954 34592 17960 34604
rect 17525 34591 17960 34592
rect 17479 34585 17960 34591
rect 17512 34564 17960 34585
rect 17221 34555 17279 34561
rect 17954 34552 17960 34564
rect 18012 34592 18018 34604
rect 18800 34592 18828 34688
rect 19996 34660 20024 34691
rect 20162 34688 20168 34740
rect 20220 34688 20226 34740
rect 20257 34731 20315 34737
rect 20257 34697 20269 34731
rect 20303 34728 20315 34731
rect 20438 34728 20444 34740
rect 20303 34700 20444 34728
rect 20303 34697 20315 34700
rect 20257 34691 20315 34697
rect 20438 34688 20444 34700
rect 20496 34688 20502 34740
rect 20533 34731 20591 34737
rect 20533 34697 20545 34731
rect 20579 34728 20591 34731
rect 20714 34728 20720 34740
rect 20579 34700 20720 34728
rect 20579 34697 20591 34700
rect 20533 34691 20591 34697
rect 20714 34688 20720 34700
rect 20772 34688 20778 34740
rect 20180 34660 20208 34688
rect 19628 34632 20024 34660
rect 20088 34632 20208 34660
rect 19628 34601 19656 34632
rect 18012 34564 18828 34592
rect 19061 34595 19119 34601
rect 18012 34552 18018 34564
rect 19061 34561 19073 34595
rect 19107 34561 19119 34595
rect 19061 34555 19119 34561
rect 19613 34595 19671 34601
rect 19613 34561 19625 34595
rect 19659 34561 19671 34595
rect 19613 34555 19671 34561
rect 19889 34595 19947 34601
rect 19889 34561 19901 34595
rect 19935 34592 19947 34595
rect 20088 34592 20116 34632
rect 20806 34620 20812 34672
rect 20864 34660 20870 34672
rect 21177 34663 21235 34669
rect 21177 34660 21189 34663
rect 20864 34632 21189 34660
rect 20864 34620 20870 34632
rect 21177 34629 21189 34632
rect 21223 34629 21235 34663
rect 21177 34623 21235 34629
rect 19935 34564 20116 34592
rect 19935 34561 19947 34564
rect 19889 34555 19947 34561
rect 8680 34496 9062 34524
rect 8680 34465 8708 34496
rect 8665 34459 8723 34465
rect 8665 34425 8677 34459
rect 8711 34425 8723 34459
rect 8665 34419 8723 34425
rect 10505 34459 10563 34465
rect 10505 34425 10517 34459
rect 10551 34456 10563 34459
rect 10594 34456 10600 34468
rect 10551 34428 10600 34456
rect 10551 34425 10563 34428
rect 10505 34419 10563 34425
rect 10594 34416 10600 34428
rect 10652 34456 10658 34468
rect 12636 34456 12664 34552
rect 19076 34456 19104 34555
rect 20162 34552 20168 34604
rect 20220 34552 20226 34604
rect 20438 34552 20444 34604
rect 20496 34552 20502 34604
rect 20717 34595 20775 34601
rect 20717 34561 20729 34595
rect 20763 34592 20775 34595
rect 20898 34592 20904 34604
rect 20763 34564 20904 34592
rect 20763 34561 20775 34564
rect 20717 34555 20775 34561
rect 20898 34552 20904 34564
rect 20956 34552 20962 34604
rect 20993 34595 21051 34601
rect 20993 34561 21005 34595
rect 21039 34592 21051 34595
rect 22278 34592 22284 34604
rect 21039 34564 22284 34592
rect 21039 34561 21051 34564
rect 20993 34555 21051 34561
rect 22278 34552 22284 34564
rect 22336 34552 22342 34604
rect 21358 34524 21364 34536
rect 19444 34496 21364 34524
rect 19444 34465 19472 34496
rect 21358 34484 21364 34496
rect 21416 34484 21422 34536
rect 10652 34428 12664 34456
rect 13740 34428 14136 34456
rect 10652 34416 10658 34428
rect 8478 34388 8484 34400
rect 7668 34360 8484 34388
rect 8478 34348 8484 34360
rect 8536 34348 8542 34400
rect 11054 34348 11060 34400
rect 11112 34388 11118 34400
rect 13740 34388 13768 34428
rect 11112 34360 13768 34388
rect 11112 34348 11118 34360
rect 13814 34348 13820 34400
rect 13872 34388 13878 34400
rect 14001 34391 14059 34397
rect 14001 34388 14013 34391
rect 13872 34360 14013 34388
rect 13872 34348 13878 34360
rect 14001 34357 14013 34360
rect 14047 34357 14059 34391
rect 14108 34388 14136 34428
rect 15304 34428 16252 34456
rect 15304 34388 15332 34428
rect 16224 34400 16252 34428
rect 17880 34428 19104 34456
rect 19429 34459 19487 34465
rect 14108 34360 15332 34388
rect 14001 34351 14059 34357
rect 15378 34348 15384 34400
rect 15436 34348 15442 34400
rect 16206 34348 16212 34400
rect 16264 34388 16270 34400
rect 17880 34388 17908 34428
rect 19429 34425 19441 34459
rect 19475 34425 19487 34459
rect 19429 34419 19487 34425
rect 16264 34360 17908 34388
rect 16264 34348 16270 34360
rect 17954 34348 17960 34400
rect 18012 34388 18018 34400
rect 18233 34391 18291 34397
rect 18233 34388 18245 34391
rect 18012 34360 18245 34388
rect 18012 34348 18018 34360
rect 18233 34357 18245 34360
rect 18279 34388 18291 34391
rect 18598 34388 18604 34400
rect 18279 34360 18604 34388
rect 18279 34357 18291 34360
rect 18233 34351 18291 34357
rect 18598 34348 18604 34360
rect 18656 34348 18662 34400
rect 20809 34391 20867 34397
rect 20809 34357 20821 34391
rect 20855 34388 20867 34391
rect 21082 34388 21088 34400
rect 20855 34360 21088 34388
rect 20855 34357 20867 34360
rect 20809 34351 20867 34357
rect 21082 34348 21088 34360
rect 21140 34348 21146 34400
rect 21450 34348 21456 34400
rect 21508 34348 21514 34400
rect 1104 34298 21896 34320
rect 1104 34246 3549 34298
rect 3601 34246 3613 34298
rect 3665 34246 3677 34298
rect 3729 34246 3741 34298
rect 3793 34246 3805 34298
rect 3857 34246 8747 34298
rect 8799 34246 8811 34298
rect 8863 34246 8875 34298
rect 8927 34246 8939 34298
rect 8991 34246 9003 34298
rect 9055 34246 13945 34298
rect 13997 34246 14009 34298
rect 14061 34246 14073 34298
rect 14125 34246 14137 34298
rect 14189 34246 14201 34298
rect 14253 34246 19143 34298
rect 19195 34246 19207 34298
rect 19259 34246 19271 34298
rect 19323 34246 19335 34298
rect 19387 34246 19399 34298
rect 19451 34246 21896 34298
rect 1104 34224 21896 34246
rect 4246 34144 4252 34196
rect 4304 34184 4310 34196
rect 7929 34187 7987 34193
rect 4304 34156 4752 34184
rect 4304 34144 4310 34156
rect 2774 34076 2780 34128
rect 2832 34116 2838 34128
rect 4522 34116 4528 34128
rect 2832 34088 4528 34116
rect 2832 34076 2838 34088
rect 4522 34076 4528 34088
rect 4580 34076 4586 34128
rect 2682 34008 2688 34060
rect 2740 34048 2746 34060
rect 3970 34048 3976 34060
rect 2740 34020 3976 34048
rect 2740 34008 2746 34020
rect 3970 34008 3976 34020
rect 4028 34008 4034 34060
rect 4724 34034 4752 34156
rect 6380 34156 7052 34184
rect 6380 34057 6408 34156
rect 6365 34051 6423 34057
rect 6365 34017 6377 34051
rect 6411 34017 6423 34051
rect 6365 34011 6423 34017
rect 7024 33992 7052 34156
rect 7929 34153 7941 34187
rect 7975 34184 7987 34187
rect 8110 34184 8116 34196
rect 7975 34156 8116 34184
rect 7975 34153 7987 34156
rect 7929 34147 7987 34153
rect 8110 34144 8116 34156
rect 8168 34144 8174 34196
rect 9582 34144 9588 34196
rect 9640 34184 9646 34196
rect 10321 34187 10379 34193
rect 10321 34184 10333 34187
rect 9640 34156 10333 34184
rect 9640 34144 9646 34156
rect 10321 34153 10333 34156
rect 10367 34153 10379 34187
rect 11054 34184 11060 34196
rect 10321 34147 10379 34153
rect 10612 34156 11060 34184
rect 7558 34076 7564 34128
rect 7616 34116 7622 34128
rect 8754 34116 8760 34128
rect 7616 34088 8760 34116
rect 7616 34076 7622 34088
rect 8754 34076 8760 34088
rect 8812 34076 8818 34128
rect 10612 34116 10640 34156
rect 11054 34144 11060 34156
rect 11112 34144 11118 34196
rect 12158 34144 12164 34196
rect 12216 34184 12222 34196
rect 13906 34184 13912 34196
rect 12216 34156 13912 34184
rect 12216 34144 12222 34156
rect 13906 34144 13912 34156
rect 13964 34144 13970 34196
rect 15194 34144 15200 34196
rect 15252 34184 15258 34196
rect 18049 34187 18107 34193
rect 15252 34156 16344 34184
rect 15252 34144 15258 34156
rect 9968 34088 10640 34116
rect 7374 34008 7380 34060
rect 7432 34048 7438 34060
rect 8021 34051 8079 34057
rect 8021 34048 8033 34051
rect 7432 34020 8033 34048
rect 7432 34008 7438 34020
rect 8021 34017 8033 34020
rect 8067 34017 8079 34051
rect 8021 34011 8079 34017
rect 8110 34008 8116 34060
rect 8168 34008 8174 34060
rect 9030 34008 9036 34060
rect 9088 34048 9094 34060
rect 9309 34051 9367 34057
rect 9309 34048 9321 34051
rect 9088 34020 9321 34048
rect 9088 34008 9094 34020
rect 9309 34017 9321 34020
rect 9355 34017 9367 34051
rect 9309 34011 9367 34017
rect 1581 33983 1639 33989
rect 1581 33949 1593 33983
rect 1627 33949 1639 33983
rect 1581 33943 1639 33949
rect 1839 33953 1897 33959
rect 1596 33844 1624 33943
rect 1839 33919 1851 33953
rect 1885 33950 1897 33953
rect 1885 33924 1900 33950
rect 2958 33940 2964 33992
rect 3016 33940 3022 33992
rect 3237 33983 3295 33989
rect 3237 33949 3249 33983
rect 3283 33949 3295 33983
rect 3237 33943 3295 33949
rect 1839 33913 1860 33919
rect 1854 33872 1860 33913
rect 1912 33872 1918 33924
rect 2406 33844 2412 33856
rect 1596 33816 2412 33844
rect 2406 33804 2412 33816
rect 2464 33804 2470 33856
rect 2590 33804 2596 33856
rect 2648 33804 2654 33856
rect 3252 33844 3280 33943
rect 3326 33940 3332 33992
rect 3384 33980 3390 33992
rect 3789 33983 3847 33989
rect 3789 33980 3801 33983
rect 3384 33952 3801 33980
rect 3384 33940 3390 33952
rect 3789 33949 3801 33952
rect 3835 33949 3847 33983
rect 3789 33943 3847 33949
rect 5074 33940 5080 33992
rect 5132 33980 5138 33992
rect 5169 33983 5227 33989
rect 5169 33980 5181 33983
rect 5132 33952 5181 33980
rect 5132 33940 5138 33952
rect 5169 33949 5181 33952
rect 5215 33949 5227 33983
rect 5169 33943 5227 33949
rect 5261 33983 5319 33989
rect 5261 33949 5273 33983
rect 5307 33980 5319 33983
rect 5442 33980 5448 33992
rect 5307 33952 5448 33980
rect 5307 33949 5319 33952
rect 5261 33943 5319 33949
rect 5442 33940 5448 33952
rect 5500 33940 5506 33992
rect 5629 33983 5687 33989
rect 5629 33949 5641 33983
rect 5675 33980 5687 33983
rect 5994 33980 6000 33992
rect 5675 33952 6000 33980
rect 5675 33949 5687 33952
rect 5629 33943 5687 33949
rect 5994 33940 6000 33952
rect 6052 33940 6058 33992
rect 6546 33940 6552 33992
rect 6604 33980 6610 33992
rect 6639 33983 6697 33989
rect 6639 33980 6651 33983
rect 6604 33952 6651 33980
rect 6604 33940 6610 33952
rect 6639 33949 6651 33952
rect 6685 33949 6697 33983
rect 6639 33943 6697 33949
rect 7006 33940 7012 33992
rect 7064 33940 7070 33992
rect 7098 33940 7104 33992
rect 7156 33980 7162 33992
rect 7745 33983 7803 33989
rect 7745 33980 7757 33983
rect 7156 33952 7757 33980
rect 7156 33940 7162 33952
rect 7745 33949 7757 33952
rect 7791 33949 7803 33983
rect 7745 33943 7803 33949
rect 7837 33983 7895 33989
rect 7837 33949 7849 33983
rect 7883 33949 7895 33983
rect 8128 33980 8156 34008
rect 9551 33983 9609 33989
rect 9551 33980 9563 33983
rect 8128 33952 9563 33980
rect 7837 33943 7895 33949
rect 9551 33949 9563 33952
rect 9597 33980 9609 33983
rect 9968 33980 9996 34088
rect 16316 34060 16344 34156
rect 18049 34153 18061 34187
rect 18095 34184 18107 34187
rect 18230 34184 18236 34196
rect 18095 34156 18236 34184
rect 18095 34153 18107 34156
rect 18049 34147 18107 34153
rect 18230 34144 18236 34156
rect 18288 34144 18294 34196
rect 19245 34187 19303 34193
rect 19245 34153 19257 34187
rect 19291 34184 19303 34187
rect 20438 34184 20444 34196
rect 19291 34156 20444 34184
rect 19291 34153 19303 34156
rect 19245 34147 19303 34153
rect 20438 34144 20444 34156
rect 20496 34144 20502 34196
rect 21174 34144 21180 34196
rect 21232 34144 21238 34196
rect 17957 34119 18015 34125
rect 17957 34085 17969 34119
rect 18003 34085 18015 34119
rect 18877 34119 18935 34125
rect 18877 34116 18889 34119
rect 17957 34079 18015 34085
rect 18156 34088 18889 34116
rect 10686 34008 10692 34060
rect 10744 34008 10750 34060
rect 13170 34008 13176 34060
rect 13228 34048 13234 34060
rect 14274 34048 14280 34060
rect 13228 34020 14280 34048
rect 13228 34008 13234 34020
rect 14274 34008 14280 34020
rect 14332 34008 14338 34060
rect 16298 34008 16304 34060
rect 16356 34008 16362 34060
rect 17972 34048 18000 34079
rect 17788 34020 18000 34048
rect 9597 33952 9996 33980
rect 9597 33949 9609 33952
rect 9551 33943 9609 33949
rect 4065 33915 4123 33921
rect 4065 33881 4077 33915
rect 4111 33912 4123 33915
rect 4338 33912 4344 33924
rect 4111 33884 4344 33912
rect 4111 33881 4123 33884
rect 4065 33875 4123 33881
rect 4338 33872 4344 33884
rect 4396 33872 4402 33924
rect 4798 33872 4804 33924
rect 4856 33912 4862 33924
rect 4893 33915 4951 33921
rect 4893 33912 4905 33915
rect 4856 33884 4905 33912
rect 4856 33872 4862 33884
rect 4893 33881 4905 33884
rect 4939 33912 4951 33915
rect 7852 33912 7880 33943
rect 10410 33940 10416 33992
rect 10468 33980 10474 33992
rect 10963 33983 11021 33989
rect 10963 33980 10975 33983
rect 10468 33952 10975 33980
rect 10468 33940 10474 33952
rect 10963 33949 10975 33952
rect 11009 33980 11021 33983
rect 11009 33952 13124 33980
rect 11009 33949 11021 33952
rect 10963 33943 11021 33949
rect 4939 33884 5210 33912
rect 4939 33881 4951 33884
rect 4893 33875 4951 33881
rect 5182 33856 5210 33884
rect 5276 33884 6224 33912
rect 5276 33856 5304 33884
rect 4982 33844 4988 33856
rect 3252 33816 4988 33844
rect 4982 33804 4988 33816
rect 5040 33804 5046 33856
rect 5166 33804 5172 33856
rect 5224 33804 5230 33856
rect 5258 33804 5264 33856
rect 5316 33804 5322 33856
rect 5997 33847 6055 33853
rect 5997 33813 6009 33847
rect 6043 33844 6055 33847
rect 6086 33844 6092 33856
rect 6043 33816 6092 33844
rect 6043 33813 6055 33816
rect 5997 33807 6055 33813
rect 6086 33804 6092 33816
rect 6144 33804 6150 33856
rect 6196 33853 6224 33884
rect 6656 33884 7880 33912
rect 6656 33856 6684 33884
rect 8018 33872 8024 33924
rect 8076 33912 8082 33924
rect 12894 33912 12900 33924
rect 8076 33884 12900 33912
rect 8076 33872 8082 33884
rect 12894 33872 12900 33884
rect 12952 33872 12958 33924
rect 13096 33912 13124 33952
rect 14550 33940 14556 33992
rect 14608 33980 14614 33992
rect 14734 33980 14740 33992
rect 14608 33952 14740 33980
rect 14608 33940 14614 33952
rect 14734 33940 14740 33952
rect 14792 33980 14798 33992
rect 14921 33983 14979 33989
rect 14921 33980 14933 33983
rect 14792 33952 14933 33980
rect 14792 33940 14798 33952
rect 14921 33949 14933 33952
rect 14967 33949 14979 33983
rect 14921 33943 14979 33949
rect 15195 33983 15253 33989
rect 15195 33949 15207 33983
rect 15241 33980 15253 33983
rect 15241 33952 15332 33980
rect 15241 33949 15253 33952
rect 15195 33943 15253 33949
rect 15304 33924 15332 33952
rect 13096 33884 13584 33912
rect 13556 33856 13584 33884
rect 15286 33872 15292 33924
rect 15344 33872 15350 33924
rect 16568 33915 16626 33921
rect 16568 33881 16580 33915
rect 16614 33912 16626 33915
rect 16942 33912 16948 33924
rect 16614 33884 16948 33912
rect 16614 33881 16626 33884
rect 16568 33875 16626 33881
rect 16942 33872 16948 33884
rect 17000 33872 17006 33924
rect 17788 33912 17816 34020
rect 18046 34008 18052 34060
rect 18104 34008 18110 34060
rect 18156 34057 18184 34088
rect 18877 34085 18889 34088
rect 18923 34085 18935 34119
rect 18877 34079 18935 34085
rect 19981 34119 20039 34125
rect 19981 34085 19993 34119
rect 20027 34116 20039 34119
rect 21192 34116 21220 34144
rect 20027 34088 21220 34116
rect 20027 34085 20039 34088
rect 19981 34079 20039 34085
rect 18141 34051 18199 34057
rect 18141 34017 18153 34051
rect 18187 34017 18199 34051
rect 18141 34011 18199 34017
rect 18598 34008 18604 34060
rect 18656 34048 18662 34060
rect 21450 34048 21456 34060
rect 18656 34020 18828 34048
rect 18656 34008 18662 34020
rect 17865 33983 17923 33989
rect 17865 33949 17877 33983
rect 17911 33980 17923 33983
rect 17954 33980 17960 33992
rect 17911 33952 17960 33980
rect 17911 33949 17923 33952
rect 17865 33943 17923 33949
rect 17954 33940 17960 33952
rect 18012 33940 18018 33992
rect 18064 33980 18092 34008
rect 18800 33989 18828 34020
rect 21192 34020 21456 34048
rect 18233 33983 18291 33989
rect 18233 33980 18245 33983
rect 18064 33952 18245 33980
rect 18233 33949 18245 33952
rect 18279 33949 18291 33983
rect 18693 33983 18751 33989
rect 18693 33980 18705 33983
rect 18233 33943 18291 33949
rect 18430 33952 18705 33980
rect 18325 33915 18383 33921
rect 18325 33912 18337 33915
rect 17788 33884 18337 33912
rect 18325 33881 18337 33884
rect 18371 33881 18383 33915
rect 18325 33875 18383 33881
rect 6181 33847 6239 33853
rect 6181 33813 6193 33847
rect 6227 33813 6239 33847
rect 6181 33807 6239 33813
rect 6638 33804 6644 33856
rect 6696 33804 6702 33856
rect 6914 33804 6920 33856
rect 6972 33844 6978 33856
rect 7377 33847 7435 33853
rect 7377 33844 7389 33847
rect 6972 33816 7389 33844
rect 6972 33804 6978 33816
rect 7377 33813 7389 33816
rect 7423 33813 7435 33847
rect 7377 33807 7435 33813
rect 9306 33804 9312 33856
rect 9364 33844 9370 33856
rect 9582 33844 9588 33856
rect 9364 33816 9588 33844
rect 9364 33804 9370 33816
rect 9582 33804 9588 33816
rect 9640 33804 9646 33856
rect 10962 33804 10968 33856
rect 11020 33844 11026 33856
rect 11701 33847 11759 33853
rect 11701 33844 11713 33847
rect 11020 33816 11713 33844
rect 11020 33804 11026 33816
rect 11701 33813 11713 33816
rect 11747 33813 11759 33847
rect 11701 33807 11759 33813
rect 13538 33804 13544 33856
rect 13596 33804 13602 33856
rect 15930 33804 15936 33856
rect 15988 33804 15994 33856
rect 17681 33847 17739 33853
rect 17681 33813 17693 33847
rect 17727 33844 17739 33847
rect 18430 33844 18458 33952
rect 18693 33949 18705 33952
rect 18739 33949 18751 33983
rect 18693 33943 18751 33949
rect 18785 33983 18843 33989
rect 18785 33949 18797 33983
rect 18831 33949 18843 33983
rect 18785 33943 18843 33949
rect 18969 33983 19027 33989
rect 18969 33949 18981 33983
rect 19015 33949 19027 33983
rect 18969 33943 19027 33949
rect 18984 33912 19012 33943
rect 19426 33940 19432 33992
rect 19484 33940 19490 33992
rect 19886 33940 19892 33992
rect 19944 33940 19950 33992
rect 20165 33983 20223 33989
rect 20165 33949 20177 33983
rect 20211 33949 20223 33983
rect 20165 33943 20223 33949
rect 18524 33884 19012 33912
rect 18524 33853 18552 33884
rect 19150 33872 19156 33924
rect 19208 33912 19214 33924
rect 20180 33912 20208 33943
rect 20346 33940 20352 33992
rect 20404 33940 20410 33992
rect 20622 33940 20628 33992
rect 20680 33940 20686 33992
rect 20714 33940 20720 33992
rect 20772 33980 20778 33992
rect 21192 33989 21220 34020
rect 21450 34008 21456 34020
rect 21508 34008 21514 34060
rect 20809 33983 20867 33989
rect 20809 33980 20821 33983
rect 20772 33952 20821 33980
rect 20772 33940 20778 33952
rect 20809 33949 20821 33952
rect 20855 33949 20867 33983
rect 20809 33943 20867 33949
rect 21177 33983 21235 33989
rect 21177 33949 21189 33983
rect 21223 33949 21235 33983
rect 21177 33943 21235 33949
rect 21266 33940 21272 33992
rect 21324 33940 21330 33992
rect 19208 33884 20208 33912
rect 19208 33872 19214 33884
rect 20254 33872 20260 33924
rect 20312 33912 20318 33924
rect 20530 33912 20536 33924
rect 20312 33884 20536 33912
rect 20312 33872 20318 33884
rect 20530 33872 20536 33884
rect 20588 33872 20594 33924
rect 17727 33816 18458 33844
rect 18509 33847 18567 33853
rect 17727 33813 17739 33816
rect 17681 33807 17739 33813
rect 18509 33813 18521 33847
rect 18555 33813 18567 33847
rect 18509 33807 18567 33813
rect 19702 33804 19708 33856
rect 19760 33804 19766 33856
rect 20441 33847 20499 33853
rect 20441 33813 20453 33847
rect 20487 33844 20499 33847
rect 20714 33844 20720 33856
rect 20487 33816 20720 33844
rect 20487 33813 20499 33816
rect 20441 33807 20499 33813
rect 20714 33804 20720 33816
rect 20772 33804 20778 33856
rect 20806 33804 20812 33856
rect 20864 33804 20870 33856
rect 20993 33847 21051 33853
rect 20993 33813 21005 33847
rect 21039 33844 21051 33847
rect 21266 33844 21272 33856
rect 21039 33816 21272 33844
rect 21039 33813 21051 33816
rect 20993 33807 21051 33813
rect 21266 33804 21272 33816
rect 21324 33804 21330 33856
rect 21453 33847 21511 33853
rect 21453 33813 21465 33847
rect 21499 33844 21511 33847
rect 22186 33844 22192 33856
rect 21499 33816 22192 33844
rect 21499 33813 21511 33816
rect 21453 33807 21511 33813
rect 22186 33804 22192 33816
rect 22244 33804 22250 33856
rect 1104 33754 22056 33776
rect 1104 33702 6148 33754
rect 6200 33702 6212 33754
rect 6264 33702 6276 33754
rect 6328 33702 6340 33754
rect 6392 33702 6404 33754
rect 6456 33702 11346 33754
rect 11398 33702 11410 33754
rect 11462 33702 11474 33754
rect 11526 33702 11538 33754
rect 11590 33702 11602 33754
rect 11654 33702 16544 33754
rect 16596 33702 16608 33754
rect 16660 33702 16672 33754
rect 16724 33702 16736 33754
rect 16788 33702 16800 33754
rect 16852 33702 21742 33754
rect 21794 33702 21806 33754
rect 21858 33702 21870 33754
rect 21922 33702 21934 33754
rect 21986 33702 21998 33754
rect 22050 33702 22056 33754
rect 1104 33680 22056 33702
rect 4157 33643 4215 33649
rect 3160 33612 4090 33640
rect 2774 33532 2780 33584
rect 2832 33572 2838 33584
rect 3160 33581 3188 33612
rect 2869 33575 2927 33581
rect 2869 33572 2881 33575
rect 2832 33544 2881 33572
rect 2832 33532 2838 33544
rect 2869 33541 2881 33544
rect 2915 33541 2927 33575
rect 2869 33535 2927 33541
rect 3145 33575 3203 33581
rect 3145 33541 3157 33575
rect 3191 33541 3203 33575
rect 3145 33535 3203 33541
rect 3878 33532 3884 33584
rect 3936 33572 3942 33584
rect 3973 33575 4031 33581
rect 3973 33572 3985 33575
rect 3936 33544 3985 33572
rect 3936 33532 3942 33544
rect 3973 33541 3985 33544
rect 4019 33541 4031 33575
rect 4062 33572 4090 33612
rect 4157 33609 4169 33643
rect 4203 33640 4215 33643
rect 15378 33640 15384 33652
rect 4203 33612 13308 33640
rect 4203 33609 4215 33612
rect 4157 33603 4215 33609
rect 4062 33544 5028 33572
rect 3973 33535 4031 33541
rect 1394 33464 1400 33516
rect 1452 33464 1458 33516
rect 1946 33464 1952 33516
rect 2004 33464 2010 33516
rect 3234 33464 3240 33516
rect 3292 33464 3298 33516
rect 3605 33507 3663 33513
rect 3605 33473 3617 33507
rect 3651 33504 3663 33507
rect 3651 33476 4016 33504
rect 3651 33473 3663 33476
rect 3605 33467 3663 33473
rect 2872 33448 2924 33454
rect 3988 33448 4016 33476
rect 4798 33464 4804 33516
rect 4856 33504 4862 33516
rect 4891 33507 4949 33513
rect 4891 33504 4903 33507
rect 4856 33476 4903 33504
rect 4856 33464 4862 33476
rect 4891 33473 4903 33476
rect 4937 33473 4949 33507
rect 5000 33504 5028 33544
rect 5074 33532 5080 33584
rect 5132 33572 5138 33584
rect 5534 33572 5540 33584
rect 5132 33544 5540 33572
rect 5132 33532 5138 33544
rect 5534 33532 5540 33544
rect 5592 33532 5598 33584
rect 6730 33532 6736 33584
rect 6788 33572 6794 33584
rect 6788 33544 8156 33572
rect 6788 33532 6794 33544
rect 5902 33504 5908 33516
rect 5000 33476 5908 33504
rect 4891 33467 4949 33473
rect 5902 33464 5908 33476
rect 5960 33464 5966 33516
rect 7467 33507 7525 33513
rect 7467 33473 7479 33507
rect 7513 33504 7525 33507
rect 8018 33504 8024 33516
rect 7513 33476 8024 33504
rect 7513 33473 7525 33476
rect 7467 33467 7525 33473
rect 8018 33464 8024 33476
rect 8076 33464 8082 33516
rect 8128 33504 8156 33544
rect 9674 33532 9680 33584
rect 9732 33572 9738 33584
rect 10689 33575 10747 33581
rect 10689 33572 10701 33575
rect 9732 33544 10701 33572
rect 9732 33532 9738 33544
rect 10689 33541 10701 33544
rect 10735 33572 10747 33575
rect 10870 33572 10876 33584
rect 10735 33544 10876 33572
rect 10735 33541 10747 33544
rect 10689 33535 10747 33541
rect 10870 33532 10876 33544
rect 10928 33532 10934 33584
rect 11054 33532 11060 33584
rect 11112 33532 11118 33584
rect 11241 33575 11299 33581
rect 11241 33541 11253 33575
rect 11287 33572 11299 33575
rect 12066 33572 12072 33584
rect 11287 33544 12072 33572
rect 11287 33541 11299 33544
rect 11241 33535 11299 33541
rect 12066 33532 12072 33544
rect 12124 33532 12130 33584
rect 13078 33532 13084 33584
rect 13136 33572 13142 33584
rect 13173 33575 13231 33581
rect 13173 33572 13185 33575
rect 13136 33544 13185 33572
rect 13136 33532 13142 33544
rect 13173 33541 13185 33544
rect 13219 33541 13231 33575
rect 13173 33535 13231 33541
rect 9307 33507 9365 33513
rect 9307 33504 9319 33507
rect 8128 33476 9319 33504
rect 9307 33473 9319 33476
rect 9353 33504 9365 33507
rect 10410 33504 10416 33516
rect 9353 33476 10416 33504
rect 9353 33473 9365 33476
rect 9307 33467 9365 33473
rect 10410 33464 10416 33476
rect 10468 33464 10474 33516
rect 10778 33464 10784 33516
rect 10836 33464 10842 33516
rect 11072 33504 11100 33532
rect 11440 33504 11560 33514
rect 11759 33507 11817 33513
rect 11759 33504 11771 33507
rect 11072 33486 11771 33504
rect 11072 33476 11468 33486
rect 11532 33476 11771 33486
rect 11759 33473 11771 33476
rect 11805 33473 11817 33507
rect 13280 33504 13308 33612
rect 13556 33612 15384 33640
rect 13354 33532 13360 33584
rect 13412 33572 13418 33584
rect 13556 33581 13584 33612
rect 15378 33600 15384 33612
rect 15436 33600 15442 33652
rect 16669 33643 16727 33649
rect 16669 33609 16681 33643
rect 16715 33609 16727 33643
rect 16669 33603 16727 33609
rect 17037 33643 17095 33649
rect 17037 33609 17049 33643
rect 17083 33640 17095 33643
rect 17126 33640 17132 33652
rect 17083 33612 17132 33640
rect 17083 33609 17095 33612
rect 17037 33603 17095 33609
rect 13449 33575 13507 33581
rect 13449 33572 13461 33575
rect 13412 33544 13461 33572
rect 13412 33532 13418 33544
rect 13449 33541 13461 33544
rect 13495 33541 13507 33575
rect 13449 33535 13507 33541
rect 13541 33575 13599 33581
rect 13541 33541 13553 33575
rect 13587 33541 13599 33575
rect 13541 33535 13599 33541
rect 13722 33532 13728 33584
rect 13780 33572 13786 33584
rect 13909 33575 13967 33581
rect 13909 33572 13921 33575
rect 13780 33544 13921 33572
rect 13780 33532 13786 33544
rect 13909 33541 13921 33544
rect 13955 33541 13967 33575
rect 13909 33535 13967 33541
rect 14274 33532 14280 33584
rect 14332 33532 14338 33584
rect 14550 33532 14556 33584
rect 14608 33572 14614 33584
rect 14608 33544 14688 33572
rect 14608 33532 14614 33544
rect 14660 33513 14688 33544
rect 15010 33532 15016 33584
rect 15068 33572 15074 33584
rect 16574 33572 16580 33584
rect 15068 33544 16580 33572
rect 15068 33532 15074 33544
rect 16574 33532 16580 33544
rect 16632 33532 16638 33584
rect 16684 33572 16712 33603
rect 17126 33600 17132 33612
rect 17184 33600 17190 33652
rect 19150 33600 19156 33652
rect 19208 33600 19214 33652
rect 19702 33600 19708 33652
rect 19760 33600 19766 33652
rect 19886 33600 19892 33652
rect 19944 33640 19950 33652
rect 19981 33643 20039 33649
rect 19981 33640 19993 33643
rect 19944 33612 19993 33640
rect 19944 33600 19950 33612
rect 19981 33609 19993 33612
rect 20027 33609 20039 33643
rect 19981 33603 20039 33609
rect 19720 33572 19748 33600
rect 20441 33575 20499 33581
rect 20441 33572 20453 33575
rect 16684 33544 17356 33572
rect 19720 33544 20453 33572
rect 14645 33507 14703 33513
rect 13280 33476 14596 33504
rect 11759 33467 11817 33473
rect 1673 33439 1731 33445
rect 1673 33405 1685 33439
rect 1719 33436 1731 33439
rect 2038 33436 2044 33448
rect 1719 33408 2044 33436
rect 1719 33405 1731 33408
rect 1673 33399 1731 33405
rect 2038 33396 2044 33408
rect 2096 33396 2102 33448
rect 2222 33396 2228 33448
rect 2280 33396 2286 33448
rect 3970 33396 3976 33448
rect 4028 33396 4034 33448
rect 4246 33396 4252 33448
rect 4304 33436 4310 33448
rect 4617 33439 4675 33445
rect 4617 33436 4629 33439
rect 4304 33408 4629 33436
rect 4304 33396 4310 33408
rect 4617 33405 4629 33408
rect 4663 33405 4675 33439
rect 4617 33399 4675 33405
rect 2872 33390 2924 33396
rect 4632 33300 4660 33399
rect 5350 33396 5356 33448
rect 5408 33436 5414 33448
rect 6730 33436 6736 33448
rect 5408 33408 6736 33436
rect 5408 33396 5414 33408
rect 6730 33396 6736 33408
rect 6788 33436 6794 33448
rect 7193 33439 7251 33445
rect 7193 33436 7205 33439
rect 6788 33408 7205 33436
rect 6788 33396 6794 33408
rect 7193 33405 7205 33408
rect 7239 33405 7251 33439
rect 7193 33399 7251 33405
rect 8478 33396 8484 33448
rect 8536 33436 8542 33448
rect 9030 33436 9036 33448
rect 8536 33408 9036 33436
rect 8536 33396 8542 33408
rect 9030 33396 9036 33408
rect 9088 33396 9094 33448
rect 9766 33396 9772 33448
rect 9824 33436 9830 33448
rect 9950 33436 9956 33448
rect 9824 33408 9956 33436
rect 9824 33396 9830 33408
rect 9950 33396 9956 33408
rect 10008 33396 10014 33448
rect 10796 33436 10824 33464
rect 11146 33436 11152 33448
rect 10796 33408 11152 33436
rect 11146 33396 11152 33408
rect 11204 33396 11210 33448
rect 11422 33396 11428 33448
rect 11480 33436 11486 33448
rect 11517 33439 11575 33445
rect 11517 33436 11529 33439
rect 11480 33408 11529 33436
rect 11480 33396 11486 33408
rect 11517 33405 11529 33408
rect 11563 33405 11575 33439
rect 11517 33399 11575 33405
rect 13814 33396 13820 33448
rect 13872 33396 13878 33448
rect 14458 33396 14464 33448
rect 14516 33396 14522 33448
rect 7006 33368 7012 33380
rect 5276 33340 7012 33368
rect 5276 33300 5304 33340
rect 7006 33328 7012 33340
rect 7064 33328 7070 33380
rect 4632 33272 5304 33300
rect 5626 33260 5632 33312
rect 5684 33260 5690 33312
rect 5810 33260 5816 33312
rect 5868 33300 5874 33312
rect 6914 33300 6920 33312
rect 5868 33272 6920 33300
rect 5868 33260 5874 33272
rect 6914 33260 6920 33272
rect 6972 33260 6978 33312
rect 7098 33260 7104 33312
rect 7156 33300 7162 33312
rect 8205 33303 8263 33309
rect 8205 33300 8217 33303
rect 7156 33272 8217 33300
rect 7156 33260 7162 33272
rect 8205 33269 8217 33272
rect 8251 33269 8263 33303
rect 8205 33263 8263 33269
rect 9766 33260 9772 33312
rect 9824 33300 9830 33312
rect 10045 33303 10103 33309
rect 10045 33300 10057 33303
rect 9824 33272 10057 33300
rect 9824 33260 9830 33272
rect 10045 33269 10057 33272
rect 10091 33269 10103 33303
rect 10045 33263 10103 33269
rect 10778 33260 10784 33312
rect 10836 33260 10842 33312
rect 11238 33260 11244 33312
rect 11296 33300 11302 33312
rect 12529 33303 12587 33309
rect 12529 33300 12541 33303
rect 11296 33272 12541 33300
rect 11296 33260 11302 33272
rect 12529 33269 12541 33272
rect 12575 33269 12587 33303
rect 12529 33263 12587 33269
rect 12618 33260 12624 33312
rect 12676 33300 12682 33312
rect 12802 33300 12808 33312
rect 12676 33272 12808 33300
rect 12676 33260 12682 33272
rect 12802 33260 12808 33272
rect 12860 33300 12866 33312
rect 12986 33300 12992 33312
rect 12860 33272 12992 33300
rect 12860 33260 12866 33272
rect 12986 33260 12992 33272
rect 13044 33260 13050 33312
rect 14476 33309 14504 33396
rect 14461 33303 14519 33309
rect 14461 33269 14473 33303
rect 14507 33269 14519 33303
rect 14568 33300 14596 33476
rect 14645 33473 14657 33507
rect 14691 33473 14703 33507
rect 14645 33467 14703 33473
rect 14919 33507 14977 33513
rect 14919 33473 14931 33507
rect 14965 33504 14977 33507
rect 15838 33504 15844 33516
rect 14965 33476 15844 33504
rect 14965 33473 14977 33476
rect 14919 33467 14977 33473
rect 15838 33464 15844 33476
rect 15896 33464 15902 33516
rect 16853 33507 16911 33513
rect 16853 33473 16865 33507
rect 16899 33473 16911 33507
rect 16853 33467 16911 33473
rect 16758 33436 16764 33448
rect 15580 33408 16764 33436
rect 15580 33300 15608 33408
rect 16758 33396 16764 33408
rect 16816 33436 16822 33448
rect 16868 33436 16896 33467
rect 17218 33464 17224 33516
rect 17276 33464 17282 33516
rect 17328 33513 17356 33544
rect 20441 33541 20453 33544
rect 20487 33541 20499 33575
rect 20441 33535 20499 33541
rect 20990 33532 20996 33584
rect 21048 33532 21054 33584
rect 17313 33507 17371 33513
rect 17313 33473 17325 33507
rect 17359 33473 17371 33507
rect 17313 33467 17371 33473
rect 19334 33464 19340 33516
rect 19392 33464 19398 33516
rect 19702 33464 19708 33516
rect 19760 33504 19766 33516
rect 19889 33507 19947 33513
rect 19889 33504 19901 33507
rect 19760 33476 19901 33504
rect 19760 33464 19766 33476
rect 19889 33473 19901 33476
rect 19935 33473 19947 33507
rect 19889 33467 19947 33473
rect 20165 33507 20223 33513
rect 20165 33473 20177 33507
rect 20211 33473 20223 33507
rect 20165 33467 20223 33473
rect 16816 33408 16896 33436
rect 16816 33396 16822 33408
rect 18874 33396 18880 33448
rect 18932 33436 18938 33448
rect 20180 33436 20208 33467
rect 20346 33464 20352 33516
rect 20404 33464 20410 33516
rect 18932 33408 20208 33436
rect 18932 33396 18938 33408
rect 16574 33328 16580 33380
rect 16632 33368 16638 33380
rect 17126 33368 17132 33380
rect 16632 33340 17132 33368
rect 16632 33328 16638 33340
rect 17126 33328 17132 33340
rect 17184 33328 17190 33380
rect 19705 33371 19763 33377
rect 19705 33337 19717 33371
rect 19751 33368 19763 33371
rect 20364 33368 20392 33464
rect 19751 33340 20392 33368
rect 19751 33337 19763 33340
rect 19705 33331 19763 33337
rect 14568 33272 15608 33300
rect 14461 33263 14519 33269
rect 15654 33260 15660 33312
rect 15712 33260 15718 33312
rect 17405 33303 17463 33309
rect 17405 33269 17417 33303
rect 17451 33300 17463 33303
rect 18046 33300 18052 33312
rect 17451 33272 18052 33300
rect 17451 33269 17463 33272
rect 17405 33263 17463 33269
rect 18046 33260 18052 33272
rect 18104 33260 18110 33312
rect 19886 33260 19892 33312
rect 19944 33300 19950 33312
rect 20438 33300 20444 33312
rect 19944 33272 20444 33300
rect 19944 33260 19950 33272
rect 20438 33260 20444 33272
rect 20496 33260 20502 33312
rect 20717 33303 20775 33309
rect 20717 33269 20729 33303
rect 20763 33300 20775 33303
rect 21174 33300 21180 33312
rect 20763 33272 21180 33300
rect 20763 33269 20775 33272
rect 20717 33263 20775 33269
rect 21174 33260 21180 33272
rect 21232 33260 21238 33312
rect 21266 33260 21272 33312
rect 21324 33260 21330 33312
rect 1104 33210 21896 33232
rect 1104 33158 3549 33210
rect 3601 33158 3613 33210
rect 3665 33158 3677 33210
rect 3729 33158 3741 33210
rect 3793 33158 3805 33210
rect 3857 33158 8747 33210
rect 8799 33158 8811 33210
rect 8863 33158 8875 33210
rect 8927 33158 8939 33210
rect 8991 33158 9003 33210
rect 9055 33158 13945 33210
rect 13997 33158 14009 33210
rect 14061 33158 14073 33210
rect 14125 33158 14137 33210
rect 14189 33158 14201 33210
rect 14253 33158 19143 33210
rect 19195 33158 19207 33210
rect 19259 33158 19271 33210
rect 19323 33158 19335 33210
rect 19387 33158 19399 33210
rect 19451 33158 21896 33210
rect 1104 33136 21896 33158
rect 2406 33056 2412 33108
rect 2464 33096 2470 33108
rect 2464 33068 3002 33096
rect 2464 33056 2470 33068
rect 2974 33028 3002 33068
rect 3234 33056 3240 33108
rect 3292 33096 3298 33108
rect 3329 33099 3387 33105
rect 3329 33096 3341 33099
rect 3292 33068 3341 33096
rect 3292 33056 3298 33068
rect 3329 33065 3341 33068
rect 3375 33065 3387 33099
rect 3329 33059 3387 33065
rect 3804 33068 4476 33096
rect 3804 33028 3832 33068
rect 2974 33000 3832 33028
rect 4448 33028 4476 33068
rect 4890 33056 4896 33108
rect 4948 33096 4954 33108
rect 5074 33096 5080 33108
rect 4948 33068 5080 33096
rect 4948 33056 4954 33068
rect 5074 33056 5080 33068
rect 5132 33056 5138 33108
rect 6638 33056 6644 33108
rect 6696 33096 6702 33108
rect 7009 33099 7067 33105
rect 7009 33096 7021 33099
rect 6696 33068 7021 33096
rect 6696 33056 6702 33068
rect 7009 33065 7021 33068
rect 7055 33065 7067 33099
rect 7009 33059 7067 33065
rect 7285 33099 7343 33105
rect 7285 33065 7297 33099
rect 7331 33096 7343 33099
rect 7374 33096 7380 33108
rect 7331 33068 7380 33096
rect 7331 33065 7343 33068
rect 7285 33059 7343 33065
rect 7374 33056 7380 33068
rect 7432 33056 7438 33108
rect 7484 33068 8156 33096
rect 5350 33028 5356 33040
rect 4448 33000 5356 33028
rect 1118 32920 1124 32972
rect 1176 32960 1182 32972
rect 1578 32960 1584 32972
rect 1176 32932 1584 32960
rect 1176 32920 1182 32932
rect 1578 32920 1584 32932
rect 1636 32920 1642 32972
rect 2130 32920 2136 32972
rect 2188 32960 2194 32972
rect 3804 32969 3832 33000
rect 5350 32988 5356 33000
rect 5408 32988 5414 33040
rect 6733 33031 6791 33037
rect 6733 32997 6745 33031
rect 6779 32997 6791 33031
rect 6733 32991 6791 32997
rect 2317 32963 2375 32969
rect 2317 32960 2329 32963
rect 2188 32932 2329 32960
rect 2188 32920 2194 32932
rect 2317 32929 2329 32932
rect 2363 32929 2375 32963
rect 2317 32923 2375 32929
rect 3789 32963 3847 32969
rect 3789 32929 3801 32963
rect 3835 32929 3847 32963
rect 3789 32923 3847 32929
rect 5626 32920 5632 32972
rect 5684 32920 5690 32972
rect 2591 32895 2649 32901
rect 2591 32861 2603 32895
rect 2637 32892 2649 32895
rect 2637 32864 3832 32892
rect 2637 32861 2649 32864
rect 2591 32855 2649 32861
rect 3804 32836 3832 32864
rect 4047 32865 4105 32871
rect 1486 32784 1492 32836
rect 1544 32784 1550 32836
rect 1673 32827 1731 32833
rect 1673 32793 1685 32827
rect 1719 32824 1731 32827
rect 1762 32824 1768 32836
rect 1719 32796 1768 32824
rect 1719 32793 1731 32796
rect 1673 32787 1731 32793
rect 1762 32784 1768 32796
rect 1820 32784 1826 32836
rect 3786 32784 3792 32836
rect 3844 32784 3850 32836
rect 4047 32831 4059 32865
rect 4093 32862 4105 32865
rect 4093 32831 4108 32862
rect 5534 32852 5540 32904
rect 5592 32892 5598 32904
rect 5592 32864 5764 32892
rect 5592 32852 5598 32864
rect 4047 32825 4108 32831
rect 4080 32768 4108 32825
rect 5166 32784 5172 32836
rect 5224 32784 5230 32836
rect 5350 32784 5356 32836
rect 5408 32824 5414 32836
rect 5736 32833 5764 32864
rect 5810 32852 5816 32904
rect 5868 32852 5874 32904
rect 6748 32892 6776 32991
rect 7484 32969 7512 33068
rect 7469 32963 7527 32969
rect 7469 32960 7481 32963
rect 7024 32932 7481 32960
rect 5920 32864 6776 32892
rect 5721 32827 5779 32833
rect 5408 32796 5580 32824
rect 5408 32784 5414 32796
rect 382 32716 388 32768
rect 440 32756 446 32768
rect 3142 32756 3148 32768
rect 440 32728 3148 32756
rect 440 32716 446 32728
rect 3142 32716 3148 32728
rect 3200 32716 3206 32768
rect 4062 32716 4068 32768
rect 4120 32716 4126 32768
rect 4801 32759 4859 32765
rect 4801 32725 4813 32759
rect 4847 32756 4859 32759
rect 4890 32756 4896 32768
rect 4847 32728 4896 32756
rect 4847 32725 4859 32728
rect 4801 32719 4859 32725
rect 4890 32716 4896 32728
rect 4948 32716 4954 32768
rect 5184 32756 5212 32784
rect 5442 32756 5448 32768
rect 5184 32728 5448 32756
rect 5442 32716 5448 32728
rect 5500 32716 5506 32768
rect 5552 32756 5580 32796
rect 5721 32793 5733 32827
rect 5767 32793 5779 32827
rect 5721 32787 5779 32793
rect 5920 32756 5948 32864
rect 6914 32852 6920 32904
rect 6972 32852 6978 32904
rect 5994 32784 6000 32836
rect 6052 32824 6058 32836
rect 6181 32827 6239 32833
rect 6181 32824 6193 32827
rect 6052 32796 6193 32824
rect 6052 32784 6058 32796
rect 6181 32793 6193 32796
rect 6227 32793 6239 32827
rect 6181 32787 6239 32793
rect 5552 32728 5948 32756
rect 6546 32716 6552 32768
rect 6604 32716 6610 32768
rect 6730 32716 6736 32768
rect 6788 32756 6794 32768
rect 7024 32756 7052 32932
rect 7469 32929 7481 32932
rect 7515 32929 7527 32963
rect 8128 32960 8156 33068
rect 8386 33056 8392 33108
rect 8444 33096 8450 33108
rect 12345 33099 12403 33105
rect 8444 33068 10364 33096
rect 8444 33056 8450 33068
rect 8478 32960 8484 32972
rect 8128 32932 8484 32960
rect 7469 32923 7527 32929
rect 8478 32920 8484 32932
rect 8536 32960 8542 32972
rect 8846 32960 8852 32972
rect 8536 32932 8852 32960
rect 8536 32920 8542 32932
rect 8846 32920 8852 32932
rect 8904 32960 8910 32972
rect 9033 32963 9091 32969
rect 9033 32960 9045 32963
rect 8904 32932 9045 32960
rect 8904 32920 8910 32932
rect 9033 32929 9045 32932
rect 9079 32929 9091 32963
rect 9033 32923 9091 32929
rect 7098 32852 7104 32904
rect 7156 32892 7162 32904
rect 7193 32895 7251 32901
rect 7193 32892 7205 32895
rect 7156 32864 7205 32892
rect 7156 32852 7162 32864
rect 7193 32861 7205 32864
rect 7239 32861 7251 32895
rect 7193 32855 7251 32861
rect 7374 32852 7380 32904
rect 7432 32852 7438 32904
rect 7711 32895 7769 32901
rect 7711 32892 7723 32895
rect 7576 32864 7723 32892
rect 7576 32836 7604 32864
rect 7711 32861 7723 32864
rect 7757 32892 7769 32895
rect 8386 32892 8392 32904
rect 7757 32864 8392 32892
rect 7757 32861 7769 32864
rect 7711 32855 7769 32861
rect 8386 32852 8392 32864
rect 8444 32852 8450 32904
rect 9291 32865 9349 32871
rect 7558 32784 7564 32836
rect 7616 32784 7622 32836
rect 9291 32831 9303 32865
rect 9337 32862 9349 32865
rect 9337 32836 9352 32862
rect 9291 32825 9312 32831
rect 9306 32784 9312 32825
rect 9364 32784 9370 32836
rect 10336 32824 10364 33068
rect 12345 33065 12357 33099
rect 12391 33096 12403 33099
rect 15654 33096 15660 33108
rect 12391 33068 14596 33096
rect 12391 33065 12403 33068
rect 12345 33059 12403 33065
rect 10962 32920 10968 32972
rect 11020 32920 11026 32972
rect 12544 32904 12572 33068
rect 14568 33040 14596 33068
rect 15212 33068 15660 33096
rect 14550 32988 14556 33040
rect 14608 32988 14614 33040
rect 15212 33037 15240 33068
rect 15654 33056 15660 33068
rect 15712 33056 15718 33108
rect 15746 33056 15752 33108
rect 15804 33096 15810 33108
rect 17494 33096 17500 33108
rect 15804 33068 17500 33096
rect 15804 33056 15810 33068
rect 17494 33056 17500 33068
rect 17552 33096 17558 33108
rect 17954 33096 17960 33108
rect 17552 33068 17960 33096
rect 17552 33056 17558 33068
rect 17954 33056 17960 33068
rect 18012 33056 18018 33108
rect 18046 33056 18052 33108
rect 18104 33056 18110 33108
rect 18138 33056 18144 33108
rect 18196 33096 18202 33108
rect 18196 33068 18828 33096
rect 18196 33056 18202 33068
rect 15197 33031 15255 33037
rect 15197 32997 15209 33031
rect 15243 32997 15255 33031
rect 15197 32991 15255 32997
rect 17865 33031 17923 33037
rect 17865 32997 17877 33031
rect 17911 33028 17923 33031
rect 18322 33028 18328 33040
rect 17911 33000 18328 33028
rect 17911 32997 17923 33000
rect 17865 32991 17923 32997
rect 18322 32988 18328 33000
rect 18380 32988 18386 33040
rect 18693 33031 18751 33037
rect 18693 33028 18705 33031
rect 18432 33000 18705 33028
rect 12618 32920 12624 32972
rect 12676 32920 12682 32972
rect 15590 32963 15648 32969
rect 15590 32960 15602 32963
rect 13262 32932 15602 32960
rect 10870 32852 10876 32904
rect 10928 32852 10934 32904
rect 11238 32852 11244 32904
rect 11296 32852 11302 32904
rect 11698 32852 11704 32904
rect 11756 32901 11762 32904
rect 11756 32895 11773 32901
rect 11761 32861 11773 32895
rect 11756 32855 11773 32861
rect 11756 32852 11762 32855
rect 12526 32852 12532 32904
rect 12584 32852 12590 32904
rect 13262 32892 13290 32932
rect 15590 32929 15602 32932
rect 15636 32929 15648 32963
rect 15590 32923 15648 32929
rect 15749 32963 15807 32969
rect 15749 32929 15761 32963
rect 15795 32960 15807 32963
rect 15930 32960 15936 32972
rect 15795 32932 15936 32960
rect 15795 32929 15807 32932
rect 15749 32923 15807 32929
rect 15930 32920 15936 32932
rect 15988 32920 15994 32972
rect 16298 32920 16304 32972
rect 16356 32960 16362 32972
rect 16485 32963 16543 32969
rect 16485 32960 16497 32963
rect 16356 32932 16497 32960
rect 16356 32920 16362 32932
rect 16485 32929 16497 32932
rect 16531 32929 16543 32963
rect 18138 32960 18144 32972
rect 16485 32923 16543 32929
rect 17880 32932 18144 32960
rect 12879 32865 12937 32871
rect 12879 32862 12891 32865
rect 10965 32827 11023 32833
rect 10336 32796 10916 32824
rect 6788 32728 7052 32756
rect 6788 32716 6794 32728
rect 7098 32716 7104 32768
rect 7156 32756 7162 32768
rect 7926 32756 7932 32768
rect 7156 32728 7932 32756
rect 7156 32716 7162 32728
rect 7926 32716 7932 32728
rect 7984 32716 7990 32768
rect 8478 32716 8484 32768
rect 8536 32716 8542 32768
rect 10042 32716 10048 32768
rect 10100 32716 10106 32768
rect 10597 32759 10655 32765
rect 10597 32725 10609 32759
rect 10643 32756 10655 32759
rect 10778 32756 10784 32768
rect 10643 32728 10784 32756
rect 10643 32725 10655 32728
rect 10597 32719 10655 32725
rect 10778 32716 10784 32728
rect 10836 32716 10842 32768
rect 10888 32756 10916 32796
rect 10965 32793 10977 32827
rect 11011 32824 11023 32827
rect 11256 32824 11284 32852
rect 11011 32796 11284 32824
rect 11333 32827 11391 32833
rect 11011 32793 11023 32796
rect 10965 32787 11023 32793
rect 11333 32793 11345 32827
rect 11379 32824 11391 32827
rect 12544 32824 12572 32852
rect 12820 32834 12891 32862
rect 12820 32824 12848 32834
rect 12879 32831 12891 32834
rect 12925 32831 12937 32865
rect 12879 32825 12937 32831
rect 13004 32864 13290 32892
rect 11379 32796 12480 32824
rect 12544 32796 12848 32824
rect 11379 32793 11391 32796
rect 11333 32787 11391 32793
rect 11885 32759 11943 32765
rect 11885 32756 11897 32759
rect 10888 32728 11897 32756
rect 11885 32725 11897 32728
rect 11931 32725 11943 32759
rect 12452 32756 12480 32796
rect 12526 32756 12532 32768
rect 12452 32728 12532 32756
rect 11885 32719 11943 32725
rect 12526 32716 12532 32728
rect 12584 32716 12590 32768
rect 12618 32716 12624 32768
rect 12676 32756 12682 32768
rect 13004 32756 13032 32864
rect 14366 32852 14372 32904
rect 14424 32892 14430 32904
rect 14553 32895 14611 32901
rect 14553 32892 14565 32895
rect 14424 32864 14565 32892
rect 14424 32852 14430 32864
rect 14553 32861 14565 32864
rect 14599 32861 14611 32895
rect 14553 32855 14611 32861
rect 14737 32895 14795 32901
rect 14737 32861 14749 32895
rect 14783 32861 14795 32895
rect 14737 32855 14795 32861
rect 14274 32784 14280 32836
rect 14332 32824 14338 32836
rect 14752 32824 14780 32855
rect 15470 32852 15476 32904
rect 15528 32852 15534 32904
rect 16393 32895 16451 32901
rect 16393 32861 16405 32895
rect 16439 32892 16451 32895
rect 17880 32892 17908 32932
rect 18138 32920 18144 32932
rect 18196 32920 18202 32972
rect 18233 32963 18291 32969
rect 18233 32929 18245 32963
rect 18279 32960 18291 32963
rect 18432 32960 18460 33000
rect 18693 32997 18705 33000
rect 18739 32997 18751 33031
rect 18693 32991 18751 32997
rect 18279 32932 18460 32960
rect 18800 32960 18828 33068
rect 18874 33056 18880 33108
rect 18932 33056 18938 33108
rect 20806 33056 20812 33108
rect 20864 33056 20870 33108
rect 20622 32988 20628 33040
rect 20680 32988 20686 33040
rect 18800 32932 19380 32960
rect 18279 32929 18291 32932
rect 18233 32923 18291 32929
rect 16439 32864 17908 32892
rect 17957 32895 18015 32901
rect 16439 32861 16451 32864
rect 16393 32855 16451 32861
rect 17957 32861 17969 32895
rect 18003 32861 18015 32895
rect 17957 32855 18015 32861
rect 16758 32833 16764 32836
rect 16752 32824 16764 32833
rect 14332 32796 14780 32824
rect 16719 32796 16764 32824
rect 14332 32784 14338 32796
rect 16752 32787 16764 32796
rect 16758 32784 16764 32787
rect 16816 32784 16822 32836
rect 17972 32824 18000 32855
rect 18322 32852 18328 32904
rect 18380 32892 18386 32904
rect 18509 32895 18567 32901
rect 18509 32892 18521 32895
rect 18380 32864 18521 32892
rect 18380 32852 18386 32864
rect 18509 32861 18521 32864
rect 18555 32861 18567 32895
rect 18601 32895 18659 32901
rect 18601 32892 18613 32895
rect 18509 32855 18567 32861
rect 18598 32861 18613 32892
rect 18647 32861 18659 32895
rect 18785 32895 18843 32901
rect 18785 32892 18797 32895
rect 18598 32855 18659 32861
rect 18708 32864 18797 32892
rect 18598 32824 18626 32855
rect 17880 32796 18626 32824
rect 17880 32768 17908 32796
rect 12676 32728 13032 32756
rect 12676 32716 12682 32728
rect 13354 32716 13360 32768
rect 13412 32756 13418 32768
rect 13633 32759 13691 32765
rect 13633 32756 13645 32759
rect 13412 32728 13645 32756
rect 13412 32716 13418 32728
rect 13633 32725 13645 32728
rect 13679 32725 13691 32759
rect 13633 32719 13691 32725
rect 17862 32716 17868 32768
rect 17920 32716 17926 32768
rect 18230 32716 18236 32768
rect 18288 32716 18294 32768
rect 18325 32759 18383 32765
rect 18325 32725 18337 32759
rect 18371 32756 18383 32759
rect 18708 32756 18736 32864
rect 18785 32861 18797 32864
rect 18831 32861 18843 32895
rect 18785 32855 18843 32861
rect 18874 32852 18880 32904
rect 18932 32892 18938 32904
rect 19061 32895 19119 32901
rect 19061 32892 19073 32895
rect 18932 32864 19073 32892
rect 18932 32852 18938 32864
rect 19061 32861 19073 32864
rect 19107 32861 19119 32895
rect 19061 32855 19119 32861
rect 19150 32852 19156 32904
rect 19208 32892 19214 32904
rect 19245 32895 19303 32901
rect 19245 32892 19257 32895
rect 19208 32864 19257 32892
rect 19208 32852 19214 32864
rect 19245 32861 19257 32864
rect 19291 32861 19303 32895
rect 19352 32892 19380 32932
rect 20640 32892 20668 32988
rect 20824 32960 20852 33056
rect 21085 33031 21143 33037
rect 21085 32997 21097 33031
rect 21131 33028 21143 33031
rect 21634 33028 21640 33040
rect 21131 33000 21640 33028
rect 21131 32997 21143 33000
rect 21085 32991 21143 32997
rect 21634 32988 21640 33000
rect 21692 32988 21698 33040
rect 20993 32963 21051 32969
rect 20993 32960 21005 32963
rect 20824 32932 21005 32960
rect 20993 32929 21005 32932
rect 21039 32929 21051 32963
rect 20993 32923 21051 32929
rect 22830 32920 22836 32972
rect 22888 32920 22894 32972
rect 20717 32895 20775 32901
rect 20717 32892 20729 32895
rect 19352 32864 19555 32892
rect 20640 32864 20729 32892
rect 19245 32855 19303 32861
rect 19527 32833 19555 32864
rect 20717 32861 20729 32864
rect 20763 32861 20775 32895
rect 20717 32855 20775 32861
rect 20806 32852 20812 32904
rect 20864 32852 20870 32904
rect 20898 32852 20904 32904
rect 20956 32852 20962 32904
rect 21174 32852 21180 32904
rect 21232 32892 21238 32904
rect 21269 32895 21327 32901
rect 21269 32892 21281 32895
rect 21232 32864 21281 32892
rect 21232 32852 21238 32864
rect 21269 32861 21281 32864
rect 21315 32861 21327 32895
rect 21269 32855 21327 32861
rect 21542 32852 21548 32904
rect 21600 32852 21606 32904
rect 22848 32892 22876 32920
rect 22848 32864 22968 32892
rect 19512 32827 19570 32833
rect 19512 32793 19524 32827
rect 19558 32824 19570 32827
rect 19702 32824 19708 32836
rect 19558 32796 19708 32824
rect 19558 32793 19570 32796
rect 19512 32787 19570 32793
rect 19702 32784 19708 32796
rect 19760 32784 19766 32836
rect 18371 32728 18736 32756
rect 18371 32725 18383 32728
rect 18325 32719 18383 32725
rect 18782 32716 18788 32768
rect 18840 32756 18846 32768
rect 19978 32756 19984 32768
rect 18840 32728 19984 32756
rect 18840 32716 18846 32728
rect 19978 32716 19984 32728
rect 20036 32716 20042 32768
rect 20625 32759 20683 32765
rect 20625 32725 20637 32759
rect 20671 32756 20683 32759
rect 20916 32756 20944 32852
rect 22830 32824 22836 32836
rect 21008 32796 22836 32824
rect 21008 32765 21036 32796
rect 22830 32784 22836 32796
rect 22888 32784 22894 32836
rect 20671 32728 20944 32756
rect 20993 32759 21051 32765
rect 20671 32725 20683 32728
rect 20625 32719 20683 32725
rect 20993 32725 21005 32759
rect 21039 32725 21051 32759
rect 20993 32719 21051 32725
rect 21358 32716 21364 32768
rect 21416 32716 21422 32768
rect 1104 32666 22056 32688
rect 1104 32614 6148 32666
rect 6200 32614 6212 32666
rect 6264 32614 6276 32666
rect 6328 32614 6340 32666
rect 6392 32614 6404 32666
rect 6456 32614 11346 32666
rect 11398 32614 11410 32666
rect 11462 32614 11474 32666
rect 11526 32614 11538 32666
rect 11590 32614 11602 32666
rect 11654 32614 16544 32666
rect 16596 32614 16608 32666
rect 16660 32614 16672 32666
rect 16724 32614 16736 32666
rect 16788 32614 16800 32666
rect 16852 32614 21742 32666
rect 21794 32614 21806 32666
rect 21858 32614 21870 32666
rect 21922 32614 21934 32666
rect 21986 32614 21998 32666
rect 22050 32614 22056 32666
rect 1104 32592 22056 32614
rect 2774 32512 2780 32564
rect 2832 32552 2838 32564
rect 3142 32552 3148 32564
rect 2832 32524 3148 32552
rect 2832 32512 2838 32524
rect 3142 32512 3148 32524
rect 3200 32512 3206 32564
rect 4154 32512 4160 32564
rect 4212 32552 4218 32564
rect 4706 32552 4712 32564
rect 4212 32524 4712 32552
rect 4212 32512 4218 32524
rect 4706 32512 4712 32524
rect 4764 32512 4770 32564
rect 5810 32512 5816 32564
rect 5868 32512 5874 32564
rect 6365 32555 6423 32561
rect 6365 32521 6377 32555
rect 6411 32552 6423 32555
rect 6914 32552 6920 32564
rect 6411 32524 6920 32552
rect 6411 32521 6423 32524
rect 6365 32515 6423 32521
rect 6914 32512 6920 32524
rect 6972 32512 6978 32564
rect 7009 32555 7067 32561
rect 7009 32521 7021 32555
rect 7055 32552 7067 32555
rect 7374 32552 7380 32564
rect 7055 32524 7380 32552
rect 7055 32521 7067 32524
rect 7009 32515 7067 32521
rect 7374 32512 7380 32524
rect 7432 32512 7438 32564
rect 8938 32552 8944 32564
rect 7484 32524 8944 32552
rect 750 32444 756 32496
rect 808 32484 814 32496
rect 808 32456 2774 32484
rect 808 32444 814 32456
rect 1823 32419 1881 32425
rect 1823 32416 1835 32419
rect 1320 32388 1835 32416
rect 1320 32212 1348 32388
rect 1823 32385 1835 32388
rect 1869 32416 1881 32419
rect 2314 32416 2320 32428
rect 1869 32388 2320 32416
rect 1869 32385 1881 32388
rect 1823 32379 1881 32385
rect 2314 32376 2320 32388
rect 2372 32376 2378 32428
rect 2746 32416 2774 32456
rect 3234 32444 3240 32496
rect 3292 32444 3298 32496
rect 3878 32484 3884 32496
rect 3712 32456 3884 32484
rect 3712 32425 3740 32456
rect 3878 32444 3884 32456
rect 3936 32444 3942 32496
rect 5828 32484 5856 32512
rect 6730 32484 6736 32496
rect 5828 32456 6736 32484
rect 6730 32444 6736 32456
rect 6788 32444 6794 32496
rect 2961 32419 3019 32425
rect 2961 32416 2973 32419
rect 2746 32388 2973 32416
rect 2961 32385 2973 32388
rect 3007 32385 3019 32419
rect 2961 32379 3019 32385
rect 3697 32419 3755 32425
rect 3697 32385 3709 32419
rect 3743 32385 3755 32419
rect 3697 32379 3755 32385
rect 5537 32419 5595 32425
rect 5537 32385 5549 32419
rect 5583 32416 5595 32419
rect 6549 32419 6607 32425
rect 6549 32416 6561 32419
rect 5583 32388 6561 32416
rect 5583 32385 5595 32388
rect 5537 32379 5595 32385
rect 6549 32385 6561 32388
rect 6595 32385 6607 32419
rect 6549 32379 6607 32385
rect 7190 32376 7196 32428
rect 7248 32376 7254 32428
rect 7285 32419 7343 32425
rect 7285 32385 7297 32419
rect 7331 32416 7343 32419
rect 7374 32416 7380 32438
rect 7331 32388 7380 32416
rect 7331 32385 7343 32388
rect 7374 32386 7380 32388
rect 7432 32416 7438 32438
rect 7484 32416 7512 32524
rect 8938 32512 8944 32524
rect 8996 32512 9002 32564
rect 9048 32524 9260 32552
rect 9048 32496 9076 32524
rect 9030 32444 9036 32496
rect 9088 32444 9094 32496
rect 9125 32487 9183 32493
rect 9125 32453 9137 32487
rect 9171 32453 9183 32487
rect 9232 32484 9260 32524
rect 9306 32512 9312 32564
rect 9364 32552 9370 32564
rect 10962 32552 10968 32564
rect 9364 32524 10968 32552
rect 9364 32512 9370 32524
rect 10962 32512 10968 32524
rect 11020 32512 11026 32564
rect 11241 32555 11299 32561
rect 11241 32521 11253 32555
rect 11287 32552 11299 32555
rect 11790 32552 11796 32564
rect 11287 32524 11796 32552
rect 11287 32521 11299 32524
rect 11241 32515 11299 32521
rect 11790 32512 11796 32524
rect 11848 32512 11854 32564
rect 12526 32512 12532 32564
rect 12584 32552 12590 32564
rect 13078 32552 13084 32564
rect 12584 32524 13084 32552
rect 12584 32512 12590 32524
rect 13078 32512 13084 32524
rect 13136 32512 13142 32564
rect 13446 32512 13452 32564
rect 13504 32552 13510 32564
rect 13906 32552 13912 32564
rect 13504 32524 13912 32552
rect 13504 32512 13510 32524
rect 13906 32512 13912 32524
rect 13964 32552 13970 32564
rect 15930 32552 15936 32564
rect 13964 32524 15936 32552
rect 13964 32512 13970 32524
rect 15930 32512 15936 32524
rect 15988 32512 15994 32564
rect 17862 32512 17868 32564
rect 17920 32512 17926 32564
rect 18969 32555 19027 32561
rect 18969 32521 18981 32555
rect 19015 32552 19027 32555
rect 19015 32524 20576 32552
rect 19015 32521 19027 32524
rect 18969 32515 19027 32521
rect 9401 32487 9459 32493
rect 9401 32484 9413 32487
rect 9232 32456 9413 32484
rect 9125 32447 9183 32453
rect 9401 32453 9413 32456
rect 9447 32453 9459 32487
rect 9401 32447 9459 32453
rect 9493 32487 9551 32493
rect 9493 32453 9505 32487
rect 9539 32484 9551 32487
rect 9766 32484 9772 32496
rect 9539 32456 9772 32484
rect 9539 32453 9551 32456
rect 9493 32447 9551 32453
rect 7432 32388 7512 32416
rect 7432 32386 7438 32388
rect 7285 32379 7343 32385
rect 1394 32308 1400 32360
rect 1452 32348 1458 32360
rect 1581 32351 1639 32357
rect 1581 32348 1593 32351
rect 1452 32320 1593 32348
rect 1452 32308 1458 32320
rect 1581 32317 1593 32320
rect 1627 32317 1639 32351
rect 1581 32311 1639 32317
rect 2590 32308 2596 32360
rect 2648 32308 2654 32360
rect 3326 32308 3332 32360
rect 3384 32348 3390 32360
rect 3881 32351 3939 32357
rect 3881 32348 3893 32351
rect 3384 32320 3893 32348
rect 3384 32308 3390 32320
rect 3881 32317 3893 32320
rect 3927 32317 3939 32351
rect 4617 32351 4675 32357
rect 4617 32348 4629 32351
rect 3881 32311 3939 32317
rect 4448 32320 4629 32348
rect 2608 32280 2636 32308
rect 4246 32280 4252 32292
rect 2608 32252 4252 32280
rect 4246 32240 4252 32252
rect 4304 32280 4310 32292
rect 4341 32283 4399 32289
rect 4341 32280 4353 32283
rect 4304 32252 4353 32280
rect 4304 32240 4310 32252
rect 4341 32249 4353 32252
rect 4387 32249 4399 32283
rect 4341 32243 4399 32249
rect 1578 32212 1584 32224
rect 1320 32184 1584 32212
rect 1578 32172 1584 32184
rect 1636 32172 1642 32224
rect 2593 32215 2651 32221
rect 2593 32181 2605 32215
rect 2639 32212 2651 32215
rect 2958 32212 2964 32224
rect 2639 32184 2964 32212
rect 2639 32181 2651 32184
rect 2593 32175 2651 32181
rect 2958 32172 2964 32184
rect 3016 32172 3022 32224
rect 4448 32212 4476 32320
rect 4617 32317 4629 32320
rect 4663 32317 4675 32351
rect 4617 32311 4675 32317
rect 4706 32308 4712 32360
rect 4764 32357 4770 32360
rect 4764 32351 4813 32357
rect 4764 32317 4767 32351
rect 4801 32317 4813 32351
rect 4764 32311 4813 32317
rect 4764 32308 4770 32311
rect 4890 32308 4896 32360
rect 4948 32348 4954 32360
rect 6178 32348 6184 32360
rect 4948 32320 6184 32348
rect 4948 32308 4954 32320
rect 6178 32308 6184 32320
rect 6236 32308 6242 32360
rect 7006 32308 7012 32360
rect 7064 32348 7070 32360
rect 7300 32348 7328 32379
rect 7558 32376 7564 32428
rect 7616 32416 7622 32428
rect 9140 32416 9168 32447
rect 9766 32444 9772 32456
rect 9824 32444 9830 32496
rect 10226 32444 10232 32496
rect 10284 32444 10290 32496
rect 10410 32444 10416 32496
rect 10468 32484 10474 32496
rect 10468 32456 17170 32484
rect 10468 32444 10474 32456
rect 9674 32416 9680 32428
rect 7616 32388 7659 32416
rect 9140 32388 9680 32416
rect 7616 32376 7622 32388
rect 9674 32376 9680 32388
rect 9732 32376 9738 32428
rect 9861 32419 9919 32425
rect 9861 32385 9873 32419
rect 9907 32416 9919 32419
rect 10686 32416 10692 32428
rect 9907 32388 10692 32416
rect 9907 32385 9919 32388
rect 9861 32379 9919 32385
rect 10686 32376 10692 32388
rect 10744 32376 10750 32428
rect 11054 32376 11060 32428
rect 11112 32376 11118 32428
rect 11330 32376 11336 32428
rect 11388 32416 11394 32428
rect 12621 32419 12679 32425
rect 12621 32416 12633 32419
rect 11388 32388 12633 32416
rect 11388 32376 11394 32388
rect 12621 32385 12633 32388
rect 12667 32416 12679 32419
rect 12802 32416 12808 32428
rect 12667 32388 12808 32416
rect 12667 32385 12679 32388
rect 12621 32379 12679 32385
rect 12802 32376 12808 32388
rect 12860 32376 12866 32428
rect 12895 32419 12953 32425
rect 12895 32385 12907 32419
rect 12941 32416 12953 32419
rect 13630 32416 13636 32428
rect 12941 32388 13636 32416
rect 12941 32385 12953 32388
rect 12895 32379 12953 32385
rect 13630 32376 13636 32388
rect 13688 32376 13694 32428
rect 13814 32376 13820 32428
rect 13872 32416 13878 32428
rect 14243 32419 14301 32425
rect 14243 32416 14255 32419
rect 13872 32388 14255 32416
rect 13872 32376 13878 32388
rect 14243 32385 14255 32388
rect 14289 32385 14301 32419
rect 14243 32379 14301 32385
rect 15470 32376 15476 32428
rect 15528 32416 15534 32428
rect 17142 32425 17170 32456
rect 17678 32444 17684 32496
rect 17736 32484 17742 32496
rect 17954 32484 17960 32496
rect 17736 32456 17960 32484
rect 17736 32444 17742 32456
rect 17954 32444 17960 32456
rect 18012 32444 18018 32496
rect 19978 32484 19984 32496
rect 19168 32456 19984 32484
rect 15657 32419 15715 32425
rect 15657 32416 15669 32419
rect 15528 32388 15669 32416
rect 15528 32376 15534 32388
rect 15657 32385 15669 32388
rect 15703 32385 15715 32419
rect 15657 32379 15715 32385
rect 17127 32419 17185 32425
rect 17127 32385 17139 32419
rect 17173 32416 17185 32419
rect 18966 32416 18972 32428
rect 17173 32388 18972 32416
rect 17173 32385 17185 32388
rect 17127 32379 17185 32385
rect 18966 32376 18972 32388
rect 19024 32376 19030 32428
rect 19168 32425 19196 32456
rect 19978 32444 19984 32456
rect 20036 32444 20042 32496
rect 20070 32444 20076 32496
rect 20128 32444 20134 32496
rect 20548 32484 20576 32524
rect 20622 32512 20628 32564
rect 20680 32512 20686 32564
rect 20806 32512 20812 32564
rect 20864 32552 20870 32564
rect 21174 32552 21180 32564
rect 20864 32524 21180 32552
rect 20864 32512 20870 32524
rect 21174 32512 21180 32524
rect 21232 32512 21238 32564
rect 20548 32456 21312 32484
rect 19153 32419 19211 32425
rect 19153 32385 19165 32419
rect 19199 32385 19211 32419
rect 19153 32379 19211 32385
rect 19426 32376 19432 32428
rect 19484 32376 19490 32428
rect 19518 32376 19524 32428
rect 19576 32376 19582 32428
rect 19610 32376 19616 32428
rect 19668 32376 19674 32428
rect 19887 32419 19945 32425
rect 19887 32385 19899 32419
rect 19933 32416 19945 32419
rect 20088 32416 20116 32444
rect 19933 32388 20116 32416
rect 19933 32385 19945 32388
rect 19887 32379 19945 32385
rect 21174 32376 21180 32428
rect 21232 32376 21238 32428
rect 21284 32425 21312 32456
rect 22278 32444 22284 32496
rect 22336 32444 22342 32496
rect 21269 32419 21327 32425
rect 21269 32385 21281 32419
rect 21315 32385 21327 32419
rect 22296 32416 22324 32444
rect 21269 32379 21327 32385
rect 21376 32388 22324 32416
rect 7064 32320 7328 32348
rect 7064 32308 7070 32320
rect 8478 32308 8484 32360
rect 8536 32348 8542 32360
rect 8536 32320 8970 32348
rect 8536 32308 8542 32320
rect 13538 32308 13544 32360
rect 13596 32348 13602 32360
rect 13832 32348 13860 32376
rect 13596 32320 13860 32348
rect 13596 32308 13602 32320
rect 13906 32308 13912 32360
rect 13964 32348 13970 32360
rect 14001 32351 14059 32357
rect 14001 32348 14013 32351
rect 13964 32320 14013 32348
rect 13964 32308 13970 32320
rect 14001 32317 14013 32320
rect 14047 32317 14059 32351
rect 14001 32311 14059 32317
rect 16853 32351 16911 32357
rect 16853 32317 16865 32351
rect 16899 32317 16911 32351
rect 16853 32311 16911 32317
rect 5902 32240 5908 32292
rect 5960 32240 5966 32292
rect 8846 32240 8852 32292
rect 8904 32240 8910 32292
rect 10410 32240 10416 32292
rect 10468 32240 10474 32292
rect 10520 32252 11100 32280
rect 5920 32212 5948 32240
rect 4448 32184 5948 32212
rect 5994 32172 6000 32224
rect 6052 32212 6058 32224
rect 6638 32212 6644 32224
rect 6052 32184 6644 32212
rect 6052 32172 6058 32184
rect 6638 32172 6644 32184
rect 6696 32172 6702 32224
rect 8018 32172 8024 32224
rect 8076 32212 8082 32224
rect 8297 32215 8355 32221
rect 8297 32212 8309 32215
rect 8076 32184 8309 32212
rect 8076 32172 8082 32184
rect 8297 32181 8309 32184
rect 8343 32181 8355 32215
rect 8297 32175 8355 32181
rect 8570 32172 8576 32224
rect 8628 32212 8634 32224
rect 8864 32212 8892 32240
rect 8628 32184 8892 32212
rect 8628 32172 8634 32184
rect 10318 32172 10324 32224
rect 10376 32212 10382 32224
rect 10520 32212 10548 32252
rect 10376 32184 10548 32212
rect 10376 32172 10382 32184
rect 10686 32172 10692 32224
rect 10744 32212 10750 32224
rect 10965 32215 11023 32221
rect 10965 32212 10977 32215
rect 10744 32184 10977 32212
rect 10744 32172 10750 32184
rect 10965 32181 10977 32184
rect 11011 32181 11023 32215
rect 11072 32212 11100 32252
rect 11238 32240 11244 32292
rect 11296 32280 11302 32292
rect 11790 32280 11796 32292
rect 11296 32252 11796 32280
rect 11296 32240 11302 32252
rect 11790 32240 11796 32252
rect 11848 32240 11854 32292
rect 13278 32252 13766 32280
rect 13278 32212 13306 32252
rect 11072 32184 13306 32212
rect 10965 32175 11023 32181
rect 13630 32172 13636 32224
rect 13688 32172 13694 32224
rect 13738 32212 13766 32252
rect 15654 32240 15660 32292
rect 15712 32280 15718 32292
rect 15712 32252 16528 32280
rect 15712 32240 15718 32252
rect 16500 32224 16528 32252
rect 16868 32224 16896 32311
rect 18782 32308 18788 32360
rect 18840 32348 18846 32360
rect 19536 32348 19564 32376
rect 21376 32348 21404 32388
rect 18840 32320 19564 32348
rect 20272 32320 21404 32348
rect 18840 32308 18846 32320
rect 14366 32212 14372 32224
rect 13738 32184 14372 32212
rect 14366 32172 14372 32184
rect 14424 32172 14430 32224
rect 15010 32172 15016 32224
rect 15068 32172 15074 32224
rect 15746 32172 15752 32224
rect 15804 32212 15810 32224
rect 16206 32212 16212 32224
rect 15804 32184 16212 32212
rect 15804 32172 15810 32184
rect 16206 32172 16212 32184
rect 16264 32172 16270 32224
rect 16482 32172 16488 32224
rect 16540 32172 16546 32224
rect 16850 32172 16856 32224
rect 16908 32212 16914 32224
rect 17126 32212 17132 32224
rect 16908 32184 17132 32212
rect 16908 32172 16914 32184
rect 17126 32172 17132 32184
rect 17184 32212 17190 32224
rect 17954 32212 17960 32224
rect 17184 32184 17960 32212
rect 17184 32172 17190 32184
rect 17954 32172 17960 32184
rect 18012 32172 18018 32224
rect 19245 32215 19303 32221
rect 19245 32181 19257 32215
rect 19291 32212 19303 32215
rect 19702 32212 19708 32224
rect 19291 32184 19708 32212
rect 19291 32181 19303 32184
rect 19245 32175 19303 32181
rect 19702 32172 19708 32184
rect 19760 32172 19766 32224
rect 19886 32172 19892 32224
rect 19944 32212 19950 32224
rect 20272 32212 20300 32320
rect 21450 32308 21456 32360
rect 21508 32308 21514 32360
rect 22278 32308 22284 32360
rect 22336 32348 22342 32360
rect 22738 32348 22744 32360
rect 22336 32320 22744 32348
rect 22336 32308 22342 32320
rect 22738 32308 22744 32320
rect 22796 32308 22802 32360
rect 21468 32280 21496 32308
rect 20916 32252 21496 32280
rect 20916 32224 20944 32252
rect 22830 32240 22836 32292
rect 22888 32240 22894 32292
rect 19944 32184 20300 32212
rect 19944 32172 19950 32184
rect 20898 32172 20904 32224
rect 20956 32172 20962 32224
rect 20990 32172 20996 32224
rect 21048 32172 21054 32224
rect 21450 32172 21456 32224
rect 21508 32172 21514 32224
rect 1104 32122 21896 32144
rect 1104 32070 3549 32122
rect 3601 32070 3613 32122
rect 3665 32070 3677 32122
rect 3729 32070 3741 32122
rect 3793 32070 3805 32122
rect 3857 32070 8747 32122
rect 8799 32070 8811 32122
rect 8863 32070 8875 32122
rect 8927 32070 8939 32122
rect 8991 32070 9003 32122
rect 9055 32070 13945 32122
rect 13997 32070 14009 32122
rect 14061 32070 14073 32122
rect 14125 32070 14137 32122
rect 14189 32070 14201 32122
rect 14253 32070 19143 32122
rect 19195 32070 19207 32122
rect 19259 32070 19271 32122
rect 19323 32070 19335 32122
rect 19387 32070 19399 32122
rect 19451 32070 21896 32122
rect 22848 32088 22876 32240
rect 1104 32048 21896 32070
rect 22830 32036 22836 32088
rect 22888 32036 22894 32088
rect 2406 32008 2412 32020
rect 1964 31980 2412 32008
rect 1964 31881 1992 31980
rect 2406 31968 2412 31980
rect 2464 32008 2470 32020
rect 3326 32008 3332 32020
rect 2464 31980 3332 32008
rect 2464 31968 2470 31980
rect 3326 31968 3332 31980
rect 3384 31968 3390 32020
rect 5166 31968 5172 32020
rect 5224 31968 5230 32020
rect 5534 31968 5540 32020
rect 5592 32008 5598 32020
rect 6825 32011 6883 32017
rect 5592 31980 6776 32008
rect 5592 31968 5598 31980
rect 5184 31940 5212 31968
rect 6748 31940 6776 31980
rect 6825 31977 6837 32011
rect 6871 32008 6883 32011
rect 7190 32008 7196 32020
rect 6871 31980 7196 32008
rect 6871 31977 6883 31980
rect 6825 31971 6883 31977
rect 7190 31968 7196 31980
rect 7248 31968 7254 32020
rect 7576 31980 8294 32008
rect 7576 31940 7604 31980
rect 2056 31912 2542 31940
rect 5184 31912 5672 31940
rect 6748 31912 7604 31940
rect 1949 31875 2007 31881
rect 1949 31841 1961 31875
rect 1995 31841 2007 31875
rect 1949 31835 2007 31841
rect 1394 31764 1400 31816
rect 1452 31764 1458 31816
rect 1762 31764 1768 31816
rect 1820 31764 1826 31816
rect 1854 31764 1860 31816
rect 1912 31804 1918 31816
rect 2056 31804 2084 31912
rect 2406 31832 2412 31884
rect 2464 31832 2470 31884
rect 2514 31872 2542 31912
rect 2514 31844 2728 31872
rect 2700 31813 2728 31844
rect 2774 31832 2780 31884
rect 2832 31881 2838 31884
rect 2832 31875 2860 31881
rect 2848 31841 2860 31875
rect 2832 31835 2860 31841
rect 3605 31875 3663 31881
rect 3605 31841 3617 31875
rect 3651 31872 3663 31875
rect 3651 31844 4200 31872
rect 3651 31841 3663 31844
rect 3605 31835 3663 31841
rect 2832 31832 2838 31835
rect 1912 31776 2084 31804
rect 2685 31807 2743 31813
rect 1912 31764 1918 31776
rect 2685 31773 2697 31807
rect 2731 31773 2743 31807
rect 2685 31767 2743 31773
rect 2958 31764 2964 31816
rect 3016 31764 3022 31816
rect 3786 31764 3792 31816
rect 3844 31764 3850 31816
rect 4062 31764 4068 31816
rect 4120 31764 4126 31816
rect 4172 31804 4200 31844
rect 4890 31832 4896 31884
rect 4948 31872 4954 31884
rect 4985 31875 5043 31881
rect 4985 31872 4997 31875
rect 4948 31844 4997 31872
rect 4948 31832 4954 31844
rect 4985 31841 4997 31844
rect 5031 31841 5043 31875
rect 4985 31835 5043 31841
rect 5258 31832 5264 31884
rect 5316 31832 5322 31884
rect 5644 31881 5672 31912
rect 5629 31875 5687 31881
rect 5629 31841 5641 31875
rect 5675 31841 5687 31875
rect 5629 31835 5687 31841
rect 5718 31832 5724 31884
rect 5776 31872 5782 31884
rect 5905 31875 5963 31881
rect 5905 31872 5917 31875
rect 5776 31844 5917 31872
rect 5776 31832 5782 31844
rect 5905 31841 5917 31844
rect 5951 31841 5963 31875
rect 5905 31835 5963 31841
rect 5994 31832 6000 31884
rect 6052 31881 6058 31884
rect 6052 31875 6080 31881
rect 6068 31841 6080 31875
rect 6052 31835 6080 31841
rect 6052 31832 6058 31835
rect 7374 31832 7380 31884
rect 7432 31872 7438 31884
rect 7469 31875 7527 31881
rect 7469 31872 7481 31875
rect 7432 31844 7481 31872
rect 7432 31832 7438 31844
rect 7469 31841 7481 31844
rect 7515 31841 7527 31875
rect 8266 31872 8294 31980
rect 10042 31968 10048 32020
rect 10100 32008 10106 32020
rect 10100 31980 10456 32008
rect 10100 31968 10106 31980
rect 10428 31949 10456 31980
rect 10870 31968 10876 32020
rect 10928 32008 10934 32020
rect 15010 32008 15016 32020
rect 10928 31980 11652 32008
rect 10928 31968 10934 31980
rect 10413 31943 10471 31949
rect 10413 31909 10425 31943
rect 10459 31909 10471 31943
rect 10413 31903 10471 31909
rect 9582 31872 9588 31884
rect 8266 31844 9588 31872
rect 7469 31835 7527 31841
rect 4430 31804 4436 31816
rect 4172 31776 4436 31804
rect 4430 31764 4436 31776
rect 4488 31764 4494 31816
rect 4522 31764 4528 31816
rect 4580 31764 4586 31816
rect 4706 31764 4712 31816
rect 4764 31764 4770 31816
rect 5169 31807 5227 31813
rect 5169 31773 5181 31807
rect 5215 31804 5227 31807
rect 5276 31804 5304 31832
rect 5215 31776 5304 31804
rect 5215 31773 5227 31776
rect 5169 31767 5227 31773
rect 4540 31736 4568 31764
rect 5184 31736 5212 31767
rect 6178 31764 6184 31816
rect 6236 31764 6242 31816
rect 4540 31708 5212 31736
rect 7484 31736 7512 31835
rect 9582 31832 9588 31844
rect 9640 31872 9646 31884
rect 9769 31875 9827 31881
rect 9769 31872 9781 31875
rect 9640 31844 9781 31872
rect 9640 31832 9646 31844
rect 9769 31841 9781 31844
rect 9815 31872 9827 31875
rect 10318 31872 10324 31884
rect 9815 31844 10324 31872
rect 9815 31841 9827 31844
rect 9769 31835 9827 31841
rect 10318 31832 10324 31844
rect 10376 31832 10382 31884
rect 10686 31832 10692 31884
rect 10744 31832 10750 31884
rect 10827 31875 10885 31881
rect 10827 31841 10839 31875
rect 10873 31872 10885 31875
rect 11146 31872 11152 31884
rect 10873 31844 11152 31872
rect 10873 31841 10885 31844
rect 10827 31835 10885 31841
rect 11146 31832 11152 31844
rect 11204 31832 11210 31884
rect 7743 31807 7801 31813
rect 7743 31773 7755 31807
rect 7789 31804 7801 31807
rect 8478 31804 8484 31816
rect 7789 31776 8484 31804
rect 7789 31773 7801 31776
rect 7743 31767 7801 31773
rect 8478 31764 8484 31776
rect 8536 31764 8542 31816
rect 9950 31764 9956 31816
rect 10008 31764 10014 31816
rect 10962 31764 10968 31816
rect 11020 31764 11026 31816
rect 11624 31813 11652 31980
rect 14752 31980 15016 32008
rect 13817 31943 13875 31949
rect 13817 31909 13829 31943
rect 13863 31940 13875 31943
rect 13906 31940 13912 31952
rect 13863 31912 13912 31940
rect 13863 31909 13875 31912
rect 13817 31903 13875 31909
rect 13906 31900 13912 31912
rect 13964 31900 13970 31952
rect 14752 31949 14780 31980
rect 15010 31968 15016 31980
rect 15068 31968 15074 32020
rect 16482 31968 16488 32020
rect 16540 32008 16546 32020
rect 17037 32011 17095 32017
rect 17037 32008 17049 32011
rect 16540 31980 17049 32008
rect 16540 31968 16546 31980
rect 17037 31977 17049 31980
rect 17083 31977 17095 32011
rect 18874 32008 18880 32020
rect 17037 31971 17095 31977
rect 17926 31980 18880 32008
rect 14737 31943 14795 31949
rect 14737 31909 14749 31943
rect 14783 31909 14795 31943
rect 14737 31903 14795 31909
rect 15930 31900 15936 31952
rect 15988 31940 15994 31952
rect 15988 31912 16068 31940
rect 15988 31900 15994 31912
rect 13354 31832 13360 31884
rect 13412 31832 13418 31884
rect 13630 31832 13636 31884
rect 13688 31832 13694 31884
rect 14274 31872 14280 31884
rect 14016 31844 14280 31872
rect 11609 31807 11667 31813
rect 11609 31773 11621 31807
rect 11655 31804 11667 31807
rect 12618 31804 12624 31816
rect 11655 31776 12624 31804
rect 11655 31773 11667 31776
rect 11609 31767 11667 31773
rect 12618 31764 12624 31776
rect 12676 31804 12682 31816
rect 12805 31807 12863 31813
rect 12805 31804 12817 31807
rect 12676 31776 12817 31804
rect 12676 31764 12682 31776
rect 12805 31773 12817 31776
rect 12851 31773 12863 31807
rect 12805 31767 12863 31773
rect 12897 31807 12955 31813
rect 12897 31773 12909 31807
rect 12943 31804 12955 31807
rect 13648 31804 13676 31832
rect 12943 31776 13676 31804
rect 12943 31773 12955 31776
rect 12897 31767 12955 31773
rect 7650 31736 7656 31748
rect 7484 31708 7656 31736
rect 7650 31696 7656 31708
rect 7708 31696 7714 31748
rect 7926 31696 7932 31748
rect 7984 31736 7990 31748
rect 9306 31736 9312 31748
rect 7984 31708 9312 31736
rect 7984 31696 7990 31708
rect 9306 31696 9312 31708
rect 9364 31736 9370 31748
rect 13265 31739 13323 31745
rect 9364 31708 9996 31736
rect 9364 31696 9370 31708
rect 1581 31671 1639 31677
rect 1581 31637 1593 31671
rect 1627 31668 1639 31671
rect 1854 31668 1860 31680
rect 1627 31640 1860 31668
rect 1627 31637 1639 31640
rect 1581 31631 1639 31637
rect 1854 31628 1860 31640
rect 1912 31668 1918 31680
rect 4154 31668 4160 31680
rect 1912 31640 4160 31668
rect 1912 31628 1918 31640
rect 4154 31628 4160 31640
rect 4212 31628 4218 31680
rect 4246 31628 4252 31680
rect 4304 31668 4310 31680
rect 4525 31671 4583 31677
rect 4525 31668 4537 31671
rect 4304 31640 4537 31668
rect 4304 31628 4310 31640
rect 4525 31637 4537 31640
rect 4571 31637 4583 31671
rect 4525 31631 4583 31637
rect 4706 31628 4712 31680
rect 4764 31668 4770 31680
rect 4890 31668 4896 31680
rect 4764 31640 4896 31668
rect 4764 31628 4770 31640
rect 4890 31628 4896 31640
rect 4948 31668 4954 31680
rect 5350 31668 5356 31680
rect 4948 31640 5356 31668
rect 4948 31628 4954 31640
rect 5350 31628 5356 31640
rect 5408 31628 5414 31680
rect 5994 31628 6000 31680
rect 6052 31668 6058 31680
rect 6270 31668 6276 31680
rect 6052 31640 6276 31668
rect 6052 31628 6058 31640
rect 6270 31628 6276 31640
rect 6328 31628 6334 31680
rect 7282 31628 7288 31680
rect 7340 31668 7346 31680
rect 8202 31668 8208 31680
rect 7340 31640 8208 31668
rect 7340 31628 7346 31640
rect 8202 31628 8208 31640
rect 8260 31628 8266 31680
rect 8478 31628 8484 31680
rect 8536 31628 8542 31680
rect 8570 31628 8576 31680
rect 8628 31668 8634 31680
rect 9674 31668 9680 31680
rect 8628 31640 9680 31668
rect 8628 31628 8634 31640
rect 9674 31628 9680 31640
rect 9732 31628 9738 31680
rect 9968 31668 9996 31708
rect 13265 31705 13277 31739
rect 13311 31736 13323 31739
rect 13354 31736 13360 31748
rect 13311 31708 13360 31736
rect 13311 31705 13323 31708
rect 13265 31699 13323 31705
rect 13354 31696 13360 31708
rect 13412 31696 13418 31748
rect 13538 31696 13544 31748
rect 13596 31736 13602 31748
rect 13633 31739 13691 31745
rect 13633 31736 13645 31739
rect 13596 31708 13645 31736
rect 13596 31696 13602 31708
rect 13633 31705 13645 31708
rect 13679 31736 13691 31739
rect 14016 31736 14044 31844
rect 14274 31832 14280 31844
rect 14332 31832 14338 31884
rect 15013 31875 15071 31881
rect 15013 31872 15025 31875
rect 14382 31844 15025 31872
rect 14090 31764 14096 31816
rect 14148 31764 14154 31816
rect 14382 31804 14410 31844
rect 15013 31841 15025 31844
rect 15059 31841 15071 31875
rect 15013 31835 15071 31841
rect 15289 31875 15347 31881
rect 15289 31841 15301 31875
rect 15335 31872 15347 31875
rect 15654 31872 15660 31884
rect 15335 31844 15660 31872
rect 15335 31841 15347 31844
rect 15289 31835 15347 31841
rect 15654 31832 15660 31844
rect 15712 31832 15718 31884
rect 16040 31881 16068 31912
rect 16025 31875 16083 31881
rect 16025 31841 16037 31875
rect 16071 31841 16083 31875
rect 16025 31835 16083 31841
rect 17218 31832 17224 31884
rect 17276 31872 17282 31884
rect 17926 31872 17954 31980
rect 18874 31968 18880 31980
rect 18932 31968 18938 32020
rect 19245 32011 19303 32017
rect 19245 31977 19257 32011
rect 19291 32008 19303 32011
rect 19886 32008 19892 32020
rect 19291 31980 19892 32008
rect 19291 31977 19303 31980
rect 19245 31971 19303 31977
rect 19886 31968 19892 31980
rect 19944 31968 19950 32020
rect 19978 31968 19984 32020
rect 20036 31968 20042 32020
rect 20257 32011 20315 32017
rect 20257 31977 20269 32011
rect 20303 32008 20315 32011
rect 21542 32008 21548 32020
rect 20303 31980 21548 32008
rect 20303 31977 20315 31980
rect 20257 31971 20315 31977
rect 21542 31968 21548 31980
rect 21600 31968 21606 32020
rect 18141 31943 18199 31949
rect 18141 31909 18153 31943
rect 18187 31940 18199 31943
rect 18693 31943 18751 31949
rect 18187 31912 18644 31940
rect 18187 31909 18199 31912
rect 18141 31903 18199 31909
rect 17276 31844 17954 31872
rect 17276 31832 17282 31844
rect 14200 31776 14410 31804
rect 13679 31708 14044 31736
rect 13679 31705 13691 31708
rect 13633 31699 13691 31705
rect 10226 31668 10232 31680
rect 9968 31640 10232 31668
rect 10226 31628 10232 31640
rect 10284 31628 10290 31680
rect 10778 31628 10784 31680
rect 10836 31668 10842 31680
rect 12158 31668 12164 31680
rect 10836 31640 12164 31668
rect 10836 31628 10842 31640
rect 12158 31628 12164 31640
rect 12216 31668 12222 31680
rect 12529 31671 12587 31677
rect 12529 31668 12541 31671
rect 12216 31640 12541 31668
rect 12216 31628 12222 31640
rect 12529 31637 12541 31640
rect 12575 31668 12587 31671
rect 14200 31668 14228 31776
rect 15102 31764 15108 31816
rect 15160 31813 15166 31816
rect 15160 31807 15188 31813
rect 15176 31773 15188 31807
rect 15160 31767 15188 31773
rect 15933 31807 15991 31813
rect 15933 31773 15945 31807
rect 15979 31804 15991 31807
rect 15979 31776 16013 31804
rect 15979 31773 15991 31776
rect 15933 31767 15991 31773
rect 15160 31764 15166 31767
rect 15948 31736 15976 31767
rect 16206 31764 16212 31816
rect 16264 31804 16270 31816
rect 16299 31807 16357 31813
rect 16299 31804 16311 31807
rect 16264 31776 16311 31804
rect 16264 31764 16270 31776
rect 16299 31773 16311 31776
rect 16345 31773 16357 31807
rect 16942 31804 16948 31816
rect 16299 31767 16357 31773
rect 16408 31776 16948 31804
rect 16408 31736 16436 31776
rect 16942 31764 16948 31776
rect 17000 31764 17006 31816
rect 18322 31764 18328 31816
rect 18380 31764 18386 31816
rect 18616 31813 18644 31912
rect 18693 31909 18705 31943
rect 18739 31909 18751 31943
rect 18693 31903 18751 31909
rect 19613 31943 19671 31949
rect 19613 31909 19625 31943
rect 19659 31940 19671 31943
rect 20898 31940 20904 31952
rect 19659 31912 20904 31940
rect 19659 31909 19671 31912
rect 19613 31903 19671 31909
rect 18708 31872 18736 31903
rect 20898 31900 20904 31912
rect 20956 31900 20962 31952
rect 18708 31844 19472 31872
rect 18417 31807 18475 31813
rect 18417 31773 18429 31807
rect 18463 31773 18475 31807
rect 18417 31767 18475 31773
rect 18601 31807 18659 31813
rect 18601 31773 18613 31807
rect 18647 31773 18659 31807
rect 18601 31767 18659 31773
rect 18877 31807 18935 31813
rect 18877 31773 18889 31807
rect 18923 31804 18935 31807
rect 18966 31804 18972 31816
rect 18923 31776 18972 31804
rect 18923 31773 18935 31776
rect 18877 31767 18935 31773
rect 18432 31736 18460 31767
rect 18966 31764 18972 31776
rect 19024 31764 19030 31816
rect 19444 31813 19472 31844
rect 19702 31832 19708 31884
rect 19760 31872 19766 31884
rect 19760 31844 20208 31872
rect 19760 31832 19766 31844
rect 19429 31807 19487 31813
rect 19429 31773 19441 31807
rect 19475 31773 19487 31807
rect 19429 31767 19487 31773
rect 19794 31764 19800 31816
rect 19852 31764 19858 31816
rect 20180 31813 20208 31844
rect 20714 31832 20720 31884
rect 20772 31832 20778 31884
rect 22940 31816 22968 32864
rect 20165 31807 20223 31813
rect 20165 31773 20177 31807
rect 20211 31773 20223 31807
rect 20165 31767 20223 31773
rect 20438 31764 20444 31816
rect 20496 31764 20502 31816
rect 20625 31807 20683 31813
rect 20625 31773 20637 31807
rect 20671 31773 20683 31807
rect 20625 31767 20683 31773
rect 15948 31708 16436 31736
rect 18156 31708 18460 31736
rect 18156 31680 18184 31708
rect 19702 31696 19708 31748
rect 19760 31736 19766 31748
rect 20640 31736 20668 31767
rect 21082 31764 21088 31816
rect 21140 31804 21146 31816
rect 21177 31807 21235 31813
rect 21177 31804 21189 31807
rect 21140 31776 21189 31804
rect 21140 31764 21146 31776
rect 21177 31773 21189 31776
rect 21223 31773 21235 31807
rect 21177 31767 21235 31773
rect 22554 31736 22560 31766
rect 19760 31708 20668 31736
rect 20732 31714 22560 31736
rect 22612 31714 22618 31766
rect 22922 31764 22928 31816
rect 22980 31764 22986 31816
rect 20732 31708 22600 31714
rect 19760 31696 19766 31708
rect 12575 31640 14228 31668
rect 12575 31637 12587 31640
rect 12529 31631 12587 31637
rect 14826 31628 14832 31680
rect 14884 31668 14890 31680
rect 15562 31668 15568 31680
rect 14884 31640 15568 31668
rect 14884 31628 14890 31640
rect 15562 31628 15568 31640
rect 15620 31628 15626 31680
rect 18138 31628 18144 31680
rect 18196 31628 18202 31680
rect 18506 31628 18512 31680
rect 18564 31628 18570 31680
rect 20070 31628 20076 31680
rect 20128 31668 20134 31680
rect 20732 31668 20760 31708
rect 20128 31640 20760 31668
rect 21453 31671 21511 31677
rect 20128 31628 20134 31640
rect 21453 31637 21465 31671
rect 21499 31668 21511 31671
rect 22186 31668 22192 31680
rect 21499 31640 22192 31668
rect 21499 31637 21511 31640
rect 21453 31631 21511 31637
rect 22186 31628 22192 31640
rect 22244 31628 22250 31680
rect 1104 31578 22056 31600
rect 1104 31526 6148 31578
rect 6200 31526 6212 31578
rect 6264 31526 6276 31578
rect 6328 31526 6340 31578
rect 6392 31526 6404 31578
rect 6456 31526 11346 31578
rect 11398 31526 11410 31578
rect 11462 31526 11474 31578
rect 11526 31526 11538 31578
rect 11590 31526 11602 31578
rect 11654 31526 16544 31578
rect 16596 31526 16608 31578
rect 16660 31526 16672 31578
rect 16724 31526 16736 31578
rect 16788 31526 16800 31578
rect 16852 31526 21742 31578
rect 21794 31526 21806 31578
rect 21858 31526 21870 31578
rect 21922 31526 21934 31578
rect 21986 31526 21998 31578
rect 22050 31526 22056 31578
rect 1104 31504 22056 31526
rect 2406 31424 2412 31476
rect 2464 31424 2470 31476
rect 2774 31424 2780 31476
rect 2832 31464 2838 31476
rect 2832 31436 3280 31464
rect 2832 31424 2838 31436
rect 1302 31356 1308 31408
rect 1360 31396 1366 31408
rect 1486 31396 1492 31408
rect 1360 31368 1492 31396
rect 1360 31356 1366 31368
rect 1412 31337 1440 31368
rect 1486 31356 1492 31368
rect 1544 31356 1550 31408
rect 2130 31356 2136 31408
rect 2188 31396 2194 31408
rect 2590 31396 2596 31408
rect 2188 31368 2596 31396
rect 2188 31356 2194 31368
rect 2590 31356 2596 31368
rect 2648 31396 2654 31408
rect 2648 31368 3154 31396
rect 2648 31356 2654 31368
rect 1397 31331 1455 31337
rect 1397 31297 1409 31331
rect 1443 31297 1455 31331
rect 1397 31291 1455 31297
rect 1671 31331 1729 31337
rect 1671 31297 1683 31331
rect 1717 31328 1729 31331
rect 2038 31328 2044 31340
rect 1717 31300 2044 31328
rect 1717 31297 1729 31300
rect 1671 31291 1729 31297
rect 2038 31288 2044 31300
rect 2096 31328 2102 31340
rect 2498 31328 2504 31340
rect 2096 31300 2504 31328
rect 2096 31288 2102 31300
rect 2498 31288 2504 31300
rect 2556 31288 2562 31340
rect 2682 31288 2688 31340
rect 2740 31328 2746 31340
rect 2774 31328 2780 31340
rect 2740 31300 2780 31328
rect 2740 31288 2746 31300
rect 2774 31288 2780 31300
rect 2832 31288 2838 31340
rect 3126 31337 3154 31368
rect 3111 31331 3169 31337
rect 3111 31297 3123 31331
rect 3157 31297 3169 31331
rect 3252 31328 3280 31436
rect 3326 31424 3332 31476
rect 3384 31464 3390 31476
rect 6454 31464 6460 31476
rect 3384 31436 6460 31464
rect 3384 31424 3390 31436
rect 6454 31424 6460 31436
rect 6512 31424 6518 31476
rect 7374 31424 7380 31476
rect 7432 31464 7438 31476
rect 10781 31467 10839 31473
rect 7432 31436 10732 31464
rect 7432 31424 7438 31436
rect 6730 31396 6736 31408
rect 4908 31368 6736 31396
rect 4908 31337 4936 31368
rect 6730 31356 6736 31368
rect 6788 31396 6794 31408
rect 9125 31399 9183 31405
rect 6788 31368 7052 31396
rect 6788 31356 6794 31368
rect 7024 31340 7052 31368
rect 9125 31365 9137 31399
rect 9171 31396 9183 31399
rect 10410 31396 10416 31408
rect 9171 31368 10416 31396
rect 9171 31365 9183 31368
rect 9125 31359 9183 31365
rect 10410 31356 10416 31368
rect 10468 31356 10474 31408
rect 10704 31396 10732 31436
rect 10781 31433 10793 31467
rect 10827 31464 10839 31467
rect 10962 31464 10968 31476
rect 10827 31436 10968 31464
rect 10827 31433 10839 31436
rect 10781 31427 10839 31433
rect 10962 31424 10968 31436
rect 11020 31424 11026 31476
rect 16114 31464 16120 31476
rect 11898 31436 16120 31464
rect 10704 31368 11742 31396
rect 11714 31358 11742 31368
rect 11775 31361 11833 31367
rect 11775 31358 11787 31361
rect 4249 31331 4307 31337
rect 4249 31328 4261 31331
rect 3252 31300 4261 31328
rect 3111 31291 3169 31297
rect 4249 31297 4261 31300
rect 4295 31297 4307 31331
rect 4249 31291 4307 31297
rect 4893 31331 4951 31337
rect 4893 31297 4905 31331
rect 4939 31297 4951 31331
rect 4893 31291 4951 31297
rect 5167 31331 5225 31337
rect 5167 31297 5179 31331
rect 5213 31328 5225 31331
rect 5258 31328 5264 31340
rect 5213 31300 5264 31328
rect 5213 31297 5225 31300
rect 5167 31291 5225 31297
rect 2866 31220 2872 31272
rect 2924 31220 2930 31272
rect 4430 31220 4436 31272
rect 4488 31220 4494 31272
rect 4908 31192 4936 31291
rect 5258 31288 5264 31300
rect 5316 31288 5322 31340
rect 5718 31288 5724 31340
rect 5776 31328 5782 31340
rect 5902 31328 5908 31340
rect 5776 31300 5908 31328
rect 5776 31288 5782 31300
rect 5902 31288 5908 31300
rect 5960 31288 5966 31340
rect 6365 31331 6423 31337
rect 6365 31297 6377 31331
rect 6411 31297 6423 31331
rect 6365 31291 6423 31297
rect 6380 31192 6408 31291
rect 6454 31288 6460 31340
rect 6512 31288 6518 31340
rect 7006 31288 7012 31340
rect 7064 31288 7070 31340
rect 7190 31288 7196 31340
rect 7248 31328 7254 31340
rect 7469 31331 7527 31337
rect 7469 31328 7481 31331
rect 7248 31300 7481 31328
rect 7248 31288 7254 31300
rect 7469 31297 7481 31300
rect 7515 31297 7527 31331
rect 7469 31291 7527 31297
rect 8478 31288 8484 31340
rect 8536 31288 8542 31340
rect 9769 31331 9827 31337
rect 9769 31297 9781 31331
rect 9815 31297 9827 31331
rect 10042 31328 10048 31340
rect 10003 31300 10048 31328
rect 9769 31291 9827 31297
rect 6472 31260 6500 31288
rect 6822 31260 6828 31272
rect 6472 31232 6828 31260
rect 6822 31220 6828 31232
rect 6880 31260 6886 31272
rect 7285 31263 7343 31269
rect 7285 31260 7297 31263
rect 6880 31232 7297 31260
rect 6880 31220 6886 31232
rect 7285 31229 7297 31232
rect 7331 31229 7343 31263
rect 7285 31223 7343 31229
rect 7926 31220 7932 31272
rect 7984 31220 7990 31272
rect 8202 31220 8208 31272
rect 8260 31220 8266 31272
rect 8343 31263 8401 31269
rect 8343 31229 8355 31263
rect 8389 31260 8401 31263
rect 8389 31232 8892 31260
rect 8389 31229 8401 31232
rect 8343 31223 8401 31229
rect 7558 31192 7564 31204
rect 3526 31164 4936 31192
rect 5552 31164 6408 31192
rect 6472 31164 7564 31192
rect 1486 31084 1492 31136
rect 1544 31124 1550 31136
rect 3526 31124 3554 31164
rect 1544 31096 3554 31124
rect 1544 31084 1550 31096
rect 3878 31084 3884 31136
rect 3936 31084 3942 31136
rect 4062 31084 4068 31136
rect 4120 31124 4126 31136
rect 5552 31124 5580 31164
rect 4120 31096 5580 31124
rect 4120 31084 4126 31096
rect 5902 31084 5908 31136
rect 5960 31084 5966 31136
rect 6086 31084 6092 31136
rect 6144 31124 6150 31136
rect 6472 31124 6500 31164
rect 7558 31152 7564 31164
rect 7616 31152 7622 31204
rect 6144 31096 6500 31124
rect 6549 31127 6607 31133
rect 6144 31084 6150 31096
rect 6549 31093 6561 31127
rect 6595 31124 6607 31127
rect 8018 31124 8024 31136
rect 6595 31096 8024 31124
rect 6595 31093 6607 31096
rect 6549 31087 6607 31093
rect 8018 31084 8024 31096
rect 8076 31084 8082 31136
rect 8478 31084 8484 31136
rect 8536 31124 8542 31136
rect 8864 31124 8892 31232
rect 9674 31220 9680 31272
rect 9732 31260 9738 31272
rect 9784 31260 9812 31291
rect 10042 31288 10048 31300
rect 10100 31288 10106 31340
rect 11238 31288 11244 31340
rect 11296 31288 11302 31340
rect 11714 31330 11787 31358
rect 11775 31327 11787 31330
rect 11821 31358 11833 31361
rect 11898 31358 11926 31436
rect 16114 31424 16120 31436
rect 16172 31464 16178 31476
rect 17218 31464 17224 31476
rect 16172 31436 17224 31464
rect 16172 31424 16178 31436
rect 17218 31424 17224 31436
rect 17276 31424 17282 31476
rect 18049 31467 18107 31473
rect 18049 31433 18061 31467
rect 18095 31464 18107 31467
rect 18322 31464 18328 31476
rect 18095 31436 18328 31464
rect 18095 31433 18107 31436
rect 18049 31427 18107 31433
rect 18322 31424 18328 31436
rect 18380 31424 18386 31476
rect 19613 31467 19671 31473
rect 18430 31436 19334 31464
rect 11821 31330 11926 31358
rect 13556 31368 14854 31396
rect 13556 31340 13584 31368
rect 12897 31331 12955 31337
rect 11821 31327 11833 31330
rect 12897 31328 12909 31331
rect 11775 31321 11833 31327
rect 12176 31300 12909 31328
rect 9732 31232 9812 31260
rect 9732 31220 9738 31232
rect 10870 31220 10876 31272
rect 10928 31260 10934 31272
rect 11256 31260 11284 31288
rect 11517 31263 11575 31269
rect 11517 31260 11529 31263
rect 10928 31232 11529 31260
rect 10928 31220 10934 31232
rect 11517 31229 11529 31232
rect 11563 31229 11575 31263
rect 11517 31223 11575 31229
rect 8536 31096 8892 31124
rect 8536 31084 8542 31096
rect 11882 31084 11888 31136
rect 11940 31124 11946 31136
rect 12176 31124 12204 31300
rect 12897 31297 12909 31300
rect 12943 31297 12955 31331
rect 12897 31291 12955 31297
rect 13078 31288 13084 31340
rect 13136 31288 13142 31340
rect 13538 31288 13544 31340
rect 13596 31288 13602 31340
rect 14703 31331 14761 31337
rect 14703 31328 14715 31331
rect 13648 31300 14715 31328
rect 12250 31220 12256 31272
rect 12308 31260 12314 31272
rect 13648 31260 13676 31300
rect 14703 31297 14715 31300
rect 14749 31297 14761 31331
rect 14826 31328 14854 31368
rect 15286 31356 15292 31408
rect 15344 31396 15350 31408
rect 18430 31396 18458 31436
rect 15344 31368 18458 31396
rect 15344 31356 15350 31368
rect 18598 31356 18604 31408
rect 18656 31356 18662 31408
rect 19306 31396 19334 31436
rect 19613 31433 19625 31467
rect 19659 31464 19671 31467
rect 19702 31464 19708 31476
rect 19659 31436 19708 31464
rect 19659 31433 19671 31436
rect 19613 31427 19671 31433
rect 19702 31424 19708 31436
rect 19760 31424 19766 31476
rect 19889 31467 19947 31473
rect 19889 31433 19901 31467
rect 19935 31464 19947 31467
rect 20438 31464 20444 31476
rect 19935 31436 20444 31464
rect 19935 31433 19947 31436
rect 19889 31427 19947 31433
rect 20438 31424 20444 31436
rect 20496 31424 20502 31476
rect 21174 31424 21180 31476
rect 21232 31424 21238 31476
rect 19306 31368 20116 31396
rect 14826 31300 16252 31328
rect 14703 31291 14761 31297
rect 12308 31232 13676 31260
rect 14461 31263 14519 31269
rect 12308 31220 12314 31232
rect 14461 31229 14473 31263
rect 14507 31229 14519 31263
rect 14461 31223 14519 31229
rect 14476 31192 14504 31223
rect 15194 31220 15200 31272
rect 15252 31220 15258 31272
rect 16224 31260 16252 31300
rect 16298 31288 16304 31340
rect 16356 31328 16362 31340
rect 16669 31331 16727 31337
rect 16669 31328 16681 31331
rect 16356 31300 16681 31328
rect 16356 31288 16362 31300
rect 16669 31297 16681 31300
rect 16715 31297 16727 31331
rect 16925 31331 16983 31337
rect 16925 31328 16937 31331
rect 16669 31291 16727 31297
rect 16767 31300 16937 31328
rect 16767 31260 16795 31300
rect 16925 31297 16937 31300
rect 16971 31328 16983 31331
rect 17218 31328 17224 31340
rect 16971 31300 17224 31328
rect 16971 31297 16983 31300
rect 16925 31291 16983 31297
rect 17218 31288 17224 31300
rect 17276 31288 17282 31340
rect 17954 31288 17960 31340
rect 18012 31328 18018 31340
rect 18141 31331 18199 31337
rect 18141 31328 18153 31331
rect 18012 31300 18153 31328
rect 18012 31288 18018 31300
rect 18141 31297 18153 31300
rect 18187 31297 18199 31331
rect 18141 31291 18199 31297
rect 18415 31331 18473 31337
rect 18415 31297 18427 31331
rect 18461 31326 18473 31331
rect 18616 31328 18644 31356
rect 18598 31326 18644 31328
rect 18461 31300 18644 31326
rect 18461 31298 18626 31300
rect 18461 31297 18473 31298
rect 18415 31291 18473 31297
rect 18874 31288 18880 31340
rect 18932 31328 18938 31340
rect 19702 31328 19708 31340
rect 18932 31300 19708 31328
rect 18932 31288 18938 31300
rect 19702 31288 19708 31300
rect 19760 31328 19766 31340
rect 20088 31337 20116 31368
rect 19797 31331 19855 31337
rect 19797 31328 19809 31331
rect 19760 31300 19809 31328
rect 19760 31288 19766 31300
rect 19797 31297 19809 31300
rect 19843 31297 19855 31331
rect 19797 31291 19855 31297
rect 20073 31331 20131 31337
rect 20073 31297 20085 31331
rect 20119 31297 20131 31331
rect 20073 31291 20131 31297
rect 20533 31331 20591 31337
rect 20533 31297 20545 31331
rect 20579 31297 20591 31331
rect 20533 31291 20591 31297
rect 16224 31232 16795 31260
rect 18966 31220 18972 31272
rect 19024 31260 19030 31272
rect 20548 31260 20576 31291
rect 20622 31288 20628 31340
rect 20680 31328 20686 31340
rect 20993 31331 21051 31337
rect 20993 31328 21005 31331
rect 20680 31300 21005 31328
rect 20680 31288 20686 31300
rect 20993 31297 21005 31300
rect 21039 31297 21051 31331
rect 20993 31291 21051 31297
rect 19024 31232 20576 31260
rect 19024 31220 19030 31232
rect 14476 31164 14565 31192
rect 12529 31127 12587 31133
rect 12529 31124 12541 31127
rect 11940 31096 12541 31124
rect 11940 31084 11946 31096
rect 12529 31093 12541 31096
rect 12575 31093 12587 31127
rect 12529 31087 12587 31093
rect 12986 31084 12992 31136
rect 13044 31084 13050 31136
rect 14537 31124 14565 31164
rect 14734 31124 14740 31136
rect 14537 31096 14740 31124
rect 14734 31084 14740 31096
rect 14792 31124 14798 31136
rect 15212 31124 15240 31220
rect 18138 31152 18144 31204
rect 18196 31152 18202 31204
rect 20349 31195 20407 31201
rect 20349 31161 20361 31195
rect 20395 31192 20407 31195
rect 21192 31192 21220 31424
rect 21266 31288 21272 31340
rect 21324 31288 21330 31340
rect 20395 31164 21220 31192
rect 20395 31161 20407 31164
rect 20349 31155 20407 31161
rect 14792 31096 15240 31124
rect 14792 31084 14798 31096
rect 15470 31084 15476 31136
rect 15528 31084 15534 31136
rect 18156 31124 18184 31152
rect 19153 31127 19211 31133
rect 19153 31124 19165 31127
rect 18156 31096 19165 31124
rect 19153 31093 19165 31096
rect 19199 31093 19211 31127
rect 19153 31087 19211 31093
rect 20809 31127 20867 31133
rect 20809 31093 20821 31127
rect 20855 31124 20867 31127
rect 21082 31124 21088 31136
rect 20855 31096 21088 31124
rect 20855 31093 20867 31096
rect 20809 31087 20867 31093
rect 21082 31084 21088 31096
rect 21140 31084 21146 31136
rect 21450 31084 21456 31136
rect 21508 31084 21514 31136
rect 1104 31034 21896 31056
rect 1104 30982 3549 31034
rect 3601 30982 3613 31034
rect 3665 30982 3677 31034
rect 3729 30982 3741 31034
rect 3793 30982 3805 31034
rect 3857 30982 8747 31034
rect 8799 30982 8811 31034
rect 8863 30982 8875 31034
rect 8927 30982 8939 31034
rect 8991 30982 9003 31034
rect 9055 30982 13945 31034
rect 13997 30982 14009 31034
rect 14061 30982 14073 31034
rect 14125 30982 14137 31034
rect 14189 30982 14201 31034
rect 14253 30982 19143 31034
rect 19195 30982 19207 31034
rect 19259 30982 19271 31034
rect 19323 30982 19335 31034
rect 19387 30982 19399 31034
rect 19451 30982 21896 31034
rect 1104 30960 21896 30982
rect 1486 30880 1492 30932
rect 1544 30880 1550 30932
rect 2406 30880 2412 30932
rect 2464 30920 2470 30932
rect 5350 30920 5356 30932
rect 2464 30892 5356 30920
rect 2464 30880 2470 30892
rect 5350 30880 5356 30892
rect 5408 30880 5414 30932
rect 8202 30880 8208 30932
rect 8260 30920 8266 30932
rect 8481 30923 8539 30929
rect 8481 30920 8493 30923
rect 8260 30892 8493 30920
rect 8260 30880 8266 30892
rect 8481 30889 8493 30892
rect 8527 30889 8539 30923
rect 8481 30883 8539 30889
rect 10042 30880 10048 30932
rect 10100 30880 10106 30932
rect 11054 30880 11060 30932
rect 11112 30920 11118 30932
rect 11885 30923 11943 30929
rect 11885 30920 11897 30923
rect 11112 30892 11897 30920
rect 11112 30880 11118 30892
rect 11885 30889 11897 30892
rect 11931 30889 11943 30923
rect 12986 30920 12992 30932
rect 11885 30883 11943 30889
rect 12360 30892 12992 30920
rect 1504 30852 1532 30880
rect 1412 30824 1532 30852
rect 1412 30793 1440 30824
rect 2958 30812 2964 30864
rect 3016 30852 3022 30864
rect 3418 30852 3424 30864
rect 3016 30824 3424 30852
rect 3016 30812 3022 30824
rect 3418 30812 3424 30824
rect 3476 30812 3482 30864
rect 3878 30812 3884 30864
rect 3936 30852 3942 30864
rect 4433 30855 4491 30861
rect 4433 30852 4445 30855
rect 3936 30824 4445 30852
rect 3936 30812 3942 30824
rect 4433 30821 4445 30824
rect 4479 30821 4491 30855
rect 10060 30852 10088 30880
rect 12250 30852 12256 30864
rect 10060 30824 12256 30852
rect 4433 30815 4491 30821
rect 12250 30812 12256 30824
rect 12308 30812 12314 30864
rect 5908 30796 5960 30802
rect 1397 30787 1455 30793
rect 1397 30753 1409 30787
rect 1443 30753 1455 30787
rect 3234 30784 3240 30796
rect 1397 30747 1455 30753
rect 2148 30756 3240 30784
rect 2148 30728 2176 30756
rect 3234 30744 3240 30756
rect 3292 30784 3298 30796
rect 3973 30787 4031 30793
rect 3973 30784 3985 30787
rect 3292 30756 3985 30784
rect 3292 30744 3298 30756
rect 3973 30753 3985 30756
rect 4019 30753 4031 30787
rect 3973 30747 4031 30753
rect 4154 30744 4160 30796
rect 4212 30784 4218 30796
rect 4826 30787 4884 30793
rect 4826 30784 4838 30787
rect 4212 30756 4838 30784
rect 4212 30744 4218 30756
rect 4826 30753 4838 30756
rect 4872 30784 4884 30787
rect 5350 30784 5356 30796
rect 4872 30756 5356 30784
rect 4872 30753 4884 30756
rect 4826 30747 4884 30753
rect 5350 30744 5356 30756
rect 5408 30744 5414 30796
rect 8018 30744 8024 30796
rect 8076 30784 8082 30796
rect 9398 30784 9404 30796
rect 8076 30756 9404 30784
rect 8076 30744 8082 30756
rect 9398 30744 9404 30756
rect 9456 30744 9462 30796
rect 11882 30784 11888 30796
rect 11716 30756 11888 30784
rect 5908 30738 5960 30744
rect 1118 30676 1124 30728
rect 1176 30716 1182 30728
rect 1639 30719 1697 30725
rect 1639 30716 1651 30719
rect 1176 30688 1651 30716
rect 1176 30676 1182 30688
rect 1639 30685 1651 30688
rect 1685 30716 1697 30719
rect 1685 30688 2084 30716
rect 1685 30685 1697 30688
rect 1639 30679 1697 30685
rect 2056 30648 2084 30688
rect 2130 30676 2136 30728
rect 2188 30676 2194 30728
rect 2774 30676 2780 30728
rect 2832 30676 2838 30728
rect 2866 30676 2872 30728
rect 2924 30716 2930 30728
rect 3053 30719 3111 30725
rect 3053 30716 3065 30719
rect 2924 30688 3065 30716
rect 2924 30676 2930 30688
rect 3053 30685 3065 30688
rect 3099 30685 3111 30719
rect 3053 30679 3111 30685
rect 3418 30676 3424 30728
rect 3476 30716 3482 30728
rect 3786 30716 3792 30728
rect 3476 30688 3792 30716
rect 3476 30676 3482 30688
rect 3786 30676 3792 30688
rect 3844 30676 3850 30728
rect 4706 30676 4712 30728
rect 4764 30676 4770 30728
rect 4982 30676 4988 30728
rect 5040 30676 5046 30728
rect 6638 30716 6644 30728
rect 6104 30688 6644 30716
rect 6104 30657 6132 30688
rect 6638 30676 6644 30688
rect 6696 30676 6702 30728
rect 6748 30716 6960 30718
rect 7374 30716 7380 30728
rect 6748 30690 7380 30716
rect 5629 30651 5687 30657
rect 2056 30620 4016 30648
rect 2314 30540 2320 30592
rect 2372 30580 2378 30592
rect 2409 30583 2467 30589
rect 2409 30580 2421 30583
rect 2372 30552 2421 30580
rect 2372 30540 2378 30552
rect 2409 30549 2421 30552
rect 2455 30549 2467 30583
rect 2409 30543 2467 30549
rect 2682 30540 2688 30592
rect 2740 30580 2746 30592
rect 2866 30580 2872 30592
rect 2740 30552 2872 30580
rect 2740 30540 2746 30552
rect 2866 30540 2872 30552
rect 2924 30540 2930 30592
rect 3988 30580 4016 30620
rect 5629 30617 5641 30651
rect 5675 30617 5687 30651
rect 5629 30611 5687 30617
rect 6089 30651 6147 30657
rect 6089 30617 6101 30651
rect 6135 30617 6147 30651
rect 6089 30611 6147 30617
rect 4246 30580 4252 30592
rect 3988 30552 4252 30580
rect 4246 30540 4252 30552
rect 4304 30540 4310 30592
rect 4890 30540 4896 30592
rect 4948 30580 4954 30592
rect 5258 30580 5264 30592
rect 4948 30552 5264 30580
rect 4948 30540 4954 30552
rect 5258 30540 5264 30552
rect 5316 30540 5322 30592
rect 5644 30580 5672 30611
rect 6362 30608 6368 30660
rect 6420 30608 6426 30660
rect 6457 30651 6515 30657
rect 6457 30617 6469 30651
rect 6503 30648 6515 30651
rect 6748 30648 6776 30690
rect 6932 30688 7380 30690
rect 7374 30676 7380 30688
rect 7432 30676 7438 30728
rect 11716 30725 11744 30756
rect 11882 30744 11888 30756
rect 11940 30744 11946 30796
rect 11977 30787 12035 30793
rect 11977 30753 11989 30787
rect 12023 30784 12035 30787
rect 12360 30784 12388 30892
rect 12986 30880 12992 30892
rect 13044 30880 13050 30932
rect 13078 30880 13084 30932
rect 13136 30880 13142 30932
rect 13262 30880 13268 30932
rect 13320 30920 13326 30932
rect 15102 30920 15108 30932
rect 13320 30892 15108 30920
rect 13320 30880 13326 30892
rect 15102 30880 15108 30892
rect 15160 30880 15166 30932
rect 16022 30880 16028 30932
rect 16080 30920 16086 30932
rect 18322 30920 18328 30932
rect 16080 30892 18328 30920
rect 16080 30880 16086 30892
rect 18322 30880 18328 30892
rect 18380 30880 18386 30932
rect 18506 30880 18512 30932
rect 18564 30880 18570 30932
rect 20625 30923 20683 30929
rect 18616 30892 20576 30920
rect 12437 30855 12495 30861
rect 12437 30821 12449 30855
rect 12483 30821 12495 30855
rect 12437 30815 12495 30821
rect 12713 30855 12771 30861
rect 12713 30821 12725 30855
rect 12759 30852 12771 30855
rect 13096 30852 13124 30880
rect 12759 30824 13124 30852
rect 17037 30855 17095 30861
rect 12759 30821 12771 30824
rect 12713 30815 12771 30821
rect 17037 30821 17049 30855
rect 17083 30821 17095 30855
rect 17037 30815 17095 30821
rect 17405 30855 17463 30861
rect 17405 30821 17417 30855
rect 17451 30821 17463 30855
rect 17405 30815 17463 30821
rect 12023 30756 12388 30784
rect 12023 30753 12035 30756
rect 11977 30747 12035 30753
rect 11701 30719 11759 30725
rect 11701 30685 11713 30719
rect 11747 30685 11759 30719
rect 11701 30679 11759 30685
rect 11793 30719 11851 30725
rect 11793 30685 11805 30719
rect 11839 30685 11851 30719
rect 11793 30679 11851 30685
rect 12161 30719 12219 30725
rect 12161 30685 12173 30719
rect 12207 30716 12219 30719
rect 12452 30716 12480 30815
rect 13446 30744 13452 30796
rect 13504 30784 13510 30796
rect 14093 30787 14151 30793
rect 14093 30784 14105 30787
rect 13504 30756 14105 30784
rect 13504 30744 13510 30756
rect 14093 30753 14105 30756
rect 14139 30753 14151 30787
rect 14093 30747 14151 30753
rect 12207 30688 12480 30716
rect 12207 30685 12219 30688
rect 12161 30679 12219 30685
rect 6503 30620 6776 30648
rect 6503 30617 6515 30620
rect 6457 30611 6515 30617
rect 6822 30608 6828 30660
rect 6880 30608 6886 30660
rect 11808 30648 11836 30679
rect 12618 30676 12624 30728
rect 12676 30676 12682 30728
rect 12894 30676 12900 30728
rect 12952 30676 12958 30728
rect 14335 30719 14393 30725
rect 14335 30716 14347 30719
rect 14200 30688 14347 30716
rect 14200 30660 14228 30688
rect 14335 30685 14347 30688
rect 14381 30716 14393 30719
rect 15286 30716 15292 30728
rect 14381 30688 15292 30716
rect 14381 30685 14393 30688
rect 14335 30679 14393 30685
rect 15286 30676 15292 30688
rect 15344 30676 15350 30728
rect 15657 30719 15715 30725
rect 15657 30685 15669 30719
rect 15703 30716 15715 30719
rect 16298 30716 16304 30728
rect 15703 30688 16304 30716
rect 15703 30685 15715 30688
rect 15657 30679 15715 30685
rect 16298 30676 16304 30688
rect 16356 30676 16362 30728
rect 17052 30716 17080 30815
rect 17420 30784 17448 30815
rect 17865 30787 17923 30793
rect 17420 30756 17816 30784
rect 17788 30725 17816 30756
rect 17865 30753 17877 30787
rect 17911 30784 17923 30787
rect 18233 30787 18291 30793
rect 18233 30784 18245 30787
rect 17911 30756 18245 30784
rect 17911 30753 17923 30756
rect 17865 30747 17923 30753
rect 18233 30753 18245 30756
rect 18279 30753 18291 30787
rect 18233 30747 18291 30753
rect 18417 30787 18475 30793
rect 18417 30753 18429 30787
rect 18463 30784 18475 30787
rect 18524 30784 18552 30880
rect 18463 30756 18552 30784
rect 18463 30753 18475 30756
rect 18417 30747 18475 30753
rect 17313 30719 17371 30725
rect 17313 30716 17325 30719
rect 17052 30688 17325 30716
rect 17313 30685 17325 30688
rect 17359 30685 17371 30719
rect 17313 30679 17371 30685
rect 17589 30719 17647 30725
rect 17589 30685 17601 30719
rect 17635 30685 17647 30719
rect 17589 30679 17647 30685
rect 17773 30719 17831 30725
rect 17773 30685 17785 30719
rect 17819 30685 17831 30719
rect 17773 30679 17831 30685
rect 12253 30651 12311 30657
rect 12253 30648 12265 30651
rect 7116 30620 9674 30648
rect 11808 30620 12265 30648
rect 7116 30580 7144 30620
rect 5644 30552 7144 30580
rect 7190 30540 7196 30592
rect 7248 30540 7254 30592
rect 7377 30583 7435 30589
rect 7377 30549 7389 30583
rect 7423 30580 7435 30583
rect 7926 30580 7932 30592
rect 7423 30552 7932 30580
rect 7423 30549 7435 30552
rect 7377 30543 7435 30549
rect 7926 30540 7932 30552
rect 7984 30540 7990 30592
rect 9646 30580 9674 30620
rect 12253 30617 12265 30620
rect 12299 30617 12311 30651
rect 12253 30611 12311 30617
rect 14182 30608 14188 30660
rect 14240 30608 14246 30660
rect 15924 30651 15982 30657
rect 15924 30617 15936 30651
rect 15970 30648 15982 30651
rect 16206 30648 16212 30660
rect 15970 30620 16212 30648
rect 15970 30617 15982 30620
rect 15924 30611 15982 30617
rect 16206 30608 16212 30620
rect 16264 30608 16270 30660
rect 17218 30608 17224 30660
rect 17276 30648 17282 30660
rect 17604 30648 17632 30679
rect 18138 30676 18144 30728
rect 18196 30676 18202 30728
rect 18616 30716 18644 30892
rect 20548 30852 20576 30892
rect 20625 30889 20637 30923
rect 20671 30920 20683 30923
rect 20806 30920 20812 30932
rect 20671 30892 20812 30920
rect 20671 30889 20683 30892
rect 20625 30883 20683 30889
rect 20806 30880 20812 30892
rect 20864 30880 20870 30932
rect 21358 30852 21364 30864
rect 20548 30824 21364 30852
rect 21358 30812 21364 30824
rect 21416 30812 21422 30864
rect 22278 30744 22284 30796
rect 22336 30784 22342 30796
rect 22554 30784 22560 30796
rect 22336 30756 22560 30784
rect 22336 30744 22342 30756
rect 22554 30744 22560 30756
rect 22612 30744 22618 30796
rect 18432 30688 18644 30716
rect 18693 30719 18751 30725
rect 17276 30620 17632 30648
rect 17276 30608 17282 30620
rect 13538 30580 13544 30592
rect 9646 30552 13544 30580
rect 13538 30540 13544 30552
rect 13596 30540 13602 30592
rect 14458 30540 14464 30592
rect 14516 30580 14522 30592
rect 15105 30583 15163 30589
rect 15105 30580 15117 30583
rect 14516 30552 15117 30580
rect 14516 30540 14522 30552
rect 15105 30549 15117 30552
rect 15151 30549 15163 30583
rect 15105 30543 15163 30549
rect 16022 30540 16028 30592
rect 16080 30580 16086 30592
rect 18432 30589 18460 30688
rect 18693 30685 18705 30719
rect 18739 30716 18751 30719
rect 18874 30716 18880 30728
rect 18739 30688 18880 30716
rect 18739 30685 18751 30688
rect 18693 30679 18751 30685
rect 18874 30676 18880 30688
rect 18932 30676 18938 30728
rect 19150 30676 19156 30728
rect 19208 30716 19214 30728
rect 19245 30719 19303 30725
rect 19245 30716 19257 30719
rect 19208 30688 19257 30716
rect 19208 30676 19214 30688
rect 19245 30685 19257 30688
rect 19291 30685 19303 30719
rect 19245 30679 19303 30685
rect 19794 30676 19800 30728
rect 19852 30676 19858 30728
rect 20898 30676 20904 30728
rect 20956 30716 20962 30728
rect 20993 30719 21051 30725
rect 20993 30716 21005 30719
rect 20956 30688 21005 30716
rect 20956 30676 20962 30688
rect 20993 30685 21005 30688
rect 21039 30685 21051 30719
rect 20993 30679 21051 30685
rect 21174 30676 21180 30728
rect 21232 30676 21238 30728
rect 18782 30608 18788 30660
rect 18840 30648 18846 30660
rect 19058 30648 19064 30660
rect 18840 30620 19064 30648
rect 18840 30608 18846 30620
rect 19058 30608 19064 30620
rect 19116 30608 19122 30660
rect 19512 30651 19570 30657
rect 19512 30617 19524 30651
rect 19558 30648 19570 30651
rect 19702 30648 19708 30660
rect 19558 30620 19708 30648
rect 19558 30617 19570 30620
rect 19512 30611 19570 30617
rect 19702 30608 19708 30620
rect 19760 30608 19766 30660
rect 17129 30583 17187 30589
rect 17129 30580 17141 30583
rect 16080 30552 17141 30580
rect 16080 30540 16086 30552
rect 17129 30549 17141 30552
rect 17175 30549 17187 30583
rect 17129 30543 17187 30549
rect 18417 30583 18475 30589
rect 18417 30549 18429 30583
rect 18463 30549 18475 30583
rect 18417 30543 18475 30549
rect 18509 30583 18567 30589
rect 18509 30549 18521 30583
rect 18555 30580 18567 30583
rect 19812 30580 19840 30676
rect 21545 30651 21603 30657
rect 21545 30617 21557 30651
rect 21591 30648 21603 30651
rect 22278 30648 22284 30660
rect 21591 30620 22284 30648
rect 21591 30617 21603 30620
rect 21545 30611 21603 30617
rect 22278 30608 22284 30620
rect 22336 30608 22342 30660
rect 18555 30552 19840 30580
rect 18555 30549 18567 30552
rect 18509 30543 18567 30549
rect 20806 30540 20812 30592
rect 20864 30540 20870 30592
rect 1104 30490 22056 30512
rect 1104 30438 6148 30490
rect 6200 30438 6212 30490
rect 6264 30438 6276 30490
rect 6328 30438 6340 30490
rect 6392 30438 6404 30490
rect 6456 30438 11346 30490
rect 11398 30438 11410 30490
rect 11462 30438 11474 30490
rect 11526 30438 11538 30490
rect 11590 30438 11602 30490
rect 11654 30438 16544 30490
rect 16596 30438 16608 30490
rect 16660 30438 16672 30490
rect 16724 30438 16736 30490
rect 16788 30438 16800 30490
rect 16852 30438 21742 30490
rect 21794 30438 21806 30490
rect 21858 30438 21870 30490
rect 21922 30438 21934 30490
rect 21986 30438 21998 30490
rect 22050 30438 22056 30490
rect 1104 30416 22056 30438
rect 1762 30336 1768 30388
rect 1820 30376 1826 30388
rect 3237 30379 3295 30385
rect 3237 30376 3249 30379
rect 1820 30348 3249 30376
rect 1820 30336 1826 30348
rect 3237 30345 3249 30348
rect 3283 30376 3295 30379
rect 3970 30376 3976 30388
rect 3283 30348 3976 30376
rect 3283 30345 3295 30348
rect 3237 30339 3295 30345
rect 3970 30336 3976 30348
rect 4028 30336 4034 30388
rect 4341 30379 4399 30385
rect 4341 30345 4353 30379
rect 4387 30376 4399 30379
rect 4982 30376 4988 30388
rect 4387 30348 4988 30376
rect 4387 30345 4399 30348
rect 4341 30339 4399 30345
rect 4982 30336 4988 30348
rect 5040 30336 5046 30388
rect 5902 30336 5908 30388
rect 5960 30336 5966 30388
rect 6086 30336 6092 30388
rect 6144 30376 6150 30388
rect 7190 30376 7196 30388
rect 6144 30348 7196 30376
rect 6144 30336 6150 30348
rect 7190 30336 7196 30348
rect 7248 30336 7254 30388
rect 7374 30336 7380 30388
rect 7432 30336 7438 30388
rect 7650 30336 7656 30388
rect 7708 30376 7714 30388
rect 10042 30376 10048 30388
rect 7708 30348 10048 30376
rect 7708 30336 7714 30348
rect 10042 30336 10048 30348
rect 10100 30336 10106 30388
rect 12618 30336 12624 30388
rect 12676 30376 12682 30388
rect 13357 30379 13415 30385
rect 13357 30376 13369 30379
rect 12676 30348 13369 30376
rect 12676 30336 12682 30348
rect 13357 30345 13369 30348
rect 13403 30345 13415 30379
rect 13357 30339 13415 30345
rect 13814 30336 13820 30388
rect 13872 30376 13878 30388
rect 14642 30376 14648 30388
rect 13872 30348 14648 30376
rect 13872 30336 13878 30348
rect 14642 30336 14648 30348
rect 14700 30336 14706 30388
rect 15838 30376 15844 30388
rect 15028 30348 15844 30376
rect 1946 30279 1952 30320
rect 1931 30273 1952 30279
rect 1394 30200 1400 30252
rect 1452 30200 1458 30252
rect 1486 30200 1492 30252
rect 1544 30240 1550 30252
rect 1673 30243 1731 30249
rect 1673 30240 1685 30243
rect 1544 30212 1685 30240
rect 1544 30200 1550 30212
rect 1673 30209 1685 30212
rect 1719 30209 1731 30243
rect 1931 30239 1943 30273
rect 2004 30268 2010 30320
rect 2406 30268 2412 30320
rect 2464 30308 2470 30320
rect 3878 30308 3884 30320
rect 2464 30280 3884 30308
rect 2464 30268 2470 30280
rect 3878 30268 3884 30280
rect 3936 30268 3942 30320
rect 5810 30308 5816 30320
rect 4908 30280 5816 30308
rect 1977 30242 1990 30268
rect 3053 30243 3111 30249
rect 1977 30239 1989 30242
rect 1931 30233 1989 30239
rect 1673 30203 1731 30209
rect 3053 30209 3065 30243
rect 3099 30240 3111 30243
rect 3234 30240 3240 30252
rect 3099 30212 3240 30240
rect 3099 30209 3111 30212
rect 3053 30203 3111 30209
rect 3234 30200 3240 30212
rect 3292 30200 3298 30252
rect 3602 30200 3608 30252
rect 3660 30240 3666 30252
rect 4154 30240 4160 30252
rect 3660 30212 4160 30240
rect 3660 30200 3666 30212
rect 4154 30200 4160 30212
rect 4212 30200 4218 30252
rect 4908 30184 4936 30280
rect 5810 30268 5816 30280
rect 5868 30268 5874 30320
rect 5166 30240 5172 30252
rect 5127 30212 5172 30240
rect 5166 30200 5172 30212
rect 5224 30200 5230 30252
rect 5920 30240 5948 30336
rect 9030 30308 9036 30320
rect 8956 30280 9036 30308
rect 8956 30264 8984 30280
rect 9030 30268 9036 30280
rect 9088 30308 9094 30320
rect 10686 30308 10692 30320
rect 9088 30280 10692 30308
rect 9088 30268 9094 30280
rect 10686 30268 10692 30280
rect 10744 30268 10750 30320
rect 8830 30259 8984 30264
rect 8815 30253 8984 30259
rect 6623 30243 6681 30249
rect 6623 30240 6635 30243
rect 5920 30212 6635 30240
rect 6623 30209 6635 30212
rect 6669 30209 6681 30243
rect 6623 30203 6681 30209
rect 7098 30200 7104 30252
rect 7156 30240 7162 30252
rect 8573 30243 8631 30249
rect 8573 30240 8585 30243
rect 7156 30212 8585 30240
rect 7156 30200 7162 30212
rect 8573 30209 8585 30212
rect 8619 30209 8631 30243
rect 8815 30219 8827 30253
rect 8861 30236 8984 30253
rect 8861 30219 8873 30236
rect 8815 30213 8873 30219
rect 8573 30203 8631 30209
rect 9214 30200 9220 30252
rect 9272 30240 9278 30252
rect 11606 30240 11612 30252
rect 9272 30212 11612 30240
rect 9272 30200 9278 30212
rect 11606 30200 11612 30212
rect 11664 30200 11670 30252
rect 12434 30200 12440 30252
rect 12492 30200 12498 30252
rect 13446 30200 13452 30252
rect 13504 30200 13510 30252
rect 13630 30200 13636 30252
rect 13688 30240 13694 30252
rect 13723 30243 13781 30249
rect 13723 30240 13735 30243
rect 13688 30212 13735 30240
rect 13688 30200 13694 30212
rect 13723 30209 13735 30212
rect 13769 30240 13781 30243
rect 15028 30240 15056 30348
rect 15838 30336 15844 30348
rect 15896 30376 15902 30388
rect 15896 30348 16611 30376
rect 15896 30336 15902 30348
rect 15194 30268 15200 30320
rect 15252 30268 15258 30320
rect 16022 30268 16028 30320
rect 16080 30308 16086 30320
rect 16583 30308 16611 30348
rect 17586 30336 17592 30388
rect 17644 30376 17650 30388
rect 18782 30376 18788 30388
rect 17644 30348 18788 30376
rect 17644 30336 17650 30348
rect 18782 30336 18788 30348
rect 18840 30336 18846 30388
rect 18966 30336 18972 30388
rect 19024 30376 19030 30388
rect 19245 30379 19303 30385
rect 19245 30376 19257 30379
rect 19024 30348 19257 30376
rect 19024 30336 19030 30348
rect 19245 30345 19257 30348
rect 19291 30345 19303 30379
rect 19245 30339 19303 30345
rect 20438 30336 20444 30388
rect 20496 30376 20502 30388
rect 22646 30376 22652 30388
rect 20496 30348 22652 30376
rect 20496 30336 20502 30348
rect 22646 30336 22652 30348
rect 22704 30336 22710 30388
rect 16080 30280 16528 30308
rect 16583 30280 19104 30308
rect 16080 30268 16086 30280
rect 13769 30212 15056 30240
rect 15103 30243 15161 30249
rect 13769 30209 13781 30212
rect 13723 30203 13781 30209
rect 15103 30209 15115 30243
rect 15149 30240 15161 30243
rect 15212 30240 15240 30268
rect 16500 30249 16528 30280
rect 15149 30212 15240 30240
rect 16301 30243 16359 30249
rect 15149 30209 15161 30212
rect 15103 30203 15161 30209
rect 16301 30209 16313 30243
rect 16347 30209 16359 30243
rect 16301 30203 16359 30209
rect 16485 30243 16543 30249
rect 16485 30209 16497 30243
rect 16531 30209 16543 30243
rect 16485 30203 16543 30209
rect 16669 30243 16727 30249
rect 16669 30209 16681 30243
rect 16715 30240 16727 30243
rect 16850 30240 16856 30252
rect 16715 30212 16856 30240
rect 16715 30209 16727 30212
rect 16669 30203 16727 30209
rect 2866 30132 2872 30184
rect 2924 30172 2930 30184
rect 3329 30175 3387 30181
rect 3329 30172 3341 30175
rect 2924 30144 3341 30172
rect 2924 30132 2930 30144
rect 3329 30141 3341 30144
rect 3375 30141 3387 30175
rect 3329 30135 3387 30141
rect 4890 30132 4896 30184
rect 4948 30132 4954 30184
rect 6362 30132 6368 30184
rect 6420 30132 6426 30184
rect 11238 30132 11244 30184
rect 11296 30172 11302 30184
rect 11517 30175 11575 30181
rect 11517 30172 11529 30175
rect 11296 30144 11529 30172
rect 11296 30132 11302 30144
rect 11517 30141 11529 30144
rect 11563 30141 11575 30175
rect 11517 30135 11575 30141
rect 11698 30132 11704 30184
rect 11756 30172 11762 30184
rect 11882 30172 11888 30184
rect 11756 30144 11888 30172
rect 11756 30132 11762 30144
rect 11882 30132 11888 30144
rect 11940 30132 11946 30184
rect 12554 30175 12612 30181
rect 12554 30172 12566 30175
rect 12268 30144 12566 30172
rect 1581 30107 1639 30113
rect 1581 30073 1593 30107
rect 1627 30073 1639 30107
rect 1581 30067 1639 30073
rect 2608 30076 3464 30104
rect 1596 30036 1624 30067
rect 2608 30036 2636 30076
rect 1596 30008 2636 30036
rect 2682 29996 2688 30048
rect 2740 29996 2746 30048
rect 3050 29996 3056 30048
rect 3108 30036 3114 30048
rect 3326 30036 3332 30048
rect 3108 30008 3332 30036
rect 3108 29996 3114 30008
rect 3326 29996 3332 30008
rect 3384 29996 3390 30048
rect 3436 30036 3464 30076
rect 5828 30076 6500 30104
rect 5828 30036 5856 30076
rect 3436 30008 5856 30036
rect 5902 29996 5908 30048
rect 5960 29996 5966 30048
rect 6472 30036 6500 30076
rect 9398 30064 9404 30116
rect 9456 30104 9462 30116
rect 9456 30076 11376 30104
rect 9456 30064 9462 30076
rect 7834 30036 7840 30048
rect 6472 30008 7840 30036
rect 7834 29996 7840 30008
rect 7892 29996 7898 30048
rect 8570 29996 8576 30048
rect 8628 30036 8634 30048
rect 9585 30039 9643 30045
rect 9585 30036 9597 30039
rect 8628 30008 9597 30036
rect 8628 29996 8634 30008
rect 9585 30005 9597 30008
rect 9631 30005 9643 30039
rect 11348 30036 11376 30076
rect 11606 30064 11612 30116
rect 11664 30104 11670 30116
rect 12161 30107 12219 30113
rect 12161 30104 12173 30107
rect 11664 30076 12173 30104
rect 11664 30064 11670 30076
rect 12161 30073 12173 30076
rect 12207 30073 12219 30107
rect 12161 30067 12219 30073
rect 12268 30036 12296 30144
rect 12554 30141 12566 30144
rect 12600 30141 12612 30175
rect 12554 30135 12612 30141
rect 12710 30132 12716 30184
rect 12768 30132 12774 30184
rect 13078 30132 13084 30184
rect 13136 30172 13142 30184
rect 13464 30172 13492 30200
rect 13136 30144 13492 30172
rect 13136 30132 13142 30144
rect 14734 30132 14740 30184
rect 14792 30172 14798 30184
rect 14829 30175 14887 30181
rect 14829 30172 14841 30175
rect 14792 30144 14841 30172
rect 14792 30132 14798 30144
rect 14829 30141 14841 30144
rect 14875 30141 14887 30175
rect 14829 30135 14887 30141
rect 16316 30104 16344 30203
rect 16850 30200 16856 30212
rect 16908 30200 16914 30252
rect 16943 30243 17001 30249
rect 16943 30209 16955 30243
rect 16989 30240 17001 30243
rect 17494 30240 17500 30252
rect 16989 30212 17500 30240
rect 16989 30209 17001 30212
rect 16943 30203 17001 30209
rect 17494 30200 17500 30212
rect 17552 30200 17558 30252
rect 18969 30243 19027 30249
rect 18969 30209 18981 30243
rect 19015 30209 19027 30243
rect 18969 30203 19027 30209
rect 18984 30104 19012 30203
rect 19076 30172 19104 30280
rect 19168 30280 20944 30308
rect 19168 30249 19196 30280
rect 19153 30243 19211 30249
rect 19153 30209 19165 30243
rect 19199 30209 19211 30243
rect 19153 30203 19211 30209
rect 19429 30243 19487 30249
rect 19429 30209 19441 30243
rect 19475 30209 19487 30243
rect 19429 30203 19487 30209
rect 19444 30172 19472 30203
rect 19518 30200 19524 30252
rect 19576 30200 19582 30252
rect 19794 30240 19800 30252
rect 19755 30212 19800 30240
rect 19794 30200 19800 30212
rect 19852 30200 19858 30252
rect 20916 30240 20944 30280
rect 20990 30268 20996 30320
rect 21048 30308 21054 30320
rect 21177 30311 21235 30317
rect 21177 30308 21189 30311
rect 21048 30280 21189 30308
rect 21048 30268 21054 30280
rect 21177 30277 21189 30280
rect 21223 30277 21235 30311
rect 21177 30271 21235 30277
rect 21634 30240 21640 30252
rect 20916 30212 21640 30240
rect 21634 30200 21640 30212
rect 21692 30200 21698 30252
rect 19076 30144 19472 30172
rect 16316 30076 16804 30104
rect 18984 30076 19656 30104
rect 16776 30048 16804 30076
rect 13354 30036 13360 30048
rect 11348 30008 13360 30036
rect 9585 29999 9643 30005
rect 13354 29996 13360 30008
rect 13412 29996 13418 30048
rect 13814 29996 13820 30048
rect 13872 30036 13878 30048
rect 14461 30039 14519 30045
rect 14461 30036 14473 30039
rect 13872 30008 14473 30036
rect 13872 29996 13878 30008
rect 14461 30005 14473 30008
rect 14507 30005 14519 30039
rect 14461 29999 14519 30005
rect 15838 29996 15844 30048
rect 15896 29996 15902 30048
rect 16390 29996 16396 30048
rect 16448 29996 16454 30048
rect 16758 29996 16764 30048
rect 16816 30036 16822 30048
rect 17681 30039 17739 30045
rect 17681 30036 17693 30039
rect 16816 30008 17693 30036
rect 16816 29996 16822 30008
rect 17681 30005 17693 30008
rect 17727 30005 17739 30039
rect 17681 29999 17739 30005
rect 19058 29996 19064 30048
rect 19116 29996 19122 30048
rect 19628 30036 19656 30076
rect 20533 30039 20591 30045
rect 20533 30036 20545 30039
rect 19628 30008 20545 30036
rect 20533 30005 20545 30008
rect 20579 30036 20591 30039
rect 20990 30036 20996 30048
rect 20579 30008 20996 30036
rect 20579 30005 20591 30008
rect 20533 29999 20591 30005
rect 20990 29996 20996 30008
rect 21048 29996 21054 30048
rect 21450 29996 21456 30048
rect 21508 29996 21514 30048
rect 1104 29946 21896 29968
rect 1104 29894 3549 29946
rect 3601 29894 3613 29946
rect 3665 29894 3677 29946
rect 3729 29894 3741 29946
rect 3793 29894 3805 29946
rect 3857 29894 8747 29946
rect 8799 29894 8811 29946
rect 8863 29894 8875 29946
rect 8927 29894 8939 29946
rect 8991 29894 9003 29946
rect 9055 29894 13945 29946
rect 13997 29894 14009 29946
rect 14061 29894 14073 29946
rect 14125 29894 14137 29946
rect 14189 29894 14201 29946
rect 14253 29894 19143 29946
rect 19195 29894 19207 29946
rect 19259 29894 19271 29946
rect 19323 29894 19335 29946
rect 19387 29894 19399 29946
rect 19451 29894 21896 29946
rect 1104 29872 21896 29894
rect 4154 29792 4160 29844
rect 4212 29832 4218 29844
rect 5166 29832 5172 29844
rect 4212 29804 5172 29832
rect 4212 29792 4218 29804
rect 5166 29792 5172 29804
rect 5224 29792 5230 29844
rect 7834 29792 7840 29844
rect 7892 29832 7898 29844
rect 9214 29832 9220 29844
rect 7892 29804 9220 29832
rect 7892 29792 7898 29804
rect 9214 29792 9220 29804
rect 9272 29792 9278 29844
rect 10962 29832 10968 29844
rect 9876 29804 10968 29832
rect 4614 29724 4620 29776
rect 4672 29724 4678 29776
rect 6730 29724 6736 29776
rect 6788 29764 6794 29776
rect 7466 29764 7472 29776
rect 6788 29736 7472 29764
rect 6788 29724 6794 29736
rect 7466 29724 7472 29736
rect 7524 29724 7530 29776
rect 9876 29764 9904 29804
rect 10962 29792 10968 29804
rect 11020 29792 11026 29844
rect 12250 29792 12256 29844
rect 12308 29832 12314 29844
rect 12308 29804 12756 29832
rect 12308 29792 12314 29804
rect 8266 29736 9904 29764
rect 10781 29767 10839 29773
rect 2314 29656 2320 29708
rect 2372 29656 2378 29708
rect 4525 29699 4583 29705
rect 4525 29665 4537 29699
rect 4571 29696 4583 29699
rect 4632 29696 4660 29724
rect 4571 29668 4660 29696
rect 4571 29665 4583 29668
rect 4525 29659 4583 29665
rect 750 29588 756 29640
rect 808 29628 814 29640
rect 1489 29631 1547 29637
rect 1489 29628 1501 29631
rect 808 29600 1501 29628
rect 808 29588 814 29600
rect 1489 29597 1501 29600
rect 1535 29597 1547 29631
rect 1489 29591 1547 29597
rect 2409 29631 2467 29637
rect 2409 29597 2421 29631
rect 2455 29628 2467 29631
rect 2682 29628 2688 29640
rect 2455 29600 2688 29628
rect 2455 29597 2467 29600
rect 2409 29591 2467 29597
rect 2682 29588 2688 29600
rect 2740 29588 2746 29640
rect 2777 29631 2835 29637
rect 2777 29597 2789 29631
rect 2823 29628 2835 29631
rect 2958 29628 2964 29640
rect 2823 29600 2964 29628
rect 2823 29597 2835 29600
rect 2777 29591 2835 29597
rect 2958 29588 2964 29600
rect 3016 29628 3022 29640
rect 3016 29600 3464 29628
rect 3016 29588 3022 29600
rect 1670 29520 1676 29572
rect 1728 29520 1734 29572
rect 1854 29520 1860 29572
rect 1912 29560 1918 29572
rect 2041 29563 2099 29569
rect 2041 29560 2053 29563
rect 1912 29532 2053 29560
rect 1912 29520 1918 29532
rect 2041 29529 2053 29532
rect 2087 29529 2099 29563
rect 2041 29523 2099 29529
rect 2317 29563 2375 29569
rect 2317 29529 2329 29563
rect 2363 29560 2375 29563
rect 2498 29560 2504 29572
rect 2363 29532 2504 29560
rect 2363 29529 2375 29532
rect 2317 29523 2375 29529
rect 2498 29520 2504 29532
rect 2556 29520 2562 29572
rect 3436 29560 3464 29600
rect 3510 29588 3516 29640
rect 3568 29628 3574 29640
rect 4249 29631 4307 29637
rect 4249 29628 4261 29631
rect 3568 29600 4261 29628
rect 3568 29588 3574 29600
rect 4249 29597 4261 29600
rect 4295 29597 4307 29631
rect 4632 29628 4660 29668
rect 5902 29656 5908 29708
rect 5960 29656 5966 29708
rect 7098 29656 7104 29708
rect 7156 29696 7162 29708
rect 8266 29696 8294 29736
rect 10781 29733 10793 29767
rect 10827 29764 10839 29767
rect 11606 29764 11612 29776
rect 10827 29736 11612 29764
rect 10827 29733 10839 29736
rect 10781 29727 10839 29733
rect 11606 29724 11612 29736
rect 11664 29764 11670 29776
rect 11773 29767 11831 29773
rect 11773 29764 11785 29767
rect 11664 29736 11785 29764
rect 11664 29724 11670 29736
rect 11773 29733 11785 29736
rect 11819 29733 11831 29767
rect 12728 29764 12756 29804
rect 12894 29792 12900 29844
rect 12952 29832 12958 29844
rect 12989 29835 13047 29841
rect 12989 29832 13001 29835
rect 12952 29804 13001 29832
rect 12952 29792 12958 29804
rect 12989 29801 13001 29804
rect 13035 29801 13047 29835
rect 15838 29832 15844 29844
rect 12989 29795 13047 29801
rect 14752 29804 15844 29832
rect 14752 29773 14780 29804
rect 15838 29792 15844 29804
rect 15896 29792 15902 29844
rect 16390 29792 16396 29844
rect 16448 29792 16454 29844
rect 18322 29792 18328 29844
rect 18380 29832 18386 29844
rect 18506 29832 18512 29844
rect 18380 29804 18512 29832
rect 18380 29792 18386 29804
rect 18506 29792 18512 29804
rect 18564 29792 18570 29844
rect 19058 29792 19064 29844
rect 19116 29792 19122 29844
rect 20073 29835 20131 29841
rect 20073 29801 20085 29835
rect 20119 29832 20131 29835
rect 20622 29832 20628 29844
rect 20119 29804 20628 29832
rect 20119 29801 20131 29804
rect 20073 29795 20131 29801
rect 20622 29792 20628 29804
rect 20680 29792 20686 29844
rect 20714 29792 20720 29844
rect 20772 29832 20778 29844
rect 20993 29835 21051 29841
rect 20993 29832 21005 29835
rect 20772 29804 21005 29832
rect 20772 29792 20778 29804
rect 20993 29801 21005 29804
rect 21039 29801 21051 29835
rect 20993 29795 21051 29801
rect 14737 29767 14795 29773
rect 12728 29736 14410 29764
rect 11773 29727 11831 29733
rect 12912 29708 12940 29736
rect 7156 29668 7512 29696
rect 7156 29656 7162 29668
rect 7374 29628 7380 29640
rect 4632 29600 7380 29628
rect 4249 29591 4307 29597
rect 7374 29588 7380 29600
rect 7432 29588 7438 29640
rect 7484 29637 7512 29668
rect 8128 29668 8294 29696
rect 7469 29631 7527 29637
rect 7469 29597 7481 29631
rect 7515 29597 7527 29631
rect 7711 29631 7769 29637
rect 7711 29628 7723 29631
rect 7469 29591 7527 29597
rect 7574 29600 7723 29628
rect 7574 29572 7602 29600
rect 7711 29597 7723 29600
rect 7757 29597 7769 29631
rect 7711 29591 7769 29597
rect 7834 29588 7840 29640
rect 7892 29628 7898 29640
rect 8128 29628 8156 29668
rect 9030 29656 9036 29708
rect 9088 29696 9094 29708
rect 9490 29696 9496 29708
rect 9088 29668 9496 29696
rect 9088 29656 9094 29668
rect 9490 29656 9496 29668
rect 9548 29656 9554 29708
rect 10594 29656 10600 29708
rect 10652 29696 10658 29708
rect 10652 29668 11284 29696
rect 10652 29656 10658 29668
rect 7892 29600 8156 29628
rect 7892 29588 7898 29600
rect 8294 29588 8300 29640
rect 8352 29628 8358 29640
rect 9214 29628 9220 29640
rect 8352 29600 9220 29628
rect 8352 29588 8358 29600
rect 9214 29588 9220 29600
rect 9272 29588 9278 29640
rect 9769 29631 9827 29637
rect 9769 29597 9781 29631
rect 9815 29597 9827 29631
rect 9769 29591 9827 29597
rect 10043 29631 10101 29637
rect 10043 29597 10055 29631
rect 10089 29628 10101 29631
rect 10134 29628 10140 29640
rect 10089 29600 10140 29628
rect 10089 29597 10101 29600
rect 10043 29591 10101 29597
rect 4154 29560 4160 29572
rect 3068 29532 3372 29560
rect 3436 29532 4160 29560
rect 1762 29452 1768 29504
rect 1820 29492 1826 29504
rect 3068 29492 3096 29532
rect 1820 29464 3096 29492
rect 3145 29495 3203 29501
rect 1820 29452 1826 29464
rect 3145 29461 3157 29495
rect 3191 29492 3203 29495
rect 3234 29492 3240 29504
rect 3191 29464 3240 29492
rect 3191 29461 3203 29464
rect 3145 29455 3203 29461
rect 3234 29452 3240 29464
rect 3292 29452 3298 29504
rect 3344 29501 3372 29532
rect 4154 29520 4160 29532
rect 4212 29520 4218 29572
rect 5353 29563 5411 29569
rect 5353 29529 5365 29563
rect 5399 29560 5411 29563
rect 5442 29560 5448 29572
rect 5399 29532 5448 29560
rect 5399 29529 5411 29532
rect 5353 29523 5411 29529
rect 5442 29520 5448 29532
rect 5500 29520 5506 29572
rect 5626 29520 5632 29572
rect 5684 29520 5690 29572
rect 5718 29520 5724 29572
rect 5776 29520 5782 29572
rect 5994 29520 6000 29572
rect 6052 29560 6058 29572
rect 6089 29563 6147 29569
rect 6089 29560 6101 29563
rect 6052 29532 6101 29560
rect 6052 29520 6058 29532
rect 6089 29529 6101 29532
rect 6135 29560 6147 29563
rect 6546 29560 6552 29572
rect 6135 29532 6552 29560
rect 6135 29529 6147 29532
rect 6089 29523 6147 29529
rect 6546 29520 6552 29532
rect 6604 29520 6610 29572
rect 6822 29520 6828 29572
rect 6880 29560 6886 29572
rect 7190 29560 7196 29572
rect 6880 29532 7196 29560
rect 6880 29520 6886 29532
rect 7190 29520 7196 29532
rect 7248 29520 7254 29572
rect 7558 29520 7564 29572
rect 7616 29520 7622 29572
rect 9784 29560 9812 29591
rect 10134 29588 10140 29600
rect 10192 29588 10198 29640
rect 10870 29588 10876 29640
rect 10928 29588 10934 29640
rect 11149 29631 11207 29637
rect 11149 29597 11161 29631
rect 11195 29597 11207 29631
rect 11256 29628 11284 29668
rect 11330 29656 11336 29708
rect 11388 29656 11394 29708
rect 12069 29699 12127 29705
rect 12069 29696 12081 29699
rect 11440 29668 12081 29696
rect 11440 29628 11468 29668
rect 12069 29665 12081 29668
rect 12115 29665 12127 29699
rect 12069 29659 12127 29665
rect 12158 29656 12164 29708
rect 12216 29705 12222 29708
rect 12216 29699 12265 29705
rect 12216 29665 12219 29699
rect 12253 29665 12265 29699
rect 12710 29696 12716 29708
rect 12216 29659 12265 29665
rect 12360 29668 12716 29696
rect 12216 29656 12222 29659
rect 12360 29637 12388 29668
rect 12710 29656 12716 29668
rect 12768 29656 12774 29708
rect 12894 29656 12900 29708
rect 12952 29656 12958 29708
rect 13906 29656 13912 29708
rect 13964 29696 13970 29708
rect 14182 29696 14188 29708
rect 13964 29668 14188 29696
rect 13964 29656 13970 29668
rect 14182 29656 14188 29668
rect 14240 29696 14246 29708
rect 14277 29699 14335 29705
rect 14277 29696 14289 29699
rect 14240 29668 14289 29696
rect 14240 29656 14246 29668
rect 14277 29665 14289 29668
rect 14323 29665 14335 29699
rect 14382 29696 14410 29736
rect 14737 29733 14749 29767
rect 14783 29733 14795 29767
rect 14737 29727 14795 29733
rect 16025 29767 16083 29773
rect 16025 29733 16037 29767
rect 16071 29733 16083 29767
rect 16025 29727 16083 29733
rect 15289 29699 15347 29705
rect 14382 29668 15056 29696
rect 14277 29659 14335 29665
rect 11256 29600 11468 29628
rect 12345 29631 12403 29637
rect 11149 29591 11207 29597
rect 12345 29597 12357 29631
rect 12391 29597 12403 29631
rect 12345 29591 12403 29597
rect 10888 29560 10916 29588
rect 7668 29532 9628 29560
rect 9784 29532 10916 29560
rect 3329 29495 3387 29501
rect 3329 29461 3341 29495
rect 3375 29461 3387 29495
rect 3329 29455 3387 29461
rect 5902 29452 5908 29504
rect 5960 29492 5966 29504
rect 6454 29492 6460 29504
rect 5960 29464 6460 29492
rect 5960 29452 5966 29464
rect 6454 29452 6460 29464
rect 6512 29452 6518 29504
rect 6638 29452 6644 29504
rect 6696 29452 6702 29504
rect 7374 29452 7380 29504
rect 7432 29492 7438 29504
rect 7668 29492 7696 29532
rect 7432 29464 7696 29492
rect 7432 29452 7438 29464
rect 8110 29452 8116 29504
rect 8168 29492 8174 29504
rect 8481 29495 8539 29501
rect 8481 29492 8493 29495
rect 8168 29464 8493 29492
rect 8168 29452 8174 29464
rect 8481 29461 8493 29464
rect 8527 29461 8539 29495
rect 9600 29492 9628 29532
rect 10042 29492 10048 29504
rect 9600 29464 10048 29492
rect 8481 29455 8539 29461
rect 10042 29452 10048 29464
rect 10100 29452 10106 29504
rect 11164 29492 11192 29591
rect 13262 29588 13268 29640
rect 13320 29628 13326 29640
rect 15028 29637 15056 29668
rect 15289 29665 15301 29699
rect 15335 29696 15347 29699
rect 15470 29696 15476 29708
rect 15335 29668 15476 29696
rect 15335 29665 15347 29668
rect 15289 29659 15347 29665
rect 15470 29656 15476 29668
rect 15528 29656 15534 29708
rect 16040 29696 16068 29727
rect 16408 29696 16436 29792
rect 16669 29767 16727 29773
rect 16669 29733 16681 29767
rect 16715 29764 16727 29767
rect 16945 29767 17003 29773
rect 16945 29764 16957 29767
rect 16715 29736 16957 29764
rect 16715 29733 16727 29736
rect 16669 29727 16727 29733
rect 16945 29733 16957 29736
rect 16991 29733 17003 29767
rect 16945 29727 17003 29733
rect 17129 29699 17187 29705
rect 17129 29696 17141 29699
rect 16040 29668 16344 29696
rect 16408 29668 17141 29696
rect 14093 29631 14151 29637
rect 14093 29628 14105 29631
rect 13320 29600 14105 29628
rect 13320 29588 13326 29600
rect 14093 29597 14105 29600
rect 14139 29628 14151 29631
rect 15013 29631 15071 29637
rect 14139 29600 14228 29628
rect 14139 29597 14151 29600
rect 14093 29591 14151 29597
rect 14200 29504 14228 29600
rect 15013 29597 15025 29631
rect 15059 29597 15071 29631
rect 15013 29591 15071 29597
rect 15102 29588 15108 29640
rect 15160 29637 15166 29640
rect 15160 29631 15188 29637
rect 15176 29597 15188 29631
rect 15160 29591 15188 29597
rect 15933 29631 15991 29637
rect 15933 29597 15945 29631
rect 15979 29628 15991 29631
rect 15979 29600 16160 29628
rect 15979 29597 15991 29600
rect 15933 29591 15991 29597
rect 15160 29588 15166 29591
rect 13998 29492 14004 29504
rect 11164 29464 14004 29492
rect 13998 29452 14004 29464
rect 14056 29452 14062 29504
rect 14182 29452 14188 29504
rect 14240 29492 14246 29504
rect 15010 29492 15016 29504
rect 14240 29464 15016 29492
rect 14240 29452 14246 29464
rect 15010 29452 15016 29464
rect 15068 29452 15074 29504
rect 16132 29492 16160 29600
rect 16206 29588 16212 29640
rect 16264 29588 16270 29640
rect 16316 29628 16344 29668
rect 17129 29665 17141 29668
rect 17175 29665 17187 29699
rect 17129 29659 17187 29665
rect 18046 29656 18052 29708
rect 18104 29696 18110 29708
rect 18322 29696 18328 29708
rect 18104 29668 18328 29696
rect 18104 29656 18110 29668
rect 18322 29656 18328 29668
rect 18380 29656 18386 29708
rect 19076 29696 19104 29792
rect 20349 29767 20407 29773
rect 20349 29733 20361 29767
rect 20395 29764 20407 29767
rect 20898 29764 20904 29776
rect 20395 29736 20904 29764
rect 20395 29733 20407 29736
rect 20349 29727 20407 29733
rect 20898 29724 20904 29736
rect 20956 29724 20962 29776
rect 21177 29699 21235 29705
rect 21177 29696 21189 29699
rect 19076 29668 21189 29696
rect 21177 29665 21189 29668
rect 21223 29665 21235 29699
rect 21177 29659 21235 29665
rect 16577 29631 16635 29637
rect 16577 29628 16589 29631
rect 16316 29600 16589 29628
rect 16577 29597 16589 29600
rect 16623 29597 16635 29631
rect 16577 29591 16635 29597
rect 16758 29588 16764 29640
rect 16816 29628 16822 29640
rect 16853 29631 16911 29637
rect 16853 29628 16865 29631
rect 16816 29600 16865 29628
rect 16816 29588 16822 29600
rect 16853 29597 16865 29600
rect 16899 29597 16911 29631
rect 17405 29631 17463 29637
rect 17405 29628 17417 29631
rect 16853 29591 16911 29597
rect 17052 29600 17417 29628
rect 17052 29504 17080 29600
rect 17405 29597 17417 29600
rect 17451 29597 17463 29631
rect 17405 29591 17463 29597
rect 18138 29588 18144 29640
rect 18196 29588 18202 29640
rect 19978 29588 19984 29640
rect 20036 29588 20042 29640
rect 20257 29631 20315 29637
rect 20257 29597 20269 29631
rect 20303 29597 20315 29631
rect 20257 29591 20315 29597
rect 19702 29560 19708 29572
rect 17144 29532 19708 29560
rect 17034 29492 17040 29504
rect 16132 29464 17040 29492
rect 17034 29452 17040 29464
rect 17092 29452 17098 29504
rect 17144 29501 17172 29532
rect 19702 29520 19708 29532
rect 19760 29520 19766 29572
rect 20272 29560 20300 29591
rect 20530 29588 20536 29640
rect 20588 29588 20594 29640
rect 20809 29631 20867 29637
rect 20809 29597 20821 29631
rect 20855 29597 20867 29631
rect 20809 29591 20867 29597
rect 20901 29631 20959 29637
rect 20901 29597 20913 29631
rect 20947 29628 20959 29631
rect 20990 29628 20996 29640
rect 20947 29600 20996 29628
rect 20947 29597 20959 29600
rect 20901 29591 20959 29597
rect 19812 29532 20300 29560
rect 17129 29495 17187 29501
rect 17129 29461 17141 29495
rect 17175 29461 17187 29495
rect 17129 29455 17187 29461
rect 17218 29452 17224 29504
rect 17276 29452 17282 29504
rect 17954 29452 17960 29504
rect 18012 29452 18018 29504
rect 19812 29501 19840 29532
rect 20438 29520 20444 29572
rect 20496 29560 20502 29572
rect 20824 29560 20852 29591
rect 20990 29588 20996 29600
rect 21048 29588 21054 29640
rect 21082 29588 21088 29640
rect 21140 29628 21146 29640
rect 21269 29631 21327 29637
rect 21269 29628 21281 29631
rect 21140 29600 21281 29628
rect 21140 29588 21146 29600
rect 21269 29597 21281 29600
rect 21315 29597 21327 29631
rect 21269 29591 21327 29597
rect 20496 29532 20852 29560
rect 20496 29520 20502 29532
rect 19797 29495 19855 29501
rect 19797 29461 19809 29495
rect 19843 29461 19855 29495
rect 19797 29455 19855 29461
rect 20625 29495 20683 29501
rect 20625 29461 20637 29495
rect 20671 29492 20683 29495
rect 20990 29492 20996 29504
rect 20671 29464 20996 29492
rect 20671 29461 20683 29464
rect 20625 29455 20683 29461
rect 20990 29452 20996 29464
rect 21048 29452 21054 29504
rect 21174 29452 21180 29504
rect 21232 29452 21238 29504
rect 21453 29495 21511 29501
rect 21453 29461 21465 29495
rect 21499 29492 21511 29495
rect 22186 29492 22192 29504
rect 21499 29464 22192 29492
rect 21499 29461 21511 29464
rect 21453 29455 21511 29461
rect 22186 29452 22192 29464
rect 22244 29452 22250 29504
rect 1104 29402 22056 29424
rect 1104 29350 6148 29402
rect 6200 29350 6212 29402
rect 6264 29350 6276 29402
rect 6328 29350 6340 29402
rect 6392 29350 6404 29402
rect 6456 29350 11346 29402
rect 11398 29350 11410 29402
rect 11462 29350 11474 29402
rect 11526 29350 11538 29402
rect 11590 29350 11602 29402
rect 11654 29350 16544 29402
rect 16596 29350 16608 29402
rect 16660 29350 16672 29402
rect 16724 29350 16736 29402
rect 16788 29350 16800 29402
rect 16852 29350 21742 29402
rect 21794 29350 21806 29402
rect 21858 29350 21870 29402
rect 21922 29350 21934 29402
rect 21986 29350 21998 29402
rect 22050 29350 22056 29402
rect 1104 29328 22056 29350
rect 14 29248 20 29300
rect 72 29288 78 29300
rect 2590 29288 2596 29300
rect 72 29260 2596 29288
rect 72 29248 78 29260
rect 2590 29248 2596 29260
rect 2648 29248 2654 29300
rect 3142 29248 3148 29300
rect 3200 29248 3206 29300
rect 5718 29248 5724 29300
rect 5776 29288 5782 29300
rect 5905 29291 5963 29297
rect 5905 29288 5917 29291
rect 5776 29260 5917 29288
rect 5776 29248 5782 29260
rect 5905 29257 5917 29260
rect 5951 29257 5963 29291
rect 5905 29251 5963 29257
rect 6012 29260 11818 29288
rect 2038 29180 2044 29232
rect 2096 29180 2102 29232
rect 2406 29180 2412 29232
rect 2464 29220 2470 29232
rect 2866 29220 2872 29232
rect 2464 29192 2872 29220
rect 2464 29180 2470 29192
rect 2866 29180 2872 29192
rect 2924 29180 2930 29232
rect 6012 29220 6040 29260
rect 3436 29192 6040 29220
rect 1855 29155 1913 29161
rect 1855 29121 1867 29155
rect 1901 29152 1913 29155
rect 2056 29152 2084 29180
rect 1901 29124 2912 29152
rect 1901 29121 1913 29124
rect 1855 29115 1913 29121
rect 1302 29044 1308 29096
rect 1360 29084 1366 29096
rect 1581 29087 1639 29093
rect 1581 29084 1593 29087
rect 1360 29056 1593 29084
rect 1360 29044 1366 29056
rect 1581 29053 1593 29056
rect 1627 29053 1639 29087
rect 2884 29084 2912 29124
rect 2958 29112 2964 29164
rect 3016 29112 3022 29164
rect 3436 29152 3464 29192
rect 9214 29180 9220 29232
rect 9272 29180 9278 29232
rect 9423 29180 9429 29232
rect 9481 29229 9487 29232
rect 9481 29223 9505 29229
rect 9493 29189 9505 29223
rect 9481 29183 9505 29189
rect 9769 29223 9827 29229
rect 9769 29189 9781 29223
rect 9815 29220 9827 29223
rect 10597 29223 10655 29229
rect 9815 29192 10548 29220
rect 9815 29189 9827 29192
rect 9769 29183 9827 29189
rect 9481 29180 9487 29183
rect 3068 29124 3464 29152
rect 3511 29155 3569 29161
rect 3068 29084 3096 29124
rect 3511 29121 3523 29155
rect 3557 29152 3569 29155
rect 4614 29152 4620 29164
rect 3557 29124 4620 29152
rect 3557 29121 3569 29124
rect 3511 29115 3569 29121
rect 4614 29112 4620 29124
rect 4672 29112 4678 29164
rect 4890 29112 4896 29164
rect 4948 29112 4954 29164
rect 5166 29152 5172 29164
rect 5127 29124 5172 29152
rect 5166 29112 5172 29124
rect 5224 29112 5230 29164
rect 7374 29112 7380 29164
rect 7432 29112 7438 29164
rect 8478 29161 8484 29164
rect 8435 29155 8484 29161
rect 8435 29121 8447 29155
rect 8481 29121 8484 29155
rect 8435 29115 8484 29121
rect 8478 29112 8484 29115
rect 8536 29112 8542 29164
rect 8570 29112 8576 29164
rect 8628 29112 8634 29164
rect 9784 29152 9812 29183
rect 9232 29124 9812 29152
rect 9861 29155 9919 29161
rect 2884 29056 3096 29084
rect 3237 29087 3295 29093
rect 1581 29047 1639 29053
rect 3237 29053 3249 29087
rect 3283 29053 3295 29087
rect 3237 29047 3295 29053
rect 7561 29087 7619 29093
rect 7561 29053 7573 29087
rect 7607 29053 7619 29087
rect 7561 29047 7619 29053
rect 8021 29087 8079 29093
rect 8021 29053 8033 29087
rect 8067 29084 8079 29087
rect 8110 29084 8116 29096
rect 8067 29056 8116 29084
rect 8067 29053 8079 29056
rect 8021 29047 8079 29053
rect 1596 28948 1624 29047
rect 2314 28976 2320 29028
rect 2372 29016 2378 29028
rect 3142 29016 3148 29028
rect 2372 28988 3148 29016
rect 2372 28976 2378 28988
rect 3142 28976 3148 28988
rect 3200 29016 3206 29028
rect 3252 29016 3280 29047
rect 3200 28988 3280 29016
rect 3200 28976 3206 28988
rect 4062 28976 4068 29028
rect 4120 29016 4126 29028
rect 4249 29019 4307 29025
rect 4249 29016 4261 29019
rect 4120 28988 4261 29016
rect 4120 28976 4126 28988
rect 4249 28985 4261 28988
rect 4295 28985 4307 29019
rect 7576 29016 7604 29047
rect 8110 29044 8116 29056
rect 8168 29044 8174 29096
rect 8297 29087 8355 29093
rect 8297 29053 8309 29087
rect 8343 29084 8355 29087
rect 9232 29084 9260 29124
rect 9861 29121 9873 29155
rect 9907 29152 9919 29155
rect 10134 29152 10140 29164
rect 9907 29124 10140 29152
rect 9907 29121 9919 29124
rect 9861 29115 9919 29121
rect 10134 29112 10140 29124
rect 10192 29112 10198 29164
rect 10226 29112 10232 29164
rect 10284 29112 10290 29164
rect 10520 29152 10548 29192
rect 10597 29189 10609 29223
rect 10643 29220 10655 29223
rect 10962 29220 10968 29232
rect 10643 29192 10968 29220
rect 10643 29189 10655 29192
rect 10597 29183 10655 29189
rect 10962 29180 10968 29192
rect 11020 29180 11026 29232
rect 10520 29124 10640 29152
rect 10612 29096 10640 29124
rect 10870 29112 10876 29164
rect 10928 29152 10934 29164
rect 11790 29161 11818 29260
rect 11882 29248 11888 29300
rect 11940 29288 11946 29300
rect 12342 29288 12348 29300
rect 11940 29260 12348 29288
rect 11940 29248 11946 29260
rect 12342 29248 12348 29260
rect 12400 29248 12406 29300
rect 12529 29291 12587 29297
rect 12529 29257 12541 29291
rect 12575 29288 12587 29291
rect 12710 29288 12716 29300
rect 12575 29260 12716 29288
rect 12575 29257 12587 29260
rect 12529 29251 12587 29257
rect 12710 29248 12716 29260
rect 12768 29248 12774 29300
rect 13262 29248 13268 29300
rect 13320 29288 13326 29300
rect 14274 29288 14280 29300
rect 13320 29260 14280 29288
rect 13320 29248 13326 29260
rect 14274 29248 14280 29260
rect 14332 29248 14338 29300
rect 14734 29248 14740 29300
rect 14792 29288 14798 29300
rect 15105 29291 15163 29297
rect 14792 29260 15056 29288
rect 14792 29248 14798 29260
rect 15028 29220 15056 29260
rect 15105 29257 15117 29291
rect 15151 29288 15163 29291
rect 16206 29288 16212 29300
rect 15151 29260 16212 29288
rect 15151 29257 15163 29260
rect 15105 29251 15163 29257
rect 16206 29248 16212 29260
rect 16264 29248 16270 29300
rect 17034 29248 17040 29300
rect 17092 29248 17098 29300
rect 18049 29291 18107 29297
rect 18049 29257 18061 29291
rect 18095 29288 18107 29291
rect 18138 29288 18144 29300
rect 18095 29260 18144 29288
rect 18095 29257 18107 29260
rect 18049 29251 18107 29257
rect 18138 29248 18144 29260
rect 18196 29248 18202 29300
rect 18506 29248 18512 29300
rect 18564 29288 18570 29300
rect 19981 29291 20039 29297
rect 18564 29260 19104 29288
rect 18564 29248 18570 29260
rect 16022 29220 16028 29232
rect 15028 29192 16028 29220
rect 11517 29155 11575 29161
rect 11517 29152 11529 29155
rect 10928 29124 11529 29152
rect 10928 29112 10934 29124
rect 11517 29121 11529 29124
rect 11563 29121 11575 29155
rect 11790 29155 11849 29161
rect 11790 29124 11803 29155
rect 11517 29115 11575 29121
rect 11791 29121 11803 29124
rect 11837 29152 11849 29155
rect 11837 29124 13584 29152
rect 11837 29121 11849 29124
rect 11791 29115 11849 29121
rect 8343 29056 9260 29084
rect 8343 29053 8355 29056
rect 8297 29047 8355 29053
rect 9398 29044 9404 29096
rect 9456 29044 9462 29096
rect 10594 29044 10600 29096
rect 10652 29084 10658 29096
rect 10652 29056 11560 29084
rect 10652 29044 10658 29056
rect 7834 29016 7840 29028
rect 7576 28988 7840 29016
rect 4249 28979 4307 28985
rect 7834 28976 7840 28988
rect 7892 28976 7898 29028
rect 9030 28976 9036 29028
rect 9088 29016 9094 29028
rect 9214 29016 9220 29028
rect 9088 28988 9220 29016
rect 9088 28976 9094 28988
rect 9214 28976 9220 28988
rect 9272 28976 9278 29028
rect 10778 28976 10784 29028
rect 10836 28976 10842 29028
rect 11532 29016 11560 29056
rect 12250 29044 12256 29096
rect 12308 29044 12314 29096
rect 13262 29044 13268 29096
rect 13320 29044 13326 29096
rect 13449 29087 13507 29093
rect 13449 29053 13461 29087
rect 13495 29053 13507 29087
rect 13449 29047 13507 29053
rect 12268 29016 12296 29044
rect 13464 29016 13492 29047
rect 11532 28988 11652 29016
rect 12268 28988 13492 29016
rect 13556 29016 13584 29124
rect 14274 29112 14280 29164
rect 14332 29161 14338 29164
rect 14332 29155 14360 29161
rect 14348 29121 14360 29155
rect 14332 29115 14360 29121
rect 14332 29112 14338 29115
rect 14458 29112 14464 29164
rect 14516 29112 14522 29164
rect 15028 29152 15056 29192
rect 16022 29180 16028 29192
rect 16080 29180 16086 29232
rect 15197 29155 15255 29161
rect 15197 29152 15209 29155
rect 15028 29124 15209 29152
rect 15197 29121 15209 29124
rect 15243 29121 15255 29155
rect 15197 29115 15255 29121
rect 15471 29155 15529 29161
rect 15471 29121 15483 29155
rect 15517 29152 15529 29155
rect 15930 29152 15936 29164
rect 15517 29124 15936 29152
rect 15517 29121 15529 29124
rect 15471 29115 15529 29121
rect 15930 29112 15936 29124
rect 15988 29112 15994 29164
rect 16298 29112 16304 29164
rect 16356 29152 16362 29164
rect 16666 29152 16672 29164
rect 16356 29124 16672 29152
rect 16356 29112 16362 29124
rect 16666 29112 16672 29124
rect 16724 29112 16730 29164
rect 16936 29155 16994 29161
rect 16936 29121 16948 29155
rect 16982 29152 16994 29155
rect 17052 29152 17080 29248
rect 18966 29180 18972 29232
rect 19024 29180 19030 29232
rect 16982 29124 17080 29152
rect 16982 29121 16994 29124
rect 16936 29115 16994 29121
rect 17494 29112 17500 29164
rect 17552 29152 17558 29164
rect 18046 29152 18052 29164
rect 17552 29124 18052 29152
rect 17552 29112 17558 29124
rect 18046 29112 18052 29124
rect 18104 29152 18110 29164
rect 18325 29155 18383 29161
rect 18325 29152 18337 29155
rect 18104 29124 18337 29152
rect 18104 29112 18110 29124
rect 18325 29121 18337 29124
rect 18371 29121 18383 29155
rect 18325 29115 18383 29121
rect 18506 29112 18512 29164
rect 18564 29152 18570 29164
rect 18599 29155 18657 29161
rect 18599 29152 18611 29155
rect 18564 29124 18611 29152
rect 18564 29112 18570 29124
rect 18599 29121 18611 29124
rect 18645 29152 18657 29155
rect 18984 29152 19012 29180
rect 18645 29124 19012 29152
rect 19076 29152 19104 29260
rect 19981 29257 19993 29291
rect 20027 29257 20039 29291
rect 19981 29251 20039 29257
rect 19996 29220 20024 29251
rect 20438 29248 20444 29300
rect 20496 29248 20502 29300
rect 20530 29248 20536 29300
rect 20588 29288 20594 29300
rect 20717 29291 20775 29297
rect 20717 29288 20729 29291
rect 20588 29260 20729 29288
rect 20588 29248 20594 29260
rect 20717 29257 20729 29260
rect 20763 29257 20775 29291
rect 20717 29251 20775 29257
rect 19996 29192 20668 29220
rect 19978 29152 19984 29164
rect 19076 29124 19984 29152
rect 18645 29121 18657 29124
rect 18599 29115 18657 29121
rect 19978 29112 19984 29124
rect 20036 29112 20042 29164
rect 20162 29112 20168 29164
rect 20220 29112 20226 29164
rect 20640 29161 20668 29192
rect 20806 29180 20812 29232
rect 20864 29220 20870 29232
rect 21177 29223 21235 29229
rect 21177 29220 21189 29223
rect 20864 29192 21189 29220
rect 20864 29180 20870 29192
rect 21177 29189 21189 29192
rect 21223 29189 21235 29223
rect 21177 29183 21235 29189
rect 20625 29155 20683 29161
rect 20625 29121 20637 29155
rect 20671 29121 20683 29155
rect 20625 29115 20683 29121
rect 20901 29155 20959 29161
rect 20901 29121 20913 29155
rect 20947 29152 20959 29155
rect 21266 29152 21272 29164
rect 20947 29124 21272 29152
rect 20947 29121 20959 29124
rect 20901 29115 20959 29121
rect 21266 29112 21272 29124
rect 21324 29112 21330 29164
rect 13906 29044 13912 29096
rect 13964 29044 13970 29096
rect 13998 29044 14004 29096
rect 14056 29084 14062 29096
rect 14185 29087 14243 29093
rect 14185 29084 14197 29087
rect 14056 29056 14197 29084
rect 14056 29044 14062 29056
rect 14185 29053 14197 29056
rect 14231 29053 14243 29087
rect 19518 29084 19524 29096
rect 14185 29047 14243 29053
rect 18984 29056 19524 29084
rect 13556 28988 13952 29016
rect 1854 28948 1860 28960
rect 1596 28920 1860 28948
rect 1854 28908 1860 28920
rect 1912 28948 1918 28960
rect 2406 28948 2412 28960
rect 1912 28920 2412 28948
rect 1912 28908 1918 28920
rect 2406 28908 2412 28920
rect 2464 28908 2470 28960
rect 2593 28951 2651 28957
rect 2593 28917 2605 28951
rect 2639 28948 2651 28951
rect 2682 28948 2688 28960
rect 2639 28920 2688 28948
rect 2639 28917 2651 28920
rect 2593 28911 2651 28917
rect 2682 28908 2688 28920
rect 2740 28908 2746 28960
rect 3326 28908 3332 28960
rect 3384 28948 3390 28960
rect 8478 28948 8484 28960
rect 3384 28920 8484 28948
rect 3384 28908 3390 28920
rect 8478 28908 8484 28920
rect 8536 28908 8542 28960
rect 10686 28908 10692 28960
rect 10744 28948 10750 28960
rect 11514 28948 11520 28960
rect 10744 28920 11520 28948
rect 10744 28908 10750 28920
rect 11514 28908 11520 28920
rect 11572 28908 11578 28960
rect 11624 28948 11652 28988
rect 13464 28960 13492 28988
rect 12434 28948 12440 28960
rect 11624 28920 12440 28948
rect 12434 28908 12440 28920
rect 12492 28908 12498 28960
rect 13446 28908 13452 28960
rect 13504 28908 13510 28960
rect 13924 28948 13952 28988
rect 15856 28988 16712 29016
rect 15856 28948 15884 28988
rect 13924 28920 15884 28948
rect 16206 28908 16212 28960
rect 16264 28908 16270 28960
rect 16684 28948 16712 28988
rect 17602 28988 18460 29016
rect 17602 28948 17630 28988
rect 16684 28920 17630 28948
rect 18432 28948 18460 28988
rect 18984 28948 19012 29056
rect 19518 29044 19524 29056
rect 19576 29044 19582 29096
rect 19702 29044 19708 29096
rect 19760 29084 19766 29096
rect 22186 29084 22192 29096
rect 19760 29056 22192 29084
rect 19760 29044 19766 29056
rect 22186 29044 22192 29056
rect 22244 29044 22250 29096
rect 18432 28920 19012 28948
rect 19337 28951 19395 28957
rect 19337 28917 19349 28951
rect 19383 28948 19395 28951
rect 19518 28948 19524 28960
rect 19383 28920 19524 28948
rect 19383 28917 19395 28920
rect 19337 28911 19395 28917
rect 19518 28908 19524 28920
rect 19576 28908 19582 28960
rect 21450 28908 21456 28960
rect 21508 28908 21514 28960
rect 1104 28858 21896 28880
rect 1104 28806 3549 28858
rect 3601 28806 3613 28858
rect 3665 28806 3677 28858
rect 3729 28806 3741 28858
rect 3793 28806 3805 28858
rect 3857 28806 8747 28858
rect 8799 28806 8811 28858
rect 8863 28806 8875 28858
rect 8927 28806 8939 28858
rect 8991 28806 9003 28858
rect 9055 28806 13945 28858
rect 13997 28806 14009 28858
rect 14061 28806 14073 28858
rect 14125 28806 14137 28858
rect 14189 28806 14201 28858
rect 14253 28806 19143 28858
rect 19195 28806 19207 28858
rect 19259 28806 19271 28858
rect 19323 28806 19335 28858
rect 19387 28806 19399 28858
rect 19451 28806 21896 28858
rect 1104 28784 21896 28806
rect 1581 28747 1639 28753
rect 1581 28713 1593 28747
rect 1627 28744 1639 28747
rect 3326 28744 3332 28756
rect 1627 28716 3332 28744
rect 1627 28713 1639 28716
rect 1581 28707 1639 28713
rect 3326 28704 3332 28716
rect 3384 28704 3390 28756
rect 3786 28704 3792 28756
rect 3844 28744 3850 28756
rect 3844 28716 5304 28744
rect 3844 28704 3850 28716
rect 1854 28636 1860 28688
rect 1912 28676 1918 28688
rect 5166 28676 5172 28688
rect 1912 28648 2268 28676
rect 1912 28636 1918 28648
rect 2240 28617 2268 28648
rect 5092 28648 5172 28676
rect 2225 28611 2283 28617
rect 1596 28580 2176 28608
rect 1596 28552 1624 28580
rect 750 28500 756 28552
rect 808 28540 814 28552
rect 1489 28543 1547 28549
rect 1489 28540 1501 28543
rect 808 28512 1501 28540
rect 808 28500 814 28512
rect 1489 28509 1501 28512
rect 1535 28509 1547 28543
rect 1489 28503 1547 28509
rect 1578 28500 1584 28552
rect 1636 28500 1642 28552
rect 1762 28500 1768 28552
rect 1820 28500 1826 28552
rect 2148 28540 2176 28580
rect 2225 28577 2237 28611
rect 2271 28577 2283 28611
rect 2225 28571 2283 28577
rect 3142 28568 3148 28620
rect 3200 28608 3206 28620
rect 3881 28611 3939 28617
rect 3881 28608 3893 28611
rect 3200 28580 3893 28608
rect 3200 28568 3206 28580
rect 3881 28577 3893 28580
rect 3927 28577 3939 28611
rect 3881 28571 3939 28577
rect 2498 28549 2504 28552
rect 2467 28543 2504 28549
rect 2467 28540 2479 28543
rect 2148 28512 2479 28540
rect 2467 28509 2479 28512
rect 2467 28503 2504 28509
rect 2498 28500 2504 28503
rect 2556 28500 2562 28552
rect 2866 28500 2872 28552
rect 2924 28540 2930 28552
rect 4123 28543 4181 28549
rect 4123 28540 4135 28543
rect 2924 28512 4135 28540
rect 2924 28500 2930 28512
rect 4123 28509 4135 28512
rect 4169 28540 4181 28543
rect 5092 28540 5120 28648
rect 5166 28636 5172 28648
rect 5224 28636 5230 28688
rect 5276 28617 5304 28716
rect 5368 28716 10362 28744
rect 5261 28611 5319 28617
rect 5261 28577 5273 28611
rect 5307 28577 5319 28611
rect 5261 28571 5319 28577
rect 4169 28512 5120 28540
rect 4169 28509 4181 28512
rect 4123 28503 4181 28509
rect 5166 28500 5172 28552
rect 5224 28540 5230 28552
rect 5368 28540 5396 28716
rect 7834 28636 7840 28688
rect 7892 28636 7898 28688
rect 8110 28636 8116 28688
rect 8168 28636 8174 28688
rect 10334 28676 10362 28716
rect 10410 28704 10416 28756
rect 10468 28744 10474 28756
rect 10689 28747 10747 28753
rect 10689 28744 10701 28747
rect 10468 28716 10701 28744
rect 10468 28704 10474 28716
rect 10689 28713 10701 28716
rect 10735 28713 10747 28747
rect 15194 28744 15200 28756
rect 10689 28707 10747 28713
rect 10796 28716 15200 28744
rect 10796 28676 10824 28716
rect 15194 28704 15200 28716
rect 15252 28704 15258 28756
rect 15286 28704 15292 28756
rect 15344 28744 15350 28756
rect 17037 28747 17095 28753
rect 17037 28744 17049 28747
rect 15344 28716 17049 28744
rect 15344 28704 15350 28716
rect 17037 28713 17049 28716
rect 17083 28713 17095 28747
rect 18046 28744 18052 28756
rect 17037 28707 17095 28713
rect 17696 28716 18052 28744
rect 10334 28648 10824 28676
rect 12158 28636 12164 28688
rect 12216 28676 12222 28688
rect 12526 28676 12532 28688
rect 12216 28648 12532 28676
rect 12216 28636 12222 28648
rect 12526 28636 12532 28648
rect 12584 28636 12590 28688
rect 14366 28636 14372 28688
rect 14424 28676 14430 28688
rect 14424 28648 14854 28676
rect 14424 28636 14430 28648
rect 5534 28568 5540 28620
rect 5592 28568 5598 28620
rect 7852 28608 7880 28636
rect 9030 28608 9036 28620
rect 7852 28580 9036 28608
rect 9030 28568 9036 28580
rect 9088 28568 9094 28620
rect 9677 28611 9735 28617
rect 9677 28608 9689 28611
rect 9508 28580 9689 28608
rect 5224 28512 5396 28540
rect 5224 28500 5230 28512
rect 7098 28500 7104 28552
rect 7156 28500 7162 28552
rect 7282 28500 7288 28552
rect 7340 28540 7346 28552
rect 7375 28543 7433 28549
rect 7375 28540 7387 28543
rect 7340 28512 7387 28540
rect 7340 28500 7346 28512
rect 7375 28509 7387 28512
rect 7421 28540 7433 28543
rect 7834 28540 7840 28552
rect 7421 28512 7840 28540
rect 7421 28509 7433 28512
rect 7375 28503 7433 28509
rect 7834 28500 7840 28512
rect 7892 28500 7898 28552
rect 8846 28500 8852 28552
rect 8904 28540 8910 28552
rect 9508 28540 9536 28580
rect 9677 28577 9689 28580
rect 9723 28577 9735 28611
rect 9677 28571 9735 28577
rect 13446 28568 13452 28620
rect 13504 28608 13510 28620
rect 14277 28611 14335 28617
rect 14277 28608 14289 28611
rect 13504 28580 14289 28608
rect 13504 28568 13510 28580
rect 14277 28577 14289 28580
rect 14323 28577 14335 28611
rect 14277 28571 14335 28577
rect 14734 28568 14740 28620
rect 14792 28568 14798 28620
rect 14826 28608 14854 28648
rect 16942 28636 16948 28688
rect 17000 28676 17006 28688
rect 17696 28676 17724 28716
rect 18046 28704 18052 28716
rect 18104 28704 18110 28756
rect 19061 28747 19119 28753
rect 19061 28713 19073 28747
rect 19107 28744 19119 28747
rect 19107 28716 20392 28744
rect 19107 28713 19119 28716
rect 19061 28707 19119 28713
rect 17000 28648 17724 28676
rect 17000 28636 17006 28648
rect 15130 28611 15188 28617
rect 15130 28608 15142 28611
rect 14826 28580 15142 28608
rect 15130 28577 15142 28580
rect 15176 28577 15188 28611
rect 15130 28571 15188 28577
rect 15838 28568 15844 28620
rect 15896 28608 15902 28620
rect 17696 28617 17724 28648
rect 19794 28636 19800 28688
rect 19852 28676 19858 28688
rect 20162 28676 20168 28688
rect 19852 28648 20168 28676
rect 19852 28636 19858 28648
rect 20162 28636 20168 28648
rect 20220 28636 20226 28688
rect 15933 28611 15991 28617
rect 15933 28608 15945 28611
rect 15896 28580 15945 28608
rect 15896 28568 15902 28580
rect 15933 28577 15945 28580
rect 15979 28577 15991 28611
rect 15933 28571 15991 28577
rect 17681 28611 17739 28617
rect 17681 28577 17693 28611
rect 17727 28577 17739 28611
rect 19521 28611 19579 28617
rect 17681 28571 17739 28577
rect 19168 28580 19472 28608
rect 8904 28512 9536 28540
rect 9919 28543 9977 28549
rect 8904 28500 8910 28512
rect 9919 28509 9931 28543
rect 9965 28540 9977 28543
rect 9965 28510 9996 28540
rect 9965 28509 10070 28510
rect 9919 28503 10070 28509
rect 1854 28472 1860 28484
rect 1596 28444 1860 28472
rect 1596 28416 1624 28444
rect 1854 28432 1860 28444
rect 1912 28432 1918 28484
rect 9306 28472 9312 28484
rect 1964 28444 9312 28472
rect 1578 28364 1584 28416
rect 1636 28364 1642 28416
rect 1964 28413 1992 28444
rect 9306 28432 9312 28444
rect 9364 28432 9370 28484
rect 9968 28482 10070 28503
rect 11054 28500 11060 28552
rect 11112 28540 11118 28552
rect 11425 28543 11483 28549
rect 11425 28540 11437 28543
rect 11112 28512 11437 28540
rect 11112 28500 11118 28512
rect 11425 28509 11437 28512
rect 11471 28509 11483 28543
rect 11425 28503 11483 28509
rect 11606 28500 11612 28552
rect 11664 28540 11670 28552
rect 11699 28543 11757 28549
rect 11699 28540 11711 28543
rect 11664 28512 11711 28540
rect 11664 28500 11670 28512
rect 11699 28509 11711 28512
rect 11745 28540 11757 28543
rect 13998 28540 14004 28552
rect 11745 28512 14004 28540
rect 11745 28509 11757 28512
rect 11699 28503 11757 28509
rect 13998 28500 14004 28512
rect 14056 28500 14062 28552
rect 14093 28543 14151 28549
rect 14093 28509 14105 28543
rect 14139 28509 14151 28543
rect 14093 28503 14151 28509
rect 10042 28472 10070 28482
rect 10134 28472 10140 28484
rect 10042 28444 10140 28472
rect 10134 28432 10140 28444
rect 10192 28432 10198 28484
rect 13262 28432 13268 28484
rect 13320 28472 13326 28484
rect 14108 28472 14136 28503
rect 15010 28500 15016 28552
rect 15068 28500 15074 28552
rect 15286 28500 15292 28552
rect 15344 28500 15350 28552
rect 16022 28500 16028 28552
rect 16080 28500 16086 28552
rect 16206 28500 16212 28552
rect 16264 28540 16270 28552
rect 16299 28543 16357 28549
rect 16299 28540 16311 28543
rect 16264 28512 16311 28540
rect 16264 28500 16270 28512
rect 16299 28509 16311 28512
rect 16345 28509 16357 28543
rect 16299 28503 16357 28509
rect 17218 28500 17224 28552
rect 17276 28540 17282 28552
rect 17405 28543 17463 28549
rect 17405 28540 17417 28543
rect 17276 28512 17417 28540
rect 17276 28500 17282 28512
rect 17405 28509 17417 28512
rect 17451 28509 17463 28543
rect 19168 28540 19196 28580
rect 17405 28503 17463 28509
rect 17972 28512 19196 28540
rect 19245 28543 19303 28549
rect 17972 28481 18000 28512
rect 19245 28509 19257 28543
rect 19291 28509 19303 28543
rect 19245 28503 19303 28509
rect 17926 28475 18000 28481
rect 17926 28472 17938 28475
rect 13320 28444 14136 28472
rect 15948 28444 16252 28472
rect 13320 28432 13326 28444
rect 1949 28407 2007 28413
rect 1949 28373 1961 28407
rect 1995 28373 2007 28407
rect 1949 28367 2007 28373
rect 2498 28364 2504 28416
rect 2556 28404 2562 28416
rect 3237 28407 3295 28413
rect 3237 28404 3249 28407
rect 2556 28376 3249 28404
rect 2556 28364 2562 28376
rect 3237 28373 3249 28376
rect 3283 28373 3295 28407
rect 3237 28367 3295 28373
rect 3694 28364 3700 28416
rect 3752 28404 3758 28416
rect 3970 28404 3976 28416
rect 3752 28376 3976 28404
rect 3752 28364 3758 28376
rect 3970 28364 3976 28376
rect 4028 28364 4034 28416
rect 4246 28364 4252 28416
rect 4304 28404 4310 28416
rect 4614 28404 4620 28416
rect 4304 28376 4620 28404
rect 4304 28364 4310 28376
rect 4614 28364 4620 28376
rect 4672 28364 4678 28416
rect 4890 28364 4896 28416
rect 4948 28364 4954 28416
rect 5534 28364 5540 28416
rect 5592 28404 5598 28416
rect 8478 28404 8484 28416
rect 5592 28376 8484 28404
rect 5592 28364 5598 28376
rect 8478 28364 8484 28376
rect 8536 28364 8542 28416
rect 8662 28364 8668 28416
rect 8720 28404 8726 28416
rect 10410 28404 10416 28416
rect 8720 28376 10416 28404
rect 8720 28364 8726 28376
rect 10410 28364 10416 28376
rect 10468 28364 10474 28416
rect 11238 28364 11244 28416
rect 11296 28404 11302 28416
rect 12250 28404 12256 28416
rect 11296 28376 12256 28404
rect 11296 28364 11302 28376
rect 12250 28364 12256 28376
rect 12308 28364 12314 28416
rect 12437 28407 12495 28413
rect 12437 28373 12449 28407
rect 12483 28404 12495 28407
rect 12618 28404 12624 28416
rect 12483 28376 12624 28404
rect 12483 28373 12495 28376
rect 12437 28367 12495 28373
rect 12618 28364 12624 28376
rect 12676 28364 12682 28416
rect 15838 28364 15844 28416
rect 15896 28404 15902 28416
rect 15948 28404 15976 28444
rect 15896 28376 15976 28404
rect 16224 28404 16252 28444
rect 16684 28444 17938 28472
rect 16684 28404 16712 28444
rect 17926 28441 17938 28444
rect 17972 28444 18000 28475
rect 19260 28472 19288 28503
rect 19334 28500 19340 28552
rect 19392 28500 19398 28552
rect 19444 28540 19472 28580
rect 19521 28577 19533 28611
rect 19567 28608 19579 28611
rect 19981 28611 20039 28617
rect 19981 28608 19993 28611
rect 19567 28580 19993 28608
rect 19567 28577 19579 28580
rect 19521 28571 19579 28577
rect 19981 28577 19993 28580
rect 20027 28577 20039 28611
rect 19981 28571 20039 28577
rect 20364 28549 20392 28716
rect 20530 28568 20536 28620
rect 20588 28608 20594 28620
rect 20588 28580 21220 28608
rect 20588 28568 20594 28580
rect 19797 28543 19855 28549
rect 19797 28540 19809 28543
rect 19444 28512 19809 28540
rect 19797 28509 19809 28512
rect 19843 28509 19855 28543
rect 19797 28503 19855 28509
rect 19889 28543 19947 28549
rect 19889 28509 19901 28543
rect 19935 28509 19947 28543
rect 19889 28503 19947 28509
rect 20073 28543 20131 28549
rect 20073 28509 20085 28543
rect 20119 28540 20131 28543
rect 20349 28543 20407 28549
rect 20119 28512 20208 28540
rect 20119 28509 20131 28512
rect 20073 28503 20131 28509
rect 19426 28472 19432 28484
rect 19260 28444 19432 28472
rect 17972 28441 17984 28444
rect 17926 28435 17984 28441
rect 19426 28432 19432 28444
rect 19484 28472 19490 28484
rect 19904 28472 19932 28503
rect 19484 28444 19932 28472
rect 19484 28432 19490 28444
rect 16224 28376 16712 28404
rect 15896 28364 15902 28376
rect 17494 28364 17500 28416
rect 17552 28364 17558 28416
rect 19518 28364 19524 28416
rect 19576 28364 19582 28416
rect 19610 28364 19616 28416
rect 19668 28364 19674 28416
rect 20180 28413 20208 28512
rect 20349 28509 20361 28543
rect 20395 28509 20407 28543
rect 20349 28503 20407 28509
rect 20622 28500 20628 28552
rect 20680 28500 20686 28552
rect 20901 28543 20959 28549
rect 20901 28509 20913 28543
rect 20947 28509 20959 28543
rect 20901 28503 20959 28509
rect 20916 28472 20944 28503
rect 20990 28500 20996 28552
rect 21048 28500 21054 28552
rect 21192 28549 21220 28580
rect 21177 28543 21235 28549
rect 21177 28509 21189 28543
rect 21223 28509 21235 28543
rect 21177 28503 21235 28509
rect 21269 28543 21327 28549
rect 21269 28509 21281 28543
rect 21315 28509 21327 28543
rect 21269 28503 21327 28509
rect 20456 28444 20944 28472
rect 21008 28472 21036 28500
rect 21284 28472 21312 28503
rect 21008 28444 21312 28472
rect 20456 28413 20484 28444
rect 20165 28407 20223 28413
rect 20165 28373 20177 28407
rect 20211 28373 20223 28407
rect 20165 28367 20223 28373
rect 20441 28407 20499 28413
rect 20441 28373 20453 28407
rect 20487 28373 20499 28407
rect 20441 28367 20499 28373
rect 20714 28364 20720 28416
rect 20772 28364 20778 28416
rect 20990 28364 20996 28416
rect 21048 28364 21054 28416
rect 21453 28407 21511 28413
rect 21453 28373 21465 28407
rect 21499 28404 21511 28407
rect 22186 28404 22192 28416
rect 21499 28376 22192 28404
rect 21499 28373 21511 28376
rect 21453 28367 21511 28373
rect 22186 28364 22192 28376
rect 22244 28364 22250 28416
rect 1104 28314 22056 28336
rect 1104 28262 6148 28314
rect 6200 28262 6212 28314
rect 6264 28262 6276 28314
rect 6328 28262 6340 28314
rect 6392 28262 6404 28314
rect 6456 28262 11346 28314
rect 11398 28262 11410 28314
rect 11462 28262 11474 28314
rect 11526 28262 11538 28314
rect 11590 28262 11602 28314
rect 11654 28262 16544 28314
rect 16596 28262 16608 28314
rect 16660 28262 16672 28314
rect 16724 28262 16736 28314
rect 16788 28262 16800 28314
rect 16852 28262 21742 28314
rect 21794 28262 21806 28314
rect 21858 28262 21870 28314
rect 21922 28262 21934 28314
rect 21986 28262 21998 28314
rect 22050 28262 22056 28314
rect 1104 28240 22056 28262
rect 2317 28203 2375 28209
rect 2317 28169 2329 28203
rect 2363 28200 2375 28203
rect 3326 28200 3332 28212
rect 2363 28172 3332 28200
rect 2363 28169 2375 28172
rect 2317 28163 2375 28169
rect 3326 28160 3332 28172
rect 3384 28160 3390 28212
rect 3605 28203 3663 28209
rect 3605 28169 3617 28203
rect 3651 28200 3663 28203
rect 5166 28200 5172 28212
rect 3651 28172 5172 28200
rect 3651 28169 3663 28172
rect 3605 28163 3663 28169
rect 5166 28160 5172 28172
rect 5224 28160 5230 28212
rect 5261 28203 5319 28209
rect 5261 28169 5273 28203
rect 5307 28200 5319 28203
rect 8938 28200 8944 28212
rect 5307 28172 8944 28200
rect 5307 28169 5319 28172
rect 5261 28163 5319 28169
rect 8938 28160 8944 28172
rect 8996 28160 9002 28212
rect 9030 28160 9036 28212
rect 9088 28200 9094 28212
rect 9088 28172 9410 28200
rect 9088 28160 9094 28172
rect 2498 28092 2504 28144
rect 2556 28132 2562 28144
rect 2685 28135 2743 28141
rect 2685 28132 2697 28135
rect 2556 28104 2697 28132
rect 2556 28092 2562 28104
rect 2685 28101 2697 28104
rect 2731 28101 2743 28135
rect 3421 28135 3479 28141
rect 2685 28095 2743 28101
rect 2792 28104 3188 28132
rect 750 28024 756 28076
rect 808 28064 814 28076
rect 1489 28067 1547 28073
rect 1489 28064 1501 28067
rect 808 28036 1501 28064
rect 808 28024 814 28036
rect 1489 28033 1501 28036
rect 1535 28033 1547 28067
rect 1489 28027 1547 28033
rect 1670 28024 1676 28076
rect 1728 28024 1734 28076
rect 1946 28024 1952 28076
rect 2004 28024 2010 28076
rect 2593 28067 2651 28073
rect 2593 28033 2605 28067
rect 2639 28064 2651 28067
rect 2792 28064 2820 28104
rect 2639 28036 2820 28064
rect 2639 28033 2651 28036
rect 2593 28027 2651 28033
rect 2866 28024 2872 28076
rect 2924 28064 2930 28076
rect 3053 28067 3111 28073
rect 3053 28064 3065 28067
rect 2924 28036 3065 28064
rect 2924 28024 2930 28036
rect 3053 28033 3065 28036
rect 3099 28033 3111 28067
rect 3160 28064 3188 28104
rect 3421 28101 3433 28135
rect 3467 28132 3479 28135
rect 3878 28132 3884 28144
rect 3467 28104 3884 28132
rect 3467 28101 3479 28104
rect 3421 28095 3479 28101
rect 3878 28092 3884 28104
rect 3936 28092 3942 28144
rect 3973 28135 4031 28141
rect 3973 28101 3985 28135
rect 4019 28101 4031 28135
rect 3973 28095 4031 28101
rect 4341 28135 4399 28141
rect 4341 28101 4353 28135
rect 4387 28132 4399 28135
rect 4890 28132 4896 28144
rect 4387 28104 4896 28132
rect 4387 28101 4399 28104
rect 4341 28095 4399 28101
rect 3602 28064 3608 28076
rect 3160 28036 3608 28064
rect 3053 28027 3111 28033
rect 3602 28024 3608 28036
rect 3660 28024 3666 28076
rect 3694 28024 3700 28076
rect 3752 28064 3758 28076
rect 3988 28064 4016 28095
rect 4890 28092 4896 28104
rect 4948 28092 4954 28144
rect 5077 28135 5135 28141
rect 5077 28101 5089 28135
rect 5123 28132 5135 28135
rect 5123 28104 5212 28132
rect 5123 28101 5135 28104
rect 5077 28095 5135 28101
rect 5184 28076 5212 28104
rect 7650 28092 7656 28144
rect 7708 28132 7714 28144
rect 7708 28104 7880 28132
rect 7708 28092 7714 28104
rect 7852 28094 7880 28104
rect 7911 28097 7969 28103
rect 7911 28094 7923 28097
rect 3752 28036 4016 28064
rect 3752 28024 3758 28036
rect 4062 28024 4068 28076
rect 4120 28024 4126 28076
rect 4249 28067 4307 28073
rect 4249 28033 4261 28067
rect 4295 28064 4307 28067
rect 4522 28064 4528 28076
rect 4295 28036 4528 28064
rect 4295 28033 4307 28036
rect 4249 28027 4307 28033
rect 4522 28024 4528 28036
rect 4580 28024 4586 28076
rect 4709 28067 4767 28073
rect 4709 28033 4721 28067
rect 4755 28064 4767 28067
rect 4798 28064 4804 28076
rect 4755 28036 4804 28064
rect 4755 28033 4767 28036
rect 4709 28027 4767 28033
rect 4798 28024 4804 28036
rect 4856 28024 4862 28076
rect 5166 28024 5172 28076
rect 5224 28024 5230 28076
rect 7852 28066 7923 28094
rect 7911 28063 7923 28066
rect 7957 28063 7969 28097
rect 8570 28092 8576 28144
rect 8628 28132 8634 28144
rect 8628 28104 9168 28132
rect 8628 28092 8634 28104
rect 7911 28057 7969 28063
rect 8846 28024 8852 28076
rect 8904 28024 8910 28076
rect 9140 28064 9168 28104
rect 9275 28077 9333 28083
rect 9275 28074 9287 28077
rect 9198 28064 9287 28074
rect 9140 28046 9287 28064
rect 9140 28036 9226 28046
rect 9275 28043 9287 28046
rect 9321 28043 9333 28077
rect 9275 28037 9333 28043
rect 9382 28064 9410 28172
rect 9582 28160 9588 28212
rect 9640 28200 9646 28212
rect 10045 28203 10103 28209
rect 10045 28200 10057 28203
rect 9640 28172 10057 28200
rect 9640 28160 9646 28172
rect 10045 28169 10057 28172
rect 10091 28169 10103 28203
rect 10045 28163 10103 28169
rect 10318 28160 10324 28212
rect 10376 28200 10382 28212
rect 10962 28200 10968 28212
rect 10376 28172 10968 28200
rect 10376 28160 10382 28172
rect 10962 28160 10968 28172
rect 11020 28160 11026 28212
rect 11808 28172 12020 28200
rect 9490 28092 9496 28144
rect 9548 28132 9554 28144
rect 11808 28132 11836 28172
rect 9548 28104 11836 28132
rect 11992 28132 12020 28172
rect 13906 28160 13912 28212
rect 13964 28200 13970 28212
rect 15654 28200 15660 28212
rect 13964 28172 15660 28200
rect 13964 28160 13970 28172
rect 15654 28160 15660 28172
rect 15712 28200 15718 28212
rect 15712 28172 16970 28200
rect 15712 28160 15718 28172
rect 15838 28132 15844 28144
rect 11992 28104 15844 28132
rect 9548 28092 9554 28104
rect 15838 28092 15844 28104
rect 15896 28092 15902 28144
rect 15930 28092 15936 28144
rect 15988 28092 15994 28144
rect 10134 28064 10140 28076
rect 9382 28036 10140 28064
rect 10134 28024 10140 28036
rect 10192 28024 10198 28076
rect 11883 28067 11941 28073
rect 11883 28033 11895 28067
rect 11929 28064 11941 28067
rect 13906 28064 13912 28076
rect 11929 28036 13912 28064
rect 11929 28033 11941 28036
rect 11883 28027 11941 28033
rect 13906 28024 13912 28036
rect 13964 28024 13970 28076
rect 14182 28024 14188 28076
rect 14240 28064 14246 28076
rect 14275 28067 14333 28073
rect 14275 28064 14287 28067
rect 14240 28036 14287 28064
rect 14240 28024 14246 28036
rect 14275 28033 14287 28036
rect 14321 28064 14333 28067
rect 14642 28064 14648 28076
rect 14321 28036 14648 28064
rect 14321 28033 14333 28036
rect 14275 28027 14333 28033
rect 14642 28024 14648 28036
rect 14700 28024 14706 28076
rect 15948 28064 15976 28092
rect 16393 28067 16451 28073
rect 16393 28064 16405 28067
rect 15948 28036 16405 28064
rect 16393 28033 16405 28036
rect 16439 28033 16451 28067
rect 16393 28027 16451 28033
rect 16853 28067 16911 28073
rect 16853 28033 16865 28067
rect 16899 28033 16911 28067
rect 16942 28064 16970 28172
rect 17034 28160 17040 28212
rect 17092 28160 17098 28212
rect 17494 28160 17500 28212
rect 17552 28200 17558 28212
rect 17552 28172 17908 28200
rect 17552 28160 17558 28172
rect 17880 28132 17908 28172
rect 17954 28160 17960 28212
rect 18012 28200 18018 28212
rect 19245 28203 19303 28209
rect 18012 28172 19104 28200
rect 18012 28160 18018 28172
rect 17880 28104 18644 28132
rect 18616 28073 18644 28104
rect 19076 28073 19104 28172
rect 19245 28169 19257 28203
rect 19291 28200 19303 28203
rect 19334 28200 19340 28212
rect 19291 28172 19340 28200
rect 19291 28169 19303 28172
rect 19245 28163 19303 28169
rect 19334 28160 19340 28172
rect 19392 28160 19398 28212
rect 19610 28160 19616 28212
rect 19668 28160 19674 28212
rect 19981 28203 20039 28209
rect 19981 28169 19993 28203
rect 20027 28169 20039 28203
rect 19981 28163 20039 28169
rect 20349 28203 20407 28209
rect 20349 28169 20361 28203
rect 20395 28200 20407 28203
rect 20530 28200 20536 28212
rect 20395 28172 20536 28200
rect 20395 28169 20407 28172
rect 20349 28163 20407 28169
rect 19628 28132 19656 28160
rect 19168 28104 19656 28132
rect 19996 28132 20024 28163
rect 20530 28160 20536 28172
rect 20588 28160 20594 28212
rect 20622 28160 20628 28212
rect 20680 28160 20686 28212
rect 20714 28160 20720 28212
rect 20772 28160 20778 28212
rect 19996 28104 20576 28132
rect 19168 28073 19196 28104
rect 17371 28067 17429 28073
rect 17371 28064 17383 28067
rect 16942 28036 17383 28064
rect 16853 28027 16911 28033
rect 17371 28033 17383 28036
rect 17417 28033 17429 28067
rect 18509 28067 18567 28073
rect 18509 28064 18521 28067
rect 17371 28027 17429 28033
rect 18156 28036 18521 28064
rect 1688 27996 1716 28024
rect 768 27968 1716 27996
rect 768 27736 796 27968
rect 2682 27956 2688 28008
rect 2740 27956 2746 28008
rect 1670 27888 1676 27940
rect 1728 27888 1734 27940
rect 3712 27928 3740 28024
rect 4080 27982 4108 28024
rect 7282 27956 7288 28008
rect 7340 27996 7346 28008
rect 7653 27999 7711 28005
rect 7653 27996 7665 27999
rect 7340 27968 7665 27996
rect 7340 27956 7346 27968
rect 7653 27965 7665 27968
rect 7699 27965 7711 27999
rect 7653 27959 7711 27965
rect 8662 27956 8668 28008
rect 8720 27996 8726 28008
rect 8864 27996 8892 28024
rect 9033 27999 9091 28005
rect 9033 27996 9045 27999
rect 8720 27968 9045 27996
rect 8720 27956 8726 27968
rect 9033 27965 9045 27968
rect 9079 27965 9091 27999
rect 9033 27959 9091 27965
rect 9766 27956 9772 28008
rect 9824 27996 9830 28008
rect 11054 27996 11060 28008
rect 9824 27968 11060 27996
rect 9824 27956 9830 27968
rect 11054 27956 11060 27968
rect 11112 27996 11118 28008
rect 11609 27999 11667 28005
rect 11609 27996 11621 27999
rect 11112 27968 11621 27996
rect 11112 27956 11118 27968
rect 11609 27965 11621 27968
rect 11655 27965 11667 27999
rect 11609 27959 11667 27965
rect 14001 27999 14059 28005
rect 14001 27965 14013 27999
rect 14047 27965 14059 27999
rect 14001 27959 14059 27965
rect 3712 27900 3924 27928
rect 3896 27872 3924 27900
rect 8478 27888 8484 27940
rect 8536 27928 8542 27940
rect 8536 27900 9168 27928
rect 8536 27888 8542 27900
rect 1765 27863 1823 27869
rect 1765 27829 1777 27863
rect 1811 27860 1823 27863
rect 2314 27860 2320 27872
rect 1811 27832 2320 27860
rect 1811 27829 1823 27832
rect 1765 27823 1823 27829
rect 2314 27820 2320 27832
rect 2372 27820 2378 27872
rect 3878 27820 3884 27872
rect 3936 27820 3942 27872
rect 5258 27820 5264 27872
rect 5316 27860 5322 27872
rect 5994 27860 6000 27872
rect 5316 27832 6000 27860
rect 5316 27820 5322 27832
rect 5994 27820 6000 27832
rect 6052 27820 6058 27872
rect 7742 27820 7748 27872
rect 7800 27860 7806 27872
rect 8665 27863 8723 27869
rect 8665 27860 8677 27863
rect 7800 27832 8677 27860
rect 7800 27820 7806 27832
rect 8665 27829 8677 27832
rect 8711 27829 8723 27863
rect 9140 27860 9168 27900
rect 11238 27860 11244 27872
rect 9140 27832 11244 27860
rect 8665 27823 8723 27829
rect 11238 27820 11244 27832
rect 11296 27820 11302 27872
rect 11882 27820 11888 27872
rect 11940 27860 11946 27872
rect 12621 27863 12679 27869
rect 12621 27860 12633 27863
rect 11940 27832 12633 27860
rect 11940 27820 11946 27832
rect 12621 27829 12633 27832
rect 12667 27829 12679 27863
rect 14016 27860 14044 27959
rect 16206 27956 16212 28008
rect 16264 27996 16270 28008
rect 16868 27996 16896 28027
rect 16264 27968 16896 27996
rect 16264 27956 16270 27968
rect 17034 27956 17040 28008
rect 17092 27996 17098 28008
rect 17129 27999 17187 28005
rect 17129 27996 17141 27999
rect 17092 27968 17141 27996
rect 17092 27956 17098 27968
rect 17129 27965 17141 27968
rect 17175 27965 17187 27999
rect 17129 27959 17187 27965
rect 15194 27888 15200 27940
rect 15252 27928 15258 27940
rect 18156 27937 18184 28036
rect 18509 28033 18521 28036
rect 18555 28033 18567 28067
rect 18509 28027 18567 28033
rect 18601 28067 18659 28073
rect 18601 28033 18613 28067
rect 18647 28033 18659 28067
rect 18877 28067 18935 28073
rect 18877 28064 18889 28067
rect 18601 28027 18659 28033
rect 18708 28036 18889 28064
rect 18524 27996 18552 28027
rect 18708 27996 18736 28036
rect 18877 28033 18889 28036
rect 18923 28033 18935 28067
rect 18877 28027 18935 28033
rect 19061 28067 19119 28073
rect 19061 28033 19073 28067
rect 19107 28033 19119 28067
rect 19061 28027 19119 28033
rect 19153 28067 19211 28073
rect 19153 28033 19165 28067
rect 19199 28033 19211 28067
rect 19153 28027 19211 28033
rect 19610 28024 19616 28076
rect 19668 28024 19674 28076
rect 19889 28067 19947 28073
rect 19889 28033 19901 28067
rect 19935 28033 19947 28067
rect 19889 28027 19947 28033
rect 18524 27968 18736 27996
rect 18785 27999 18843 28005
rect 18785 27965 18797 27999
rect 18831 27996 18843 27999
rect 18969 27999 19027 28005
rect 18969 27996 18981 27999
rect 18831 27968 18981 27996
rect 18831 27965 18843 27968
rect 18785 27959 18843 27965
rect 18969 27965 18981 27968
rect 19015 27965 19027 27999
rect 19904 27996 19932 28027
rect 20162 28024 20168 28076
rect 20220 28024 20226 28076
rect 20548 28073 20576 28104
rect 20533 28067 20591 28073
rect 20533 28033 20545 28067
rect 20579 28033 20591 28067
rect 20533 28027 20591 28033
rect 18969 27959 19027 27965
rect 19352 27968 19932 27996
rect 18141 27931 18199 27937
rect 15252 27900 16528 27928
rect 15252 27888 15258 27900
rect 14366 27860 14372 27872
rect 14016 27832 14372 27860
rect 12621 27823 12679 27829
rect 14366 27820 14372 27832
rect 14424 27820 14430 27872
rect 15013 27863 15071 27869
rect 15013 27829 15025 27863
rect 15059 27860 15071 27863
rect 15286 27860 15292 27872
rect 15059 27832 15292 27860
rect 15059 27829 15071 27832
rect 15013 27823 15071 27829
rect 15286 27820 15292 27832
rect 15344 27820 15350 27872
rect 16209 27863 16267 27869
rect 16209 27829 16221 27863
rect 16255 27860 16267 27863
rect 16390 27860 16396 27872
rect 16255 27832 16396 27860
rect 16255 27829 16267 27832
rect 16209 27823 16267 27829
rect 16390 27820 16396 27832
rect 16448 27820 16454 27872
rect 16500 27860 16528 27900
rect 18141 27897 18153 27931
rect 18187 27897 18199 27931
rect 19058 27928 19064 27940
rect 18141 27891 18199 27897
rect 18616 27900 19064 27928
rect 18616 27860 18644 27900
rect 19058 27888 19064 27900
rect 19116 27928 19122 27940
rect 19352 27928 19380 27968
rect 19116 27900 19380 27928
rect 19429 27931 19487 27937
rect 19116 27888 19122 27900
rect 19429 27897 19441 27931
rect 19475 27928 19487 27931
rect 20640 27928 20668 28160
rect 20732 28132 20760 28160
rect 20732 28104 20944 28132
rect 20806 28024 20812 28076
rect 20864 28024 20870 28076
rect 20916 28073 20944 28104
rect 20901 28067 20959 28073
rect 20901 28033 20913 28067
rect 20947 28033 20959 28067
rect 20901 28027 20959 28033
rect 21266 28024 21272 28076
rect 21324 28024 21330 28076
rect 19475 27900 20668 27928
rect 19475 27897 19487 27900
rect 19429 27891 19487 27897
rect 16500 27832 18644 27860
rect 18693 27863 18751 27869
rect 18693 27829 18705 27863
rect 18739 27860 18751 27863
rect 19610 27860 19616 27872
rect 18739 27832 19616 27860
rect 18739 27829 18751 27832
rect 18693 27823 18751 27829
rect 19610 27820 19616 27832
rect 19668 27820 19674 27872
rect 19705 27863 19763 27869
rect 19705 27829 19717 27863
rect 19751 27860 19763 27863
rect 19794 27860 19800 27872
rect 19751 27832 19800 27860
rect 19751 27829 19763 27832
rect 19705 27823 19763 27829
rect 19794 27820 19800 27832
rect 19852 27820 19858 27872
rect 20625 27863 20683 27869
rect 20625 27829 20637 27863
rect 20671 27860 20683 27863
rect 20898 27860 20904 27872
rect 20671 27832 20904 27860
rect 20671 27829 20683 27832
rect 20625 27823 20683 27829
rect 20898 27820 20904 27832
rect 20956 27820 20962 27872
rect 21082 27820 21088 27872
rect 21140 27820 21146 27872
rect 21450 27820 21456 27872
rect 21508 27820 21514 27872
rect 1104 27770 21896 27792
rect 750 27684 756 27736
rect 808 27684 814 27736
rect 1104 27718 3549 27770
rect 3601 27718 3613 27770
rect 3665 27718 3677 27770
rect 3729 27718 3741 27770
rect 3793 27718 3805 27770
rect 3857 27718 8747 27770
rect 8799 27718 8811 27770
rect 8863 27718 8875 27770
rect 8927 27718 8939 27770
rect 8991 27718 9003 27770
rect 9055 27718 13945 27770
rect 13997 27718 14009 27770
rect 14061 27718 14073 27770
rect 14125 27718 14137 27770
rect 14189 27718 14201 27770
rect 14253 27718 19143 27770
rect 19195 27718 19207 27770
rect 19259 27718 19271 27770
rect 19323 27718 19335 27770
rect 19387 27718 19399 27770
rect 19451 27718 21896 27770
rect 1104 27696 21896 27718
rect 1670 27616 1676 27668
rect 1728 27656 1734 27668
rect 1728 27628 2820 27656
rect 1728 27616 1734 27628
rect 2792 27588 2820 27628
rect 2866 27616 2872 27668
rect 2924 27656 2930 27668
rect 2924 27628 5028 27656
rect 2924 27616 2930 27628
rect 3142 27588 3148 27600
rect 2792 27560 3148 27588
rect 3142 27548 3148 27560
rect 3200 27548 3206 27600
rect 3973 27591 4031 27597
rect 3973 27557 3985 27591
rect 4019 27588 4031 27591
rect 4246 27588 4252 27600
rect 4019 27560 4252 27588
rect 4019 27557 4031 27560
rect 3973 27551 4031 27557
rect 4246 27548 4252 27560
rect 4304 27548 4310 27600
rect 5000 27588 5028 27628
rect 9122 27616 9128 27668
rect 9180 27656 9186 27668
rect 9490 27656 9496 27668
rect 9180 27628 9496 27656
rect 9180 27616 9186 27628
rect 9490 27616 9496 27628
rect 9548 27616 9554 27668
rect 14366 27656 14372 27668
rect 14108 27628 14372 27656
rect 5166 27588 5172 27600
rect 5000 27560 5172 27588
rect 5166 27548 5172 27560
rect 5224 27548 5230 27600
rect 8665 27591 8723 27597
rect 8665 27588 8677 27591
rect 8496 27560 8677 27588
rect 2240 27492 3832 27520
rect 1578 27412 1584 27464
rect 1636 27412 1642 27464
rect 1854 27452 1860 27464
rect 1815 27424 1860 27452
rect 1854 27412 1860 27424
rect 1912 27412 1918 27464
rect 1302 27344 1308 27396
rect 1360 27384 1366 27396
rect 2240 27384 2268 27492
rect 2406 27412 2412 27464
rect 2464 27452 2470 27464
rect 3804 27461 3832 27492
rect 8110 27480 8116 27532
rect 8168 27480 8174 27532
rect 2961 27455 3019 27461
rect 2961 27452 2973 27455
rect 2464 27424 2973 27452
rect 2464 27412 2470 27424
rect 2961 27421 2973 27424
rect 3007 27421 3019 27455
rect 2961 27415 3019 27421
rect 3237 27455 3295 27461
rect 3237 27421 3249 27455
rect 3283 27421 3295 27455
rect 3237 27415 3295 27421
rect 3789 27455 3847 27461
rect 3789 27421 3801 27455
rect 3835 27421 3847 27455
rect 3789 27415 3847 27421
rect 1360 27356 2268 27384
rect 1360 27344 1366 27356
rect 2498 27344 2504 27396
rect 2556 27384 2562 27396
rect 3252 27384 3280 27415
rect 4154 27412 4160 27464
rect 4212 27452 4218 27464
rect 4249 27455 4307 27461
rect 4249 27452 4261 27455
rect 4212 27424 4261 27452
rect 4212 27412 4218 27424
rect 4249 27421 4261 27424
rect 4295 27421 4307 27455
rect 4491 27455 4549 27461
rect 4491 27452 4503 27455
rect 4249 27415 4307 27421
rect 4344 27424 4503 27452
rect 2556 27356 3280 27384
rect 2556 27344 2562 27356
rect 3694 27344 3700 27396
rect 3752 27384 3758 27396
rect 4062 27384 4068 27396
rect 3752 27356 4068 27384
rect 3752 27344 3758 27356
rect 4062 27344 4068 27356
rect 4120 27384 4126 27396
rect 4344 27384 4372 27424
rect 4491 27421 4503 27424
rect 4537 27421 4549 27455
rect 4491 27415 4549 27421
rect 5534 27412 5540 27464
rect 5592 27452 5598 27464
rect 5629 27455 5687 27461
rect 5629 27452 5641 27455
rect 5592 27424 5641 27452
rect 5592 27412 5598 27424
rect 5629 27421 5641 27424
rect 5675 27421 5687 27455
rect 5629 27415 5687 27421
rect 5871 27455 5929 27461
rect 5871 27421 5883 27455
rect 5917 27452 5929 27455
rect 5994 27452 6000 27464
rect 5917 27424 6000 27452
rect 5917 27421 5929 27424
rect 5871 27415 5929 27421
rect 5994 27412 6000 27424
rect 6052 27412 6058 27464
rect 7282 27452 7288 27464
rect 6564 27424 7288 27452
rect 4120 27356 4372 27384
rect 4120 27344 4126 27356
rect 4890 27344 4896 27396
rect 4948 27384 4954 27396
rect 6564 27384 6592 27424
rect 7282 27412 7288 27424
rect 7340 27412 7346 27464
rect 7466 27412 7472 27464
rect 7524 27452 7530 27464
rect 7524 27424 7880 27452
rect 7524 27412 7530 27424
rect 7558 27384 7564 27396
rect 4948 27356 6592 27384
rect 6656 27356 7564 27384
rect 4948 27344 4954 27356
rect 2590 27276 2596 27328
rect 2648 27276 2654 27328
rect 3142 27276 3148 27328
rect 3200 27276 3206 27328
rect 3326 27276 3332 27328
rect 3384 27316 3390 27328
rect 3421 27319 3479 27325
rect 3421 27316 3433 27319
rect 3384 27288 3433 27316
rect 3384 27276 3390 27288
rect 3421 27285 3433 27288
rect 3467 27316 3479 27319
rect 4798 27316 4804 27328
rect 3467 27288 4804 27316
rect 3467 27285 3479 27288
rect 3421 27279 3479 27285
rect 4798 27276 4804 27288
rect 4856 27276 4862 27328
rect 5261 27319 5319 27325
rect 5261 27285 5273 27319
rect 5307 27316 5319 27319
rect 5994 27316 6000 27328
rect 5307 27288 6000 27316
rect 5307 27285 5319 27288
rect 5261 27279 5319 27285
rect 5994 27276 6000 27288
rect 6052 27276 6058 27328
rect 6656 27325 6684 27356
rect 7558 27344 7564 27356
rect 7616 27344 7622 27396
rect 7650 27344 7656 27396
rect 7708 27344 7714 27396
rect 7742 27344 7748 27396
rect 7800 27344 7806 27396
rect 7852 27384 7880 27424
rect 8018 27412 8024 27464
rect 8076 27452 8082 27464
rect 8496 27452 8524 27560
rect 8665 27557 8677 27560
rect 8711 27557 8723 27591
rect 8665 27551 8723 27557
rect 10965 27591 11023 27597
rect 10965 27557 10977 27591
rect 11011 27588 11023 27591
rect 11011 27560 11376 27588
rect 11011 27557 11023 27560
rect 10965 27551 11023 27557
rect 9766 27480 9772 27532
rect 9824 27520 9830 27532
rect 9953 27523 10011 27529
rect 9953 27520 9965 27523
rect 9824 27492 9965 27520
rect 9824 27480 9830 27492
rect 9953 27489 9965 27492
rect 9999 27489 10011 27523
rect 11348 27506 11376 27560
rect 14108 27529 14136 27628
rect 14366 27616 14372 27628
rect 14424 27656 14430 27668
rect 14550 27656 14556 27668
rect 14424 27628 14556 27656
rect 14424 27616 14430 27628
rect 14550 27616 14556 27628
rect 14608 27656 14614 27668
rect 16206 27656 16212 27668
rect 14608 27628 16212 27656
rect 14608 27616 14614 27628
rect 16206 27616 16212 27628
rect 16264 27616 16270 27668
rect 17034 27616 17040 27668
rect 17092 27656 17098 27668
rect 17494 27656 17500 27668
rect 17092 27628 17500 27656
rect 17092 27616 17098 27628
rect 17494 27616 17500 27628
rect 17552 27616 17558 27668
rect 17681 27659 17739 27665
rect 17681 27625 17693 27659
rect 17727 27656 17739 27659
rect 18046 27656 18052 27668
rect 17727 27628 18052 27656
rect 17727 27625 17739 27628
rect 17681 27619 17739 27625
rect 18046 27616 18052 27628
rect 18104 27616 18110 27668
rect 18138 27616 18144 27668
rect 18196 27616 18202 27668
rect 19518 27616 19524 27668
rect 19576 27656 19582 27668
rect 20714 27656 20720 27668
rect 19576 27628 20720 27656
rect 19576 27616 19582 27628
rect 20714 27616 20720 27628
rect 20772 27616 20778 27668
rect 20806 27616 20812 27668
rect 20864 27616 20870 27668
rect 17770 27588 17776 27600
rect 17512 27560 17776 27588
rect 14093 27523 14151 27529
rect 9953 27483 10011 27489
rect 14093 27489 14105 27523
rect 14139 27489 14151 27523
rect 17512 27520 17540 27560
rect 17770 27548 17776 27560
rect 17828 27588 17834 27600
rect 18156 27588 18184 27616
rect 20625 27591 20683 27597
rect 17828 27560 19288 27588
rect 17828 27548 17834 27560
rect 14093 27483 14151 27489
rect 17236 27492 17540 27520
rect 17589 27523 17647 27529
rect 8076 27424 8524 27452
rect 10227 27455 10285 27461
rect 8076 27412 8082 27424
rect 10227 27421 10239 27455
rect 10273 27452 10285 27455
rect 11606 27452 11612 27464
rect 10273 27424 11612 27452
rect 10273 27421 10285 27424
rect 10227 27415 10285 27421
rect 11606 27412 11612 27424
rect 11664 27412 11670 27464
rect 12645 27455 12703 27461
rect 11714 27424 12388 27452
rect 8113 27387 8171 27393
rect 8113 27384 8125 27387
rect 7852 27356 8125 27384
rect 8113 27353 8125 27356
rect 8159 27384 8171 27387
rect 9214 27384 9220 27396
rect 8159 27356 9220 27384
rect 8159 27353 8171 27356
rect 8113 27347 8171 27353
rect 9214 27344 9220 27356
rect 9272 27344 9278 27396
rect 9582 27344 9588 27396
rect 9640 27384 9646 27396
rect 9950 27384 9956 27396
rect 9640 27356 9956 27384
rect 9640 27344 9646 27356
rect 9950 27344 9956 27356
rect 10008 27344 10014 27396
rect 10594 27344 10600 27396
rect 10652 27384 10658 27396
rect 11714 27384 11742 27424
rect 10652 27356 11742 27384
rect 11793 27387 11851 27393
rect 10652 27344 10658 27356
rect 11793 27353 11805 27387
rect 11839 27353 11851 27387
rect 11793 27347 11851 27353
rect 6641 27319 6699 27325
rect 6641 27285 6653 27319
rect 6687 27285 6699 27319
rect 6641 27279 6699 27285
rect 7098 27276 7104 27328
rect 7156 27316 7162 27328
rect 7377 27319 7435 27325
rect 7377 27316 7389 27319
rect 7156 27288 7389 27316
rect 7156 27276 7162 27288
rect 7377 27285 7389 27288
rect 7423 27316 7435 27319
rect 8386 27316 8392 27328
rect 7423 27288 8392 27316
rect 7423 27285 7435 27288
rect 7377 27279 7435 27285
rect 8386 27276 8392 27288
rect 8444 27276 8450 27328
rect 8478 27276 8484 27328
rect 8536 27276 8542 27328
rect 9398 27276 9404 27328
rect 9456 27316 9462 27328
rect 10778 27316 10784 27328
rect 9456 27288 10784 27316
rect 9456 27276 9462 27288
rect 10778 27276 10784 27288
rect 10836 27276 10842 27328
rect 11146 27276 11152 27328
rect 11204 27316 11210 27328
rect 11517 27319 11575 27325
rect 11517 27316 11529 27319
rect 11204 27288 11529 27316
rect 11204 27276 11210 27288
rect 11517 27285 11529 27288
rect 11563 27285 11575 27319
rect 11808 27316 11836 27347
rect 11882 27344 11888 27396
rect 11940 27344 11946 27396
rect 11974 27344 11980 27396
rect 12032 27344 12038 27396
rect 12250 27344 12256 27396
rect 12308 27344 12314 27396
rect 12360 27384 12388 27424
rect 12645 27421 12657 27455
rect 12691 27452 12703 27455
rect 12986 27452 12992 27464
rect 12691 27424 12992 27452
rect 12691 27421 12703 27424
rect 12645 27415 12703 27421
rect 12986 27412 12992 27424
rect 13044 27412 13050 27464
rect 13078 27412 13084 27464
rect 13136 27452 13142 27464
rect 13262 27452 13268 27464
rect 13136 27424 13268 27452
rect 13136 27412 13142 27424
rect 13262 27412 13268 27424
rect 13320 27412 13326 27464
rect 14367 27455 14425 27461
rect 14367 27452 14379 27455
rect 13372 27424 14379 27452
rect 13372 27384 13400 27424
rect 14367 27421 14379 27424
rect 14413 27452 14425 27455
rect 15841 27455 15899 27461
rect 14413 27424 15516 27452
rect 14413 27421 14425 27424
rect 14367 27415 14425 27421
rect 12360 27356 13400 27384
rect 11992 27316 12020 27344
rect 15488 27328 15516 27424
rect 15841 27421 15853 27455
rect 15887 27452 15899 27455
rect 17236 27452 17264 27492
rect 17589 27489 17601 27523
rect 17635 27520 17647 27523
rect 18138 27520 18144 27532
rect 17635 27492 18144 27520
rect 17635 27489 17647 27492
rect 17589 27483 17647 27489
rect 18138 27480 18144 27492
rect 18196 27480 18202 27532
rect 19058 27480 19064 27532
rect 19116 27480 19122 27532
rect 19260 27529 19288 27560
rect 20625 27557 20637 27591
rect 20671 27588 20683 27591
rect 20824 27588 20852 27616
rect 20671 27560 20852 27588
rect 20671 27557 20683 27560
rect 20625 27551 20683 27557
rect 19245 27523 19303 27529
rect 19245 27489 19257 27523
rect 19291 27489 19303 27523
rect 19245 27483 19303 27489
rect 20254 27480 20260 27532
rect 20312 27520 20318 27532
rect 21634 27520 21640 27532
rect 20312 27492 21640 27520
rect 20312 27480 20318 27492
rect 21634 27480 21640 27492
rect 21692 27480 21698 27532
rect 15887 27424 17264 27452
rect 15887 27421 15899 27424
rect 15841 27415 15899 27421
rect 17310 27412 17316 27464
rect 17368 27412 17374 27464
rect 17402 27412 17408 27464
rect 17460 27412 17466 27464
rect 17865 27455 17923 27461
rect 17865 27421 17877 27455
rect 17911 27421 17923 27455
rect 19076 27452 19104 27480
rect 19501 27455 19559 27461
rect 19501 27452 19513 27455
rect 19076 27424 19513 27452
rect 17865 27415 17923 27421
rect 19501 27421 19513 27424
rect 19547 27421 19559 27455
rect 19501 27415 19559 27421
rect 15930 27344 15936 27396
rect 15988 27384 15994 27396
rect 16086 27387 16144 27393
rect 16086 27384 16098 27387
rect 15988 27356 16098 27384
rect 15988 27344 15994 27356
rect 16086 27353 16098 27356
rect 16132 27353 16144 27387
rect 17880 27384 17908 27415
rect 20990 27412 20996 27464
rect 21048 27412 21054 27464
rect 16086 27347 16144 27353
rect 17236 27356 17908 27384
rect 11808 27288 12020 27316
rect 11517 27279 11575 27285
rect 12710 27276 12716 27328
rect 12768 27316 12774 27328
rect 12805 27319 12863 27325
rect 12805 27316 12817 27319
rect 12768 27288 12817 27316
rect 12768 27276 12774 27288
rect 12805 27285 12817 27288
rect 12851 27285 12863 27319
rect 12805 27279 12863 27285
rect 14458 27276 14464 27328
rect 14516 27316 14522 27328
rect 15105 27319 15163 27325
rect 15105 27316 15117 27319
rect 14516 27288 15117 27316
rect 14516 27276 14522 27288
rect 15105 27285 15117 27288
rect 15151 27285 15163 27319
rect 15105 27279 15163 27285
rect 15470 27276 15476 27328
rect 15528 27276 15534 27328
rect 17236 27325 17264 27356
rect 19610 27344 19616 27396
rect 19668 27384 19674 27396
rect 21361 27387 21419 27393
rect 19668 27356 20944 27384
rect 19668 27344 19674 27356
rect 17221 27319 17279 27325
rect 17221 27285 17233 27319
rect 17267 27285 17279 27319
rect 17221 27279 17279 27285
rect 17589 27319 17647 27325
rect 17589 27285 17601 27319
rect 17635 27316 17647 27319
rect 20714 27316 20720 27328
rect 17635 27288 20720 27316
rect 17635 27285 17647 27288
rect 17589 27279 17647 27285
rect 20714 27276 20720 27288
rect 20772 27276 20778 27328
rect 20916 27316 20944 27356
rect 21361 27353 21373 27387
rect 21407 27384 21419 27387
rect 22186 27384 22192 27396
rect 21407 27356 22192 27384
rect 21407 27353 21419 27356
rect 21361 27347 21419 27353
rect 22186 27344 22192 27356
rect 22244 27344 22250 27396
rect 20990 27316 20996 27328
rect 20916 27288 20996 27316
rect 20990 27276 20996 27288
rect 21048 27276 21054 27328
rect 1104 27226 22056 27248
rect 1104 27174 6148 27226
rect 6200 27174 6212 27226
rect 6264 27174 6276 27226
rect 6328 27174 6340 27226
rect 6392 27174 6404 27226
rect 6456 27174 11346 27226
rect 11398 27174 11410 27226
rect 11462 27174 11474 27226
rect 11526 27174 11538 27226
rect 11590 27174 11602 27226
rect 11654 27174 16544 27226
rect 16596 27174 16608 27226
rect 16660 27174 16672 27226
rect 16724 27174 16736 27226
rect 16788 27174 16800 27226
rect 16852 27174 21742 27226
rect 21794 27174 21806 27226
rect 21858 27174 21870 27226
rect 21922 27174 21934 27226
rect 21986 27174 21998 27226
rect 22050 27174 22056 27226
rect 1104 27152 22056 27174
rect 1210 27072 1216 27124
rect 1268 27112 1274 27124
rect 2406 27112 2412 27124
rect 1268 27084 2412 27112
rect 1268 27072 1274 27084
rect 2406 27072 2412 27084
rect 2464 27072 2470 27124
rect 2498 27072 2504 27124
rect 2556 27072 2562 27124
rect 2590 27072 2596 27124
rect 2648 27072 2654 27124
rect 2682 27072 2688 27124
rect 2740 27112 2746 27124
rect 2777 27115 2835 27121
rect 2777 27112 2789 27115
rect 2740 27084 2789 27112
rect 2740 27072 2746 27084
rect 2777 27081 2789 27084
rect 2823 27081 2835 27115
rect 2777 27075 2835 27081
rect 3326 27072 3332 27124
rect 3384 27112 3390 27124
rect 3694 27112 3700 27124
rect 3384 27084 3700 27112
rect 3384 27072 3390 27084
rect 3694 27072 3700 27084
rect 3752 27072 3758 27124
rect 3970 27072 3976 27124
rect 4028 27112 4034 27124
rect 4246 27112 4252 27124
rect 4028 27084 4252 27112
rect 4028 27072 4034 27084
rect 4246 27072 4252 27084
rect 4304 27072 4310 27124
rect 5534 27112 5540 27124
rect 4344 27084 5540 27112
rect 1302 27004 1308 27056
rect 1360 27044 1366 27056
rect 2516 27044 2544 27072
rect 1360 27016 2544 27044
rect 1360 27004 1366 27016
rect 1394 26936 1400 26988
rect 1452 26936 1458 26988
rect 1486 26936 1492 26988
rect 1544 26976 1550 26988
rect 2317 26979 2375 26985
rect 2317 26976 2329 26979
rect 1544 26948 2329 26976
rect 1544 26936 1550 26948
rect 2317 26945 2329 26948
rect 2363 26945 2375 26979
rect 2317 26939 2375 26945
rect 474 26868 480 26920
rect 532 26908 538 26920
rect 1026 26908 1032 26920
rect 532 26880 1032 26908
rect 532 26868 538 26880
rect 1026 26868 1032 26880
rect 1084 26868 1090 26920
rect 1673 26911 1731 26917
rect 1673 26877 1685 26911
rect 1719 26877 1731 26911
rect 1673 26871 1731 26877
rect 1688 26840 1716 26871
rect 2038 26868 2044 26920
rect 2096 26908 2102 26920
rect 2096 26880 2452 26908
rect 2608 26894 2636 27072
rect 2746 27016 3556 27044
rect 2746 26988 2774 27016
rect 2682 26936 2688 26988
rect 2740 26948 2774 26988
rect 2740 26936 2746 26948
rect 2958 26936 2964 26988
rect 3016 26976 3022 26988
rect 3053 26979 3111 26985
rect 3053 26976 3065 26979
rect 3016 26948 3065 26976
rect 3016 26936 3022 26948
rect 3053 26945 3065 26948
rect 3099 26945 3111 26979
rect 3053 26939 3111 26945
rect 3142 26936 3148 26988
rect 3200 26936 3206 26988
rect 3528 26985 3556 27016
rect 3786 27004 3792 27056
rect 3844 27044 3850 27056
rect 3881 27047 3939 27053
rect 3881 27044 3893 27047
rect 3844 27016 3893 27044
rect 3844 27004 3850 27016
rect 3881 27013 3893 27016
rect 3927 27013 3939 27047
rect 3881 27007 3939 27013
rect 4154 27004 4160 27056
rect 4212 27044 4218 27056
rect 4344 27044 4372 27084
rect 5534 27072 5540 27084
rect 5592 27112 5598 27124
rect 10686 27112 10692 27124
rect 5592 27084 10692 27112
rect 5592 27072 5598 27084
rect 10686 27072 10692 27084
rect 10744 27072 10750 27124
rect 11146 27072 11152 27124
rect 11204 27112 11210 27124
rect 11701 27115 11759 27121
rect 11701 27112 11713 27115
rect 11204 27084 11713 27112
rect 11204 27072 11210 27084
rect 11701 27081 11713 27084
rect 11747 27081 11759 27115
rect 14826 27112 14832 27124
rect 11701 27075 11759 27081
rect 13924 27084 14832 27112
rect 5258 27044 5264 27056
rect 4212 27016 4372 27044
rect 4908 27016 5264 27044
rect 4212 27004 4218 27016
rect 3513 26979 3571 26985
rect 3513 26945 3525 26979
rect 3559 26976 3571 26979
rect 3970 26976 3976 26988
rect 3559 26948 3976 26976
rect 3559 26945 3571 26948
rect 3513 26939 3571 26945
rect 3970 26936 3976 26948
rect 4028 26936 4034 26988
rect 4908 26985 4936 27016
rect 5258 27004 5264 27016
rect 5316 27004 5322 27056
rect 5350 27004 5356 27056
rect 5408 27004 5414 27056
rect 5994 27004 6000 27056
rect 6052 27004 6058 27056
rect 8110 27004 8116 27056
rect 8168 27044 8174 27056
rect 9306 27044 9312 27056
rect 8168 27016 9312 27044
rect 8168 27004 8174 27016
rect 9306 27004 9312 27016
rect 9364 27004 9370 27056
rect 9784 27016 10088 27044
rect 4249 26979 4307 26985
rect 4249 26945 4261 26979
rect 4295 26976 4307 26979
rect 4893 26979 4951 26985
rect 4295 26948 4844 26976
rect 4295 26945 4307 26948
rect 4249 26939 4307 26945
rect 2096 26868 2102 26880
rect 1688 26812 2360 26840
rect 2332 26784 2360 26812
rect 2314 26732 2320 26784
rect 2372 26732 2378 26784
rect 2424 26772 2452 26880
rect 4062 26868 4068 26920
rect 4120 26908 4126 26920
rect 4614 26908 4620 26920
rect 4120 26880 4620 26908
rect 4120 26868 4126 26880
rect 4614 26868 4620 26880
rect 4672 26868 4678 26920
rect 2498 26800 2504 26852
rect 2556 26800 2562 26852
rect 2590 26772 2596 26784
rect 2424 26744 2596 26772
rect 2590 26732 2596 26744
rect 2648 26732 2654 26784
rect 4062 26732 4068 26784
rect 4120 26732 4126 26784
rect 4430 26732 4436 26784
rect 4488 26732 4494 26784
rect 4816 26772 4844 26948
rect 4893 26945 4905 26979
rect 4939 26945 4951 26979
rect 4893 26939 4951 26945
rect 5167 26979 5225 26985
rect 5167 26945 5179 26979
rect 5213 26976 5225 26979
rect 5368 26976 5396 27004
rect 5213 26948 5396 26976
rect 6012 26976 6040 27004
rect 9784 26988 9812 27016
rect 6012 26948 6684 26976
rect 5213 26945 5225 26948
rect 5167 26939 5225 26945
rect 5626 26868 5632 26920
rect 5684 26908 5690 26920
rect 6365 26911 6423 26917
rect 6365 26908 6377 26911
rect 5684 26880 6377 26908
rect 5684 26868 5690 26880
rect 6365 26877 6377 26880
rect 6411 26877 6423 26911
rect 6365 26871 6423 26877
rect 6546 26868 6552 26920
rect 6604 26868 6610 26920
rect 6656 26908 6684 26948
rect 7374 26936 7380 26988
rect 7432 26985 7438 26988
rect 7432 26979 7460 26985
rect 7448 26945 7460 26979
rect 7432 26939 7460 26945
rect 7432 26936 7438 26939
rect 7558 26936 7564 26988
rect 7616 26936 7622 26988
rect 8571 26979 8629 26985
rect 8571 26945 8583 26979
rect 8617 26976 8629 26979
rect 8662 26976 8668 26988
rect 8617 26948 8668 26976
rect 8617 26945 8629 26948
rect 8571 26939 8629 26945
rect 8662 26936 8668 26948
rect 8720 26936 8726 26988
rect 9677 26979 9735 26985
rect 9677 26976 9689 26979
rect 9324 26948 9689 26976
rect 7009 26911 7067 26917
rect 7009 26908 7021 26911
rect 6656 26880 7021 26908
rect 7009 26877 7021 26880
rect 7055 26877 7067 26911
rect 7009 26871 7067 26877
rect 7098 26868 7104 26920
rect 7156 26908 7162 26920
rect 7285 26911 7343 26917
rect 7285 26908 7297 26911
rect 7156 26880 7297 26908
rect 7156 26868 7162 26880
rect 7285 26877 7297 26880
rect 7331 26877 7343 26911
rect 7285 26871 7343 26877
rect 8110 26868 8116 26920
rect 8168 26908 8174 26920
rect 8285 26911 8343 26917
rect 8285 26908 8297 26911
rect 8168 26880 8297 26908
rect 8168 26868 8174 26880
rect 8266 26877 8297 26880
rect 8331 26877 8343 26911
rect 8266 26871 8343 26877
rect 8266 26840 8294 26871
rect 5552 26812 6132 26840
rect 8266 26812 8340 26840
rect 5552 26772 5580 26812
rect 4816 26744 5580 26772
rect 5905 26775 5963 26781
rect 5905 26741 5917 26775
rect 5951 26772 5963 26775
rect 5994 26772 6000 26784
rect 5951 26744 6000 26772
rect 5951 26741 5963 26744
rect 5905 26735 5963 26741
rect 5994 26732 6000 26744
rect 6052 26732 6058 26784
rect 6104 26772 6132 26812
rect 8205 26775 8263 26781
rect 8205 26772 8217 26775
rect 6104 26744 8217 26772
rect 8205 26741 8217 26744
rect 8251 26741 8263 26775
rect 8312 26772 8340 26812
rect 9324 26784 9352 26948
rect 9677 26945 9689 26948
rect 9723 26945 9735 26979
rect 9677 26939 9735 26945
rect 9766 26936 9772 26988
rect 9824 26936 9830 26988
rect 10060 26985 10088 27016
rect 10134 27004 10140 27056
rect 10192 27004 10198 27056
rect 10778 27004 10784 27056
rect 10836 27044 10842 27056
rect 11790 27044 11796 27056
rect 10836 27016 11796 27044
rect 10836 27004 10842 27016
rect 11790 27004 11796 27016
rect 11848 27004 11854 27056
rect 11974 27004 11980 27056
rect 12032 27004 12038 27056
rect 12069 27047 12127 27053
rect 12069 27013 12081 27047
rect 12115 27044 12127 27047
rect 12158 27044 12164 27056
rect 12115 27016 12164 27044
rect 12115 27013 12127 27016
rect 12069 27007 12127 27013
rect 12158 27004 12164 27016
rect 12216 27004 12222 27056
rect 12250 27004 12256 27056
rect 12308 27044 12314 27056
rect 12437 27047 12495 27053
rect 12437 27044 12449 27047
rect 12308 27016 12449 27044
rect 12308 27004 12314 27016
rect 12437 27013 12449 27016
rect 12483 27013 12495 27047
rect 12437 27007 12495 27013
rect 12618 27004 12624 27056
rect 12676 27044 12682 27056
rect 12805 27047 12863 27053
rect 12805 27044 12817 27047
rect 12676 27016 12817 27044
rect 12676 27004 12682 27016
rect 12805 27013 12817 27016
rect 12851 27044 12863 27047
rect 12986 27044 12992 27056
rect 12851 27016 12992 27044
rect 12851 27013 12863 27016
rect 12805 27007 12863 27013
rect 12986 27004 12992 27016
rect 13044 27004 13050 27056
rect 9861 26979 9919 26985
rect 9861 26945 9873 26979
rect 9907 26945 9919 26979
rect 9861 26939 9919 26945
rect 10045 26979 10103 26985
rect 10045 26945 10057 26979
rect 10091 26945 10103 26979
rect 10152 26976 10180 27004
rect 10287 26979 10345 26985
rect 10287 26976 10299 26979
rect 10152 26948 10299 26976
rect 10045 26939 10103 26945
rect 10287 26945 10299 26948
rect 10333 26945 10345 26979
rect 10287 26939 10345 26945
rect 9398 26868 9404 26920
rect 9456 26908 9462 26920
rect 9876 26908 9904 26939
rect 10686 26936 10692 26988
rect 10744 26976 10750 26988
rect 13924 26976 13952 27084
rect 14826 27072 14832 27084
rect 14884 27072 14890 27124
rect 16114 27072 16120 27124
rect 16172 27112 16178 27124
rect 16850 27112 16856 27124
rect 16172 27084 16856 27112
rect 16172 27072 16178 27084
rect 16850 27072 16856 27084
rect 16908 27072 16914 27124
rect 17310 27072 17316 27124
rect 17368 27072 17374 27124
rect 18046 27072 18052 27124
rect 18104 27072 18110 27124
rect 18138 27072 18144 27124
rect 18196 27072 18202 27124
rect 19337 27115 19395 27121
rect 19337 27081 19349 27115
rect 19383 27112 19395 27115
rect 20254 27112 20260 27124
rect 19383 27084 20260 27112
rect 19383 27081 19395 27084
rect 19337 27075 19395 27081
rect 20254 27072 20260 27084
rect 20312 27072 20318 27124
rect 21266 27072 21272 27124
rect 21324 27112 21330 27124
rect 21361 27115 21419 27121
rect 21361 27112 21373 27115
rect 21324 27084 21373 27112
rect 21324 27072 21330 27084
rect 21361 27081 21373 27084
rect 21407 27081 21419 27115
rect 21361 27075 21419 27081
rect 15654 27004 15660 27056
rect 15712 27044 15718 27056
rect 16298 27044 16304 27056
rect 15712 27016 16304 27044
rect 15712 27004 15718 27016
rect 16298 27004 16304 27016
rect 16356 27004 16362 27056
rect 10744 26948 13952 26976
rect 10744 26936 10750 26948
rect 14642 26936 14648 26988
rect 14700 26936 14706 26988
rect 15565 26979 15623 26985
rect 15565 26945 15577 26979
rect 15611 26976 15623 26979
rect 15841 26979 15899 26985
rect 15841 26976 15853 26979
rect 15611 26948 15853 26976
rect 15611 26945 15623 26948
rect 15565 26939 15623 26945
rect 15841 26945 15853 26948
rect 15887 26945 15899 26979
rect 15841 26939 15899 26945
rect 16114 26936 16120 26988
rect 16172 26936 16178 26988
rect 16209 26979 16267 26985
rect 16209 26945 16221 26979
rect 16255 26945 16267 26979
rect 16209 26939 16267 26945
rect 9456 26880 9904 26908
rect 9456 26868 9462 26880
rect 11057 26843 11115 26849
rect 11057 26809 11069 26843
rect 11103 26840 11115 26843
rect 11532 26840 11560 26894
rect 13354 26868 13360 26920
rect 13412 26908 13418 26920
rect 13630 26908 13636 26920
rect 13412 26880 13636 26908
rect 13412 26868 13418 26880
rect 13630 26868 13636 26880
rect 13688 26908 13694 26920
rect 13725 26911 13783 26917
rect 13725 26908 13737 26911
rect 13688 26880 13737 26908
rect 13688 26868 13694 26880
rect 13725 26877 13737 26880
rect 13771 26877 13783 26911
rect 13725 26871 13783 26877
rect 13909 26911 13967 26917
rect 13909 26877 13921 26911
rect 13955 26877 13967 26911
rect 13909 26871 13967 26877
rect 14369 26911 14427 26917
rect 14369 26877 14381 26911
rect 14415 26908 14427 26911
rect 14458 26908 14464 26920
rect 14415 26880 14464 26908
rect 14415 26877 14427 26880
rect 14369 26871 14427 26877
rect 13924 26840 13952 26871
rect 14458 26868 14464 26880
rect 14516 26868 14522 26920
rect 14734 26868 14740 26920
rect 14792 26917 14798 26920
rect 14792 26911 14820 26917
rect 14808 26877 14820 26911
rect 14792 26871 14820 26877
rect 14921 26911 14979 26917
rect 14921 26877 14933 26911
rect 14967 26908 14979 26911
rect 15286 26908 15292 26920
rect 14967 26880 15292 26908
rect 14967 26877 14979 26880
rect 14921 26871 14979 26877
rect 14792 26868 14798 26871
rect 15286 26868 15292 26880
rect 15344 26868 15350 26920
rect 16224 26908 16252 26939
rect 16850 26936 16856 26988
rect 16908 26976 16914 26988
rect 16943 26979 17001 26985
rect 16943 26976 16955 26979
rect 16908 26948 16955 26976
rect 16908 26936 16914 26948
rect 16943 26945 16955 26948
rect 16989 26945 17001 26979
rect 16943 26939 17001 26945
rect 17328 26976 17356 27072
rect 18064 27044 18092 27072
rect 18064 27016 18276 27044
rect 18248 26985 18276 27016
rect 19886 27015 19892 27056
rect 19871 27009 19892 27015
rect 18049 26979 18107 26985
rect 18049 26976 18061 26979
rect 17328 26948 18061 26976
rect 15948 26880 16252 26908
rect 16669 26911 16727 26917
rect 15948 26849 15976 26880
rect 16669 26877 16681 26911
rect 16715 26877 16727 26911
rect 16669 26871 16727 26877
rect 11103 26812 11560 26840
rect 13004 26812 13952 26840
rect 15933 26843 15991 26849
rect 11103 26809 11115 26812
rect 11057 26803 11115 26809
rect 13004 26784 13032 26812
rect 15933 26809 15945 26843
rect 15979 26809 15991 26843
rect 15933 26803 15991 26809
rect 8754 26772 8760 26784
rect 8312 26744 8760 26772
rect 8205 26735 8263 26741
rect 8754 26732 8760 26744
rect 8812 26732 8818 26784
rect 9306 26732 9312 26784
rect 9364 26732 9370 26784
rect 9766 26732 9772 26784
rect 9824 26732 9830 26784
rect 12986 26732 12992 26784
rect 13044 26732 13050 26784
rect 13630 26732 13636 26784
rect 13688 26772 13694 26784
rect 14734 26772 14740 26784
rect 13688 26744 14740 26772
rect 13688 26732 13694 26744
rect 14734 26732 14740 26744
rect 14792 26732 14798 26784
rect 15654 26732 15660 26784
rect 15712 26732 15718 26784
rect 15746 26732 15752 26784
rect 15804 26772 15810 26784
rect 16301 26775 16359 26781
rect 16301 26772 16313 26775
rect 15804 26744 16313 26772
rect 15804 26732 15810 26744
rect 16301 26741 16313 26744
rect 16347 26741 16359 26775
rect 16684 26772 16712 26871
rect 17328 26840 17356 26948
rect 18049 26945 18061 26948
rect 18095 26945 18107 26979
rect 18049 26939 18107 26945
rect 18233 26979 18291 26985
rect 18233 26945 18245 26979
rect 18279 26945 18291 26979
rect 18233 26939 18291 26945
rect 19521 26979 19579 26985
rect 19521 26945 19533 26979
rect 19567 26945 19579 26979
rect 19871 26975 19883 27009
rect 19944 27004 19950 27056
rect 20070 27004 20076 27056
rect 20128 27044 20134 27056
rect 20128 27016 21588 27044
rect 20128 27004 20134 27016
rect 19917 26978 19932 27004
rect 21560 26985 21588 27016
rect 20993 26979 21051 26985
rect 19917 26975 19929 26978
rect 20993 26976 21005 26979
rect 19871 26969 19929 26975
rect 19521 26939 19579 26945
rect 20640 26948 21005 26976
rect 18138 26868 18144 26920
rect 18196 26908 18202 26920
rect 19536 26908 19564 26939
rect 18196 26880 19564 26908
rect 19613 26911 19671 26917
rect 18196 26868 18202 26880
rect 19613 26877 19625 26911
rect 19659 26877 19671 26911
rect 19613 26871 19671 26877
rect 17681 26843 17739 26849
rect 17681 26840 17693 26843
rect 17328 26812 17693 26840
rect 17681 26809 17693 26812
rect 17727 26809 17739 26843
rect 17681 26803 17739 26809
rect 17034 26772 17040 26784
rect 16684 26744 17040 26772
rect 16301 26735 16359 26741
rect 17034 26732 17040 26744
rect 17092 26772 17098 26784
rect 18874 26772 18880 26784
rect 17092 26744 18880 26772
rect 17092 26732 17098 26744
rect 18874 26732 18880 26744
rect 18932 26772 18938 26784
rect 19628 26772 19656 26871
rect 20640 26852 20668 26948
rect 20993 26945 21005 26948
rect 21039 26945 21051 26979
rect 20993 26939 21051 26945
rect 21545 26979 21603 26985
rect 21545 26945 21557 26979
rect 21591 26945 21603 26979
rect 21545 26939 21603 26945
rect 21266 26868 21272 26920
rect 21324 26868 21330 26920
rect 20622 26800 20628 26852
rect 20680 26800 20686 26852
rect 18932 26744 19656 26772
rect 18932 26732 18938 26744
rect 20438 26732 20444 26784
rect 20496 26772 20502 26784
rect 21085 26775 21143 26781
rect 21085 26772 21097 26775
rect 20496 26744 21097 26772
rect 20496 26732 20502 26744
rect 21085 26741 21097 26744
rect 21131 26741 21143 26775
rect 21085 26735 21143 26741
rect 21177 26775 21235 26781
rect 21177 26741 21189 26775
rect 21223 26772 21235 26775
rect 22646 26772 22652 26784
rect 21223 26744 22652 26772
rect 21223 26741 21235 26744
rect 21177 26735 21235 26741
rect 22646 26732 22652 26744
rect 22704 26732 22710 26784
rect 1104 26682 21896 26704
rect 1104 26630 3549 26682
rect 3601 26630 3613 26682
rect 3665 26630 3677 26682
rect 3729 26630 3741 26682
rect 3793 26630 3805 26682
rect 3857 26630 8747 26682
rect 8799 26630 8811 26682
rect 8863 26630 8875 26682
rect 8927 26630 8939 26682
rect 8991 26630 9003 26682
rect 9055 26630 13945 26682
rect 13997 26630 14009 26682
rect 14061 26630 14073 26682
rect 14125 26630 14137 26682
rect 14189 26630 14201 26682
rect 14253 26630 19143 26682
rect 19195 26630 19207 26682
rect 19259 26630 19271 26682
rect 19323 26630 19335 26682
rect 19387 26630 19399 26682
rect 19451 26630 21896 26682
rect 1104 26608 21896 26630
rect 2958 26528 2964 26580
rect 3016 26528 3022 26580
rect 3142 26528 3148 26580
rect 3200 26568 3206 26580
rect 4801 26571 4859 26577
rect 4801 26568 4813 26571
rect 3200 26540 4813 26568
rect 3200 26528 3206 26540
rect 4801 26537 4813 26540
rect 4847 26537 4859 26571
rect 8478 26568 8484 26580
rect 4801 26531 4859 26537
rect 5552 26540 8484 26568
rect 2498 26500 2504 26512
rect 2148 26472 2504 26500
rect 1394 26392 1400 26444
rect 1452 26392 1458 26444
rect 1671 26367 1729 26373
rect 1671 26333 1683 26367
rect 1717 26364 1729 26367
rect 2038 26364 2044 26376
rect 1717 26336 2044 26364
rect 1717 26333 1729 26336
rect 1671 26327 1729 26333
rect 2038 26324 2044 26336
rect 2096 26364 2102 26376
rect 2148 26364 2176 26472
rect 2498 26460 2504 26472
rect 2556 26460 2562 26512
rect 3237 26503 3295 26509
rect 3237 26469 3249 26503
rect 3283 26500 3295 26503
rect 3326 26500 3332 26512
rect 3283 26472 3332 26500
rect 3283 26469 3295 26472
rect 3237 26463 3295 26469
rect 3326 26460 3332 26472
rect 3384 26460 3390 26512
rect 3418 26460 3424 26512
rect 3476 26500 3482 26512
rect 3513 26503 3571 26509
rect 3513 26500 3525 26503
rect 3476 26472 3525 26500
rect 3476 26460 3482 26472
rect 3513 26469 3525 26472
rect 3559 26469 3571 26503
rect 3513 26463 3571 26469
rect 4614 26460 4620 26512
rect 4672 26500 4678 26512
rect 4672 26472 5488 26500
rect 4672 26460 4678 26472
rect 2096 26336 2176 26364
rect 2240 26404 3832 26432
rect 2096 26324 2102 26336
rect 1578 26256 1584 26308
rect 1636 26296 1642 26308
rect 2240 26296 2268 26404
rect 2777 26367 2835 26373
rect 2777 26333 2789 26367
rect 2823 26333 2835 26367
rect 2777 26327 2835 26333
rect 1636 26268 2268 26296
rect 1636 26256 1642 26268
rect 2792 26240 2820 26327
rect 3050 26324 3056 26376
rect 3108 26324 3114 26376
rect 3326 26324 3332 26376
rect 3384 26324 3390 26376
rect 3804 26373 3832 26404
rect 3789 26367 3847 26373
rect 3789 26333 3801 26367
rect 3835 26333 3847 26367
rect 3789 26327 3847 26333
rect 4063 26367 4121 26373
rect 4063 26333 4075 26367
rect 4109 26364 4121 26367
rect 5166 26364 5172 26376
rect 4109 26336 5172 26364
rect 4109 26333 4121 26336
rect 4063 26327 4121 26333
rect 2406 26188 2412 26240
rect 2464 26188 2470 26240
rect 2774 26188 2780 26240
rect 2832 26188 2838 26240
rect 3804 26228 3832 26327
rect 5166 26324 5172 26336
rect 5224 26324 5230 26376
rect 5350 26324 5356 26376
rect 5408 26324 5414 26376
rect 5460 26364 5488 26472
rect 5552 26441 5580 26540
rect 5644 26472 6132 26500
rect 5537 26435 5595 26441
rect 5537 26401 5549 26435
rect 5583 26401 5595 26435
rect 5537 26395 5595 26401
rect 5644 26364 5672 26472
rect 5994 26392 6000 26444
rect 6052 26392 6058 26444
rect 6104 26432 6132 26472
rect 6390 26435 6448 26441
rect 6390 26432 6402 26435
rect 6104 26404 6402 26432
rect 6390 26401 6402 26404
rect 6436 26401 6448 26435
rect 6390 26395 6448 26401
rect 6549 26435 6607 26441
rect 6549 26401 6561 26435
rect 6595 26432 6607 26435
rect 6914 26432 6920 26444
rect 6595 26404 6920 26432
rect 6595 26401 6607 26404
rect 6549 26395 6607 26401
rect 6914 26392 6920 26404
rect 6972 26392 6978 26444
rect 5460 26336 5672 26364
rect 6270 26324 6276 26376
rect 6328 26324 6334 26376
rect 6638 26228 6644 26240
rect 3804 26200 6644 26228
rect 6638 26188 6644 26200
rect 6696 26188 6702 26240
rect 7190 26188 7196 26240
rect 7248 26188 7254 26240
rect 7300 26228 7328 26540
rect 8478 26528 8484 26540
rect 8536 26528 8542 26580
rect 9122 26528 9128 26580
rect 9180 26568 9186 26580
rect 9401 26571 9459 26577
rect 9401 26568 9413 26571
rect 9180 26540 9413 26568
rect 9180 26528 9186 26540
rect 9401 26537 9413 26540
rect 9447 26537 9459 26571
rect 9401 26531 9459 26537
rect 9766 26528 9772 26580
rect 9824 26528 9830 26580
rect 12526 26528 12532 26580
rect 12584 26568 12590 26580
rect 12621 26571 12679 26577
rect 12621 26568 12633 26571
rect 12584 26540 12633 26568
rect 12584 26528 12590 26540
rect 12621 26537 12633 26540
rect 12667 26568 12679 26571
rect 13630 26568 13636 26580
rect 12667 26540 13636 26568
rect 12667 26537 12679 26540
rect 12621 26531 12679 26537
rect 13630 26528 13636 26540
rect 13688 26528 13694 26580
rect 14458 26528 14464 26580
rect 14516 26528 14522 26580
rect 15010 26568 15016 26580
rect 14844 26540 15016 26568
rect 9306 26392 9312 26444
rect 9364 26392 9370 26444
rect 9784 26432 9812 26528
rect 10781 26503 10839 26509
rect 10781 26469 10793 26503
rect 10827 26500 10839 26503
rect 14476 26500 14504 26528
rect 14737 26503 14795 26509
rect 14737 26500 14749 26503
rect 10827 26472 11192 26500
rect 14476 26472 14749 26500
rect 10827 26469 10839 26472
rect 10781 26463 10839 26469
rect 9508 26404 9812 26432
rect 10704 26404 10916 26432
rect 11164 26418 11192 26472
rect 14737 26469 14749 26472
rect 14783 26469 14795 26503
rect 14737 26463 14795 26469
rect 7469 26367 7527 26373
rect 7469 26333 7481 26367
rect 7515 26333 7527 26367
rect 7469 26327 7527 26333
rect 7743 26367 7801 26373
rect 7743 26333 7755 26367
rect 7789 26364 7801 26367
rect 7834 26364 7840 26376
rect 7789 26336 7840 26364
rect 7789 26333 7801 26336
rect 7743 26327 7801 26333
rect 7484 26296 7512 26327
rect 7834 26324 7840 26336
rect 7892 26324 7898 26376
rect 8110 26324 8116 26376
rect 8168 26364 8174 26376
rect 9508 26373 9536 26404
rect 9125 26367 9183 26373
rect 9125 26364 9137 26367
rect 8168 26336 9137 26364
rect 8168 26324 8174 26336
rect 9125 26333 9137 26336
rect 9171 26333 9183 26367
rect 9125 26327 9183 26333
rect 9493 26367 9551 26373
rect 9493 26333 9505 26367
rect 9539 26333 9551 26367
rect 9493 26327 9551 26333
rect 9766 26324 9772 26376
rect 9824 26324 9830 26376
rect 9950 26324 9956 26376
rect 10008 26364 10014 26376
rect 10043 26367 10101 26373
rect 10043 26364 10055 26367
rect 10008 26336 10055 26364
rect 10008 26324 10014 26336
rect 10043 26333 10055 26336
rect 10089 26364 10101 26367
rect 10704 26364 10732 26404
rect 10888 26376 10916 26404
rect 12710 26392 12716 26444
rect 12768 26432 12774 26444
rect 14844 26432 14872 26540
rect 15010 26528 15016 26540
rect 15068 26528 15074 26580
rect 15933 26571 15991 26577
rect 15933 26537 15945 26571
rect 15979 26568 15991 26571
rect 16114 26568 16120 26580
rect 15979 26540 16120 26568
rect 15979 26537 15991 26540
rect 15933 26531 15991 26537
rect 16114 26528 16120 26540
rect 16172 26528 16178 26580
rect 17402 26528 17408 26580
rect 17460 26568 17466 26580
rect 17497 26571 17555 26577
rect 17497 26568 17509 26571
rect 17460 26540 17509 26568
rect 17460 26528 17466 26540
rect 17497 26537 17509 26540
rect 17543 26537 17555 26571
rect 17497 26531 17555 26537
rect 18230 26528 18236 26580
rect 18288 26568 18294 26580
rect 18288 26540 20024 26568
rect 18288 26528 18294 26540
rect 18325 26503 18383 26509
rect 18325 26469 18337 26503
rect 18371 26469 18383 26503
rect 18325 26463 18383 26469
rect 15194 26441 15200 26444
rect 15013 26435 15071 26441
rect 15013 26432 15025 26435
rect 12768 26404 15025 26432
rect 12768 26392 12774 26404
rect 15013 26401 15025 26404
rect 15059 26401 15071 26435
rect 15013 26395 15071 26401
rect 15151 26435 15200 26441
rect 15151 26401 15163 26435
rect 15197 26401 15200 26435
rect 15151 26395 15200 26401
rect 15194 26392 15200 26395
rect 15252 26392 15258 26444
rect 15286 26392 15292 26444
rect 15344 26392 15350 26444
rect 16025 26435 16083 26441
rect 16025 26401 16037 26435
rect 16071 26401 16083 26435
rect 18340 26432 18368 26463
rect 19996 26432 20024 26540
rect 20070 26528 20076 26580
rect 20128 26528 20134 26580
rect 20438 26528 20444 26580
rect 20496 26528 20502 26580
rect 20622 26528 20628 26580
rect 20680 26528 20686 26580
rect 20714 26528 20720 26580
rect 20772 26528 20778 26580
rect 20901 26571 20959 26577
rect 20901 26537 20913 26571
rect 20947 26568 20959 26571
rect 21266 26568 21272 26580
rect 20947 26540 21272 26568
rect 20947 26537 20959 26540
rect 20901 26531 20959 26537
rect 21266 26528 21272 26540
rect 21324 26528 21330 26580
rect 18340 26404 19288 26432
rect 19996 26404 20576 26432
rect 16025 26395 16083 26401
rect 10089 26336 10732 26364
rect 10089 26333 10101 26336
rect 10043 26327 10101 26333
rect 10778 26324 10784 26376
rect 10836 26324 10842 26376
rect 10870 26324 10876 26376
rect 10928 26324 10934 26376
rect 11701 26367 11759 26373
rect 11701 26333 11713 26367
rect 11747 26364 11759 26367
rect 13906 26364 13912 26376
rect 11747 26336 13912 26364
rect 11747 26333 11759 26336
rect 11701 26327 11759 26333
rect 13906 26324 13912 26336
rect 13964 26324 13970 26376
rect 14093 26367 14151 26373
rect 14093 26333 14105 26367
rect 14139 26364 14151 26367
rect 14182 26364 14188 26376
rect 14139 26336 14188 26364
rect 14139 26333 14151 26336
rect 14093 26327 14151 26333
rect 14182 26324 14188 26336
rect 14240 26324 14246 26376
rect 14277 26367 14335 26373
rect 14277 26333 14289 26367
rect 14323 26333 14335 26367
rect 14277 26327 14335 26333
rect 9214 26296 9220 26308
rect 7484 26268 9220 26296
rect 9214 26256 9220 26268
rect 9272 26256 9278 26308
rect 9784 26296 9812 26324
rect 10796 26296 10824 26324
rect 9784 26268 10824 26296
rect 11609 26299 11667 26305
rect 11609 26265 11621 26299
rect 11655 26296 11667 26299
rect 11974 26296 11980 26308
rect 11655 26268 11980 26296
rect 11655 26265 11667 26268
rect 11609 26259 11667 26265
rect 11974 26256 11980 26268
rect 12032 26256 12038 26308
rect 12069 26299 12127 26305
rect 12069 26265 12081 26299
rect 12115 26296 12127 26299
rect 12250 26296 12256 26308
rect 12115 26268 12256 26296
rect 12115 26265 12127 26268
rect 12069 26259 12127 26265
rect 12250 26256 12256 26268
rect 12308 26256 12314 26308
rect 12437 26299 12495 26305
rect 12437 26265 12449 26299
rect 12483 26296 12495 26299
rect 12618 26296 12624 26308
rect 12483 26268 12624 26296
rect 12483 26265 12495 26268
rect 12437 26259 12495 26265
rect 12618 26256 12624 26268
rect 12676 26256 12682 26308
rect 12986 26256 12992 26308
rect 13044 26296 13050 26308
rect 14292 26296 14320 26327
rect 13044 26268 14320 26296
rect 16040 26296 16068 26395
rect 16283 26337 16341 26343
rect 16114 26296 16120 26308
rect 16040 26268 16120 26296
rect 13044 26256 13050 26268
rect 16114 26256 16120 26268
rect 16172 26256 16178 26308
rect 16283 26303 16295 26337
rect 16329 26334 16341 26337
rect 16329 26308 16342 26334
rect 16390 26324 16396 26376
rect 16448 26364 16454 26376
rect 19260 26373 19288 26404
rect 17405 26367 17463 26373
rect 17405 26364 17417 26367
rect 16448 26336 17417 26364
rect 16448 26324 16454 26336
rect 17405 26333 17417 26336
rect 17451 26333 17463 26367
rect 17405 26327 17463 26333
rect 18509 26367 18567 26373
rect 18509 26333 18521 26367
rect 18555 26333 18567 26367
rect 18509 26327 18567 26333
rect 19245 26367 19303 26373
rect 19245 26333 19257 26367
rect 19291 26333 19303 26367
rect 19245 26327 19303 26333
rect 19337 26367 19395 26373
rect 19337 26333 19349 26367
rect 19383 26364 19395 26367
rect 19518 26364 19524 26376
rect 19383 26336 19524 26364
rect 19383 26333 19395 26336
rect 19337 26327 19395 26333
rect 16283 26297 16304 26303
rect 16298 26256 16304 26297
rect 16356 26256 16362 26308
rect 18524 26240 18552 26327
rect 19518 26324 19524 26336
rect 19576 26324 19582 26376
rect 19705 26367 19763 26373
rect 19705 26333 19717 26367
rect 19751 26333 19763 26367
rect 19705 26327 19763 26333
rect 19150 26256 19156 26308
rect 19208 26296 19214 26308
rect 19720 26296 19748 26327
rect 19794 26324 19800 26376
rect 19852 26324 19858 26376
rect 20254 26324 20260 26376
rect 20312 26324 20318 26376
rect 20349 26367 20407 26373
rect 20349 26333 20361 26367
rect 20395 26333 20407 26367
rect 20349 26327 20407 26333
rect 19208 26268 19748 26296
rect 19812 26296 19840 26324
rect 20364 26296 20392 26327
rect 19812 26268 20392 26296
rect 20548 26296 20576 26404
rect 20640 26364 20668 26528
rect 20732 26432 20760 26528
rect 20732 26404 21220 26432
rect 20809 26367 20867 26373
rect 20809 26364 20821 26367
rect 20640 26336 20821 26364
rect 20809 26333 20821 26336
rect 20855 26333 20867 26367
rect 20809 26327 20867 26333
rect 20898 26324 20904 26376
rect 20956 26364 20962 26376
rect 21192 26373 21220 26404
rect 20993 26367 21051 26373
rect 20993 26364 21005 26367
rect 20956 26336 21005 26364
rect 20956 26324 20962 26336
rect 20993 26333 21005 26336
rect 21039 26333 21051 26367
rect 20993 26327 21051 26333
rect 21177 26367 21235 26373
rect 21177 26333 21189 26367
rect 21223 26333 21235 26367
rect 21177 26327 21235 26333
rect 21266 26296 21272 26308
rect 20548 26268 21272 26296
rect 19208 26256 19214 26268
rect 21266 26256 21272 26268
rect 21324 26256 21330 26308
rect 21545 26299 21603 26305
rect 21545 26265 21557 26299
rect 21591 26296 21603 26299
rect 22278 26296 22284 26308
rect 21591 26268 22284 26296
rect 21591 26265 21603 26268
rect 21545 26259 21603 26265
rect 22278 26256 22284 26268
rect 22336 26256 22342 26308
rect 7834 26228 7840 26240
rect 7300 26200 7840 26228
rect 7834 26188 7840 26200
rect 7892 26188 7898 26240
rect 8478 26188 8484 26240
rect 8536 26188 8542 26240
rect 9306 26188 9312 26240
rect 9364 26228 9370 26240
rect 10502 26228 10508 26240
rect 9364 26200 10508 26228
rect 9364 26188 9370 26200
rect 10502 26188 10508 26200
rect 10560 26188 10566 26240
rect 11146 26188 11152 26240
rect 11204 26228 11210 26240
rect 11333 26231 11391 26237
rect 11333 26228 11345 26231
rect 11204 26200 11345 26228
rect 11204 26188 11210 26200
rect 11333 26197 11345 26200
rect 11379 26197 11391 26231
rect 11333 26191 11391 26197
rect 12158 26188 12164 26240
rect 12216 26228 12222 26240
rect 13538 26228 13544 26240
rect 12216 26200 13544 26228
rect 12216 26188 12222 26200
rect 13538 26188 13544 26200
rect 13596 26188 13602 26240
rect 16206 26188 16212 26240
rect 16264 26228 16270 26240
rect 17037 26231 17095 26237
rect 17037 26228 17049 26231
rect 16264 26200 17049 26228
rect 16264 26188 16270 26200
rect 17037 26197 17049 26200
rect 17083 26197 17095 26231
rect 17037 26191 17095 26197
rect 18506 26188 18512 26240
rect 18564 26188 18570 26240
rect 19521 26231 19579 26237
rect 19521 26197 19533 26231
rect 19567 26228 19579 26231
rect 19794 26228 19800 26240
rect 19567 26200 19800 26228
rect 19567 26197 19579 26200
rect 19521 26191 19579 26197
rect 19794 26188 19800 26200
rect 19852 26188 19858 26240
rect 1104 26138 22056 26160
rect 1104 26086 6148 26138
rect 6200 26086 6212 26138
rect 6264 26086 6276 26138
rect 6328 26086 6340 26138
rect 6392 26086 6404 26138
rect 6456 26086 11346 26138
rect 11398 26086 11410 26138
rect 11462 26086 11474 26138
rect 11526 26086 11538 26138
rect 11590 26086 11602 26138
rect 11654 26086 16544 26138
rect 16596 26086 16608 26138
rect 16660 26086 16672 26138
rect 16724 26086 16736 26138
rect 16788 26086 16800 26138
rect 16852 26086 21742 26138
rect 21794 26086 21806 26138
rect 21858 26086 21870 26138
rect 21922 26086 21934 26138
rect 21986 26086 21998 26138
rect 22050 26086 22056 26138
rect 1104 26064 22056 26086
rect 1397 26027 1455 26033
rect 1397 25993 1409 26027
rect 1443 26024 1455 26027
rect 3878 26024 3884 26036
rect 1443 25996 3884 26024
rect 1443 25993 1455 25996
rect 1397 25987 1455 25993
rect 3878 25984 3884 25996
rect 3936 26024 3942 26036
rect 4341 26027 4399 26033
rect 4341 26024 4353 26027
rect 3936 25996 4353 26024
rect 3936 25984 3942 25996
rect 4341 25993 4353 25996
rect 4387 26024 4399 26027
rect 5350 26024 5356 26036
rect 4387 25996 5356 26024
rect 4387 25993 4399 25996
rect 4341 25987 4399 25993
rect 5350 25984 5356 25996
rect 5408 25984 5414 26036
rect 7190 25984 7196 26036
rect 7248 25984 7254 26036
rect 7282 25984 7288 26036
rect 7340 26024 7346 26036
rect 8202 26024 8208 26036
rect 7340 25996 8208 26024
rect 7340 25984 7346 25996
rect 8202 25984 8208 25996
rect 8260 25984 8266 26036
rect 10689 26027 10747 26033
rect 10689 26024 10701 26027
rect 8588 25996 10701 26024
rect 2222 25956 2228 25968
rect 1688 25928 2228 25956
rect 1578 25848 1584 25900
rect 1636 25848 1642 25900
rect 1688 25897 1716 25928
rect 2222 25916 2228 25928
rect 2280 25916 2286 25968
rect 2314 25916 2320 25968
rect 2372 25956 2378 25968
rect 3237 25959 3295 25965
rect 3237 25956 3249 25959
rect 2372 25928 3249 25956
rect 2372 25916 2378 25928
rect 3237 25925 3249 25928
rect 3283 25925 3295 25959
rect 3237 25919 3295 25925
rect 3326 25916 3332 25968
rect 3384 25956 3390 25968
rect 3605 25959 3663 25965
rect 3605 25956 3617 25959
rect 3384 25928 3617 25956
rect 3384 25916 3390 25928
rect 3605 25925 3617 25928
rect 3651 25925 3663 25959
rect 3605 25919 3663 25925
rect 3970 25916 3976 25968
rect 4028 25916 4034 25968
rect 7208 25956 7236 25984
rect 6564 25928 7236 25956
rect 1673 25891 1731 25897
rect 1673 25857 1685 25891
rect 1719 25857 1731 25891
rect 1673 25851 1731 25857
rect 1947 25891 2005 25897
rect 1947 25857 1959 25891
rect 1993 25888 2005 25891
rect 2038 25888 2044 25900
rect 1993 25860 2044 25888
rect 1993 25857 2005 25860
rect 1947 25851 2005 25857
rect 2038 25848 2044 25860
rect 2096 25848 2102 25900
rect 3510 25848 3516 25900
rect 3568 25848 3574 25900
rect 6564 25897 6592 25928
rect 8386 25916 8392 25968
rect 8444 25956 8450 25968
rect 8588 25965 8616 25996
rect 10689 25993 10701 25996
rect 10735 25993 10747 26027
rect 10689 25987 10747 25993
rect 10870 25984 10876 26036
rect 10928 26024 10934 26036
rect 10928 25996 13860 26024
rect 10928 25984 10934 25996
rect 8481 25959 8539 25965
rect 8481 25956 8493 25959
rect 8444 25928 8493 25956
rect 8444 25916 8450 25928
rect 8481 25925 8493 25928
rect 8527 25925 8539 25959
rect 8481 25919 8539 25925
rect 8573 25959 8631 25965
rect 8573 25925 8585 25959
rect 8619 25925 8631 25959
rect 8573 25919 8631 25925
rect 8662 25916 8668 25968
rect 8720 25956 8726 25968
rect 8941 25959 8999 25965
rect 8941 25956 8953 25959
rect 8720 25928 8953 25956
rect 8720 25916 8726 25928
rect 8941 25925 8953 25928
rect 8987 25925 8999 25959
rect 8941 25919 8999 25925
rect 9309 25959 9367 25965
rect 9309 25925 9321 25959
rect 9355 25925 9367 25959
rect 13262 25956 13268 25968
rect 9309 25919 9367 25925
rect 9692 25928 13268 25956
rect 6549 25891 6607 25897
rect 6549 25857 6561 25891
rect 6595 25857 6607 25891
rect 6549 25851 6607 25857
rect 6915 25891 6973 25897
rect 6915 25857 6927 25891
rect 6961 25888 6973 25891
rect 7742 25888 7748 25900
rect 6961 25860 7748 25888
rect 6961 25857 6973 25860
rect 6915 25851 6973 25857
rect 7742 25848 7748 25860
rect 7800 25848 7806 25900
rect 7834 25848 7840 25900
rect 7892 25888 7898 25900
rect 9324 25888 9352 25919
rect 9692 25897 9720 25928
rect 13262 25916 13268 25928
rect 13320 25956 13326 25968
rect 13832 25956 13860 25996
rect 13906 25984 13912 26036
rect 13964 25984 13970 26036
rect 14642 25984 14648 26036
rect 14700 25984 14706 26036
rect 15654 25984 15660 26036
rect 15712 26024 15718 26036
rect 15712 25996 16436 26024
rect 15712 25984 15718 25996
rect 14660 25956 14688 25984
rect 13320 25928 13774 25956
rect 13832 25928 14688 25956
rect 16025 25959 16083 25965
rect 13320 25916 13326 25928
rect 7892 25860 9352 25888
rect 9677 25891 9735 25897
rect 7892 25848 7898 25860
rect 9677 25857 9689 25891
rect 9723 25857 9735 25891
rect 9677 25851 9735 25857
rect 9858 25848 9864 25900
rect 9916 25888 9922 25900
rect 9951 25891 10009 25897
rect 9951 25888 9963 25891
rect 9916 25860 9963 25888
rect 9916 25848 9922 25860
rect 9951 25857 9963 25860
rect 9997 25888 10009 25891
rect 10594 25888 10600 25900
rect 9997 25860 10600 25888
rect 9997 25857 10009 25860
rect 9951 25851 10009 25857
rect 10594 25848 10600 25860
rect 10652 25848 10658 25900
rect 11054 25848 11060 25900
rect 11112 25888 11118 25900
rect 11238 25888 11244 25900
rect 11112 25860 11244 25888
rect 11112 25848 11118 25860
rect 11238 25848 11244 25860
rect 11296 25888 11302 25900
rect 11517 25891 11575 25897
rect 11517 25888 11529 25891
rect 11296 25860 11529 25888
rect 11296 25848 11302 25860
rect 11517 25857 11529 25860
rect 11563 25857 11575 25891
rect 11517 25851 11575 25857
rect 11791 25891 11849 25897
rect 11791 25857 11803 25891
rect 11837 25888 11849 25891
rect 12158 25888 12164 25900
rect 11837 25860 12164 25888
rect 11837 25857 11849 25860
rect 11791 25851 11849 25857
rect 12158 25848 12164 25860
rect 12216 25848 12222 25900
rect 13171 25891 13229 25897
rect 13171 25857 13183 25891
rect 13217 25888 13229 25891
rect 13630 25888 13636 25900
rect 13217 25860 13636 25888
rect 13217 25857 13229 25860
rect 13171 25851 13229 25857
rect 13630 25848 13636 25860
rect 13688 25848 13694 25900
rect 13746 25888 13774 25928
rect 16025 25925 16037 25959
rect 16071 25956 16083 25959
rect 16301 25959 16359 25965
rect 16301 25956 16313 25959
rect 16071 25928 16313 25956
rect 16071 25925 16083 25928
rect 16025 25919 16083 25925
rect 16301 25925 16313 25928
rect 16347 25925 16359 25959
rect 16301 25919 16359 25925
rect 14918 25888 14924 25900
rect 13746 25860 14924 25888
rect 14918 25848 14924 25860
rect 14976 25848 14982 25900
rect 15286 25848 15292 25900
rect 15344 25848 15350 25900
rect 15657 25891 15715 25897
rect 15657 25857 15669 25891
rect 15703 25888 15715 25891
rect 15746 25888 15752 25900
rect 15703 25860 15752 25888
rect 15703 25857 15715 25860
rect 15657 25851 15715 25857
rect 15746 25848 15752 25860
rect 15804 25848 15810 25900
rect 15841 25891 15899 25897
rect 15841 25857 15853 25891
rect 15887 25888 15899 25891
rect 16206 25888 16212 25900
rect 15887 25860 16212 25888
rect 15887 25857 15899 25860
rect 15841 25851 15899 25857
rect 16206 25848 16212 25860
rect 16264 25848 16270 25900
rect 16408 25897 16436 25996
rect 17034 25984 17040 26036
rect 17092 26024 17098 26036
rect 18598 26024 18604 26036
rect 17092 25996 18604 26024
rect 17092 25984 17098 25996
rect 18598 25984 18604 25996
rect 18656 25984 18662 26036
rect 19150 25984 19156 26036
rect 19208 25984 19214 26036
rect 19702 26024 19708 26036
rect 19536 25996 19708 26024
rect 19536 25927 19564 25996
rect 19702 25984 19708 25996
rect 19760 25984 19766 26036
rect 19503 25921 19564 25927
rect 16393 25891 16451 25897
rect 16393 25857 16405 25891
rect 16439 25857 16451 25891
rect 16393 25851 16451 25857
rect 17770 25848 17776 25900
rect 17828 25848 17834 25900
rect 18029 25891 18087 25897
rect 18029 25888 18041 25891
rect 17878 25860 18041 25888
rect 2685 25687 2743 25693
rect 2685 25653 2697 25687
rect 2731 25684 2743 25687
rect 3068 25684 3096 25806
rect 6638 25780 6644 25832
rect 6696 25780 6702 25832
rect 4522 25712 4528 25764
rect 4580 25712 4586 25764
rect 7653 25755 7711 25761
rect 7653 25721 7665 25755
rect 7699 25752 7711 25755
rect 8036 25752 8064 25806
rect 12894 25780 12900 25832
rect 12952 25780 12958 25832
rect 15304 25820 15332 25848
rect 17878 25820 17906 25860
rect 18029 25857 18041 25860
rect 18075 25888 18087 25891
rect 18506 25888 18512 25900
rect 18075 25860 18512 25888
rect 18075 25857 18087 25860
rect 18029 25851 18087 25857
rect 18506 25848 18512 25860
rect 18564 25848 18570 25900
rect 19503 25887 19515 25921
rect 19549 25890 19564 25921
rect 19610 25916 19616 25968
rect 19668 25956 19674 25968
rect 19668 25928 21312 25956
rect 19668 25916 19674 25928
rect 19549 25887 19561 25890
rect 19503 25881 19561 25887
rect 20898 25848 20904 25900
rect 20956 25848 20962 25900
rect 21284 25897 21312 25928
rect 20993 25891 21051 25897
rect 20993 25857 21005 25891
rect 21039 25857 21051 25891
rect 20993 25851 21051 25857
rect 21269 25891 21327 25897
rect 21269 25857 21281 25891
rect 21315 25857 21327 25891
rect 21269 25851 21327 25857
rect 15304 25792 17906 25820
rect 18874 25780 18880 25832
rect 18932 25820 18938 25832
rect 19245 25823 19303 25829
rect 19245 25820 19257 25823
rect 18932 25792 19257 25820
rect 18932 25780 18938 25792
rect 19245 25789 19257 25792
rect 19291 25789 19303 25823
rect 19245 25783 19303 25789
rect 20070 25780 20076 25832
rect 20128 25820 20134 25832
rect 21008 25820 21036 25851
rect 20128 25792 21036 25820
rect 20128 25780 20134 25792
rect 12802 25752 12808 25764
rect 7699 25724 8064 25752
rect 12406 25724 12808 25752
rect 7699 25721 7711 25724
rect 7653 25715 7711 25721
rect 2731 25656 3096 25684
rect 6365 25687 6423 25693
rect 2731 25653 2743 25656
rect 2685 25647 2743 25653
rect 6365 25653 6377 25687
rect 6411 25684 6423 25687
rect 7098 25684 7104 25696
rect 6411 25656 7104 25684
rect 6411 25653 6423 25656
rect 6365 25647 6423 25653
rect 7098 25644 7104 25656
rect 7156 25644 7162 25696
rect 9493 25687 9551 25693
rect 9493 25653 9505 25687
rect 9539 25684 9551 25687
rect 9582 25684 9588 25696
rect 9539 25656 9588 25684
rect 9539 25653 9551 25656
rect 9493 25647 9551 25653
rect 9582 25644 9588 25656
rect 9640 25644 9646 25696
rect 10778 25644 10784 25696
rect 10836 25684 10842 25696
rect 12406 25684 12434 25724
rect 12802 25712 12808 25724
rect 12860 25712 12866 25764
rect 10836 25656 12434 25684
rect 10836 25644 10842 25656
rect 12526 25644 12532 25696
rect 12584 25644 12590 25696
rect 12912 25684 12940 25780
rect 13262 25684 13268 25696
rect 12912 25656 13268 25684
rect 13262 25644 13268 25656
rect 13320 25644 13326 25696
rect 15930 25644 15936 25696
rect 15988 25644 15994 25696
rect 17678 25644 17684 25696
rect 17736 25684 17742 25696
rect 18690 25684 18696 25696
rect 17736 25656 18696 25684
rect 17736 25644 17742 25656
rect 18690 25644 18696 25656
rect 18748 25644 18754 25696
rect 19702 25644 19708 25696
rect 19760 25684 19766 25696
rect 20257 25687 20315 25693
rect 20257 25684 20269 25687
rect 19760 25656 20269 25684
rect 19760 25644 19766 25656
rect 20257 25653 20269 25656
rect 20303 25653 20315 25687
rect 20257 25647 20315 25653
rect 20714 25644 20720 25696
rect 20772 25644 20778 25696
rect 21082 25644 21088 25696
rect 21140 25644 21146 25696
rect 21450 25644 21456 25696
rect 21508 25644 21514 25696
rect 1104 25594 21896 25616
rect 1104 25542 3549 25594
rect 3601 25542 3613 25594
rect 3665 25542 3677 25594
rect 3729 25542 3741 25594
rect 3793 25542 3805 25594
rect 3857 25542 8747 25594
rect 8799 25542 8811 25594
rect 8863 25542 8875 25594
rect 8927 25542 8939 25594
rect 8991 25542 9003 25594
rect 9055 25542 13945 25594
rect 13997 25542 14009 25594
rect 14061 25542 14073 25594
rect 14125 25542 14137 25594
rect 14189 25542 14201 25594
rect 14253 25542 19143 25594
rect 19195 25542 19207 25594
rect 19259 25542 19271 25594
rect 19323 25542 19335 25594
rect 19387 25542 19399 25594
rect 19451 25542 21896 25594
rect 1104 25520 21896 25542
rect 2130 25440 2136 25492
rect 2188 25440 2194 25492
rect 3326 25440 3332 25492
rect 3384 25440 3390 25492
rect 6730 25480 6736 25492
rect 3988 25452 6736 25480
rect 1670 25304 1676 25356
rect 1728 25304 1734 25356
rect 1394 25236 1400 25288
rect 1452 25236 1458 25288
rect 2148 25276 2176 25440
rect 3988 25421 4016 25452
rect 6730 25440 6736 25452
rect 6788 25440 6794 25492
rect 7098 25440 7104 25492
rect 7156 25480 7162 25492
rect 7156 25452 8064 25480
rect 7156 25440 7162 25452
rect 3973 25415 4031 25421
rect 3973 25381 3985 25415
rect 4019 25381 4031 25415
rect 3973 25375 4031 25381
rect 5994 25372 6000 25424
rect 6052 25412 6058 25424
rect 6365 25415 6423 25421
rect 6365 25412 6377 25415
rect 6052 25384 6377 25412
rect 6052 25372 6058 25384
rect 6365 25381 6377 25384
rect 6411 25381 6423 25415
rect 6365 25375 6423 25381
rect 2222 25304 2228 25356
rect 2280 25344 2286 25356
rect 2317 25347 2375 25353
rect 2317 25344 2329 25347
rect 2280 25316 2329 25344
rect 2280 25304 2286 25316
rect 2317 25313 2329 25316
rect 2363 25313 2375 25347
rect 2317 25307 2375 25313
rect 5902 25304 5908 25356
rect 5960 25304 5966 25356
rect 6086 25304 6092 25356
rect 6144 25344 6150 25356
rect 6641 25347 6699 25353
rect 6641 25344 6653 25347
rect 6144 25316 6653 25344
rect 6144 25304 6150 25316
rect 6641 25313 6653 25316
rect 6687 25313 6699 25347
rect 6641 25307 6699 25313
rect 6779 25347 6837 25353
rect 6779 25313 6791 25347
rect 6825 25344 6837 25347
rect 6825 25316 7512 25344
rect 6825 25313 6837 25316
rect 6779 25307 6837 25313
rect 2498 25276 2504 25288
rect 2148 25248 2504 25276
rect 2498 25236 2504 25248
rect 2556 25285 2562 25288
rect 2556 25279 2617 25285
rect 2556 25245 2571 25279
rect 2605 25245 2617 25279
rect 2556 25239 2617 25245
rect 2556 25236 2562 25239
rect 3234 25236 3240 25288
rect 3292 25276 3298 25288
rect 3789 25279 3847 25285
rect 3789 25276 3801 25279
rect 3292 25248 3801 25276
rect 3292 25236 3298 25248
rect 3789 25245 3801 25248
rect 3835 25245 3847 25279
rect 3789 25239 3847 25245
rect 4341 25279 4399 25285
rect 4341 25245 4353 25279
rect 4387 25245 4399 25279
rect 4341 25239 4399 25245
rect 4615 25279 4673 25285
rect 4615 25245 4627 25279
rect 4661 25245 4673 25279
rect 4615 25239 4673 25245
rect 4356 25140 4384 25239
rect 4522 25168 4528 25220
rect 4580 25208 4586 25220
rect 4630 25208 4658 25239
rect 5350 25236 5356 25288
rect 5408 25236 5414 25288
rect 5626 25236 5632 25288
rect 5684 25276 5690 25288
rect 5721 25279 5779 25285
rect 5721 25276 5733 25279
rect 5684 25248 5733 25276
rect 5684 25236 5690 25248
rect 5721 25245 5733 25248
rect 5767 25245 5779 25279
rect 5721 25239 5779 25245
rect 6914 25236 6920 25288
rect 6972 25236 6978 25288
rect 5368 25208 5396 25236
rect 4580 25180 4658 25208
rect 4706 25180 5396 25208
rect 7484 25208 7512 25316
rect 8036 25285 8064 25452
rect 8110 25440 8116 25492
rect 8168 25440 8174 25492
rect 8478 25440 8484 25492
rect 8536 25440 8542 25492
rect 9122 25440 9128 25492
rect 9180 25480 9186 25492
rect 9180 25452 9720 25480
rect 9180 25440 9186 25452
rect 8496 25412 8524 25440
rect 9585 25415 9643 25421
rect 9585 25412 9597 25415
rect 8496 25384 9597 25412
rect 9585 25381 9597 25384
rect 9631 25381 9643 25415
rect 9585 25375 9643 25381
rect 8202 25304 8208 25356
rect 8260 25304 8266 25356
rect 8662 25304 8668 25356
rect 8720 25344 8726 25356
rect 9125 25347 9183 25353
rect 9125 25344 9137 25347
rect 8720 25316 9137 25344
rect 8720 25304 8726 25316
rect 9125 25313 9137 25316
rect 9171 25313 9183 25347
rect 9692 25344 9720 25452
rect 10778 25440 10784 25492
rect 10836 25440 10842 25492
rect 12802 25440 12808 25492
rect 12860 25480 12866 25492
rect 12860 25452 19012 25480
rect 12860 25440 12866 25452
rect 18693 25415 18751 25421
rect 18693 25381 18705 25415
rect 18739 25381 18751 25415
rect 18693 25375 18751 25381
rect 12532 25356 12584 25362
rect 9978 25347 10036 25353
rect 9978 25344 9990 25347
rect 9692 25316 9990 25344
rect 9125 25307 9183 25313
rect 9978 25313 9990 25316
rect 10024 25313 10036 25347
rect 9978 25307 10036 25313
rect 7561 25279 7619 25285
rect 7561 25245 7573 25279
rect 7607 25276 7619 25279
rect 7929 25279 7987 25285
rect 7929 25276 7941 25279
rect 7607 25248 7941 25276
rect 7607 25245 7619 25248
rect 7561 25239 7619 25245
rect 7929 25245 7941 25248
rect 7975 25245 7987 25279
rect 7929 25239 7987 25245
rect 8021 25279 8079 25285
rect 8021 25245 8033 25279
rect 8067 25245 8079 25279
rect 8220 25276 8248 25304
rect 12532 25298 12584 25304
rect 8941 25279 8999 25285
rect 8941 25276 8953 25279
rect 8220 25248 8953 25276
rect 8021 25239 8079 25245
rect 8941 25245 8953 25248
rect 8987 25245 8999 25279
rect 8941 25239 8999 25245
rect 9858 25236 9864 25288
rect 9916 25236 9922 25288
rect 10134 25236 10140 25288
rect 10192 25236 10198 25288
rect 11793 25279 11851 25285
rect 11793 25245 11805 25279
rect 11839 25276 11851 25279
rect 11974 25276 11980 25288
rect 11839 25248 11980 25276
rect 11839 25245 11851 25248
rect 11793 25239 11851 25245
rect 11974 25236 11980 25248
rect 12032 25236 12038 25288
rect 12342 25236 12348 25288
rect 12400 25276 12406 25288
rect 12802 25276 12808 25288
rect 12400 25270 12480 25276
rect 12636 25270 12808 25276
rect 12400 25248 12808 25270
rect 12400 25236 12406 25248
rect 12452 25242 12664 25248
rect 12802 25236 12808 25248
rect 12860 25236 12866 25288
rect 14093 25279 14151 25285
rect 14093 25245 14105 25279
rect 14139 25276 14151 25279
rect 14826 25276 14832 25288
rect 14139 25248 14832 25276
rect 14139 25245 14151 25248
rect 14093 25239 14151 25245
rect 14826 25236 14832 25248
rect 14884 25236 14890 25288
rect 15010 25236 15016 25288
rect 15068 25276 15074 25288
rect 15105 25279 15163 25285
rect 15105 25276 15117 25279
rect 15068 25248 15117 25276
rect 15068 25236 15074 25248
rect 15105 25245 15117 25248
rect 15151 25245 15163 25279
rect 15378 25276 15384 25288
rect 15339 25248 15384 25276
rect 15105 25239 15163 25245
rect 8386 25208 8392 25220
rect 7484 25180 8392 25208
rect 4580 25168 4586 25180
rect 4706 25140 4734 25180
rect 8386 25168 8392 25180
rect 8444 25208 8450 25220
rect 8662 25208 8668 25220
rect 8444 25180 8668 25208
rect 8444 25168 8450 25180
rect 8662 25168 8668 25180
rect 8720 25168 8726 25220
rect 11882 25168 11888 25220
rect 11940 25168 11946 25220
rect 12250 25168 12256 25220
rect 12308 25168 12314 25220
rect 15120 25208 15148 25239
rect 15378 25236 15384 25248
rect 15436 25236 15442 25288
rect 16485 25279 16543 25285
rect 16485 25245 16497 25279
rect 16531 25245 16543 25279
rect 18049 25279 18107 25285
rect 18049 25276 18061 25279
rect 16485 25239 16543 25245
rect 16743 25249 16801 25255
rect 16022 25208 16028 25220
rect 15120 25180 16028 25208
rect 16022 25168 16028 25180
rect 16080 25208 16086 25220
rect 16500 25208 16528 25239
rect 16743 25215 16755 25249
rect 16789 25215 16801 25249
rect 16743 25209 16801 25215
rect 17420 25248 18061 25276
rect 16080 25180 16528 25208
rect 16080 25168 16086 25180
rect 4356 25112 4734 25140
rect 5353 25143 5411 25149
rect 5353 25109 5365 25143
rect 5399 25140 5411 25143
rect 6914 25140 6920 25152
rect 5399 25112 6920 25140
rect 5399 25109 5411 25112
rect 5353 25103 5411 25109
rect 6914 25100 6920 25112
rect 6972 25100 6978 25152
rect 7745 25143 7803 25149
rect 7745 25109 7757 25143
rect 7791 25140 7803 25143
rect 9398 25140 9404 25152
rect 7791 25112 9404 25140
rect 7791 25109 7803 25112
rect 7745 25103 7803 25109
rect 9398 25100 9404 25112
rect 9456 25100 9462 25152
rect 11146 25100 11152 25152
rect 11204 25140 11210 25152
rect 11517 25143 11575 25149
rect 11517 25140 11529 25143
rect 11204 25112 11529 25140
rect 11204 25100 11210 25112
rect 11517 25109 11529 25112
rect 11563 25140 11575 25143
rect 12342 25140 12348 25152
rect 11563 25112 12348 25140
rect 11563 25109 11575 25112
rect 11517 25103 11575 25109
rect 12342 25100 12348 25112
rect 12400 25100 12406 25152
rect 12618 25100 12624 25152
rect 12676 25100 12682 25152
rect 12805 25143 12863 25149
rect 12805 25109 12817 25143
rect 12851 25140 12863 25143
rect 13354 25140 13360 25152
rect 12851 25112 13360 25140
rect 12851 25109 12863 25112
rect 12805 25103 12863 25109
rect 13354 25100 13360 25112
rect 13412 25100 13418 25152
rect 14185 25143 14243 25149
rect 14185 25109 14197 25143
rect 14231 25140 14243 25143
rect 14274 25140 14280 25152
rect 14231 25112 14280 25140
rect 14231 25109 14243 25112
rect 14185 25103 14243 25109
rect 14274 25100 14280 25112
rect 14332 25100 14338 25152
rect 14918 25100 14924 25152
rect 14976 25140 14982 25152
rect 15838 25140 15844 25152
rect 14976 25112 15844 25140
rect 14976 25100 14982 25112
rect 15838 25100 15844 25112
rect 15896 25100 15902 25152
rect 16114 25100 16120 25152
rect 16172 25100 16178 25152
rect 16758 25140 16786 25209
rect 17420 25152 17448 25248
rect 18049 25245 18061 25248
rect 18095 25245 18107 25279
rect 18049 25239 18107 25245
rect 18417 25279 18475 25285
rect 18417 25245 18429 25279
rect 18463 25276 18475 25279
rect 18506 25276 18512 25288
rect 18463 25248 18512 25276
rect 18463 25245 18475 25248
rect 18417 25239 18475 25245
rect 18506 25236 18512 25248
rect 18564 25236 18570 25288
rect 18601 25279 18659 25285
rect 18601 25245 18613 25279
rect 18647 25276 18659 25279
rect 18708 25276 18736 25375
rect 18647 25248 18736 25276
rect 18647 25245 18659 25248
rect 18601 25239 18659 25245
rect 18874 25236 18880 25288
rect 18932 25236 18938 25288
rect 18984 25276 19012 25452
rect 19518 25440 19524 25492
rect 19576 25440 19582 25492
rect 19610 25440 19616 25492
rect 19668 25440 19674 25492
rect 19702 25440 19708 25492
rect 19760 25440 19766 25492
rect 19794 25440 19800 25492
rect 19852 25440 19858 25492
rect 20070 25440 20076 25492
rect 20128 25440 20134 25492
rect 20714 25440 20720 25492
rect 20772 25440 20778 25492
rect 19720 25412 19748 25440
rect 19628 25384 19748 25412
rect 19812 25412 19840 25440
rect 19812 25384 20024 25412
rect 19429 25279 19487 25285
rect 18984 25248 19380 25276
rect 18966 25208 18972 25220
rect 17880 25180 18972 25208
rect 17034 25140 17040 25152
rect 16758 25112 17040 25140
rect 17034 25100 17040 25112
rect 17092 25100 17098 25152
rect 17402 25100 17408 25152
rect 17460 25100 17466 25152
rect 17494 25100 17500 25152
rect 17552 25100 17558 25152
rect 17880 25149 17908 25180
rect 18966 25168 18972 25180
rect 19024 25168 19030 25220
rect 19352 25208 19380 25248
rect 19429 25245 19441 25279
rect 19475 25276 19487 25279
rect 19628 25276 19656 25384
rect 19705 25347 19763 25353
rect 19705 25313 19717 25347
rect 19751 25344 19763 25347
rect 19889 25347 19947 25353
rect 19889 25344 19901 25347
rect 19751 25316 19901 25344
rect 19751 25313 19763 25316
rect 19705 25307 19763 25313
rect 19889 25313 19901 25316
rect 19935 25313 19947 25347
rect 19889 25307 19947 25313
rect 19996 25285 20024 25384
rect 20530 25344 20536 25356
rect 20364 25316 20536 25344
rect 19797 25279 19855 25285
rect 19797 25276 19809 25279
rect 19475 25248 19809 25276
rect 19475 25245 19487 25248
rect 19429 25239 19487 25245
rect 19797 25245 19809 25248
rect 19843 25245 19855 25279
rect 19797 25239 19855 25245
rect 19981 25279 20039 25285
rect 19981 25245 19993 25279
rect 20027 25245 20039 25279
rect 19981 25239 20039 25245
rect 20257 25279 20315 25285
rect 20257 25245 20269 25279
rect 20303 25245 20315 25279
rect 20257 25239 20315 25245
rect 19886 25208 19892 25220
rect 19352 25180 19892 25208
rect 19886 25168 19892 25180
rect 19944 25208 19950 25220
rect 20272 25208 20300 25239
rect 19944 25180 20300 25208
rect 19944 25168 19950 25180
rect 17865 25143 17923 25149
rect 17865 25109 17877 25143
rect 17911 25109 17923 25143
rect 17865 25103 17923 25109
rect 18598 25100 18604 25152
rect 18656 25100 18662 25152
rect 19702 25100 19708 25152
rect 19760 25140 19766 25152
rect 20364 25140 20392 25316
rect 20530 25304 20536 25316
rect 20588 25304 20594 25356
rect 20438 25236 20444 25288
rect 20496 25236 20502 25288
rect 20625 25279 20683 25285
rect 20625 25245 20637 25279
rect 20671 25276 20683 25279
rect 20732 25276 20760 25440
rect 20671 25248 20760 25276
rect 20901 25279 20959 25285
rect 20671 25245 20683 25248
rect 20625 25239 20683 25245
rect 20901 25245 20913 25279
rect 20947 25245 20959 25279
rect 20901 25239 20959 25245
rect 21177 25279 21235 25285
rect 21177 25245 21189 25279
rect 21223 25276 21235 25279
rect 21266 25276 21272 25288
rect 21223 25248 21272 25276
rect 21223 25245 21235 25248
rect 21177 25239 21235 25245
rect 20530 25168 20536 25220
rect 20588 25208 20594 25220
rect 20916 25208 20944 25239
rect 21266 25236 21272 25248
rect 21324 25236 21330 25288
rect 20588 25180 20944 25208
rect 21545 25211 21603 25217
rect 20588 25168 20594 25180
rect 21545 25177 21557 25211
rect 21591 25208 21603 25211
rect 22278 25208 22284 25220
rect 21591 25180 22284 25208
rect 21591 25177 21603 25180
rect 21545 25171 21603 25177
rect 22278 25168 22284 25180
rect 22336 25168 22342 25220
rect 19760 25112 20392 25140
rect 19760 25100 19766 25112
rect 20622 25100 20628 25152
rect 20680 25100 20686 25152
rect 20714 25100 20720 25152
rect 20772 25100 20778 25152
rect 14 25032 20 25084
rect 72 25072 78 25084
rect 290 25072 296 25084
rect 72 25044 296 25072
rect 72 25032 78 25044
rect 290 25032 296 25044
rect 348 25032 354 25084
rect 1104 25050 22056 25072
rect 1104 24998 6148 25050
rect 6200 24998 6212 25050
rect 6264 24998 6276 25050
rect 6328 24998 6340 25050
rect 6392 24998 6404 25050
rect 6456 24998 11346 25050
rect 11398 24998 11410 25050
rect 11462 24998 11474 25050
rect 11526 24998 11538 25050
rect 11590 24998 11602 25050
rect 11654 24998 16544 25050
rect 16596 24998 16608 25050
rect 16660 24998 16672 25050
rect 16724 24998 16736 25050
rect 16788 24998 16800 25050
rect 16852 24998 21742 25050
rect 21794 24998 21806 25050
rect 21858 24998 21870 25050
rect 21922 24998 21934 25050
rect 21986 24998 21998 25050
rect 22050 24998 22056 25050
rect 1104 24976 22056 24998
rect 1397 24939 1455 24945
rect 1397 24905 1409 24939
rect 1443 24936 1455 24939
rect 2866 24936 2872 24948
rect 1443 24908 2872 24936
rect 1443 24905 1455 24908
rect 1397 24899 1455 24905
rect 2866 24896 2872 24908
rect 2924 24896 2930 24948
rect 4062 24896 4068 24948
rect 4120 24936 4126 24948
rect 4982 24936 4988 24948
rect 4120 24908 4988 24936
rect 4120 24896 4126 24908
rect 4982 24896 4988 24908
rect 5040 24896 5046 24948
rect 5442 24896 5448 24948
rect 5500 24936 5506 24948
rect 5994 24936 6000 24948
rect 5500 24908 6000 24936
rect 5500 24896 5506 24908
rect 5994 24896 6000 24908
rect 6052 24896 6058 24948
rect 8110 24936 8116 24948
rect 6104 24908 8116 24936
rect 1854 24828 1860 24880
rect 1912 24828 1918 24880
rect 2130 24828 2136 24880
rect 2188 24828 2194 24880
rect 2961 24871 3019 24877
rect 2961 24837 2973 24871
rect 3007 24868 3019 24871
rect 3326 24868 3332 24880
rect 3007 24840 3332 24868
rect 3007 24837 3019 24840
rect 2961 24831 3019 24837
rect 3326 24828 3332 24840
rect 3384 24828 3390 24880
rect 4522 24828 4528 24880
rect 4580 24828 4586 24880
rect 5902 24828 5908 24880
rect 5960 24868 5966 24880
rect 6104 24868 6132 24908
rect 8110 24896 8116 24908
rect 8168 24936 8174 24948
rect 9858 24936 9864 24948
rect 8168 24908 9864 24936
rect 8168 24896 8174 24908
rect 9858 24896 9864 24908
rect 9916 24896 9922 24948
rect 10134 24896 10140 24948
rect 10192 24936 10198 24948
rect 10597 24939 10655 24945
rect 10597 24936 10609 24939
rect 10192 24908 10609 24936
rect 10192 24896 10198 24908
rect 10597 24905 10609 24908
rect 10643 24905 10655 24939
rect 10597 24899 10655 24905
rect 11882 24896 11888 24948
rect 11940 24936 11946 24948
rect 12529 24939 12587 24945
rect 12529 24936 12541 24939
rect 11940 24908 12541 24936
rect 11940 24896 11946 24908
rect 12529 24905 12541 24908
rect 12575 24905 12587 24939
rect 14366 24936 14372 24948
rect 12529 24899 12587 24905
rect 13464 24908 14372 24936
rect 5960 24840 6132 24868
rect 5960 24828 5966 24840
rect 6546 24828 6552 24880
rect 6604 24828 6610 24880
rect 9490 24828 9496 24880
rect 9548 24828 9554 24880
rect 10778 24828 10784 24880
rect 10836 24868 10842 24880
rect 12434 24868 12440 24880
rect 10836 24840 12440 24868
rect 10836 24828 10842 24840
rect 12434 24828 12440 24840
rect 12492 24828 12498 24880
rect 842 24760 848 24812
rect 900 24800 906 24812
rect 1581 24803 1639 24809
rect 1581 24800 1593 24803
rect 900 24772 1593 24800
rect 900 24760 906 24772
rect 1581 24769 1593 24772
rect 1627 24769 1639 24803
rect 1581 24763 1639 24769
rect 2225 24803 2283 24809
rect 2225 24769 2237 24803
rect 2271 24800 2283 24803
rect 2498 24800 2504 24812
rect 2271 24772 2504 24800
rect 2271 24769 2283 24772
rect 2225 24763 2283 24769
rect 2498 24760 2504 24772
rect 2556 24760 2562 24812
rect 2593 24803 2651 24809
rect 2593 24769 2605 24803
rect 2639 24800 2651 24803
rect 3418 24800 3424 24812
rect 2639 24772 3424 24800
rect 2639 24769 2651 24772
rect 2593 24763 2651 24769
rect 3418 24760 3424 24772
rect 3476 24760 3482 24812
rect 4540 24800 4568 24828
rect 4707 24803 4765 24809
rect 4707 24800 4719 24803
rect 4540 24772 4719 24800
rect 4707 24769 4719 24772
rect 4753 24800 4765 24803
rect 6564 24800 6592 24828
rect 4753 24772 6592 24800
rect 4753 24769 4765 24772
rect 4707 24763 4765 24769
rect 6822 24760 6828 24812
rect 6880 24760 6886 24812
rect 7282 24760 7288 24812
rect 7340 24800 7346 24812
rect 8754 24809 8760 24812
rect 7653 24803 7711 24809
rect 7653 24800 7665 24803
rect 7340 24772 7665 24800
rect 7340 24760 7346 24772
rect 7653 24769 7665 24772
rect 7699 24769 7711 24803
rect 7653 24763 7711 24769
rect 8711 24803 8760 24809
rect 8711 24769 8723 24803
rect 8757 24769 8760 24803
rect 8711 24763 8760 24769
rect 8754 24760 8760 24763
rect 8812 24760 8818 24812
rect 9508 24800 9536 24828
rect 13464 24819 13492 24908
rect 14366 24896 14372 24908
rect 14424 24896 14430 24948
rect 18138 24936 18144 24948
rect 15394 24908 18144 24936
rect 13814 24828 13820 24880
rect 13872 24868 13878 24880
rect 13872 24840 15148 24868
rect 13872 24828 13878 24840
rect 13447 24813 13505 24819
rect 13447 24812 13459 24813
rect 13493 24812 13505 24813
rect 9859 24803 9917 24809
rect 9859 24800 9871 24803
rect 9508 24772 9871 24800
rect 9859 24769 9871 24772
rect 9905 24800 9917 24803
rect 10502 24800 10508 24812
rect 9905 24772 10508 24800
rect 9905 24769 9917 24772
rect 9859 24763 9917 24769
rect 10502 24760 10508 24772
rect 10560 24760 10566 24812
rect 11238 24760 11244 24812
rect 11296 24760 11302 24812
rect 11791 24803 11849 24809
rect 11791 24769 11803 24803
rect 11837 24800 11849 24803
rect 12526 24800 12532 24812
rect 11837 24772 12532 24800
rect 11837 24769 11849 24772
rect 11791 24763 11849 24769
rect 12526 24760 12532 24772
rect 12584 24760 12590 24812
rect 12986 24760 12992 24812
rect 13044 24800 13050 24812
rect 13446 24800 13452 24812
rect 13044 24772 13452 24800
rect 13044 24760 13050 24772
rect 13446 24760 13452 24772
rect 13504 24760 13510 24812
rect 14553 24803 14611 24809
rect 14553 24800 14565 24803
rect 14200 24772 14565 24800
rect 2406 24692 2412 24744
rect 2464 24692 2470 24744
rect 3878 24692 3884 24744
rect 3936 24732 3942 24744
rect 4433 24735 4491 24741
rect 4433 24732 4445 24735
rect 3936 24704 4445 24732
rect 3936 24692 3942 24704
rect 4433 24701 4445 24704
rect 4479 24701 4491 24735
rect 4433 24695 4491 24701
rect 5718 24664 5724 24676
rect 5368 24636 5724 24664
rect 3145 24599 3203 24605
rect 3145 24565 3157 24599
rect 3191 24596 3203 24599
rect 3602 24596 3608 24608
rect 3191 24568 3608 24596
rect 3191 24565 3203 24568
rect 3145 24559 3203 24565
rect 3602 24556 3608 24568
rect 3660 24556 3666 24608
rect 4338 24556 4344 24608
rect 4396 24596 4402 24608
rect 5368 24596 5396 24636
rect 5718 24624 5724 24636
rect 5776 24624 5782 24676
rect 6840 24664 6868 24760
rect 7374 24692 7380 24744
rect 7432 24732 7438 24744
rect 7834 24732 7840 24744
rect 7432 24704 7840 24732
rect 7432 24692 7438 24704
rect 7834 24692 7840 24704
rect 7892 24692 7898 24744
rect 8573 24735 8631 24741
rect 8573 24732 8585 24735
rect 7926 24704 8585 24732
rect 7098 24664 7104 24676
rect 6840 24636 7104 24664
rect 7098 24624 7104 24636
rect 7156 24664 7162 24676
rect 7926 24664 7954 24704
rect 8573 24701 8585 24704
rect 8619 24701 8631 24735
rect 8573 24695 8631 24701
rect 8849 24735 8907 24741
rect 8849 24701 8861 24735
rect 8895 24732 8907 24735
rect 9030 24732 9036 24744
rect 8895 24704 9036 24732
rect 8895 24701 8907 24704
rect 8849 24695 8907 24701
rect 9030 24692 9036 24704
rect 9088 24692 9094 24744
rect 9214 24692 9220 24744
rect 9272 24732 9278 24744
rect 9585 24735 9643 24741
rect 9585 24732 9597 24735
rect 9272 24704 9597 24732
rect 9272 24692 9278 24704
rect 9585 24701 9597 24704
rect 9631 24701 9643 24735
rect 9585 24695 9643 24701
rect 11256 24732 11284 24760
rect 11517 24735 11575 24741
rect 11517 24732 11529 24735
rect 11256 24704 11529 24732
rect 7156 24636 7954 24664
rect 7156 24624 7162 24636
rect 8294 24624 8300 24676
rect 8352 24624 8358 24676
rect 4396 24568 5396 24596
rect 5445 24599 5503 24605
rect 4396 24556 4402 24568
rect 5445 24565 5457 24599
rect 5491 24596 5503 24599
rect 5626 24596 5632 24608
rect 5491 24568 5632 24596
rect 5491 24565 5503 24568
rect 5445 24559 5503 24565
rect 5626 24556 5632 24568
rect 5684 24556 5690 24608
rect 8386 24556 8392 24608
rect 8444 24596 8450 24608
rect 9232 24596 9260 24692
rect 9398 24624 9404 24676
rect 9456 24664 9462 24676
rect 11256 24664 11284 24704
rect 11517 24701 11529 24704
rect 11563 24701 11575 24735
rect 11517 24695 11575 24701
rect 13173 24735 13231 24741
rect 13173 24701 13185 24735
rect 13219 24701 13231 24735
rect 13173 24695 13231 24701
rect 9456 24636 9674 24664
rect 9456 24624 9462 24636
rect 8444 24568 9260 24596
rect 8444 24556 8450 24568
rect 9490 24556 9496 24608
rect 9548 24556 9554 24608
rect 9646 24596 9674 24636
rect 10242 24636 11284 24664
rect 10242 24596 10270 24636
rect 13188 24608 13216 24695
rect 14200 24673 14228 24772
rect 14553 24769 14565 24772
rect 14599 24769 14611 24803
rect 14553 24763 14611 24769
rect 14734 24760 14740 24812
rect 14792 24760 14798 24812
rect 14918 24760 14924 24812
rect 14976 24800 14982 24812
rect 15013 24803 15071 24809
rect 15013 24800 15025 24803
rect 14976 24772 15025 24800
rect 14976 24760 14982 24772
rect 15013 24769 15025 24772
rect 15059 24769 15071 24803
rect 15120 24800 15148 24840
rect 15271 24833 15329 24839
rect 15271 24800 15283 24833
rect 15120 24799 15283 24800
rect 15317 24830 15329 24833
rect 15317 24800 15330 24830
rect 15394 24800 15422 24908
rect 18138 24896 18144 24908
rect 18196 24896 18202 24948
rect 18693 24939 18751 24945
rect 18693 24905 18705 24939
rect 18739 24936 18751 24939
rect 18874 24936 18880 24948
rect 18739 24908 18880 24936
rect 18739 24905 18751 24908
rect 18693 24899 18751 24905
rect 18874 24896 18880 24908
rect 18932 24896 18938 24948
rect 19518 24896 19524 24948
rect 19576 24936 19582 24948
rect 20714 24936 20720 24948
rect 19576 24908 20720 24936
rect 19576 24896 19582 24908
rect 20714 24896 20720 24908
rect 20772 24896 20778 24948
rect 20898 24896 20904 24948
rect 20956 24936 20962 24948
rect 20993 24939 21051 24945
rect 20993 24936 21005 24939
rect 20956 24908 21005 24936
rect 20956 24896 20962 24908
rect 20993 24905 21005 24908
rect 21039 24905 21051 24939
rect 20993 24899 21051 24905
rect 22002 24896 22008 24948
rect 22060 24936 22066 24948
rect 22186 24936 22192 24948
rect 22060 24908 22192 24936
rect 22060 24896 22066 24908
rect 22186 24896 22192 24908
rect 22244 24896 22250 24948
rect 17770 24868 17776 24880
rect 17328 24840 17776 24868
rect 17328 24809 17356 24840
rect 17770 24828 17776 24840
rect 17828 24868 17834 24880
rect 19886 24877 19892 24880
rect 19880 24868 19892 24877
rect 17828 24840 19334 24868
rect 19847 24840 19892 24868
rect 17828 24828 17834 24840
rect 18892 24812 18920 24840
rect 15317 24799 15422 24800
rect 15120 24772 15422 24799
rect 17313 24803 17371 24809
rect 15013 24763 15071 24769
rect 17313 24769 17325 24803
rect 17359 24769 17371 24803
rect 17313 24763 17371 24769
rect 17402 24760 17408 24812
rect 17460 24800 17466 24812
rect 17569 24803 17627 24809
rect 17569 24800 17581 24803
rect 17460 24772 17581 24800
rect 17460 24760 17466 24772
rect 17569 24769 17581 24772
rect 17615 24769 17627 24803
rect 17569 24763 17627 24769
rect 18598 24760 18604 24812
rect 18656 24760 18662 24812
rect 18690 24760 18696 24812
rect 18748 24800 18754 24812
rect 18785 24803 18843 24809
rect 18785 24800 18797 24803
rect 18748 24772 18797 24800
rect 18748 24760 18754 24772
rect 18785 24769 18797 24772
rect 18831 24769 18843 24803
rect 18785 24763 18843 24769
rect 18874 24760 18880 24812
rect 18932 24760 18938 24812
rect 18966 24760 18972 24812
rect 19024 24800 19030 24812
rect 19153 24803 19211 24809
rect 19153 24800 19165 24803
rect 19024 24772 19165 24800
rect 19024 24760 19030 24772
rect 19153 24769 19165 24772
rect 19199 24769 19211 24803
rect 19306 24800 19334 24840
rect 19880 24831 19892 24840
rect 19886 24828 19892 24831
rect 19944 24828 19950 24880
rect 20070 24828 20076 24880
rect 20128 24828 20134 24880
rect 19613 24803 19671 24809
rect 19613 24800 19625 24803
rect 19306 24772 19625 24800
rect 19153 24763 19211 24769
rect 19613 24769 19625 24772
rect 19659 24769 19671 24803
rect 20088 24800 20116 24828
rect 19613 24763 19671 24769
rect 19720 24772 20116 24800
rect 21177 24803 21235 24809
rect 18616 24732 18644 24760
rect 19061 24735 19119 24741
rect 19061 24732 19073 24735
rect 18616 24704 19073 24732
rect 19061 24701 19073 24704
rect 19107 24701 19119 24735
rect 19061 24695 19119 24701
rect 19334 24692 19340 24744
rect 19392 24732 19398 24744
rect 19720 24732 19748 24772
rect 21177 24769 21189 24803
rect 21223 24769 21235 24803
rect 21177 24763 21235 24769
rect 19392 24704 19748 24732
rect 19392 24692 19398 24704
rect 14185 24667 14243 24673
rect 14185 24633 14197 24667
rect 14231 24664 14243 24667
rect 14366 24664 14372 24676
rect 14231 24636 14372 24664
rect 14231 24633 14243 24636
rect 14185 24627 14243 24633
rect 14366 24624 14372 24636
rect 14424 24624 14430 24676
rect 18877 24667 18935 24673
rect 14476 24636 15056 24664
rect 9646 24568 10270 24596
rect 13170 24556 13176 24608
rect 13228 24596 13234 24608
rect 14476 24596 14504 24636
rect 15028 24608 15056 24636
rect 18877 24633 18889 24667
rect 18923 24664 18935 24667
rect 19245 24667 19303 24673
rect 19245 24664 19257 24667
rect 18923 24636 19257 24664
rect 18923 24633 18935 24636
rect 18877 24627 18935 24633
rect 19245 24633 19257 24636
rect 19291 24633 19303 24667
rect 19245 24627 19303 24633
rect 13228 24568 14504 24596
rect 13228 24556 13234 24568
rect 14642 24556 14648 24608
rect 14700 24556 14706 24608
rect 15010 24556 15016 24608
rect 15068 24556 15074 24608
rect 16022 24556 16028 24608
rect 16080 24556 16086 24608
rect 18969 24599 19027 24605
rect 18969 24565 18981 24599
rect 19015 24596 19027 24599
rect 21192 24596 21220 24763
rect 19015 24568 21220 24596
rect 19015 24565 19027 24568
rect 18969 24559 19027 24565
rect 21450 24556 21456 24608
rect 21508 24556 21514 24608
rect 1104 24506 21896 24528
rect 1104 24454 3549 24506
rect 3601 24454 3613 24506
rect 3665 24454 3677 24506
rect 3729 24454 3741 24506
rect 3793 24454 3805 24506
rect 3857 24454 8747 24506
rect 8799 24454 8811 24506
rect 8863 24454 8875 24506
rect 8927 24454 8939 24506
rect 8991 24454 9003 24506
rect 9055 24454 13945 24506
rect 13997 24454 14009 24506
rect 14061 24454 14073 24506
rect 14125 24454 14137 24506
rect 14189 24454 14201 24506
rect 14253 24454 19143 24506
rect 19195 24454 19207 24506
rect 19259 24454 19271 24506
rect 19323 24454 19335 24506
rect 19387 24454 19399 24506
rect 19451 24454 21896 24506
rect 1104 24432 21896 24454
rect 1581 24395 1639 24401
rect 1581 24361 1593 24395
rect 1627 24392 1639 24395
rect 1762 24392 1768 24404
rect 1627 24364 1768 24392
rect 1627 24361 1639 24364
rect 1581 24355 1639 24361
rect 1762 24352 1768 24364
rect 1820 24352 1826 24404
rect 2498 24352 2504 24404
rect 2556 24392 2562 24404
rect 2685 24395 2743 24401
rect 2685 24392 2697 24395
rect 2556 24364 2697 24392
rect 2556 24352 2562 24364
rect 2685 24361 2697 24364
rect 2731 24361 2743 24395
rect 2685 24355 2743 24361
rect 3234 24352 3240 24404
rect 3292 24392 3298 24404
rect 4246 24392 4252 24404
rect 3292 24364 4252 24392
rect 3292 24352 3298 24364
rect 4246 24352 4252 24364
rect 4304 24352 4310 24404
rect 5626 24392 5632 24404
rect 5368 24364 5632 24392
rect 1394 24284 1400 24336
rect 1452 24324 1458 24336
rect 1452 24296 1716 24324
rect 1452 24284 1458 24296
rect 1688 24265 1716 24296
rect 4982 24284 4988 24336
rect 5040 24324 5046 24336
rect 5368 24333 5396 24364
rect 5626 24352 5632 24364
rect 5684 24352 5690 24404
rect 5718 24352 5724 24404
rect 5776 24392 5782 24404
rect 8205 24395 8263 24401
rect 5776 24364 7878 24392
rect 5776 24352 5782 24364
rect 5353 24327 5411 24333
rect 5040 24296 5304 24324
rect 5040 24284 5046 24296
rect 1673 24259 1731 24265
rect 1673 24225 1685 24259
rect 1719 24225 1731 24259
rect 5276 24256 5304 24296
rect 5353 24293 5365 24327
rect 5399 24293 5411 24327
rect 5353 24287 5411 24293
rect 5767 24259 5825 24265
rect 5276 24228 5672 24256
rect 1673 24219 1731 24225
rect 750 24148 756 24200
rect 808 24188 814 24200
rect 1397 24191 1455 24197
rect 1397 24188 1409 24191
rect 808 24160 1409 24188
rect 808 24148 814 24160
rect 1397 24157 1409 24160
rect 1443 24157 1455 24191
rect 1397 24151 1455 24157
rect 1486 24148 1492 24200
rect 1544 24188 1550 24200
rect 1544 24161 1992 24188
rect 1544 24160 1943 24161
rect 1544 24148 1550 24160
rect 1931 24127 1943 24160
rect 1977 24127 1992 24161
rect 2590 24148 2596 24200
rect 2648 24188 2654 24200
rect 2648 24160 4476 24188
rect 2648 24148 2654 24160
rect 1931 24121 1992 24127
rect 1964 24120 1992 24121
rect 4338 24120 4344 24132
rect 1964 24092 4344 24120
rect 4338 24080 4344 24092
rect 4396 24080 4402 24132
rect 4448 24052 4476 24160
rect 4522 24148 4528 24200
rect 4580 24148 4586 24200
rect 4709 24191 4767 24197
rect 4709 24157 4721 24191
rect 4755 24188 4767 24191
rect 4798 24188 4804 24200
rect 4755 24160 4804 24188
rect 4755 24157 4767 24160
rect 4709 24151 4767 24157
rect 4798 24148 4804 24160
rect 4856 24148 4862 24200
rect 4890 24148 4896 24200
rect 4948 24148 4954 24200
rect 5644 24197 5672 24228
rect 5767 24225 5779 24259
rect 5813 24256 5825 24259
rect 6086 24256 6092 24268
rect 5813 24228 6092 24256
rect 5813 24225 5825 24228
rect 5767 24219 5825 24225
rect 6086 24216 6092 24228
rect 6144 24216 6150 24268
rect 7850 24256 7878 24364
rect 8205 24361 8217 24395
rect 8251 24392 8263 24395
rect 8294 24392 8300 24404
rect 8251 24364 8300 24392
rect 8251 24361 8263 24364
rect 8205 24355 8263 24361
rect 8294 24352 8300 24364
rect 8352 24352 8358 24404
rect 9490 24352 9496 24404
rect 9548 24392 9554 24404
rect 10042 24392 10048 24404
rect 9548 24364 10048 24392
rect 9548 24352 9554 24364
rect 10042 24352 10048 24364
rect 10100 24352 10106 24404
rect 12434 24392 12440 24404
rect 10152 24364 12440 24392
rect 10152 24256 10180 24364
rect 7850 24228 10180 24256
rect 11072 24228 11834 24256
rect 5629 24191 5687 24197
rect 5629 24157 5641 24191
rect 5675 24157 5687 24191
rect 5629 24151 5687 24157
rect 5902 24148 5908 24200
rect 5960 24148 5966 24200
rect 6822 24148 6828 24200
rect 6880 24188 6886 24200
rect 7193 24191 7251 24197
rect 7193 24188 7205 24191
rect 6880 24160 7205 24188
rect 6880 24148 6886 24160
rect 7193 24157 7205 24160
rect 7239 24157 7251 24191
rect 7451 24191 7509 24197
rect 7451 24188 7463 24191
rect 7450 24158 7463 24188
rect 7193 24151 7251 24157
rect 7417 24157 7463 24158
rect 7497 24157 7509 24191
rect 7417 24151 7509 24157
rect 4540 24120 4568 24148
rect 4908 24120 4936 24148
rect 7417 24130 7478 24151
rect 7558 24148 7564 24200
rect 7616 24188 7622 24200
rect 7926 24188 7932 24200
rect 7616 24160 7932 24188
rect 7616 24148 7622 24160
rect 7926 24148 7932 24160
rect 7984 24148 7990 24200
rect 10042 24148 10048 24200
rect 10100 24148 10106 24200
rect 10137 24191 10195 24197
rect 10137 24157 10149 24191
rect 10183 24157 10195 24191
rect 10137 24151 10195 24157
rect 7417 24120 7445 24130
rect 10152 24120 10180 24151
rect 10318 24148 10324 24200
rect 10376 24188 10382 24200
rect 10411 24191 10469 24197
rect 10411 24188 10423 24191
rect 10376 24160 10423 24188
rect 10376 24148 10382 24160
rect 10411 24157 10423 24160
rect 10457 24157 10469 24191
rect 10411 24151 10469 24157
rect 11072 24120 11100 24228
rect 11517 24191 11575 24197
rect 11517 24188 11529 24191
rect 4540 24092 4936 24120
rect 6472 24092 7445 24120
rect 8266 24092 11100 24120
rect 11164 24160 11529 24188
rect 6472 24052 6500 24092
rect 4448 24024 6500 24052
rect 6546 24012 6552 24064
rect 6604 24012 6610 24064
rect 7742 24012 7748 24064
rect 7800 24052 7806 24064
rect 8266 24052 8294 24092
rect 11164 24064 11192 24160
rect 11517 24157 11529 24160
rect 11563 24157 11575 24191
rect 11517 24151 11575 24157
rect 11701 24191 11759 24197
rect 11701 24157 11713 24191
rect 11747 24157 11759 24191
rect 11701 24151 11759 24157
rect 11238 24080 11244 24132
rect 11296 24120 11302 24132
rect 11716 24120 11744 24151
rect 11296 24092 11744 24120
rect 11806 24120 11834 24228
rect 12360 24188 12388 24364
rect 12434 24352 12440 24364
rect 12492 24352 12498 24404
rect 13170 24392 13176 24404
rect 12544 24364 13176 24392
rect 12544 24324 12572 24364
rect 13170 24352 13176 24364
rect 13228 24352 13234 24404
rect 14366 24352 14372 24404
rect 14424 24352 14430 24404
rect 14642 24352 14648 24404
rect 14700 24352 14706 24404
rect 14737 24395 14795 24401
rect 14737 24361 14749 24395
rect 14783 24392 14795 24395
rect 14826 24392 14832 24404
rect 14783 24364 14832 24392
rect 14783 24361 14795 24364
rect 14737 24355 14795 24361
rect 14826 24352 14832 24364
rect 14884 24352 14890 24404
rect 15470 24352 15476 24404
rect 15528 24392 15534 24404
rect 16942 24392 16948 24404
rect 15528 24364 16948 24392
rect 15528 24352 15534 24364
rect 16942 24352 16948 24364
rect 17000 24352 17006 24404
rect 17221 24395 17279 24401
rect 17221 24361 17233 24395
rect 17267 24392 17279 24395
rect 17402 24392 17408 24404
rect 17267 24364 17408 24392
rect 17267 24361 17279 24364
rect 17221 24355 17279 24361
rect 17402 24352 17408 24364
rect 17460 24352 17466 24404
rect 18601 24395 18659 24401
rect 17604 24364 18276 24392
rect 12452 24296 12572 24324
rect 12452 24265 12480 24296
rect 14384 24265 14412 24352
rect 12437 24259 12495 24265
rect 12437 24225 12449 24259
rect 12483 24225 12495 24259
rect 12437 24219 12495 24225
rect 14369 24259 14427 24265
rect 14369 24225 14381 24259
rect 14415 24225 14427 24259
rect 14369 24219 14427 24225
rect 12711 24191 12769 24197
rect 12711 24188 12723 24191
rect 12360 24160 12723 24188
rect 12711 24157 12723 24160
rect 12757 24188 12769 24191
rect 13814 24188 13820 24200
rect 12757 24160 13820 24188
rect 12757 24157 12769 24160
rect 12711 24151 12769 24157
rect 13814 24148 13820 24160
rect 13872 24148 13878 24200
rect 14274 24148 14280 24200
rect 14332 24148 14338 24200
rect 14660 24197 14688 24352
rect 16025 24327 16083 24333
rect 16025 24293 16037 24327
rect 16071 24324 16083 24327
rect 16114 24324 16120 24336
rect 16071 24296 16120 24324
rect 16071 24293 16083 24296
rect 16025 24287 16083 24293
rect 16114 24284 16120 24296
rect 16172 24284 16178 24336
rect 15565 24259 15623 24265
rect 15565 24256 15577 24259
rect 15212 24228 15577 24256
rect 15212 24200 15240 24228
rect 15565 24225 15577 24228
rect 15611 24225 15623 24259
rect 15565 24219 15623 24225
rect 16577 24259 16635 24265
rect 16577 24225 16589 24259
rect 16623 24256 16635 24259
rect 17494 24256 17500 24268
rect 16623 24228 17500 24256
rect 16623 24225 16635 24228
rect 16577 24219 16635 24225
rect 17494 24216 17500 24228
rect 17552 24216 17558 24268
rect 17604 24265 17632 24364
rect 18248 24324 18276 24364
rect 18601 24361 18613 24395
rect 18647 24392 18659 24395
rect 18690 24392 18696 24404
rect 18647 24364 18696 24392
rect 18647 24361 18659 24364
rect 18601 24355 18659 24361
rect 18690 24352 18696 24364
rect 18748 24352 18754 24404
rect 18874 24352 18880 24404
rect 18932 24392 18938 24404
rect 18932 24364 19104 24392
rect 18932 24352 18938 24364
rect 18248 24296 19012 24324
rect 18984 24268 19012 24296
rect 19076 24268 19104 24364
rect 20530 24352 20536 24404
rect 20588 24352 20594 24404
rect 20622 24352 20628 24404
rect 20680 24352 20686 24404
rect 20809 24395 20867 24401
rect 20809 24361 20821 24395
rect 20855 24392 20867 24395
rect 21082 24392 21088 24404
rect 20855 24364 21088 24392
rect 20855 24361 20867 24364
rect 20809 24355 20867 24361
rect 21082 24352 21088 24364
rect 21140 24352 21146 24404
rect 17589 24259 17647 24265
rect 17589 24225 17601 24259
rect 17635 24225 17647 24259
rect 17589 24219 17647 24225
rect 18966 24216 18972 24268
rect 19024 24216 19030 24268
rect 19058 24216 19064 24268
rect 19116 24256 19122 24268
rect 19245 24259 19303 24265
rect 19245 24256 19257 24259
rect 19116 24228 19257 24256
rect 19116 24216 19122 24228
rect 19245 24225 19257 24228
rect 19291 24225 19303 24259
rect 19245 24219 19303 24225
rect 14645 24191 14703 24197
rect 14645 24157 14657 24191
rect 14691 24157 14703 24191
rect 14645 24151 14703 24157
rect 14918 24148 14924 24200
rect 14976 24148 14982 24200
rect 15194 24148 15200 24200
rect 15252 24148 15258 24200
rect 15286 24148 15292 24200
rect 15344 24188 15350 24200
rect 15381 24191 15439 24197
rect 15381 24188 15393 24191
rect 15344 24160 15393 24188
rect 15344 24148 15350 24160
rect 15381 24157 15393 24160
rect 15427 24157 15439 24191
rect 15381 24151 15439 24157
rect 16298 24148 16304 24200
rect 16356 24148 16362 24200
rect 16390 24148 16396 24200
rect 16448 24197 16454 24200
rect 16448 24191 16476 24197
rect 16464 24157 16476 24191
rect 16448 24151 16476 24157
rect 17847 24161 17905 24167
rect 16448 24148 16454 24151
rect 14366 24120 14372 24132
rect 11806 24092 14372 24120
rect 11296 24080 11302 24092
rect 14366 24080 14372 24092
rect 14424 24080 14430 24132
rect 14553 24123 14611 24129
rect 14553 24089 14565 24123
rect 14599 24120 14611 24123
rect 14826 24120 14832 24132
rect 14599 24092 14832 24120
rect 14599 24089 14611 24092
rect 14553 24083 14611 24089
rect 14826 24080 14832 24092
rect 14884 24080 14890 24132
rect 17494 24080 17500 24132
rect 17552 24120 17558 24132
rect 17678 24120 17684 24132
rect 17552 24092 17684 24120
rect 17552 24080 17558 24092
rect 17678 24080 17684 24092
rect 17736 24080 17742 24132
rect 17847 24127 17859 24161
rect 17893 24158 17905 24161
rect 17893 24132 17906 24158
rect 18874 24148 18880 24200
rect 18932 24188 18938 24200
rect 18932 24160 19748 24188
rect 18932 24148 18938 24160
rect 19720 24132 19748 24160
rect 17847 24121 17868 24127
rect 17862 24080 17868 24121
rect 17920 24120 17926 24132
rect 18046 24120 18052 24132
rect 17920 24092 18052 24120
rect 17920 24080 17926 24092
rect 18046 24080 18052 24092
rect 18104 24080 18110 24132
rect 19334 24080 19340 24132
rect 19392 24120 19398 24132
rect 19490 24123 19548 24129
rect 19490 24120 19502 24123
rect 19392 24092 19502 24120
rect 19392 24080 19398 24092
rect 19490 24089 19502 24092
rect 19536 24089 19548 24123
rect 19490 24083 19548 24089
rect 19702 24080 19708 24132
rect 19760 24120 19766 24132
rect 19886 24120 19892 24132
rect 19760 24092 19892 24120
rect 19760 24080 19766 24092
rect 19886 24080 19892 24092
rect 19944 24080 19950 24132
rect 7800 24024 8294 24052
rect 7800 24012 7806 24024
rect 9858 24012 9864 24064
rect 9916 24012 9922 24064
rect 10134 24012 10140 24064
rect 10192 24052 10198 24064
rect 10870 24052 10876 24064
rect 10192 24024 10876 24052
rect 10192 24012 10198 24024
rect 10870 24012 10876 24024
rect 10928 24012 10934 24064
rect 11146 24012 11152 24064
rect 11204 24012 11210 24064
rect 11698 24012 11704 24064
rect 11756 24012 11762 24064
rect 13446 24012 13452 24064
rect 13504 24012 13510 24064
rect 13814 24012 13820 24064
rect 13872 24052 13878 24064
rect 14642 24052 14648 24064
rect 13872 24024 14648 24052
rect 13872 24012 13878 24024
rect 14642 24012 14648 24024
rect 14700 24052 14706 24064
rect 16298 24052 16304 24064
rect 14700 24024 16304 24052
rect 14700 24012 14706 24024
rect 16298 24012 16304 24024
rect 16356 24012 16362 24064
rect 17310 24012 17316 24064
rect 17368 24052 17374 24064
rect 20162 24052 20168 24064
rect 17368 24024 20168 24052
rect 17368 24012 17374 24024
rect 20162 24012 20168 24024
rect 20220 24012 20226 24064
rect 20548 24052 20576 24352
rect 20640 24256 20668 24352
rect 20993 24259 21051 24265
rect 20993 24256 21005 24259
rect 20640 24228 21005 24256
rect 20993 24225 21005 24228
rect 21039 24225 21051 24259
rect 20993 24219 21051 24225
rect 20622 24148 20628 24200
rect 20680 24188 20686 24200
rect 20717 24191 20775 24197
rect 20717 24188 20729 24191
rect 20680 24160 20729 24188
rect 20680 24148 20686 24160
rect 20717 24157 20729 24160
rect 20763 24157 20775 24191
rect 20717 24151 20775 24157
rect 20898 24148 20904 24200
rect 20956 24188 20962 24200
rect 21269 24191 21327 24197
rect 21269 24188 21281 24191
rect 20956 24160 21281 24188
rect 20956 24148 20962 24160
rect 21269 24157 21281 24160
rect 21315 24157 21327 24191
rect 21269 24151 21327 24157
rect 21082 24080 21088 24132
rect 21140 24120 21146 24132
rect 21542 24120 21548 24132
rect 21140 24092 21548 24120
rect 21140 24080 21146 24092
rect 21542 24080 21548 24092
rect 21600 24080 21606 24132
rect 20625 24055 20683 24061
rect 20625 24052 20637 24055
rect 20548 24024 20637 24052
rect 20625 24021 20637 24024
rect 20671 24021 20683 24055
rect 20625 24015 20683 24021
rect 20990 24012 20996 24064
rect 21048 24012 21054 24064
rect 21453 24055 21511 24061
rect 21453 24021 21465 24055
rect 21499 24052 21511 24055
rect 22186 24052 22192 24064
rect 21499 24024 22192 24052
rect 21499 24021 21511 24024
rect 21453 24015 21511 24021
rect 22186 24012 22192 24024
rect 22244 24012 22250 24064
rect 1104 23962 22056 23984
rect 1104 23910 6148 23962
rect 6200 23910 6212 23962
rect 6264 23910 6276 23962
rect 6328 23910 6340 23962
rect 6392 23910 6404 23962
rect 6456 23910 11346 23962
rect 11398 23910 11410 23962
rect 11462 23910 11474 23962
rect 11526 23910 11538 23962
rect 11590 23910 11602 23962
rect 11654 23910 16544 23962
rect 16596 23910 16608 23962
rect 16660 23910 16672 23962
rect 16724 23910 16736 23962
rect 16788 23910 16800 23962
rect 16852 23910 21742 23962
rect 21794 23910 21806 23962
rect 21858 23910 21870 23962
rect 21922 23910 21934 23962
rect 21986 23910 21998 23962
rect 22050 23910 22056 23962
rect 1104 23888 22056 23910
rect 5920 23820 9536 23848
rect 5350 23740 5356 23792
rect 5408 23780 5414 23792
rect 5920 23780 5948 23820
rect 5408 23752 5948 23780
rect 5408 23740 5414 23752
rect 1394 23672 1400 23724
rect 1452 23672 1458 23724
rect 1671 23715 1729 23721
rect 1671 23681 1683 23715
rect 1717 23712 1729 23715
rect 1762 23712 1768 23724
rect 1717 23684 1768 23712
rect 1717 23681 1729 23684
rect 1671 23675 1729 23681
rect 1762 23672 1768 23684
rect 1820 23672 1826 23724
rect 3878 23672 3884 23724
rect 3936 23712 3942 23724
rect 4893 23715 4951 23721
rect 4893 23712 4905 23715
rect 3936 23684 4905 23712
rect 3936 23672 3942 23684
rect 4893 23681 4905 23684
rect 4939 23681 4951 23715
rect 5166 23712 5172 23724
rect 5127 23684 5172 23712
rect 4893 23675 4951 23681
rect 5166 23672 5172 23684
rect 5224 23672 5230 23724
rect 6546 23672 6552 23724
rect 6604 23712 6610 23724
rect 7009 23715 7067 23721
rect 7009 23712 7021 23715
rect 6604 23684 7021 23712
rect 6604 23672 6610 23684
rect 7009 23681 7021 23684
rect 7055 23681 7067 23715
rect 7009 23675 7067 23681
rect 7377 23715 7435 23721
rect 7377 23681 7389 23715
rect 7423 23681 7435 23715
rect 7377 23675 7435 23681
rect 2774 23604 2780 23656
rect 2832 23604 2838 23656
rect 3053 23647 3111 23653
rect 3053 23613 3065 23647
rect 3099 23644 3111 23647
rect 3970 23644 3976 23656
rect 3099 23616 3976 23644
rect 3099 23613 3111 23616
rect 3053 23607 3111 23613
rect 3970 23604 3976 23616
rect 4028 23604 4034 23656
rect 7392 23644 7420 23675
rect 7466 23672 7472 23724
rect 7524 23672 7530 23724
rect 7558 23672 7564 23724
rect 7616 23712 7622 23724
rect 7929 23715 7987 23721
rect 7929 23712 7941 23715
rect 7616 23684 7941 23712
rect 7616 23672 7622 23684
rect 7929 23681 7941 23684
rect 7975 23712 7987 23715
rect 8110 23712 8116 23724
rect 7975 23684 8116 23712
rect 7975 23681 7987 23684
rect 7929 23675 7987 23681
rect 8110 23672 8116 23684
rect 8168 23672 8174 23724
rect 6840 23616 7420 23644
rect 7484 23644 7512 23672
rect 7745 23647 7803 23653
rect 7745 23644 7757 23647
rect 7484 23616 7757 23644
rect 4430 23576 4436 23588
rect 2056 23548 4436 23576
rect 658 23468 664 23520
rect 716 23508 722 23520
rect 2056 23508 2084 23548
rect 4430 23536 4436 23548
rect 4488 23536 4494 23588
rect 6840 23585 6868 23616
rect 7745 23613 7757 23616
rect 7791 23613 7803 23647
rect 7745 23607 7803 23613
rect 8018 23604 8024 23656
rect 8076 23604 8082 23656
rect 8294 23604 8300 23656
rect 8352 23644 8358 23656
rect 8389 23647 8447 23653
rect 8389 23644 8401 23647
rect 8352 23616 8401 23644
rect 8352 23604 8358 23616
rect 8389 23613 8401 23616
rect 8435 23613 8447 23647
rect 8665 23647 8723 23653
rect 8665 23644 8677 23647
rect 8389 23607 8447 23613
rect 8496 23616 8677 23644
rect 6825 23579 6883 23585
rect 6825 23545 6837 23579
rect 6871 23545 6883 23579
rect 8036 23576 8064 23604
rect 8496 23576 8524 23616
rect 8665 23613 8677 23616
rect 8711 23613 8723 23647
rect 8665 23607 8723 23613
rect 8754 23604 8760 23656
rect 8812 23653 8818 23656
rect 8812 23647 8840 23653
rect 8828 23613 8840 23647
rect 8812 23607 8840 23613
rect 8941 23647 8999 23653
rect 8941 23613 8953 23647
rect 8987 23644 8999 23647
rect 9122 23644 9128 23656
rect 8987 23616 9128 23644
rect 8987 23613 8999 23616
rect 8941 23607 8999 23613
rect 8812 23604 8818 23607
rect 9122 23604 9128 23616
rect 9180 23604 9186 23656
rect 9508 23644 9536 23820
rect 9858 23808 9864 23860
rect 9916 23808 9922 23860
rect 10962 23808 10968 23860
rect 11020 23848 11026 23860
rect 11606 23848 11612 23860
rect 11020 23820 11612 23848
rect 11020 23808 11026 23820
rect 11606 23808 11612 23820
rect 11664 23808 11670 23860
rect 11698 23808 11704 23860
rect 11756 23808 11762 23860
rect 11882 23808 11888 23860
rect 11940 23848 11946 23860
rect 12802 23848 12808 23860
rect 11940 23820 12808 23848
rect 11940 23808 11946 23820
rect 12802 23808 12808 23820
rect 12860 23808 12866 23860
rect 14737 23851 14795 23857
rect 12912 23820 14688 23848
rect 9876 23780 9904 23808
rect 11333 23783 11391 23789
rect 9876 23752 10548 23780
rect 10520 23721 10548 23752
rect 11333 23749 11345 23783
rect 11379 23780 11391 23783
rect 11716 23780 11744 23808
rect 12912 23792 12940 23820
rect 12710 23780 12716 23792
rect 11379 23752 11744 23780
rect 12544 23752 12716 23780
rect 11379 23749 11391 23752
rect 11333 23743 11391 23749
rect 9585 23715 9643 23721
rect 9585 23681 9597 23715
rect 9631 23712 9643 23715
rect 10413 23715 10471 23721
rect 10413 23712 10425 23715
rect 9631 23684 10425 23712
rect 9631 23681 9643 23684
rect 9585 23675 9643 23681
rect 10413 23681 10425 23684
rect 10459 23681 10471 23715
rect 10413 23675 10471 23681
rect 10505 23715 10563 23721
rect 10505 23681 10517 23715
rect 10551 23681 10563 23715
rect 10505 23675 10563 23681
rect 10597 23715 10655 23721
rect 10597 23681 10609 23715
rect 10643 23712 10655 23715
rect 10965 23715 11023 23721
rect 10965 23712 10977 23715
rect 10643 23684 10977 23712
rect 10643 23681 10655 23684
rect 10597 23675 10655 23681
rect 10965 23681 10977 23684
rect 11011 23681 11023 23715
rect 10965 23675 11023 23681
rect 11149 23715 11207 23721
rect 11149 23681 11161 23715
rect 11195 23712 11207 23715
rect 11238 23712 11244 23724
rect 11195 23684 11244 23712
rect 11195 23681 11207 23684
rect 11149 23675 11207 23681
rect 11238 23672 11244 23684
rect 11296 23672 11302 23724
rect 11698 23672 11704 23724
rect 11756 23712 11762 23724
rect 11974 23712 11980 23724
rect 11756 23684 11980 23712
rect 11756 23672 11762 23684
rect 11974 23672 11980 23684
rect 12032 23672 12038 23724
rect 12544 23644 12572 23752
rect 12710 23740 12716 23752
rect 12768 23740 12774 23792
rect 12894 23740 12900 23792
rect 12952 23740 12958 23792
rect 14660 23780 14688 23820
rect 14737 23817 14749 23851
rect 14783 23848 14795 23851
rect 14918 23848 14924 23860
rect 14783 23820 14924 23848
rect 14783 23817 14795 23820
rect 14737 23811 14795 23817
rect 14918 23808 14924 23820
rect 14976 23808 14982 23860
rect 19337 23851 19395 23857
rect 19337 23817 19349 23851
rect 19383 23848 19395 23851
rect 19383 23820 20576 23848
rect 19383 23817 19395 23820
rect 19337 23811 19395 23817
rect 15194 23780 15200 23792
rect 14660 23752 15200 23780
rect 15194 23740 15200 23752
rect 15252 23740 15258 23792
rect 19153 23783 19211 23789
rect 19153 23749 19165 23783
rect 19199 23780 19211 23783
rect 20548 23780 20576 23820
rect 20622 23808 20628 23860
rect 20680 23808 20686 23860
rect 19199 23752 20300 23780
rect 20548 23752 21404 23780
rect 19199 23749 19211 23752
rect 19153 23743 19211 23749
rect 12618 23672 12624 23724
rect 12676 23712 12682 23724
rect 12676 23684 13318 23712
rect 12676 23672 12682 23684
rect 9508 23616 12572 23644
rect 12894 23604 12900 23656
rect 12952 23604 12958 23656
rect 13081 23647 13139 23653
rect 13081 23613 13093 23647
rect 13127 23613 13139 23647
rect 13081 23607 13139 23613
rect 6825 23539 6883 23545
rect 6930 23548 8524 23576
rect 716 23480 2084 23508
rect 716 23468 722 23480
rect 2314 23468 2320 23520
rect 2372 23508 2378 23520
rect 2409 23511 2467 23517
rect 2409 23508 2421 23511
rect 2372 23480 2421 23508
rect 2372 23468 2378 23480
rect 2409 23477 2421 23480
rect 2455 23477 2467 23511
rect 2409 23471 2467 23477
rect 5902 23468 5908 23520
rect 5960 23508 5966 23520
rect 6454 23508 6460 23520
rect 5960 23480 6460 23508
rect 5960 23468 5966 23480
rect 6454 23468 6460 23480
rect 6512 23468 6518 23520
rect 6546 23468 6552 23520
rect 6604 23508 6610 23520
rect 6930 23508 6958 23548
rect 9582 23536 9588 23588
rect 9640 23576 9646 23588
rect 10502 23576 10508 23588
rect 9640 23548 10508 23576
rect 9640 23536 9646 23548
rect 10502 23536 10508 23548
rect 10560 23536 10566 23588
rect 10962 23536 10968 23588
rect 11020 23576 11026 23588
rect 11020 23548 11558 23576
rect 11020 23536 11026 23548
rect 6604 23480 6958 23508
rect 6604 23468 6610 23480
rect 7466 23468 7472 23520
rect 7524 23468 7530 23520
rect 7650 23468 7656 23520
rect 7708 23508 7714 23520
rect 8754 23508 8760 23520
rect 7708 23480 8760 23508
rect 7708 23468 7714 23480
rect 8754 23468 8760 23480
rect 8812 23468 8818 23520
rect 10229 23511 10287 23517
rect 10229 23477 10241 23511
rect 10275 23508 10287 23511
rect 11146 23508 11152 23520
rect 10275 23480 11152 23508
rect 10275 23477 10287 23480
rect 10229 23471 10287 23477
rect 11146 23468 11152 23480
rect 11204 23468 11210 23520
rect 11241 23511 11299 23517
rect 11241 23477 11253 23511
rect 11287 23508 11299 23511
rect 11422 23508 11428 23520
rect 11287 23480 11428 23508
rect 11287 23477 11299 23480
rect 11241 23471 11299 23477
rect 11422 23468 11428 23480
rect 11480 23468 11486 23520
rect 11530 23508 11558 23548
rect 11606 23536 11612 23588
rect 11664 23576 11670 23588
rect 11974 23576 11980 23588
rect 11664 23548 11980 23576
rect 11664 23536 11670 23548
rect 11974 23536 11980 23548
rect 12032 23536 12038 23588
rect 12710 23536 12716 23588
rect 12768 23576 12774 23588
rect 13096 23576 13124 23607
rect 12768 23548 13124 23576
rect 12768 23536 12774 23548
rect 13078 23508 13084 23520
rect 11530 23480 13084 23508
rect 13078 23468 13084 23480
rect 13136 23468 13142 23520
rect 13290 23508 13318 23684
rect 13814 23672 13820 23724
rect 13872 23672 13878 23724
rect 15071 23715 15129 23721
rect 15071 23712 15083 23715
rect 14752 23684 15083 23712
rect 13446 23604 13452 23656
rect 13504 23644 13510 23656
rect 13541 23647 13599 23653
rect 13541 23644 13553 23647
rect 13504 23616 13553 23644
rect 13504 23604 13510 23616
rect 13541 23613 13553 23616
rect 13587 23613 13599 23647
rect 13541 23607 13599 23613
rect 13906 23604 13912 23656
rect 13964 23653 13970 23656
rect 13964 23647 13992 23653
rect 13980 23613 13992 23647
rect 13964 23607 13992 23613
rect 14093 23647 14151 23653
rect 14093 23613 14105 23647
rect 14139 23644 14151 23647
rect 14274 23644 14280 23656
rect 14139 23616 14280 23644
rect 14139 23613 14151 23616
rect 14093 23607 14151 23613
rect 13964 23604 13970 23607
rect 14274 23604 14280 23616
rect 14332 23604 14338 23656
rect 14752 23576 14780 23684
rect 15071 23681 15083 23684
rect 15117 23712 15129 23715
rect 16911 23715 16969 23721
rect 16911 23712 16923 23715
rect 15117 23684 16923 23712
rect 15117 23681 15129 23684
rect 15071 23675 15129 23681
rect 16911 23681 16923 23684
rect 16957 23712 16969 23715
rect 17310 23712 17316 23724
rect 16957 23684 17316 23712
rect 16957 23681 16969 23684
rect 16911 23675 16969 23681
rect 17310 23672 17316 23684
rect 17368 23672 17374 23724
rect 19061 23715 19119 23721
rect 19061 23681 19073 23715
rect 19107 23681 19119 23715
rect 19061 23675 19119 23681
rect 14826 23604 14832 23656
rect 14884 23604 14890 23656
rect 15838 23604 15844 23656
rect 15896 23644 15902 23656
rect 16114 23644 16120 23656
rect 15896 23616 16120 23644
rect 15896 23604 15902 23616
rect 16114 23604 16120 23616
rect 16172 23644 16178 23656
rect 16669 23647 16727 23653
rect 16669 23644 16681 23647
rect 16172 23616 16681 23644
rect 16172 23604 16178 23616
rect 16669 23613 16681 23616
rect 16715 23613 16727 23647
rect 16669 23607 16727 23613
rect 14476 23548 14780 23576
rect 19076 23576 19104 23675
rect 19242 23672 19248 23724
rect 19300 23672 19306 23724
rect 19334 23672 19340 23724
rect 19392 23712 19398 23724
rect 19521 23715 19579 23721
rect 19521 23712 19533 23715
rect 19392 23684 19533 23712
rect 19392 23672 19398 23684
rect 19521 23681 19533 23684
rect 19567 23681 19579 23715
rect 19886 23712 19892 23724
rect 19847 23684 19892 23712
rect 19521 23675 19579 23681
rect 19886 23672 19892 23684
rect 19944 23672 19950 23724
rect 19613 23647 19671 23653
rect 19613 23613 19625 23647
rect 19659 23613 19671 23647
rect 20272 23644 20300 23752
rect 20530 23672 20536 23724
rect 20588 23712 20594 23724
rect 21376 23721 21404 23752
rect 20993 23715 21051 23721
rect 20993 23712 21005 23715
rect 20588 23684 21005 23712
rect 20588 23672 20594 23684
rect 20993 23681 21005 23684
rect 21039 23681 21051 23715
rect 20993 23675 21051 23681
rect 21361 23715 21419 23721
rect 21361 23681 21373 23715
rect 21407 23681 21419 23715
rect 21361 23675 21419 23681
rect 21269 23647 21327 23653
rect 21269 23644 21281 23647
rect 20272 23616 21281 23644
rect 19613 23607 19671 23613
rect 21269 23613 21281 23616
rect 21315 23613 21327 23647
rect 21269 23607 21327 23613
rect 19518 23576 19524 23588
rect 19076 23548 19524 23576
rect 14476 23508 14504 23548
rect 19518 23536 19524 23548
rect 19576 23536 19582 23588
rect 19628 23520 19656 23607
rect 21085 23579 21143 23585
rect 21085 23545 21097 23579
rect 21131 23576 21143 23579
rect 21453 23579 21511 23585
rect 21453 23576 21465 23579
rect 21131 23548 21465 23576
rect 21131 23545 21143 23548
rect 21085 23539 21143 23545
rect 21453 23545 21465 23548
rect 21499 23545 21511 23579
rect 21453 23539 21511 23545
rect 13290 23480 14504 23508
rect 14550 23468 14556 23520
rect 14608 23508 14614 23520
rect 15841 23511 15899 23517
rect 15841 23508 15853 23511
rect 14608 23480 15853 23508
rect 14608 23468 14614 23480
rect 15841 23477 15853 23480
rect 15887 23477 15899 23511
rect 15841 23471 15899 23477
rect 17678 23468 17684 23520
rect 17736 23468 17742 23520
rect 18966 23468 18972 23520
rect 19024 23508 19030 23520
rect 19610 23508 19616 23520
rect 19024 23480 19616 23508
rect 19024 23468 19030 23480
rect 19610 23468 19616 23480
rect 19668 23468 19674 23520
rect 20714 23468 20720 23520
rect 20772 23508 20778 23520
rect 21177 23511 21235 23517
rect 21177 23508 21189 23511
rect 20772 23480 21189 23508
rect 20772 23468 20778 23480
rect 21177 23477 21189 23480
rect 21223 23477 21235 23511
rect 21177 23471 21235 23477
rect 1104 23418 21896 23440
rect 1104 23366 3549 23418
rect 3601 23366 3613 23418
rect 3665 23366 3677 23418
rect 3729 23366 3741 23418
rect 3793 23366 3805 23418
rect 3857 23366 8747 23418
rect 8799 23366 8811 23418
rect 8863 23366 8875 23418
rect 8927 23366 8939 23418
rect 8991 23366 9003 23418
rect 9055 23366 13945 23418
rect 13997 23366 14009 23418
rect 14061 23366 14073 23418
rect 14125 23366 14137 23418
rect 14189 23366 14201 23418
rect 14253 23366 19143 23418
rect 19195 23366 19207 23418
rect 19259 23366 19271 23418
rect 19323 23366 19335 23418
rect 19387 23366 19399 23418
rect 19451 23366 21896 23418
rect 1104 23344 21896 23366
rect 1118 23264 1124 23316
rect 1176 23304 1182 23316
rect 1176 23276 3372 23304
rect 1176 23264 1182 23276
rect 3234 23196 3240 23248
rect 3292 23196 3298 23248
rect 1486 23128 1492 23180
rect 1544 23168 1550 23180
rect 1673 23171 1731 23177
rect 1673 23168 1685 23171
rect 1544 23140 1685 23168
rect 1544 23128 1550 23140
rect 1673 23137 1685 23140
rect 1719 23137 1731 23171
rect 1673 23131 1731 23137
rect 1394 23060 1400 23112
rect 1452 23060 1458 23112
rect 1854 23060 1860 23112
rect 1912 23100 1918 23112
rect 1947 23103 2005 23109
rect 1947 23100 1959 23103
rect 1912 23072 1959 23100
rect 1912 23060 1918 23072
rect 1947 23069 1959 23072
rect 1993 23100 2005 23103
rect 2682 23100 2688 23112
rect 1993 23072 2688 23100
rect 1993 23069 2005 23072
rect 1947 23063 2005 23069
rect 2682 23060 2688 23072
rect 2740 23060 2746 23112
rect 3344 23109 3372 23276
rect 3418 23264 3424 23316
rect 3476 23304 3482 23316
rect 3513 23307 3571 23313
rect 3513 23304 3525 23307
rect 3476 23276 3525 23304
rect 3476 23264 3482 23276
rect 3513 23273 3525 23276
rect 3559 23273 3571 23307
rect 3513 23267 3571 23273
rect 4798 23264 4804 23316
rect 4856 23304 4862 23316
rect 5718 23304 5724 23316
rect 4856 23276 5724 23304
rect 4856 23264 4862 23276
rect 5718 23264 5724 23276
rect 5776 23264 5782 23316
rect 5810 23264 5816 23316
rect 5868 23304 5874 23316
rect 6270 23304 6276 23316
rect 5868 23276 6276 23304
rect 5868 23264 5874 23276
rect 6270 23264 6276 23276
rect 6328 23264 6334 23316
rect 7742 23304 7748 23316
rect 7484 23276 7748 23304
rect 5626 23196 5632 23248
rect 5684 23236 5690 23248
rect 5905 23239 5963 23245
rect 5905 23236 5917 23239
rect 5684 23208 5917 23236
rect 5684 23196 5690 23208
rect 5905 23205 5917 23208
rect 5951 23205 5963 23239
rect 5905 23199 5963 23205
rect 6181 23171 6239 23177
rect 6181 23168 6193 23171
rect 5368 23140 6193 23168
rect 5368 23112 5396 23140
rect 6181 23137 6193 23140
rect 6227 23137 6239 23171
rect 6181 23131 6239 23137
rect 6270 23128 6276 23180
rect 6328 23177 6334 23180
rect 6328 23171 6356 23177
rect 6344 23137 6356 23171
rect 6328 23131 6356 23137
rect 6328 23128 6334 23131
rect 6454 23128 6460 23180
rect 6512 23128 6518 23180
rect 6822 23128 6828 23180
rect 6880 23168 6886 23180
rect 7484 23177 7512 23276
rect 7742 23264 7748 23276
rect 7800 23264 7806 23316
rect 7926 23264 7932 23316
rect 7984 23304 7990 23316
rect 8481 23307 8539 23313
rect 7984 23276 8432 23304
rect 7984 23264 7990 23276
rect 8404 23236 8432 23276
rect 8481 23273 8493 23307
rect 8527 23304 8539 23307
rect 9122 23304 9128 23316
rect 8527 23276 9128 23304
rect 8527 23273 8539 23276
rect 8481 23267 8539 23273
rect 9122 23264 9128 23276
rect 9180 23264 9186 23316
rect 9232 23276 10640 23304
rect 9232 23236 9260 23276
rect 8404 23208 9260 23236
rect 7469 23171 7527 23177
rect 7469 23168 7481 23171
rect 6880 23140 7481 23168
rect 6880 23128 6886 23140
rect 7469 23137 7481 23140
rect 7515 23137 7527 23171
rect 7469 23131 7527 23137
rect 3053 23103 3111 23109
rect 3053 23069 3065 23103
rect 3099 23069 3111 23103
rect 3053 23063 3111 23069
rect 3329 23103 3387 23109
rect 3329 23069 3341 23103
rect 3375 23069 3387 23103
rect 3329 23063 3387 23069
rect 1302 22992 1308 23044
rect 1360 23032 1366 23044
rect 3068 23032 3096 23063
rect 3418 23060 3424 23112
rect 3476 23100 3482 23112
rect 3786 23100 3792 23112
rect 3476 23072 3792 23100
rect 3476 23060 3482 23072
rect 3786 23060 3792 23072
rect 3844 23060 3850 23112
rect 3970 23060 3976 23112
rect 4028 23100 4034 23112
rect 4063 23103 4121 23109
rect 4063 23100 4075 23103
rect 4028 23072 4075 23100
rect 4028 23060 4034 23072
rect 4063 23069 4075 23072
rect 4109 23069 4121 23103
rect 4063 23063 4121 23069
rect 4706 23060 4712 23112
rect 4764 23100 4770 23112
rect 5258 23100 5264 23112
rect 4764 23072 5264 23100
rect 4764 23060 4770 23072
rect 5258 23060 5264 23072
rect 5316 23060 5322 23112
rect 5350 23060 5356 23112
rect 5408 23060 5414 23112
rect 5445 23103 5503 23109
rect 5445 23069 5457 23103
rect 5491 23069 5503 23103
rect 5445 23063 5503 23069
rect 7101 23103 7159 23109
rect 7101 23069 7113 23103
rect 7147 23100 7159 23103
rect 7377 23103 7435 23109
rect 7377 23100 7389 23103
rect 7147 23072 7389 23100
rect 7147 23069 7159 23072
rect 7101 23063 7159 23069
rect 7377 23069 7389 23072
rect 7423 23069 7435 23103
rect 7742 23100 7748 23112
rect 7703 23072 7748 23100
rect 7377 23063 7435 23069
rect 1360 23004 3096 23032
rect 1360 22992 1366 23004
rect 4614 22992 4620 23044
rect 4672 23032 4678 23044
rect 4982 23032 4988 23044
rect 4672 23004 4988 23032
rect 4672 22992 4678 23004
rect 4982 22992 4988 23004
rect 5040 23032 5046 23044
rect 5460 23032 5488 23063
rect 7742 23060 7748 23072
rect 7800 23060 7806 23112
rect 9674 23100 9680 23112
rect 8266 23072 9680 23100
rect 8266 23032 8294 23072
rect 9674 23060 9680 23072
rect 9732 23060 9738 23112
rect 9919 23103 9977 23109
rect 9919 23069 9931 23103
rect 9965 23100 9977 23103
rect 10042 23100 10048 23112
rect 9965 23072 10048 23100
rect 9965 23069 9977 23072
rect 9919 23063 9977 23069
rect 10042 23060 10048 23072
rect 10100 23060 10106 23112
rect 5040 23004 5488 23032
rect 6930 23004 8294 23032
rect 5040 22992 5046 23004
rect 1578 22924 1584 22976
rect 1636 22924 1642 22976
rect 2498 22924 2504 22976
rect 2556 22964 2562 22976
rect 2685 22967 2743 22973
rect 2685 22964 2697 22967
rect 2556 22936 2697 22964
rect 2556 22924 2562 22936
rect 2685 22933 2697 22936
rect 2731 22933 2743 22967
rect 2685 22927 2743 22933
rect 4062 22924 4068 22976
rect 4120 22964 4126 22976
rect 4338 22964 4344 22976
rect 4120 22936 4344 22964
rect 4120 22924 4126 22936
rect 4338 22924 4344 22936
rect 4396 22924 4402 22976
rect 4798 22924 4804 22976
rect 4856 22924 4862 22976
rect 5442 22924 5448 22976
rect 5500 22964 5506 22976
rect 6546 22964 6552 22976
rect 5500 22936 6552 22964
rect 5500 22924 5506 22936
rect 6546 22924 6552 22936
rect 6604 22964 6610 22976
rect 6930 22964 6958 23004
rect 9766 22992 9772 23044
rect 9824 23032 9830 23044
rect 10318 23032 10324 23044
rect 9824 23004 10324 23032
rect 9824 22992 9830 23004
rect 10318 22992 10324 23004
rect 10376 22992 10382 23044
rect 10612 23032 10640 23276
rect 10686 23264 10692 23316
rect 10744 23304 10750 23316
rect 11514 23304 11520 23316
rect 10744 23276 11520 23304
rect 10744 23264 10750 23276
rect 11072 23177 11100 23276
rect 11514 23264 11520 23276
rect 11572 23264 11578 23316
rect 12158 23304 12164 23316
rect 11714 23276 12164 23304
rect 11057 23171 11115 23177
rect 11057 23137 11069 23171
rect 11103 23137 11115 23171
rect 11057 23131 11115 23137
rect 11238 23060 11244 23112
rect 11296 23100 11302 23112
rect 11331 23103 11389 23109
rect 11331 23100 11343 23103
rect 11296 23072 11343 23100
rect 11296 23060 11302 23072
rect 11331 23069 11343 23072
rect 11377 23100 11389 23103
rect 11714 23100 11742 23276
rect 12158 23264 12164 23276
rect 12216 23264 12222 23316
rect 12268 23276 13860 23304
rect 12268 23236 12296 23276
rect 13832 23248 13860 23276
rect 14274 23264 14280 23316
rect 14332 23304 14338 23316
rect 14550 23304 14556 23316
rect 14332 23276 14556 23304
rect 14332 23264 14338 23276
rect 14550 23264 14556 23276
rect 14608 23264 14614 23316
rect 14645 23307 14703 23313
rect 14645 23273 14657 23307
rect 14691 23304 14703 23307
rect 14734 23304 14740 23316
rect 14691 23276 14740 23304
rect 14691 23273 14703 23276
rect 14645 23267 14703 23273
rect 14734 23264 14740 23276
rect 14792 23264 14798 23316
rect 16390 23304 16396 23316
rect 14844 23276 16396 23304
rect 11377 23072 11742 23100
rect 11790 23208 12296 23236
rect 11377 23069 11389 23072
rect 11331 23063 11389 23069
rect 11790 23032 11818 23208
rect 13814 23196 13820 23248
rect 13872 23236 13878 23248
rect 14844 23236 14872 23276
rect 16390 23264 16396 23276
rect 16448 23264 16454 23316
rect 19518 23304 19524 23316
rect 17236 23276 19524 23304
rect 13872 23208 14872 23236
rect 13872 23196 13878 23208
rect 16022 23196 16028 23248
rect 16080 23196 16086 23248
rect 17236 23245 17264 23276
rect 19518 23264 19524 23276
rect 19576 23264 19582 23316
rect 19610 23264 19616 23316
rect 19668 23264 19674 23316
rect 19886 23264 19892 23316
rect 19944 23304 19950 23316
rect 20530 23304 20536 23316
rect 19944 23276 20536 23304
rect 19944 23264 19950 23276
rect 20530 23264 20536 23276
rect 20588 23264 20594 23316
rect 21453 23307 21511 23313
rect 21453 23273 21465 23307
rect 21499 23304 21511 23307
rect 21542 23304 21548 23316
rect 21499 23276 21548 23304
rect 21499 23273 21511 23276
rect 21453 23267 21511 23273
rect 21542 23264 21548 23276
rect 21600 23264 21606 23316
rect 17221 23239 17279 23245
rect 17221 23205 17233 23239
rect 17267 23205 17279 23239
rect 17221 23199 17279 23205
rect 17954 23196 17960 23248
rect 18012 23236 18018 23248
rect 18506 23236 18512 23248
rect 18012 23208 18512 23236
rect 18012 23196 18018 23208
rect 18506 23196 18512 23208
rect 18564 23196 18570 23248
rect 19245 23239 19303 23245
rect 19245 23205 19257 23239
rect 19291 23205 19303 23239
rect 19628 23236 19656 23264
rect 19245 23199 19303 23205
rect 19536 23208 19656 23236
rect 12158 23128 12164 23180
rect 12216 23168 12222 23180
rect 12342 23168 12348 23180
rect 12216 23140 12348 23168
rect 12216 23128 12222 23140
rect 12342 23128 12348 23140
rect 12400 23128 12406 23180
rect 12437 23171 12495 23177
rect 12437 23137 12449 23171
rect 12483 23137 12495 23171
rect 12437 23131 12495 23137
rect 12452 23100 12480 23131
rect 15194 23128 15200 23180
rect 15252 23168 15258 23180
rect 15565 23171 15623 23177
rect 15565 23168 15577 23171
rect 15252 23140 15577 23168
rect 15252 23128 15258 23140
rect 15565 23137 15577 23140
rect 15611 23137 15623 23171
rect 15565 23131 15623 23137
rect 15746 23128 15752 23180
rect 15804 23168 15810 23180
rect 16301 23171 16359 23177
rect 16301 23168 16313 23171
rect 15804 23140 16313 23168
rect 15804 23128 15810 23140
rect 16301 23137 16313 23140
rect 16347 23137 16359 23171
rect 16301 23131 16359 23137
rect 16577 23171 16635 23177
rect 16577 23137 16589 23171
rect 16623 23168 16635 23171
rect 17678 23168 17684 23180
rect 16623 23140 17684 23168
rect 16623 23137 16635 23140
rect 16577 23131 16635 23137
rect 17678 23128 17684 23140
rect 17736 23128 17742 23180
rect 18414 23168 18420 23180
rect 17788 23140 18420 23168
rect 12452 23072 12572 23100
rect 12544 23032 12572 23072
rect 12618 23060 12624 23112
rect 12676 23100 12682 23112
rect 12711 23103 12769 23109
rect 12711 23100 12723 23103
rect 12676 23072 12723 23100
rect 12676 23060 12682 23072
rect 12711 23069 12723 23072
rect 12757 23069 12769 23103
rect 12711 23063 12769 23069
rect 12802 23060 12808 23112
rect 12860 23100 12866 23112
rect 12860 23072 14688 23100
rect 12860 23060 12866 23072
rect 14550 23032 14556 23044
rect 10612 23004 11818 23032
rect 11882 23004 14556 23032
rect 6604 22936 6958 22964
rect 7193 22967 7251 22973
rect 6604 22924 6610 22936
rect 7193 22933 7205 22967
rect 7239 22964 7251 22967
rect 8018 22964 8024 22976
rect 7239 22936 8024 22964
rect 7239 22933 7251 22936
rect 7193 22927 7251 22933
rect 8018 22924 8024 22936
rect 8076 22924 8082 22976
rect 8202 22924 8208 22976
rect 8260 22964 8266 22976
rect 9858 22964 9864 22976
rect 8260 22936 9864 22964
rect 8260 22924 8266 22936
rect 9858 22924 9864 22936
rect 9916 22924 9922 22976
rect 10686 22924 10692 22976
rect 10744 22924 10750 22976
rect 11514 22924 11520 22976
rect 11572 22964 11578 22976
rect 11882 22964 11910 23004
rect 14550 22992 14556 23004
rect 14608 22992 14614 23044
rect 11572 22936 11910 22964
rect 12069 22967 12127 22973
rect 11572 22924 11578 22936
rect 12069 22933 12081 22967
rect 12115 22964 12127 22967
rect 12618 22964 12624 22976
rect 12115 22936 12624 22964
rect 12115 22933 12127 22936
rect 12069 22927 12127 22933
rect 12618 22924 12624 22936
rect 12676 22924 12682 22976
rect 13262 22924 13268 22976
rect 13320 22964 13326 22976
rect 13449 22967 13507 22973
rect 13449 22964 13461 22967
rect 13320 22936 13461 22964
rect 13320 22924 13326 22936
rect 13449 22933 13461 22936
rect 13495 22933 13507 22967
rect 14660 22964 14688 23072
rect 14826 23060 14832 23112
rect 14884 23060 14890 23112
rect 15286 23060 15292 23112
rect 15344 23100 15350 23112
rect 15381 23103 15439 23109
rect 15381 23100 15393 23103
rect 15344 23072 15393 23100
rect 15344 23060 15350 23072
rect 15381 23069 15393 23072
rect 15427 23069 15439 23103
rect 15381 23063 15439 23069
rect 16390 23060 16396 23112
rect 16448 23109 16454 23112
rect 16448 23103 16476 23109
rect 16464 23069 16476 23103
rect 16448 23063 16476 23069
rect 16448 23060 16454 23063
rect 17494 22992 17500 23044
rect 17552 23032 17558 23044
rect 17678 23032 17684 23044
rect 17552 23004 17684 23032
rect 17552 22992 17558 23004
rect 17678 22992 17684 23004
rect 17736 22992 17742 23044
rect 17788 22964 17816 23140
rect 18414 23128 18420 23140
rect 18472 23128 18478 23180
rect 18509 23103 18567 23109
rect 18509 23100 18521 23103
rect 18156 23072 18521 23100
rect 18156 22976 18184 23072
rect 18509 23069 18521 23072
rect 18555 23069 18567 23103
rect 18509 23063 18567 23069
rect 18877 23103 18935 23109
rect 18877 23069 18889 23103
rect 18923 23069 18935 23103
rect 18877 23063 18935 23069
rect 19061 23103 19119 23109
rect 19061 23069 19073 23103
rect 19107 23100 19119 23103
rect 19260 23100 19288 23199
rect 19536 23177 19564 23208
rect 20438 23196 20444 23248
rect 20496 23236 20502 23248
rect 21174 23236 21180 23248
rect 20496 23208 21180 23236
rect 20496 23196 20502 23208
rect 21174 23196 21180 23208
rect 21232 23196 21238 23248
rect 19521 23171 19579 23177
rect 19521 23137 19533 23171
rect 19567 23137 19579 23171
rect 19521 23131 19579 23137
rect 19334 23100 19340 23112
rect 19107 23072 19288 23100
rect 19107 23069 19119 23072
rect 19061 23063 19119 23069
rect 18892 23032 18920 23063
rect 19321 23060 19340 23100
rect 19392 23060 19398 23112
rect 19886 23100 19892 23112
rect 19429 23079 19487 23085
rect 19794 23079 19892 23100
rect 19321 23032 19349 23060
rect 19429 23045 19441 23079
rect 19475 23045 19487 23079
rect 19429 23039 19487 23045
rect 19779 23073 19892 23079
rect 19779 23039 19791 23073
rect 19825 23072 19892 23073
rect 19825 23039 19837 23072
rect 19886 23060 19892 23072
rect 19944 23060 19950 23112
rect 20990 23060 20996 23112
rect 21048 23100 21054 23112
rect 21177 23103 21235 23109
rect 21177 23100 21189 23103
rect 21048 23072 21189 23100
rect 21048 23060 21054 23072
rect 21177 23069 21189 23072
rect 21223 23069 21235 23103
rect 21177 23063 21235 23069
rect 18892 23004 19349 23032
rect 19444 22976 19472 23039
rect 19779 23033 19837 23039
rect 14660 22936 17816 22964
rect 13449 22927 13507 22933
rect 18138 22924 18144 22976
rect 18196 22924 18202 22976
rect 18322 22924 18328 22976
rect 18380 22924 18386 22976
rect 19058 22924 19064 22976
rect 19116 22924 19122 22976
rect 19150 22924 19156 22976
rect 19208 22964 19214 22976
rect 19288 22964 19294 22976
rect 19208 22936 19294 22964
rect 19208 22924 19214 22936
rect 19288 22924 19294 22936
rect 19346 22924 19352 22976
rect 19426 22924 19432 22976
rect 19484 22924 19490 22976
rect 1104 22874 22056 22896
rect 1104 22822 6148 22874
rect 6200 22822 6212 22874
rect 6264 22822 6276 22874
rect 6328 22822 6340 22874
rect 6392 22822 6404 22874
rect 6456 22822 11346 22874
rect 11398 22822 11410 22874
rect 11462 22822 11474 22874
rect 11526 22822 11538 22874
rect 11590 22822 11602 22874
rect 11654 22822 16544 22874
rect 16596 22822 16608 22874
rect 16660 22822 16672 22874
rect 16724 22822 16736 22874
rect 16788 22822 16800 22874
rect 16852 22822 21742 22874
rect 21794 22822 21806 22874
rect 21858 22822 21870 22874
rect 21922 22822 21934 22874
rect 21986 22822 21998 22874
rect 22050 22822 22056 22874
rect 1104 22800 22056 22822
rect 1670 22720 1676 22772
rect 1728 22720 1734 22772
rect 2866 22720 2872 22772
rect 2924 22760 2930 22772
rect 2961 22763 3019 22769
rect 2961 22760 2973 22763
rect 2924 22732 2973 22760
rect 2924 22720 2930 22732
rect 2961 22729 2973 22732
rect 3007 22729 3019 22763
rect 2961 22723 3019 22729
rect 3050 22720 3056 22772
rect 3108 22760 3114 22772
rect 3329 22763 3387 22769
rect 3329 22760 3341 22763
rect 3108 22732 3341 22760
rect 3108 22720 3114 22732
rect 3329 22729 3341 22732
rect 3375 22729 3387 22763
rect 4798 22760 4804 22772
rect 3329 22723 3387 22729
rect 3712 22732 4804 22760
rect 2041 22695 2099 22701
rect 2041 22661 2053 22695
rect 2087 22692 2099 22695
rect 2498 22692 2504 22704
rect 2087 22664 2504 22692
rect 2087 22661 2099 22664
rect 2041 22655 2099 22661
rect 2498 22652 2504 22664
rect 2556 22652 2562 22704
rect 2774 22652 2780 22704
rect 2832 22652 2838 22704
rect 3510 22692 3516 22704
rect 2976 22664 3516 22692
rect 1946 22584 1952 22636
rect 2004 22584 2010 22636
rect 2406 22584 2412 22636
rect 2464 22584 2470 22636
rect 2976 22568 3004 22664
rect 3510 22652 3516 22664
rect 3568 22652 3574 22704
rect 3602 22652 3608 22704
rect 3660 22652 3666 22704
rect 3712 22701 3740 22732
rect 4798 22720 4804 22732
rect 4856 22720 4862 22772
rect 5902 22720 5908 22772
rect 5960 22760 5966 22772
rect 7374 22760 7380 22772
rect 5960 22732 7380 22760
rect 5960 22720 5966 22732
rect 7374 22720 7380 22732
rect 7432 22720 7438 22772
rect 7926 22720 7932 22772
rect 7984 22760 7990 22772
rect 9861 22763 9919 22769
rect 9861 22760 9873 22763
rect 7984 22732 9873 22760
rect 7984 22720 7990 22732
rect 9861 22729 9873 22732
rect 9907 22729 9919 22763
rect 10318 22760 10324 22772
rect 9861 22723 9919 22729
rect 9968 22732 10324 22760
rect 3697 22695 3755 22701
rect 3697 22661 3709 22695
rect 3743 22661 3755 22695
rect 3697 22655 3755 22661
rect 4065 22695 4123 22701
rect 4065 22661 4077 22695
rect 4111 22692 4123 22695
rect 4338 22692 4344 22704
rect 4111 22664 4344 22692
rect 4111 22661 4123 22664
rect 4065 22655 4123 22661
rect 4338 22652 4344 22664
rect 4396 22652 4402 22704
rect 4430 22652 4436 22704
rect 4488 22652 4494 22704
rect 9968 22692 9996 22732
rect 10318 22720 10324 22732
rect 10376 22720 10382 22772
rect 10502 22720 10508 22772
rect 10560 22760 10566 22772
rect 12802 22760 12808 22772
rect 10560 22732 12808 22760
rect 10560 22720 10566 22732
rect 12802 22720 12808 22732
rect 12860 22720 12866 22772
rect 14737 22763 14795 22769
rect 12912 22732 14596 22760
rect 7392 22664 9996 22692
rect 3418 22584 3424 22636
rect 3476 22624 3482 22636
rect 6822 22624 6828 22636
rect 3476 22596 6828 22624
rect 3476 22584 3482 22596
rect 6822 22584 6828 22596
rect 6880 22584 6886 22636
rect 7099 22627 7157 22633
rect 7099 22593 7111 22627
rect 7145 22624 7157 22627
rect 7392 22624 7420 22664
rect 10042 22652 10048 22704
rect 10100 22652 10106 22704
rect 10229 22695 10287 22701
rect 10229 22661 10241 22695
rect 10275 22692 10287 22695
rect 10686 22692 10692 22704
rect 10275 22664 10692 22692
rect 10275 22661 10287 22664
rect 10229 22655 10287 22661
rect 10686 22652 10692 22664
rect 10744 22652 10750 22704
rect 10870 22652 10876 22704
rect 10928 22652 10934 22704
rect 10962 22652 10968 22704
rect 11020 22652 11026 22704
rect 11790 22652 11796 22704
rect 11848 22692 11854 22704
rect 12342 22692 12348 22704
rect 11848 22664 12348 22692
rect 11848 22652 11854 22664
rect 12342 22652 12348 22664
rect 12400 22652 12406 22704
rect 7145 22596 7420 22624
rect 7145 22593 7157 22596
rect 7099 22587 7157 22593
rect 7466 22584 7472 22636
rect 7524 22624 7530 22636
rect 8573 22627 8631 22633
rect 8573 22624 8585 22627
rect 7524 22596 8585 22624
rect 7524 22584 7530 22596
rect 8573 22593 8585 22596
rect 8619 22593 8631 22627
rect 8573 22587 8631 22593
rect 8662 22584 8668 22636
rect 8720 22624 8726 22636
rect 9033 22627 9091 22633
rect 9033 22624 9045 22627
rect 8720 22596 9045 22624
rect 8720 22584 8726 22596
rect 9033 22593 9045 22596
rect 9079 22593 9091 22627
rect 9033 22587 9091 22593
rect 9490 22584 9496 22636
rect 9548 22624 9554 22636
rect 10060 22624 10088 22652
rect 10137 22627 10195 22633
rect 10137 22624 10149 22627
rect 9548 22596 10149 22624
rect 9548 22584 9554 22596
rect 10137 22593 10149 22596
rect 10183 22593 10195 22627
rect 10137 22587 10195 22593
rect 10318 22584 10324 22636
rect 10376 22624 10382 22636
rect 10502 22624 10508 22636
rect 10376 22596 10508 22624
rect 10376 22584 10382 22596
rect 10502 22584 10508 22596
rect 10560 22584 10566 22636
rect 10597 22627 10655 22633
rect 10597 22593 10609 22627
rect 10643 22624 10655 22627
rect 10888 22624 10916 22652
rect 10643 22596 10916 22624
rect 10643 22593 10655 22596
rect 10597 22587 10655 22593
rect 11238 22584 11244 22636
rect 11296 22624 11302 22636
rect 11296 22596 12204 22624
rect 11296 22584 11302 22596
rect 2314 22516 2320 22568
rect 2372 22516 2378 22568
rect 2958 22516 2964 22568
rect 3016 22516 3022 22568
rect 3878 22516 3884 22568
rect 3936 22516 3942 22568
rect 5074 22516 5080 22568
rect 5132 22516 5138 22568
rect 5442 22516 5448 22568
rect 5500 22556 5506 22568
rect 6546 22556 6552 22568
rect 5500 22528 6552 22556
rect 5500 22516 5506 22528
rect 6546 22516 6552 22528
rect 6604 22516 6610 22568
rect 8297 22559 8355 22565
rect 8297 22525 8309 22559
rect 8343 22525 8355 22559
rect 8297 22519 8355 22525
rect 4614 22448 4620 22500
rect 4672 22448 4678 22500
rect 5092 22420 5120 22516
rect 7837 22491 7895 22497
rect 7837 22457 7849 22491
rect 7883 22488 7895 22491
rect 7926 22488 7932 22500
rect 7883 22460 7932 22488
rect 7883 22457 7895 22460
rect 7837 22451 7895 22457
rect 7926 22448 7932 22460
rect 7984 22488 7990 22500
rect 8312 22488 8340 22519
rect 10042 22516 10048 22568
rect 10100 22516 10106 22568
rect 11146 22516 11152 22568
rect 11204 22556 11210 22568
rect 11204 22528 11284 22556
rect 11204 22516 11210 22528
rect 7984 22460 8340 22488
rect 7984 22448 7990 22460
rect 8478 22448 8484 22500
rect 8536 22488 8542 22500
rect 9033 22491 9091 22497
rect 9033 22488 9045 22491
rect 8536 22460 9045 22488
rect 8536 22448 8542 22460
rect 9033 22457 9045 22460
rect 9079 22457 9091 22491
rect 9033 22451 9091 22457
rect 7742 22420 7748 22432
rect 5092 22392 7748 22420
rect 7742 22380 7748 22392
rect 7800 22380 7806 22432
rect 9122 22380 9128 22432
rect 9180 22420 9186 22432
rect 9858 22420 9864 22432
rect 9180 22392 9864 22420
rect 9180 22380 9186 22392
rect 9858 22380 9864 22392
rect 9916 22380 9922 22432
rect 11146 22380 11152 22432
rect 11204 22380 11210 22432
rect 11256 22420 11284 22528
rect 12176 22488 12204 22596
rect 12802 22584 12808 22636
rect 12860 22624 12866 22636
rect 12912 22633 12940 22732
rect 14568 22692 14596 22732
rect 14737 22729 14749 22763
rect 14783 22760 14795 22763
rect 14826 22760 14832 22772
rect 14783 22732 14832 22760
rect 14783 22729 14795 22732
rect 14737 22723 14795 22729
rect 14826 22720 14832 22732
rect 14884 22720 14890 22772
rect 15746 22760 15752 22772
rect 14936 22732 15752 22760
rect 14936 22692 14964 22732
rect 15746 22720 15752 22732
rect 15804 22720 15810 22772
rect 16390 22720 16396 22772
rect 16448 22760 16454 22772
rect 18046 22760 18052 22772
rect 16448 22732 18052 22760
rect 16448 22720 16454 22732
rect 18046 22720 18052 22732
rect 18104 22720 18110 22772
rect 19058 22720 19064 22772
rect 19116 22720 19122 22772
rect 19245 22763 19303 22769
rect 19245 22729 19257 22763
rect 19291 22760 19303 22763
rect 19426 22760 19432 22772
rect 19291 22732 19432 22760
rect 19291 22729 19303 22732
rect 19245 22723 19303 22729
rect 19426 22720 19432 22732
rect 19484 22720 19490 22772
rect 20346 22720 20352 22772
rect 20404 22720 20410 22772
rect 21085 22763 21143 22769
rect 21085 22729 21097 22763
rect 21131 22760 21143 22763
rect 22186 22760 22192 22772
rect 21131 22732 22192 22760
rect 21131 22729 21143 22732
rect 21085 22723 21143 22729
rect 22186 22720 22192 22732
rect 22244 22720 22250 22772
rect 19076 22692 19104 22720
rect 19334 22692 19340 22704
rect 14568 22664 14964 22692
rect 15580 22664 18276 22692
rect 19076 22664 19340 22692
rect 15179 22657 15237 22663
rect 15179 22654 15191 22657
rect 12897 22627 12955 22633
rect 12897 22624 12909 22627
rect 12860 22596 12909 22624
rect 12860 22584 12866 22596
rect 12897 22593 12909 22596
rect 12943 22593 12955 22627
rect 12897 22587 12955 22593
rect 13078 22584 13084 22636
rect 13136 22584 13142 22636
rect 15178 22624 15191 22654
rect 14660 22623 15191 22624
rect 15225 22623 15237 22657
rect 14660 22617 15237 22623
rect 14660 22596 15206 22617
rect 13446 22516 13452 22568
rect 13504 22556 13510 22568
rect 13541 22559 13599 22565
rect 13541 22556 13553 22559
rect 13504 22528 13553 22556
rect 13504 22516 13510 22528
rect 13541 22525 13553 22528
rect 13587 22525 13599 22559
rect 13817 22559 13875 22565
rect 13817 22556 13829 22559
rect 13541 22519 13599 22525
rect 13648 22528 13829 22556
rect 13078 22488 13084 22500
rect 12176 22460 13084 22488
rect 13078 22448 13084 22460
rect 13136 22488 13142 22500
rect 13648 22488 13676 22528
rect 13817 22525 13829 22528
rect 13863 22525 13875 22559
rect 13817 22519 13875 22525
rect 13906 22516 13912 22568
rect 13964 22565 13970 22568
rect 13964 22559 13992 22565
rect 13980 22525 13992 22559
rect 13964 22519 13992 22525
rect 14093 22559 14151 22565
rect 14093 22525 14105 22559
rect 14139 22556 14151 22559
rect 14274 22556 14280 22568
rect 14139 22528 14280 22556
rect 14139 22525 14151 22528
rect 14093 22519 14151 22525
rect 13964 22516 13970 22519
rect 14274 22516 14280 22528
rect 14332 22516 14338 22568
rect 13136 22460 13676 22488
rect 13136 22448 13142 22460
rect 14660 22420 14688 22596
rect 14734 22516 14740 22568
rect 14792 22556 14798 22568
rect 14921 22559 14979 22565
rect 14921 22556 14933 22559
rect 14792 22528 14933 22556
rect 14792 22516 14798 22528
rect 14921 22525 14933 22528
rect 14967 22525 14979 22559
rect 14921 22519 14979 22525
rect 11256 22392 14688 22420
rect 15010 22380 15016 22432
rect 15068 22420 15074 22432
rect 15580 22420 15608 22664
rect 16390 22584 16396 22636
rect 16448 22624 16454 22636
rect 16942 22624 16948 22636
rect 16448 22596 16948 22624
rect 16448 22584 16454 22596
rect 16942 22584 16948 22596
rect 17000 22584 17006 22636
rect 17770 22584 17776 22636
rect 17828 22624 17834 22636
rect 18138 22633 18144 22636
rect 17865 22627 17923 22633
rect 17865 22624 17877 22627
rect 17828 22596 17877 22624
rect 17828 22584 17834 22596
rect 17865 22593 17877 22596
rect 17911 22593 17923 22627
rect 18132 22624 18144 22633
rect 18099 22596 18144 22624
rect 17865 22587 17923 22593
rect 18132 22587 18144 22596
rect 18138 22584 18144 22587
rect 18196 22584 18202 22636
rect 18248 22624 18276 22664
rect 19334 22652 19340 22664
rect 19392 22652 19398 22704
rect 20364 22692 20392 22720
rect 20364 22664 21312 22692
rect 19150 22624 19156 22636
rect 18248 22596 19156 22624
rect 19150 22584 19156 22596
rect 19208 22584 19214 22636
rect 19487 22624 19493 22646
rect 19352 22596 19493 22624
rect 19352 22565 19380 22596
rect 19487 22594 19493 22596
rect 19545 22594 19551 22646
rect 19579 22627 19637 22633
rect 19579 22593 19591 22627
rect 19625 22624 19637 22627
rect 20162 22624 20168 22636
rect 19625 22596 20168 22624
rect 19625 22593 19637 22596
rect 19579 22587 19637 22593
rect 20162 22584 20168 22596
rect 20220 22584 20226 22636
rect 20806 22584 20812 22636
rect 20864 22624 20870 22636
rect 21284 22633 21312 22664
rect 21910 22652 21916 22704
rect 21968 22692 21974 22704
rect 22738 22692 22744 22704
rect 21968 22664 22744 22692
rect 21968 22652 21974 22664
rect 22738 22652 22744 22664
rect 22796 22652 22802 22704
rect 20901 22627 20959 22633
rect 20901 22624 20913 22627
rect 20864 22596 20913 22624
rect 20864 22584 20870 22596
rect 20901 22593 20913 22596
rect 20947 22593 20959 22627
rect 20901 22587 20959 22593
rect 21269 22627 21327 22633
rect 21269 22593 21281 22627
rect 21315 22593 21327 22627
rect 21269 22587 21327 22593
rect 21726 22584 21732 22636
rect 21784 22624 21790 22636
rect 22370 22624 22376 22636
rect 21784 22596 22376 22624
rect 21784 22584 21790 22596
rect 22370 22584 22376 22596
rect 22428 22584 22434 22636
rect 19337 22559 19395 22565
rect 19337 22525 19349 22559
rect 19383 22525 19395 22559
rect 19337 22519 19395 22525
rect 21542 22516 21548 22568
rect 21600 22516 21606 22568
rect 21266 22448 21272 22500
rect 21324 22488 21330 22500
rect 21324 22460 21496 22488
rect 21324 22448 21330 22460
rect 15068 22392 15608 22420
rect 15068 22380 15074 22392
rect 15930 22380 15936 22432
rect 15988 22380 15994 22432
rect 17770 22380 17776 22432
rect 17828 22420 17834 22432
rect 18966 22420 18972 22432
rect 17828 22392 18972 22420
rect 17828 22380 17834 22392
rect 18966 22380 18972 22392
rect 19024 22380 19030 22432
rect 21358 22380 21364 22432
rect 21416 22380 21422 22432
rect 21468 22429 21496 22460
rect 21453 22423 21511 22429
rect 21453 22389 21465 22423
rect 21499 22389 21511 22423
rect 21453 22383 21511 22389
rect 1104 22330 21896 22352
rect 1104 22278 3549 22330
rect 3601 22278 3613 22330
rect 3665 22278 3677 22330
rect 3729 22278 3741 22330
rect 3793 22278 3805 22330
rect 3857 22278 8747 22330
rect 8799 22278 8811 22330
rect 8863 22278 8875 22330
rect 8927 22278 8939 22330
rect 8991 22278 9003 22330
rect 9055 22278 13945 22330
rect 13997 22278 14009 22330
rect 14061 22278 14073 22330
rect 14125 22278 14137 22330
rect 14189 22278 14201 22330
rect 14253 22278 19143 22330
rect 19195 22278 19207 22330
rect 19259 22278 19271 22330
rect 19323 22278 19335 22330
rect 19387 22278 19399 22330
rect 19451 22278 21896 22330
rect 1104 22256 21896 22278
rect 4154 22216 4160 22228
rect 1964 22188 4160 22216
rect 1964 22160 1992 22188
rect 4154 22176 4160 22188
rect 4212 22216 4218 22228
rect 4614 22216 4620 22228
rect 4212 22188 4620 22216
rect 4212 22176 4218 22188
rect 4614 22176 4620 22188
rect 4672 22176 4678 22228
rect 7374 22176 7380 22228
rect 7432 22216 7438 22228
rect 8202 22216 8208 22228
rect 7432 22188 8208 22216
rect 7432 22176 7438 22188
rect 8202 22176 8208 22188
rect 8260 22176 8266 22228
rect 9230 22188 9812 22216
rect 1946 22108 1952 22160
rect 2004 22108 2010 22160
rect 2406 22108 2412 22160
rect 2464 22148 2470 22160
rect 2777 22151 2835 22157
rect 2777 22148 2789 22151
rect 2464 22120 2789 22148
rect 2464 22108 2470 22120
rect 2777 22117 2789 22120
rect 2823 22117 2835 22151
rect 2777 22111 2835 22117
rect 474 22040 480 22092
rect 532 22080 538 22092
rect 658 22080 664 22092
rect 532 22052 664 22080
rect 532 22040 538 22052
rect 658 22040 664 22052
rect 716 22040 722 22092
rect 1394 22040 1400 22092
rect 1452 22040 1458 22092
rect 2792 22080 2820 22111
rect 3326 22108 3332 22160
rect 3384 22148 3390 22160
rect 3421 22151 3479 22157
rect 3421 22148 3433 22151
rect 3384 22120 3433 22148
rect 3384 22108 3390 22120
rect 3421 22117 3433 22120
rect 3467 22117 3479 22151
rect 3421 22111 3479 22117
rect 4246 22108 4252 22160
rect 4304 22148 4310 22160
rect 4798 22148 4804 22160
rect 4304 22120 4804 22148
rect 4304 22108 4310 22120
rect 4798 22108 4804 22120
rect 4856 22108 4862 22160
rect 6362 22108 6368 22160
rect 6420 22108 6426 22160
rect 7282 22108 7288 22160
rect 7340 22148 7346 22160
rect 8570 22148 8576 22160
rect 7340 22120 8576 22148
rect 7340 22108 7346 22120
rect 8570 22108 8576 22120
rect 8628 22108 8634 22160
rect 9230 22148 9258 22188
rect 9140 22120 9258 22148
rect 4896 22092 4948 22098
rect 1504 22052 2636 22080
rect 2792 22052 4844 22080
rect 1210 21972 1216 22024
rect 1268 22012 1274 22024
rect 1504 22012 1532 22052
rect 1268 21984 1532 22012
rect 1268 21972 1274 21984
rect 1670 21972 1676 22024
rect 1728 21972 1734 22024
rect 2314 21972 2320 22024
rect 2372 21972 2378 22024
rect 2608 22021 2636 22052
rect 2593 22015 2651 22021
rect 2593 21981 2605 22015
rect 2639 21981 2651 22015
rect 2593 21975 2651 21981
rect 3237 21991 3295 21997
rect 3237 21957 3249 21991
rect 3283 21957 3295 21991
rect 4614 21972 4620 22024
rect 4672 21972 4678 22024
rect 4816 22006 4844 22052
rect 6454 22040 6460 22092
rect 6512 22080 6518 22092
rect 6549 22083 6607 22089
rect 6549 22080 6561 22083
rect 6512 22052 6561 22080
rect 6512 22040 6518 22052
rect 6549 22049 6561 22052
rect 6595 22049 6607 22083
rect 6549 22043 6607 22049
rect 8021 22083 8079 22089
rect 8021 22049 8033 22083
rect 8067 22080 8079 22083
rect 8662 22080 8668 22092
rect 8067 22052 8668 22080
rect 8067 22049 8079 22052
rect 8021 22043 8079 22049
rect 8662 22040 8668 22052
rect 8720 22040 8726 22092
rect 9140 22089 9168 22120
rect 9125 22083 9183 22089
rect 9125 22049 9137 22083
rect 9171 22049 9183 22083
rect 9125 22043 9183 22049
rect 9784 22080 9812 22188
rect 10042 22176 10048 22228
rect 10100 22216 10106 22228
rect 10137 22219 10195 22225
rect 10137 22216 10149 22219
rect 10100 22188 10149 22216
rect 10100 22176 10106 22188
rect 10137 22185 10149 22188
rect 10183 22185 10195 22219
rect 10870 22216 10876 22228
rect 10137 22179 10195 22185
rect 10242 22188 10876 22216
rect 9858 22108 9864 22160
rect 9916 22148 9922 22160
rect 10242 22148 10270 22188
rect 10870 22176 10876 22188
rect 10928 22176 10934 22228
rect 11054 22176 11060 22228
rect 11112 22216 11118 22228
rect 12066 22216 12072 22228
rect 11112 22188 12072 22216
rect 11112 22176 11118 22188
rect 12066 22176 12072 22188
rect 12124 22176 12130 22228
rect 13814 22216 13820 22228
rect 12820 22188 13820 22216
rect 9916 22120 10270 22148
rect 9916 22108 9922 22120
rect 12618 22108 12624 22160
rect 12676 22148 12682 22160
rect 12676 22120 12756 22148
rect 12676 22108 12682 22120
rect 10594 22080 10600 22092
rect 9784 22052 10600 22080
rect 4896 22034 4948 22040
rect 9784 22024 9812 22052
rect 10594 22040 10600 22052
rect 10652 22040 10658 22092
rect 11698 22040 11704 22092
rect 11756 22080 11762 22092
rect 12728 22089 12756 22120
rect 12069 22083 12127 22089
rect 12069 22080 12081 22083
rect 11756 22052 12081 22080
rect 11756 22040 11762 22052
rect 12069 22049 12081 22052
rect 12115 22049 12127 22083
rect 12069 22043 12127 22049
rect 12713 22083 12771 22089
rect 12713 22049 12725 22083
rect 12759 22049 12771 22083
rect 12820 22080 12848 22188
rect 13814 22176 13820 22188
rect 13872 22216 13878 22228
rect 14182 22216 14188 22228
rect 13872 22188 14188 22216
rect 13872 22176 13878 22188
rect 14182 22176 14188 22188
rect 14240 22176 14246 22228
rect 14366 22176 14372 22228
rect 14424 22176 14430 22228
rect 14734 22176 14740 22228
rect 14792 22216 14798 22228
rect 15194 22216 15200 22228
rect 14792 22188 15200 22216
rect 14792 22176 14798 22188
rect 15194 22176 15200 22188
rect 15252 22216 15258 22228
rect 15252 22188 17356 22216
rect 15252 22176 15258 22188
rect 14384 22148 14412 22176
rect 13832 22120 14412 22148
rect 13832 22092 13860 22120
rect 15562 22108 15568 22160
rect 15620 22108 15626 22160
rect 15930 22108 15936 22160
rect 15988 22148 15994 22160
rect 16025 22151 16083 22157
rect 16025 22148 16037 22151
rect 15988 22120 16037 22148
rect 15988 22108 15994 22120
rect 16025 22117 16037 22120
rect 16071 22117 16083 22151
rect 16025 22111 16083 22117
rect 12989 22083 13047 22089
rect 12989 22080 13001 22083
rect 12820 22052 13001 22080
rect 12713 22043 12771 22049
rect 12989 22049 13001 22052
rect 13035 22049 13047 22083
rect 12989 22043 13047 22049
rect 13262 22040 13268 22092
rect 13320 22040 13326 22092
rect 13814 22040 13820 22092
rect 13872 22040 13878 22092
rect 15378 22040 15384 22092
rect 15436 22040 15442 22092
rect 15580 22080 15608 22108
rect 17328 22089 17356 22188
rect 17402 22176 17408 22228
rect 17460 22216 17466 22228
rect 19426 22216 19432 22228
rect 17460 22188 19432 22216
rect 17460 22176 17466 22188
rect 19426 22176 19432 22188
rect 19484 22176 19490 22228
rect 20346 22176 20352 22228
rect 20404 22216 20410 22228
rect 20404 22188 20484 22216
rect 20404 22176 20410 22188
rect 20456 22148 20484 22188
rect 21450 22176 21456 22228
rect 21508 22176 21514 22228
rect 22922 22176 22928 22228
rect 22980 22176 22986 22228
rect 22940 22148 22968 22176
rect 20456 22120 22968 22148
rect 16418 22083 16476 22089
rect 16418 22080 16430 22083
rect 15580 22052 16430 22080
rect 16418 22049 16430 22052
rect 16464 22049 16476 22083
rect 16418 22043 16476 22049
rect 16577 22083 16635 22089
rect 16577 22049 16589 22083
rect 16623 22080 16635 22083
rect 17313 22083 17371 22089
rect 16623 22052 17264 22080
rect 16623 22049 16635 22052
rect 16577 22043 16635 22049
rect 4982 22006 4988 22024
rect 4816 21978 4988 22006
rect 4982 21972 4988 21978
rect 5040 21972 5046 22024
rect 5350 21972 5356 22024
rect 5408 21972 5414 22024
rect 5445 22015 5503 22021
rect 5445 21981 5457 22015
rect 5491 22012 5503 22015
rect 6823 22015 6881 22021
rect 5491 21984 6040 22012
rect 5491 21981 5503 21984
rect 5445 21975 5503 21981
rect 750 21904 756 21956
rect 808 21944 814 21956
rect 2961 21947 3019 21953
rect 3237 21951 3295 21957
rect 2961 21944 2973 21947
rect 808 21916 2973 21944
rect 808 21904 814 21916
rect 2961 21913 2973 21916
rect 3007 21913 3019 21947
rect 2961 21907 3019 21913
rect 3252 21888 3280 21951
rect 4632 21944 4660 21972
rect 5368 21944 5396 21972
rect 5813 21947 5871 21953
rect 5813 21944 5825 21947
rect 4632 21916 5396 21944
rect 5552 21916 5825 21944
rect 2501 21879 2559 21885
rect 2501 21845 2513 21879
rect 2547 21876 2559 21879
rect 2682 21876 2688 21888
rect 2547 21848 2688 21876
rect 2547 21845 2559 21848
rect 2501 21839 2559 21845
rect 2682 21836 2688 21848
rect 2740 21836 2746 21888
rect 2866 21836 2872 21888
rect 2924 21876 2930 21888
rect 3053 21879 3111 21885
rect 3053 21876 3065 21879
rect 2924 21848 3065 21876
rect 2924 21836 2930 21848
rect 3053 21845 3065 21848
rect 3099 21845 3111 21879
rect 3053 21839 3111 21845
rect 3234 21836 3240 21888
rect 3292 21836 3298 21888
rect 4982 21836 4988 21888
rect 5040 21876 5046 21888
rect 5077 21879 5135 21885
rect 5077 21876 5089 21879
rect 5040 21848 5089 21876
rect 5040 21836 5046 21848
rect 5077 21845 5089 21848
rect 5123 21845 5135 21879
rect 5077 21839 5135 21845
rect 5350 21836 5356 21888
rect 5408 21876 5414 21888
rect 5552 21876 5580 21916
rect 5813 21913 5825 21916
rect 5859 21913 5871 21947
rect 6012 21944 6040 21984
rect 6823 21981 6835 22015
rect 6869 22012 6881 22015
rect 7742 22012 7748 22024
rect 6869 21984 7748 22012
rect 6869 21981 6881 21984
rect 6823 21975 6881 21981
rect 7742 21972 7748 21984
rect 7800 21972 7806 22024
rect 7926 21972 7932 22024
rect 7984 21972 7990 22024
rect 8113 22015 8171 22021
rect 8113 22012 8125 22015
rect 8036 21984 8125 22012
rect 8036 21956 8064 21984
rect 8113 21981 8125 21984
rect 8159 21981 8171 22015
rect 8113 21975 8171 21981
rect 8294 21972 8300 22024
rect 8352 21972 8358 22024
rect 8386 21972 8392 22024
rect 8444 22012 8450 22024
rect 9367 22015 9425 22021
rect 8956 22012 9076 22014
rect 9140 22012 9260 22014
rect 9367 22012 9379 22015
rect 8444 21986 9379 22012
rect 8444 21984 8984 21986
rect 9048 21984 9168 21986
rect 9232 21984 9379 21986
rect 8444 21972 8450 21984
rect 9367 21981 9379 21984
rect 9413 21981 9425 22015
rect 9367 21975 9425 21981
rect 9766 21972 9772 22024
rect 9824 21972 9830 22024
rect 10318 21972 10324 22024
rect 10376 22012 10382 22024
rect 10839 22015 10897 22021
rect 10839 22012 10851 22015
rect 10376 21984 10851 22012
rect 10376 21972 10382 21984
rect 10839 21981 10851 21984
rect 10885 21981 10897 22015
rect 10839 21975 10897 21981
rect 12250 21972 12256 22024
rect 12308 21972 12314 22024
rect 13078 21972 13084 22024
rect 13136 22021 13142 22024
rect 13136 22015 13164 22021
rect 13152 21981 13164 22015
rect 15194 22012 15200 22024
rect 13136 21975 13164 21981
rect 14317 21984 15200 22012
rect 13136 21972 13142 21975
rect 6012 21916 6592 21944
rect 5813 21907 5871 21913
rect 5408 21848 5580 21876
rect 5408 21836 5414 21848
rect 5626 21836 5632 21888
rect 5684 21876 5690 21888
rect 6181 21879 6239 21885
rect 6181 21876 6193 21879
rect 5684 21848 6193 21876
rect 5684 21836 5690 21848
rect 6181 21845 6193 21848
rect 6227 21845 6239 21879
rect 6564 21876 6592 21916
rect 6730 21904 6736 21956
rect 6788 21944 6794 21956
rect 6788 21916 7696 21944
rect 6788 21904 6794 21916
rect 7561 21879 7619 21885
rect 7561 21876 7573 21879
rect 6564 21848 7573 21876
rect 6181 21839 6239 21845
rect 7561 21845 7573 21848
rect 7607 21845 7619 21879
rect 7668 21876 7696 21916
rect 8018 21904 8024 21956
rect 8076 21904 8082 21956
rect 8312 21944 8340 21972
rect 8662 21944 8668 21956
rect 8312 21916 8668 21944
rect 8662 21904 8668 21916
rect 8720 21904 8726 21956
rect 14317 21944 14345 21984
rect 15194 21972 15200 21984
rect 15252 22012 15258 22024
rect 15565 22015 15623 22021
rect 15252 21984 15332 22012
rect 15252 21972 15258 21984
rect 9876 21916 12296 21944
rect 9876 21876 9904 21916
rect 7668 21848 9904 21876
rect 11609 21879 11667 21885
rect 7561 21839 7619 21845
rect 11609 21845 11621 21879
rect 11655 21876 11667 21879
rect 11698 21876 11704 21888
rect 11655 21848 11704 21876
rect 11655 21845 11667 21848
rect 11609 21839 11667 21845
rect 11698 21836 11704 21848
rect 11756 21836 11762 21888
rect 12268 21876 12296 21916
rect 13832 21916 14345 21944
rect 15304 21944 15332 21984
rect 15565 21981 15577 22015
rect 15611 21981 15623 22015
rect 15565 21975 15623 21981
rect 15580 21944 15608 21975
rect 16298 21972 16304 22024
rect 16356 21972 16362 22024
rect 17236 22012 17264 22052
rect 17313 22049 17325 22083
rect 17359 22049 17371 22083
rect 21450 22080 21456 22092
rect 17313 22043 17371 22049
rect 20916 22052 21456 22080
rect 17587 22015 17645 22021
rect 17236 21984 17448 22012
rect 15304 21916 15608 21944
rect 13832 21876 13860 21916
rect 12268 21848 13860 21876
rect 13909 21879 13967 21885
rect 13909 21845 13921 21879
rect 13955 21876 13967 21879
rect 14366 21876 14372 21888
rect 13955 21848 14372 21876
rect 13955 21845 13967 21848
rect 13909 21839 13967 21845
rect 14366 21836 14372 21848
rect 14424 21836 14430 21888
rect 17034 21836 17040 21888
rect 17092 21876 17098 21888
rect 17221 21879 17279 21885
rect 17221 21876 17233 21879
rect 17092 21848 17233 21876
rect 17092 21836 17098 21848
rect 17221 21845 17233 21848
rect 17267 21845 17279 21879
rect 17420 21876 17448 21984
rect 17587 21981 17599 22015
rect 17633 22012 17645 22015
rect 17633 21984 17724 22012
rect 17633 21981 17645 21984
rect 17587 21975 17645 21981
rect 17696 21956 17724 21984
rect 18322 21972 18328 22024
rect 18380 22012 18386 22024
rect 18877 22015 18935 22021
rect 18877 22012 18889 22015
rect 18380 21984 18889 22012
rect 18380 21972 18386 21984
rect 18877 21981 18889 21984
rect 18923 21981 18935 22015
rect 18877 21975 18935 21981
rect 18966 21972 18972 22024
rect 19024 22012 19030 22024
rect 20916 22021 20944 22052
rect 21450 22040 21456 22052
rect 21508 22040 21514 22092
rect 19429 22015 19487 22021
rect 19429 22012 19441 22015
rect 19024 21984 19441 22012
rect 19024 21972 19030 21984
rect 19429 21981 19441 21984
rect 19475 21981 19487 22015
rect 19429 21975 19487 21981
rect 20901 22015 20959 22021
rect 20901 21981 20913 22015
rect 20947 21981 20959 22015
rect 20901 21975 20959 21981
rect 21266 21972 21272 22024
rect 21324 21972 21330 22024
rect 21358 21972 21364 22024
rect 21416 21972 21422 22024
rect 21542 21972 21548 22024
rect 21600 22012 21606 22024
rect 22186 22012 22192 22024
rect 21600 21984 22192 22012
rect 21600 21972 21606 21984
rect 22186 21972 22192 21984
rect 22244 21972 22250 22024
rect 17678 21904 17684 21956
rect 17736 21904 17742 21956
rect 19696 21947 19754 21953
rect 19696 21913 19708 21947
rect 19742 21944 19754 21947
rect 20070 21944 20076 21956
rect 19742 21916 20076 21944
rect 19742 21913 19754 21916
rect 19696 21907 19754 21913
rect 20070 21904 20076 21916
rect 20128 21904 20134 21956
rect 21376 21944 21404 21972
rect 20180 21916 21404 21944
rect 18325 21879 18383 21885
rect 18325 21876 18337 21879
rect 17420 21848 18337 21876
rect 17221 21839 17279 21845
rect 18325 21845 18337 21848
rect 18371 21845 18383 21879
rect 18325 21839 18383 21845
rect 18969 21879 19027 21885
rect 18969 21845 18981 21879
rect 19015 21876 19027 21879
rect 20180 21876 20208 21916
rect 19015 21848 20208 21876
rect 20809 21879 20867 21885
rect 19015 21845 19027 21848
rect 18969 21839 19027 21845
rect 20809 21845 20821 21879
rect 20855 21876 20867 21879
rect 20990 21876 20996 21888
rect 20855 21848 20996 21876
rect 20855 21845 20867 21848
rect 20809 21839 20867 21845
rect 20990 21836 20996 21848
rect 21048 21836 21054 21888
rect 21085 21879 21143 21885
rect 21085 21845 21097 21879
rect 21131 21876 21143 21879
rect 22186 21876 22192 21888
rect 21131 21848 22192 21876
rect 21131 21845 21143 21848
rect 21085 21839 21143 21845
rect 22186 21836 22192 21848
rect 22244 21836 22250 21888
rect 1104 21786 22056 21808
rect 1104 21734 6148 21786
rect 6200 21734 6212 21786
rect 6264 21734 6276 21786
rect 6328 21734 6340 21786
rect 6392 21734 6404 21786
rect 6456 21734 11346 21786
rect 11398 21734 11410 21786
rect 11462 21734 11474 21786
rect 11526 21734 11538 21786
rect 11590 21734 11602 21786
rect 11654 21734 16544 21786
rect 16596 21734 16608 21786
rect 16660 21734 16672 21786
rect 16724 21734 16736 21786
rect 16788 21734 16800 21786
rect 16852 21734 21742 21786
rect 21794 21734 21806 21786
rect 21858 21734 21870 21786
rect 21922 21734 21934 21786
rect 21986 21734 21998 21786
rect 22050 21734 22056 21786
rect 1104 21712 22056 21734
rect 3418 21672 3424 21684
rect 2884 21644 3424 21672
rect 1670 21496 1676 21548
rect 1728 21536 1734 21548
rect 2884 21545 2912 21644
rect 3418 21632 3424 21644
rect 3476 21632 3482 21684
rect 3878 21632 3884 21684
rect 3936 21632 3942 21684
rect 4522 21632 4528 21684
rect 4580 21672 4586 21684
rect 5626 21672 5632 21684
rect 4580 21644 5632 21672
rect 4580 21632 4586 21644
rect 5626 21632 5632 21644
rect 5684 21632 5690 21684
rect 5718 21632 5724 21684
rect 5776 21672 5782 21684
rect 5813 21675 5871 21681
rect 5813 21672 5825 21675
rect 5776 21644 5825 21672
rect 5776 21632 5782 21644
rect 5813 21641 5825 21644
rect 5859 21641 5871 21675
rect 5813 21635 5871 21641
rect 7742 21632 7748 21684
rect 7800 21672 7806 21684
rect 9490 21672 9496 21684
rect 7800 21644 9496 21672
rect 7800 21632 7806 21644
rect 9490 21632 9496 21644
rect 9548 21632 9554 21684
rect 9950 21632 9956 21684
rect 10008 21632 10014 21684
rect 10226 21632 10232 21684
rect 10284 21632 10290 21684
rect 10413 21675 10471 21681
rect 10413 21641 10425 21675
rect 10459 21672 10471 21675
rect 12618 21672 12624 21684
rect 10459 21644 12624 21672
rect 10459 21641 10471 21644
rect 10413 21635 10471 21641
rect 12618 21632 12624 21644
rect 12676 21632 12682 21684
rect 12710 21632 12716 21684
rect 12768 21672 12774 21684
rect 12805 21675 12863 21681
rect 12805 21672 12817 21675
rect 12768 21644 12817 21672
rect 12768 21632 12774 21644
rect 12805 21641 12817 21644
rect 12851 21641 12863 21675
rect 12805 21635 12863 21641
rect 12894 21632 12900 21684
rect 12952 21672 12958 21684
rect 13078 21672 13084 21684
rect 12952 21644 13084 21672
rect 12952 21632 12958 21644
rect 13078 21632 13084 21644
rect 13136 21632 13142 21684
rect 15194 21632 15200 21684
rect 15252 21672 15258 21684
rect 15252 21644 16712 21672
rect 15252 21632 15258 21644
rect 4338 21604 4344 21616
rect 3068 21576 4344 21604
rect 3068 21548 3096 21576
rect 1763 21539 1821 21545
rect 1763 21536 1775 21539
rect 1728 21508 1775 21536
rect 1728 21496 1734 21508
rect 1763 21505 1775 21508
rect 1809 21505 1821 21539
rect 1763 21499 1821 21505
rect 2869 21539 2927 21545
rect 2869 21505 2881 21539
rect 2915 21505 2927 21539
rect 2869 21499 2927 21505
rect 3050 21496 3056 21548
rect 3108 21496 3114 21548
rect 3143 21539 3201 21545
rect 3143 21505 3155 21539
rect 3189 21536 3201 21539
rect 4062 21536 4068 21548
rect 3189 21508 4068 21536
rect 3189 21505 3201 21508
rect 3143 21499 3201 21505
rect 4062 21496 4068 21508
rect 4120 21496 4126 21548
rect 1210 21428 1216 21480
rect 1268 21468 1274 21480
rect 4264 21477 4292 21576
rect 4338 21564 4344 21576
rect 4396 21564 4402 21616
rect 9030 21604 9036 21616
rect 4816 21576 9036 21604
rect 4523 21549 4581 21555
rect 4523 21515 4535 21549
rect 4569 21536 4581 21549
rect 4816 21536 4844 21576
rect 9030 21564 9036 21576
rect 9088 21564 9094 21616
rect 9122 21564 9128 21616
rect 9180 21564 9186 21616
rect 9766 21570 9772 21616
rect 9600 21564 9772 21570
rect 9824 21564 9830 21616
rect 9861 21607 9919 21613
rect 9861 21573 9873 21607
rect 9907 21604 9919 21607
rect 9968 21604 9996 21632
rect 9907 21576 9996 21604
rect 9907 21573 9919 21576
rect 9861 21567 9919 21573
rect 11054 21564 11060 21616
rect 11112 21604 11118 21616
rect 11701 21607 11759 21613
rect 11701 21604 11713 21607
rect 11112 21576 11713 21604
rect 11112 21564 11118 21576
rect 11701 21573 11713 21576
rect 11747 21573 11759 21607
rect 11701 21567 11759 21573
rect 12437 21607 12495 21613
rect 12437 21573 12449 21607
rect 12483 21573 12495 21607
rect 12437 21567 12495 21573
rect 4569 21515 4844 21536
rect 4523 21509 4844 21515
rect 4538 21508 4844 21509
rect 4890 21496 4896 21548
rect 4948 21496 4954 21548
rect 7374 21496 7380 21548
rect 7432 21536 7438 21548
rect 7803 21539 7861 21545
rect 7803 21536 7815 21539
rect 7432 21508 7815 21536
rect 7432 21496 7438 21508
rect 7803 21505 7815 21508
rect 7849 21505 7861 21539
rect 7803 21499 7861 21505
rect 9398 21496 9404 21548
rect 9456 21496 9462 21548
rect 9493 21539 9551 21545
rect 9493 21505 9505 21539
rect 9539 21536 9551 21539
rect 9600 21542 9812 21564
rect 9600 21536 9628 21542
rect 9539 21508 9628 21536
rect 9539 21505 9551 21508
rect 9493 21499 9551 21505
rect 11238 21496 11244 21548
rect 11296 21536 11302 21548
rect 11977 21539 12035 21545
rect 11977 21536 11989 21539
rect 11296 21508 11989 21536
rect 11296 21496 11302 21508
rect 11977 21505 11989 21508
rect 12023 21505 12035 21539
rect 11977 21499 12035 21505
rect 12066 21496 12072 21548
rect 12124 21496 12130 21548
rect 12452 21536 12480 21567
rect 13630 21564 13636 21616
rect 13688 21604 13694 21616
rect 13688 21576 15240 21604
rect 13688 21564 13694 21576
rect 15212 21548 15240 21576
rect 13446 21536 13452 21548
rect 12452 21508 13452 21536
rect 13446 21496 13452 21508
rect 13504 21496 13510 21548
rect 15194 21496 15200 21548
rect 15252 21496 15258 21548
rect 16684 21545 16712 21644
rect 20070 21564 20076 21616
rect 20128 21604 20134 21616
rect 20622 21604 20628 21616
rect 20128 21576 20628 21604
rect 20128 21564 20134 21576
rect 20622 21564 20628 21576
rect 20680 21604 20686 21616
rect 20680 21576 21588 21604
rect 20680 21564 20686 21576
rect 19855 21549 19913 21555
rect 16669 21539 16727 21545
rect 16669 21505 16681 21539
rect 16715 21505 16727 21539
rect 16669 21499 16727 21505
rect 17586 21496 17592 21548
rect 17644 21496 17650 21548
rect 19426 21496 19432 21548
rect 19484 21536 19490 21548
rect 19855 21536 19867 21549
rect 19484 21515 19867 21536
rect 19901 21546 19913 21549
rect 19901 21515 19914 21546
rect 19484 21508 19914 21515
rect 19484 21496 19490 21508
rect 20898 21496 20904 21548
rect 20956 21536 20962 21548
rect 21560 21545 21588 21576
rect 20993 21539 21051 21545
rect 20993 21536 21005 21539
rect 20956 21508 21005 21536
rect 20956 21496 20962 21508
rect 20993 21505 21005 21508
rect 21039 21505 21051 21539
rect 20993 21499 21051 21505
rect 21545 21539 21603 21545
rect 21545 21505 21557 21539
rect 21591 21505 21603 21539
rect 21545 21499 21603 21505
rect 1489 21471 1547 21477
rect 1489 21468 1501 21471
rect 1268 21440 1501 21468
rect 1268 21428 1274 21440
rect 1489 21437 1501 21440
rect 1535 21437 1547 21471
rect 1489 21431 1547 21437
rect 4249 21471 4307 21477
rect 4249 21437 4261 21471
rect 4295 21437 4307 21471
rect 4249 21431 4307 21437
rect 4908 21400 4936 21496
rect 6914 21468 6920 21480
rect 5552 21440 6920 21468
rect 5261 21403 5319 21409
rect 5261 21400 5273 21403
rect 4908 21372 5273 21400
rect 5261 21369 5273 21372
rect 5307 21369 5319 21403
rect 5261 21363 5319 21369
rect 198 21292 204 21344
rect 256 21332 262 21344
rect 2406 21332 2412 21344
rect 256 21304 2412 21332
rect 256 21292 262 21304
rect 2406 21292 2412 21304
rect 2464 21292 2470 21344
rect 2501 21335 2559 21341
rect 2501 21301 2513 21335
rect 2547 21332 2559 21335
rect 3878 21332 3884 21344
rect 2547 21304 3884 21332
rect 2547 21301 2559 21304
rect 2501 21295 2559 21301
rect 3878 21292 3884 21304
rect 3936 21292 3942 21344
rect 4246 21292 4252 21344
rect 4304 21332 4310 21344
rect 5552 21332 5580 21440
rect 6914 21428 6920 21440
rect 6972 21428 6978 21480
rect 7558 21428 7564 21480
rect 7616 21428 7622 21480
rect 8588 21440 8970 21468
rect 4304 21304 5580 21332
rect 4304 21292 4310 21304
rect 5626 21292 5632 21344
rect 5684 21332 5690 21344
rect 5902 21332 5908 21344
rect 5684 21304 5908 21332
rect 5684 21292 5690 21304
rect 5902 21292 5908 21304
rect 5960 21292 5966 21344
rect 6178 21292 6184 21344
rect 6236 21332 6242 21344
rect 6730 21332 6736 21344
rect 6236 21304 6736 21332
rect 6236 21292 6242 21304
rect 6730 21292 6736 21304
rect 6788 21292 6794 21344
rect 7576 21332 7604 21428
rect 8588 21409 8616 21440
rect 11606 21428 11612 21480
rect 11664 21428 11670 21480
rect 16206 21468 16212 21480
rect 13740 21440 16212 21468
rect 8573 21403 8631 21409
rect 8573 21369 8585 21403
rect 8619 21369 8631 21403
rect 8573 21363 8631 21369
rect 13262 21360 13268 21412
rect 13320 21400 13326 21412
rect 13446 21400 13452 21412
rect 13320 21372 13452 21400
rect 13320 21360 13326 21372
rect 13446 21360 13452 21372
rect 13504 21360 13510 21412
rect 13740 21344 13768 21440
rect 16206 21428 16212 21440
rect 16264 21428 16270 21480
rect 16850 21428 16856 21480
rect 16908 21428 16914 21480
rect 17706 21471 17764 21477
rect 17706 21468 17718 21471
rect 16942 21440 17718 21468
rect 14458 21360 14464 21412
rect 14516 21400 14522 21412
rect 15378 21400 15384 21412
rect 14516 21372 15384 21400
rect 14516 21360 14522 21372
rect 15378 21360 15384 21372
rect 15436 21400 15442 21412
rect 16942 21400 16970 21440
rect 17706 21437 17718 21440
rect 17752 21437 17764 21471
rect 17706 21431 17764 21437
rect 17862 21428 17868 21480
rect 17920 21428 17926 21480
rect 19518 21428 19524 21480
rect 19576 21468 19582 21480
rect 19613 21471 19671 21477
rect 19613 21468 19625 21471
rect 19576 21440 19625 21468
rect 19576 21428 19582 21440
rect 19613 21437 19625 21440
rect 19659 21437 19671 21471
rect 19613 21431 19671 21437
rect 15436 21372 16970 21400
rect 17313 21403 17371 21409
rect 15436 21360 15442 21372
rect 17313 21369 17325 21403
rect 17359 21400 17371 21403
rect 17402 21400 17408 21412
rect 17359 21372 17408 21400
rect 17359 21369 17371 21372
rect 17313 21363 17371 21369
rect 17402 21360 17408 21372
rect 17460 21360 17466 21412
rect 20625 21403 20683 21409
rect 20625 21369 20637 21403
rect 20671 21400 20683 21403
rect 20916 21400 20944 21496
rect 21269 21471 21327 21477
rect 21269 21437 21281 21471
rect 21315 21468 21327 21471
rect 21358 21468 21364 21480
rect 21315 21440 21364 21468
rect 21315 21437 21327 21440
rect 21269 21431 21327 21437
rect 21358 21428 21364 21440
rect 21416 21428 21422 21480
rect 20671 21372 20944 21400
rect 20671 21369 20683 21372
rect 20625 21363 20683 21369
rect 7926 21332 7932 21344
rect 7576 21304 7932 21332
rect 7926 21292 7932 21304
rect 7984 21292 7990 21344
rect 10318 21292 10324 21344
rect 10376 21332 10382 21344
rect 10781 21335 10839 21341
rect 10781 21332 10793 21335
rect 10376 21304 10793 21332
rect 10376 21292 10382 21304
rect 10781 21301 10793 21304
rect 10827 21301 10839 21335
rect 10781 21295 10839 21301
rect 12986 21292 12992 21344
rect 13044 21292 13050 21344
rect 13722 21292 13728 21344
rect 13780 21292 13786 21344
rect 14274 21292 14280 21344
rect 14332 21332 14338 21344
rect 15746 21332 15752 21344
rect 14332 21304 15752 21332
rect 14332 21292 14338 21304
rect 15746 21292 15752 21304
rect 15804 21332 15810 21344
rect 17586 21332 17592 21344
rect 15804 21304 17592 21332
rect 15804 21292 15810 21304
rect 17586 21292 17592 21304
rect 17644 21292 17650 21344
rect 18509 21335 18567 21341
rect 18509 21301 18521 21335
rect 18555 21332 18567 21335
rect 19058 21332 19064 21344
rect 18555 21304 19064 21332
rect 18555 21301 18567 21304
rect 18509 21295 18567 21301
rect 19058 21292 19064 21304
rect 19116 21292 19122 21344
rect 20070 21292 20076 21344
rect 20128 21332 20134 21344
rect 20346 21332 20352 21344
rect 20128 21304 20352 21332
rect 20128 21292 20134 21304
rect 20346 21292 20352 21304
rect 20404 21292 20410 21344
rect 20530 21292 20536 21344
rect 20588 21332 20594 21344
rect 21085 21335 21143 21341
rect 21085 21332 21097 21335
rect 20588 21304 21097 21332
rect 20588 21292 20594 21304
rect 21085 21301 21097 21304
rect 21131 21301 21143 21335
rect 21085 21295 21143 21301
rect 21174 21292 21180 21344
rect 21232 21292 21238 21344
rect 21266 21292 21272 21344
rect 21324 21332 21330 21344
rect 21361 21335 21419 21341
rect 21361 21332 21373 21335
rect 21324 21304 21373 21332
rect 21324 21292 21330 21304
rect 21361 21301 21373 21304
rect 21407 21301 21419 21335
rect 21361 21295 21419 21301
rect 1104 21242 21896 21264
rect 1104 21190 3549 21242
rect 3601 21190 3613 21242
rect 3665 21190 3677 21242
rect 3729 21190 3741 21242
rect 3793 21190 3805 21242
rect 3857 21190 8747 21242
rect 8799 21190 8811 21242
rect 8863 21190 8875 21242
rect 8927 21190 8939 21242
rect 8991 21190 9003 21242
rect 9055 21190 13945 21242
rect 13997 21190 14009 21242
rect 14061 21190 14073 21242
rect 14125 21190 14137 21242
rect 14189 21190 14201 21242
rect 14253 21190 19143 21242
rect 19195 21190 19207 21242
rect 19259 21190 19271 21242
rect 19323 21190 19335 21242
rect 19387 21190 19399 21242
rect 19451 21190 21896 21242
rect 1104 21168 21896 21190
rect 2038 21088 2044 21140
rect 2096 21128 2102 21140
rect 2096 21100 3096 21128
rect 2096 21088 2102 21100
rect 2222 21060 2228 21072
rect 1688 21032 2228 21060
rect 750 20952 756 21004
rect 808 20992 814 21004
rect 1688 21001 1716 21032
rect 2222 21020 2228 21032
rect 2280 21020 2286 21072
rect 3068 21060 3096 21100
rect 3142 21088 3148 21140
rect 3200 21128 3206 21140
rect 3973 21131 4031 21137
rect 3973 21128 3985 21131
rect 3200 21100 3985 21128
rect 3200 21088 3206 21100
rect 3973 21097 3985 21100
rect 4019 21097 4031 21131
rect 4522 21128 4528 21140
rect 3973 21091 4031 21097
rect 4170 21100 4528 21128
rect 4170 21060 4198 21100
rect 4522 21088 4528 21100
rect 4580 21088 4586 21140
rect 5721 21131 5779 21137
rect 5721 21097 5733 21131
rect 5767 21128 5779 21131
rect 6178 21128 6184 21140
rect 5767 21100 6184 21128
rect 5767 21097 5779 21100
rect 5721 21091 5779 21097
rect 6178 21088 6184 21100
rect 6236 21088 6242 21140
rect 8110 21088 8116 21140
rect 8168 21128 8174 21140
rect 9030 21128 9036 21140
rect 8168 21100 9036 21128
rect 8168 21088 8174 21100
rect 9030 21088 9036 21100
rect 9088 21088 9094 21140
rect 9214 21088 9220 21140
rect 9272 21128 9278 21140
rect 9272 21100 9628 21128
rect 9272 21088 9278 21100
rect 3068 21032 4198 21060
rect 5077 21063 5135 21069
rect 5077 21029 5089 21063
rect 5123 21060 5135 21063
rect 9600 21060 9628 21100
rect 9766 21088 9772 21140
rect 9824 21128 9830 21140
rect 9953 21131 10011 21137
rect 9953 21128 9965 21131
rect 9824 21100 9965 21128
rect 9824 21088 9830 21100
rect 9953 21097 9965 21100
rect 9999 21097 10011 21131
rect 9953 21091 10011 21097
rect 11238 21088 11244 21140
rect 11296 21088 11302 21140
rect 12066 21088 12072 21140
rect 12124 21128 12130 21140
rect 12253 21131 12311 21137
rect 12253 21128 12265 21131
rect 12124 21100 12265 21128
rect 12124 21088 12130 21100
rect 12253 21097 12265 21100
rect 12299 21097 12311 21131
rect 12253 21091 12311 21097
rect 12618 21088 12624 21140
rect 12676 21128 12682 21140
rect 12676 21100 17356 21128
rect 12676 21088 12682 21100
rect 11256 21060 11284 21088
rect 5123 21032 6040 21060
rect 9600 21032 11284 21060
rect 5123 21029 5135 21032
rect 5077 21023 5135 21029
rect 1397 20995 1455 21001
rect 1397 20992 1409 20995
rect 808 20964 1409 20992
rect 808 20952 814 20964
rect 1397 20961 1409 20964
rect 1443 20961 1455 20995
rect 1397 20955 1455 20961
rect 1673 20995 1731 21001
rect 1673 20961 1685 20995
rect 1719 20961 1731 20995
rect 1673 20955 1731 20961
rect 5442 20952 5448 21004
rect 5500 20992 5506 21004
rect 5500 20964 5856 20992
rect 6012 20978 6040 21032
rect 15010 21020 15016 21072
rect 15068 21060 15074 21072
rect 15562 21060 15568 21072
rect 15068 21032 15568 21060
rect 15068 21020 15074 21032
rect 15562 21020 15568 21032
rect 15620 21020 15626 21072
rect 16114 21020 16120 21072
rect 16172 21020 16178 21072
rect 17328 21060 17356 21100
rect 17402 21088 17408 21140
rect 17460 21128 17466 21140
rect 17681 21131 17739 21137
rect 17681 21128 17693 21131
rect 17460 21100 17693 21128
rect 17460 21088 17466 21100
rect 17681 21097 17693 21100
rect 17727 21097 17739 21131
rect 17681 21091 17739 21097
rect 20165 21131 20223 21137
rect 20165 21097 20177 21131
rect 20211 21128 20223 21131
rect 20530 21128 20536 21140
rect 20211 21100 20536 21128
rect 20211 21097 20223 21100
rect 20165 21091 20223 21097
rect 20530 21088 20536 21100
rect 20588 21088 20594 21140
rect 20717 21131 20775 21137
rect 20717 21097 20729 21131
rect 20763 21128 20775 21131
rect 20806 21128 20812 21140
rect 20763 21100 20812 21128
rect 20763 21097 20775 21100
rect 20717 21091 20775 21097
rect 20806 21088 20812 21100
rect 20864 21088 20870 21140
rect 18782 21060 18788 21072
rect 17328 21032 18788 21060
rect 18782 21020 18788 21032
rect 18840 21020 18846 21072
rect 7742 20992 7748 21004
rect 5500 20952 5506 20964
rect 1946 20884 1952 20936
rect 2004 20924 2010 20936
rect 2317 20927 2375 20933
rect 2004 20920 2268 20924
rect 2317 20920 2329 20927
rect 2004 20896 2329 20920
rect 2004 20884 2010 20896
rect 2240 20893 2329 20896
rect 2363 20893 2375 20927
rect 2240 20892 2375 20893
rect 2317 20887 2375 20892
rect 2498 20884 2504 20936
rect 2556 20924 2562 20936
rect 2591 20927 2649 20933
rect 2591 20924 2603 20927
rect 2556 20896 2603 20924
rect 2556 20884 2562 20896
rect 2591 20893 2603 20896
rect 2637 20893 2649 20927
rect 3789 20927 3847 20933
rect 3789 20924 3801 20927
rect 2591 20887 2649 20893
rect 2746 20896 3801 20924
rect 1302 20816 1308 20868
rect 1360 20856 1366 20868
rect 2746 20856 2774 20896
rect 3789 20893 3801 20896
rect 3835 20893 3847 20927
rect 3789 20887 3847 20893
rect 4065 20927 4123 20933
rect 4065 20893 4077 20927
rect 4111 20924 4123 20927
rect 4246 20924 4252 20936
rect 4111 20896 4252 20924
rect 4111 20893 4123 20896
rect 4065 20887 4123 20893
rect 4246 20884 4252 20896
rect 4304 20884 4310 20936
rect 4339 20927 4397 20933
rect 4339 20893 4351 20927
rect 4385 20924 4397 20927
rect 5718 20924 5724 20936
rect 4385 20896 5724 20924
rect 4385 20893 4397 20896
rect 4339 20887 4397 20893
rect 5718 20884 5724 20896
rect 5776 20884 5782 20936
rect 1360 20828 2774 20856
rect 1360 20816 1366 20828
rect 2958 20816 2964 20868
rect 3016 20856 3022 20868
rect 4430 20856 4436 20868
rect 3016 20828 4436 20856
rect 3016 20816 3022 20828
rect 4430 20816 4436 20828
rect 4488 20816 4494 20868
rect 5828 20856 5856 20964
rect 7300 20964 7748 20992
rect 5902 20884 5908 20936
rect 5960 20924 5966 20936
rect 6549 20927 6607 20933
rect 6549 20924 6561 20927
rect 5960 20896 6561 20924
rect 5960 20884 5966 20896
rect 6549 20893 6561 20896
rect 6595 20893 6607 20927
rect 6549 20887 6607 20893
rect 6730 20884 6736 20936
rect 6788 20924 6794 20936
rect 6917 20927 6975 20933
rect 6917 20924 6929 20927
rect 6788 20896 6929 20924
rect 6788 20884 6794 20896
rect 6917 20893 6929 20896
rect 6963 20924 6975 20927
rect 7300 20924 7328 20964
rect 7742 20952 7748 20964
rect 7800 20952 7806 21004
rect 10042 20952 10048 21004
rect 10100 20992 10106 21004
rect 10502 20992 10508 21004
rect 10100 20964 10508 20992
rect 10100 20952 10106 20964
rect 10502 20952 10508 20964
rect 10560 20952 10566 21004
rect 13354 20952 13360 21004
rect 13412 20992 13418 21004
rect 13814 20992 13820 21004
rect 13412 20964 13820 20992
rect 13412 20952 13418 20964
rect 13814 20952 13820 20964
rect 13872 20992 13878 21004
rect 14090 20992 14096 21004
rect 13872 20964 14096 20992
rect 13872 20952 13878 20964
rect 14090 20952 14096 20964
rect 14148 20952 14154 21004
rect 16132 20992 16160 21020
rect 16669 20995 16727 21001
rect 16669 20992 16681 20995
rect 16132 20964 16681 20992
rect 16669 20961 16681 20964
rect 16715 20961 16727 20995
rect 16669 20955 16727 20961
rect 6963 20896 7328 20924
rect 6963 20893 6975 20896
rect 6917 20887 6975 20893
rect 7926 20884 7932 20936
rect 7984 20924 7990 20936
rect 8941 20927 8999 20933
rect 8941 20924 8953 20927
rect 7984 20896 8953 20924
rect 7984 20884 7990 20896
rect 8941 20893 8953 20896
rect 8987 20893 8999 20927
rect 8941 20887 8999 20893
rect 6457 20859 6515 20865
rect 5828 20828 6316 20856
rect 2130 20748 2136 20800
rect 2188 20788 2194 20800
rect 2498 20788 2504 20800
rect 2188 20760 2504 20788
rect 2188 20748 2194 20760
rect 2498 20748 2504 20760
rect 2556 20748 2562 20800
rect 2682 20748 2688 20800
rect 2740 20788 2746 20800
rect 3329 20791 3387 20797
rect 3329 20788 3341 20791
rect 2740 20760 3341 20788
rect 2740 20748 2746 20760
rect 3329 20757 3341 20760
rect 3375 20757 3387 20791
rect 3329 20751 3387 20757
rect 3418 20748 3424 20800
rect 3476 20788 3482 20800
rect 4522 20788 4528 20800
rect 3476 20760 4528 20788
rect 3476 20748 3482 20760
rect 4522 20748 4528 20760
rect 4580 20748 4586 20800
rect 4890 20748 4896 20800
rect 4948 20788 4954 20800
rect 5166 20788 5172 20800
rect 4948 20760 5172 20788
rect 4948 20748 4954 20760
rect 5166 20748 5172 20760
rect 5224 20748 5230 20800
rect 6178 20748 6184 20800
rect 6236 20748 6242 20800
rect 6288 20788 6316 20828
rect 6457 20825 6469 20859
rect 6503 20856 6515 20859
rect 6822 20856 6828 20868
rect 6503 20828 6828 20856
rect 6503 20825 6515 20828
rect 6457 20819 6515 20825
rect 6822 20816 6828 20828
rect 6880 20816 6886 20868
rect 8956 20856 8984 20887
rect 9122 20884 9128 20936
rect 9180 20924 9186 20936
rect 9215 20927 9273 20933
rect 9215 20924 9227 20927
rect 9180 20896 9227 20924
rect 9180 20884 9186 20896
rect 9215 20893 9227 20896
rect 9261 20893 9273 20927
rect 9215 20887 9273 20893
rect 9582 20884 9588 20936
rect 9640 20884 9646 20936
rect 10594 20884 10600 20936
rect 10652 20924 10658 20936
rect 11241 20927 11299 20933
rect 11241 20924 11253 20927
rect 10652 20896 11253 20924
rect 10652 20884 10658 20896
rect 11241 20893 11253 20896
rect 11287 20893 11299 20927
rect 11241 20887 11299 20893
rect 9600 20856 9628 20884
rect 6930 20828 7512 20856
rect 8956 20828 9628 20856
rect 6930 20788 6958 20828
rect 6288 20760 6958 20788
rect 7098 20748 7104 20800
rect 7156 20788 7162 20800
rect 7484 20797 7512 20828
rect 7285 20791 7343 20797
rect 7285 20788 7297 20791
rect 7156 20760 7297 20788
rect 7156 20748 7162 20760
rect 7285 20757 7297 20760
rect 7331 20757 7343 20791
rect 7285 20751 7343 20757
rect 7469 20791 7527 20797
rect 7469 20757 7481 20791
rect 7515 20757 7527 20791
rect 7469 20751 7527 20757
rect 9490 20748 9496 20800
rect 9548 20788 9554 20800
rect 10318 20788 10324 20800
rect 9548 20760 10324 20788
rect 9548 20748 9554 20760
rect 10318 20748 10324 20760
rect 10376 20748 10382 20800
rect 11256 20788 11284 20887
rect 11422 20884 11428 20936
rect 11480 20924 11486 20936
rect 11515 20927 11573 20933
rect 11515 20924 11527 20927
rect 11480 20896 11527 20924
rect 11480 20884 11486 20896
rect 11515 20893 11527 20896
rect 11561 20924 11573 20927
rect 12618 20924 12624 20936
rect 11561 20896 12624 20924
rect 11561 20893 11573 20896
rect 11515 20887 11573 20893
rect 12618 20884 12624 20896
rect 12676 20884 12682 20936
rect 14335 20927 14393 20933
rect 14335 20893 14347 20927
rect 14381 20893 14393 20927
rect 14335 20887 14393 20893
rect 11790 20816 11796 20868
rect 11848 20856 11854 20868
rect 14350 20856 14378 20887
rect 16022 20884 16028 20936
rect 16080 20884 16086 20936
rect 16117 20927 16175 20933
rect 16117 20893 16129 20927
rect 16163 20893 16175 20927
rect 16117 20887 16175 20893
rect 15657 20859 15715 20865
rect 15657 20856 15669 20859
rect 11848 20828 14412 20856
rect 11848 20816 11854 20828
rect 13906 20788 13912 20800
rect 11256 20760 13912 20788
rect 13906 20748 13912 20760
rect 13964 20748 13970 20800
rect 14384 20788 14412 20828
rect 14568 20828 15669 20856
rect 14568 20788 14596 20828
rect 15657 20825 15669 20828
rect 15703 20825 15715 20859
rect 15657 20819 15715 20825
rect 16132 20800 16160 20887
rect 16206 20884 16212 20936
rect 16264 20924 16270 20936
rect 16301 20927 16359 20933
rect 16301 20924 16313 20927
rect 16264 20896 16313 20924
rect 16264 20884 16270 20896
rect 16301 20893 16313 20896
rect 16347 20893 16359 20927
rect 16301 20887 16359 20893
rect 14384 20760 14596 20788
rect 14918 20748 14924 20800
rect 14976 20788 14982 20800
rect 15105 20791 15163 20797
rect 15105 20788 15117 20791
rect 14976 20760 15117 20788
rect 14976 20748 14982 20760
rect 15105 20757 15117 20760
rect 15151 20757 15163 20791
rect 15105 20751 15163 20757
rect 15838 20748 15844 20800
rect 15896 20748 15902 20800
rect 16114 20748 16120 20800
rect 16172 20748 16178 20800
rect 16298 20748 16304 20800
rect 16356 20748 16362 20800
rect 16684 20788 16712 20955
rect 18598 20952 18604 21004
rect 18656 20992 18662 21004
rect 20346 20992 20352 21004
rect 18656 20964 20352 20992
rect 18656 20952 18662 20964
rect 20346 20952 20352 20964
rect 20404 20952 20410 21004
rect 22646 20952 22652 21004
rect 22704 20992 22710 21004
rect 22704 20964 22968 20992
rect 22704 20952 22710 20964
rect 16943 20927 17001 20933
rect 16943 20893 16955 20927
rect 16989 20924 17001 20927
rect 17034 20924 17040 20936
rect 16989 20896 17040 20924
rect 16989 20893 17001 20896
rect 16943 20887 17001 20893
rect 17034 20884 17040 20896
rect 17092 20924 17098 20936
rect 17954 20924 17960 20936
rect 17092 20896 17960 20924
rect 17092 20884 17098 20896
rect 17954 20884 17960 20896
rect 18012 20884 18018 20936
rect 20073 20927 20131 20933
rect 20073 20893 20085 20927
rect 20119 20924 20131 20927
rect 21266 20924 21272 20936
rect 20119 20896 21272 20924
rect 20119 20893 20131 20896
rect 20073 20887 20131 20893
rect 21266 20884 21272 20896
rect 21324 20884 21330 20936
rect 17218 20816 17224 20868
rect 17276 20856 17282 20868
rect 18874 20856 18880 20868
rect 17276 20828 18880 20856
rect 17276 20816 17282 20828
rect 18874 20816 18880 20828
rect 18932 20816 18938 20868
rect 20441 20859 20499 20865
rect 20441 20825 20453 20859
rect 20487 20856 20499 20859
rect 20622 20856 20628 20868
rect 20487 20828 20628 20856
rect 20487 20825 20499 20828
rect 20441 20819 20499 20825
rect 20622 20816 20628 20828
rect 20680 20816 20686 20868
rect 20993 20859 21051 20865
rect 20993 20825 21005 20859
rect 21039 20825 21051 20859
rect 20993 20819 21051 20825
rect 21361 20859 21419 20865
rect 21361 20825 21373 20859
rect 21407 20856 21419 20859
rect 22186 20856 22192 20868
rect 21407 20828 22192 20856
rect 21407 20825 21419 20828
rect 21361 20819 21419 20825
rect 17586 20788 17592 20800
rect 16684 20760 17592 20788
rect 17586 20748 17592 20760
rect 17644 20748 17650 20800
rect 21008 20788 21036 20819
rect 22186 20816 22192 20828
rect 22244 20816 22250 20868
rect 21450 20788 21456 20800
rect 21008 20760 21456 20788
rect 21450 20748 21456 20760
rect 21508 20748 21514 20800
rect 1104 20698 22056 20720
rect 1104 20646 6148 20698
rect 6200 20646 6212 20698
rect 6264 20646 6276 20698
rect 6328 20646 6340 20698
rect 6392 20646 6404 20698
rect 6456 20646 11346 20698
rect 11398 20646 11410 20698
rect 11462 20646 11474 20698
rect 11526 20646 11538 20698
rect 11590 20646 11602 20698
rect 11654 20646 16544 20698
rect 16596 20646 16608 20698
rect 16660 20646 16672 20698
rect 16724 20646 16736 20698
rect 16788 20646 16800 20698
rect 16852 20646 21742 20698
rect 21794 20646 21806 20698
rect 21858 20646 21870 20698
rect 21922 20646 21934 20698
rect 21986 20646 21998 20698
rect 22050 20646 22056 20698
rect 22940 20664 22968 20964
rect 1104 20624 22056 20646
rect 22922 20612 22928 20664
rect 22980 20612 22986 20664
rect 934 20544 940 20596
rect 992 20584 998 20596
rect 1302 20584 1308 20596
rect 992 20556 1308 20584
rect 992 20544 998 20556
rect 1302 20544 1308 20556
rect 1360 20544 1366 20596
rect 2314 20544 2320 20596
rect 2372 20544 2378 20596
rect 3973 20587 4031 20593
rect 2424 20556 3554 20584
rect 1397 20451 1455 20457
rect 1397 20417 1409 20451
rect 1443 20448 1455 20451
rect 1486 20448 1492 20460
rect 1443 20420 1492 20448
rect 1443 20417 1455 20420
rect 1397 20411 1455 20417
rect 1486 20408 1492 20420
rect 1544 20408 1550 20460
rect 2041 20451 2099 20457
rect 2041 20417 2053 20451
rect 2087 20448 2099 20451
rect 2424 20448 2452 20556
rect 2498 20476 2504 20528
rect 2556 20516 2562 20528
rect 2593 20519 2651 20525
rect 2593 20516 2605 20519
rect 2556 20488 2605 20516
rect 2556 20476 2562 20488
rect 2593 20485 2605 20488
rect 2639 20516 2651 20519
rect 3142 20516 3148 20528
rect 2639 20488 3148 20516
rect 2639 20485 2651 20488
rect 2593 20479 2651 20485
rect 3142 20476 3148 20488
rect 3200 20476 3206 20528
rect 3326 20476 3332 20528
rect 3384 20516 3390 20528
rect 3421 20519 3479 20525
rect 3421 20516 3433 20519
rect 3384 20488 3433 20516
rect 3384 20476 3390 20488
rect 3421 20485 3433 20488
rect 3467 20485 3479 20519
rect 3526 20516 3554 20556
rect 3973 20553 3985 20587
rect 4019 20584 4031 20587
rect 4154 20584 4160 20596
rect 4019 20556 4160 20584
rect 4019 20553 4031 20556
rect 3973 20547 4031 20553
rect 4154 20544 4160 20556
rect 4212 20544 4218 20596
rect 4338 20544 4344 20596
rect 4396 20544 4402 20596
rect 4522 20544 4528 20596
rect 4580 20584 4586 20596
rect 5077 20587 5135 20593
rect 5077 20584 5089 20587
rect 4580 20556 5089 20584
rect 4580 20544 4586 20556
rect 5077 20553 5089 20556
rect 5123 20553 5135 20587
rect 6822 20584 6828 20596
rect 5077 20547 5135 20553
rect 5552 20556 6828 20584
rect 4249 20519 4307 20525
rect 4249 20516 4261 20519
rect 3526 20488 4261 20516
rect 3421 20479 3479 20485
rect 4249 20485 4261 20488
rect 4295 20485 4307 20519
rect 4356 20516 4384 20544
rect 5552 20525 5580 20556
rect 6822 20544 6828 20556
rect 6880 20544 6886 20596
rect 7926 20584 7932 20596
rect 6930 20556 7932 20584
rect 4709 20519 4767 20525
rect 4709 20516 4721 20519
rect 4356 20488 4721 20516
rect 4249 20479 4307 20485
rect 4709 20485 4721 20488
rect 4755 20485 4767 20519
rect 4709 20479 4767 20485
rect 5537 20519 5595 20525
rect 5537 20485 5549 20519
rect 5583 20485 5595 20519
rect 5537 20479 5595 20485
rect 5721 20519 5779 20525
rect 5721 20485 5733 20519
rect 5767 20516 5779 20519
rect 6454 20516 6460 20528
rect 5767 20488 6460 20516
rect 5767 20485 5779 20488
rect 5721 20479 5779 20485
rect 6454 20476 6460 20488
rect 6512 20476 6518 20528
rect 6546 20476 6552 20528
rect 6604 20516 6610 20528
rect 6730 20516 6736 20528
rect 6604 20488 6736 20516
rect 6604 20476 6610 20488
rect 6730 20476 6736 20488
rect 6788 20476 6794 20528
rect 2087 20420 2452 20448
rect 2087 20417 2099 20420
rect 2041 20411 2099 20417
rect 2682 20408 2688 20460
rect 2740 20408 2746 20460
rect 2866 20408 2872 20460
rect 2924 20448 2930 20460
rect 3053 20451 3111 20457
rect 3053 20448 3065 20451
rect 2924 20420 3065 20448
rect 2924 20408 2930 20420
rect 3053 20417 3065 20420
rect 3099 20417 3111 20451
rect 3053 20411 3111 20417
rect 4341 20451 4399 20457
rect 4341 20417 4353 20451
rect 4387 20448 4399 20451
rect 4430 20448 4436 20460
rect 4387 20420 4436 20448
rect 4387 20417 4399 20420
rect 4341 20411 4399 20417
rect 4430 20408 4436 20420
rect 4488 20408 4494 20460
rect 4522 20408 4528 20460
rect 4580 20448 4586 20460
rect 5442 20448 5448 20460
rect 4580 20420 5448 20448
rect 4580 20408 4586 20420
rect 5442 20408 5448 20420
rect 5500 20448 5506 20460
rect 6930 20448 6958 20556
rect 7926 20544 7932 20556
rect 7984 20544 7990 20596
rect 8018 20544 8024 20596
rect 8076 20584 8082 20596
rect 8076 20556 8432 20584
rect 8076 20544 8082 20556
rect 7561 20519 7619 20525
rect 7561 20485 7573 20519
rect 7607 20516 7619 20519
rect 7650 20516 7656 20528
rect 7607 20488 7656 20516
rect 7607 20485 7619 20488
rect 7561 20479 7619 20485
rect 7650 20476 7656 20488
rect 7708 20476 7714 20528
rect 7834 20476 7840 20528
rect 7892 20476 7898 20528
rect 8294 20476 8300 20528
rect 8352 20476 8358 20528
rect 8404 20516 8432 20556
rect 8570 20544 8576 20596
rect 8628 20584 8634 20596
rect 9398 20584 9404 20596
rect 8628 20556 9404 20584
rect 8628 20544 8634 20556
rect 9398 20544 9404 20556
rect 9456 20584 9462 20596
rect 12894 20584 12900 20596
rect 9456 20556 10088 20584
rect 9456 20544 9462 20556
rect 8665 20519 8723 20525
rect 8665 20516 8677 20519
rect 8404 20488 8677 20516
rect 8665 20485 8677 20488
rect 8711 20516 8723 20519
rect 9214 20516 9220 20528
rect 8711 20488 9220 20516
rect 8711 20485 8723 20488
rect 8665 20479 8723 20485
rect 9214 20476 9220 20488
rect 9272 20476 9278 20528
rect 5500 20420 6958 20448
rect 5500 20408 5506 20420
rect 7926 20408 7932 20460
rect 7984 20408 7990 20460
rect 10060 20457 10088 20556
rect 11790 20556 12900 20584
rect 11790 20487 11818 20556
rect 12894 20544 12900 20556
rect 12952 20584 12958 20596
rect 13078 20584 13084 20596
rect 12952 20556 13084 20584
rect 12952 20544 12958 20556
rect 13078 20544 13084 20556
rect 13136 20544 13142 20596
rect 13170 20544 13176 20596
rect 13228 20544 13234 20596
rect 14090 20544 14096 20596
rect 14148 20584 14154 20596
rect 14148 20556 14872 20584
rect 14148 20544 14154 20556
rect 11775 20481 11833 20487
rect 10045 20451 10103 20457
rect 10045 20417 10057 20451
rect 10091 20417 10103 20451
rect 10045 20411 10103 20417
rect 10318 20408 10324 20460
rect 10376 20448 10382 20460
rect 11422 20448 11428 20460
rect 10376 20420 11428 20448
rect 10376 20408 10382 20420
rect 11422 20408 11428 20420
rect 11480 20408 11486 20460
rect 11775 20447 11787 20481
rect 11821 20447 11833 20481
rect 11775 20441 11833 20447
rect 12802 20408 12808 20460
rect 12860 20408 12866 20460
rect 12894 20408 12900 20460
rect 12952 20448 12958 20460
rect 13188 20448 13216 20544
rect 13265 20451 13323 20457
rect 13265 20448 13277 20451
rect 12952 20420 13277 20448
rect 12952 20408 12958 20420
rect 13265 20417 13277 20420
rect 13311 20417 13323 20451
rect 14844 20448 14872 20556
rect 15562 20544 15568 20596
rect 15620 20584 15626 20596
rect 17773 20587 17831 20593
rect 15620 20556 15792 20584
rect 15620 20544 15626 20556
rect 14921 20519 14979 20525
rect 14921 20485 14933 20519
rect 14967 20516 14979 20519
rect 15654 20516 15660 20528
rect 14967 20488 15660 20516
rect 14967 20485 14979 20488
rect 14921 20479 14979 20485
rect 15654 20476 15660 20488
rect 15712 20476 15718 20528
rect 15013 20451 15071 20457
rect 15013 20448 15025 20451
rect 14844 20420 15025 20448
rect 13265 20411 13323 20417
rect 15013 20417 15025 20420
rect 15059 20417 15071 20451
rect 15013 20411 15071 20417
rect 15194 20408 15200 20460
rect 15252 20448 15258 20460
rect 15287 20451 15345 20457
rect 15287 20448 15299 20451
rect 15252 20420 15299 20448
rect 15252 20408 15258 20420
rect 15287 20417 15299 20420
rect 15333 20448 15345 20451
rect 15764 20448 15792 20556
rect 17773 20553 17785 20587
rect 17819 20584 17831 20587
rect 17862 20584 17868 20596
rect 17819 20556 17868 20584
rect 17819 20553 17831 20556
rect 17773 20547 17831 20553
rect 17862 20544 17868 20556
rect 17920 20544 17926 20596
rect 19245 20587 19303 20593
rect 19245 20553 19257 20587
rect 19291 20584 19303 20587
rect 20806 20584 20812 20596
rect 19291 20556 20812 20584
rect 19291 20553 19303 20556
rect 19245 20547 19303 20553
rect 20806 20544 20812 20556
rect 20864 20544 20870 20596
rect 21174 20544 21180 20596
rect 21232 20544 21238 20596
rect 15930 20476 15936 20528
rect 15988 20516 15994 20528
rect 21192 20516 21220 20544
rect 15988 20488 17046 20516
rect 21192 20488 21312 20516
rect 15988 20476 15994 20488
rect 17018 20457 17046 20488
rect 19779 20481 19837 20487
rect 15333 20420 15792 20448
rect 17003 20451 17061 20457
rect 15333 20417 15345 20420
rect 15287 20411 15345 20417
rect 17003 20417 17015 20451
rect 17049 20417 17061 20451
rect 17003 20411 17061 20417
rect 19429 20451 19487 20457
rect 19429 20417 19441 20451
rect 19475 20417 19487 20451
rect 19779 20447 19791 20481
rect 19825 20478 19837 20481
rect 19825 20448 19840 20478
rect 20162 20448 20168 20460
rect 19825 20447 20168 20448
rect 19779 20441 20168 20447
rect 19812 20420 20168 20441
rect 19429 20411 19487 20417
rect 2498 20340 2504 20392
rect 2556 20340 2562 20392
rect 3878 20340 3884 20392
rect 3936 20340 3942 20392
rect 5350 20340 5356 20392
rect 5408 20380 5414 20392
rect 6914 20380 6920 20392
rect 5408 20352 6920 20380
rect 5408 20340 5414 20352
rect 6914 20340 6920 20352
rect 6972 20340 6978 20392
rect 7006 20340 7012 20392
rect 7064 20340 7070 20392
rect 7098 20340 7104 20392
rect 7156 20380 7162 20392
rect 11514 20380 11520 20392
rect 7156 20352 7406 20380
rect 10704 20352 11520 20380
rect 7156 20340 7162 20352
rect 1578 20272 1584 20324
rect 1636 20272 1642 20324
rect 5718 20272 5724 20324
rect 5776 20312 5782 20324
rect 6454 20312 6460 20324
rect 5776 20284 6460 20312
rect 5776 20272 5782 20284
rect 6454 20272 6460 20284
rect 6512 20272 6518 20324
rect 6546 20272 6552 20324
rect 6604 20312 6610 20324
rect 7024 20312 7052 20340
rect 6604 20284 7052 20312
rect 6604 20272 6610 20284
rect 3510 20204 3516 20256
rect 3568 20244 3574 20256
rect 3605 20247 3663 20253
rect 3605 20244 3617 20247
rect 3568 20216 3617 20244
rect 3568 20204 3574 20216
rect 3605 20213 3617 20216
rect 3651 20213 3663 20247
rect 3605 20207 3663 20213
rect 5258 20204 5264 20256
rect 5316 20204 5322 20256
rect 6638 20204 6644 20256
rect 6696 20204 6702 20256
rect 8849 20247 8907 20253
rect 8849 20213 8861 20247
rect 8895 20244 8907 20247
rect 9122 20244 9128 20256
rect 8895 20216 9128 20244
rect 8895 20213 8907 20216
rect 8849 20207 8907 20213
rect 9122 20204 9128 20216
rect 9180 20204 9186 20256
rect 9858 20204 9864 20256
rect 9916 20244 9922 20256
rect 10704 20244 10732 20352
rect 11514 20340 11520 20352
rect 11572 20340 11578 20392
rect 12820 20380 12848 20408
rect 13081 20383 13139 20389
rect 13081 20380 13093 20383
rect 12820 20352 13093 20380
rect 13081 20349 13093 20352
rect 13127 20380 13139 20383
rect 13170 20380 13176 20392
rect 13127 20352 13176 20380
rect 13127 20349 13139 20352
rect 13081 20343 13139 20349
rect 13170 20340 13176 20352
rect 13228 20340 13234 20392
rect 14001 20383 14059 20389
rect 14001 20380 14013 20383
rect 13372 20352 14013 20380
rect 10962 20272 10968 20324
rect 11020 20312 11026 20324
rect 11330 20312 11336 20324
rect 11020 20284 11336 20312
rect 11020 20272 11026 20284
rect 11330 20272 11336 20284
rect 11388 20272 11394 20324
rect 13372 20312 13400 20352
rect 14001 20349 14013 20352
rect 14047 20349 14059 20383
rect 14001 20343 14059 20349
rect 14136 20340 14142 20392
rect 14194 20340 14200 20392
rect 14277 20383 14335 20389
rect 14277 20349 14289 20383
rect 14323 20380 14335 20383
rect 14918 20380 14924 20392
rect 14323 20352 14924 20380
rect 14323 20349 14335 20352
rect 14277 20343 14335 20349
rect 14918 20340 14924 20352
rect 14976 20340 14982 20392
rect 16761 20383 16819 20389
rect 16761 20349 16773 20383
rect 16807 20349 16819 20383
rect 16761 20343 16819 20349
rect 12406 20284 13400 20312
rect 9916 20216 10732 20244
rect 9916 20204 9922 20216
rect 11054 20204 11060 20256
rect 11112 20204 11118 20256
rect 11238 20204 11244 20256
rect 11296 20244 11302 20256
rect 12406 20244 12434 20284
rect 13722 20272 13728 20324
rect 13780 20272 13786 20324
rect 11296 20216 12434 20244
rect 12529 20247 12587 20253
rect 11296 20204 11302 20216
rect 12529 20213 12541 20247
rect 12575 20244 12587 20247
rect 12618 20244 12624 20256
rect 12575 20216 12624 20244
rect 12575 20213 12587 20216
rect 12529 20207 12587 20213
rect 12618 20204 12624 20216
rect 12676 20204 12682 20256
rect 14936 20244 14964 20340
rect 15378 20244 15384 20256
rect 14936 20216 15384 20244
rect 15378 20204 15384 20216
rect 15436 20204 15442 20256
rect 16025 20247 16083 20253
rect 16025 20213 16037 20247
rect 16071 20244 16083 20247
rect 16114 20244 16120 20256
rect 16071 20216 16120 20244
rect 16071 20213 16083 20216
rect 16025 20207 16083 20213
rect 16114 20204 16120 20216
rect 16172 20204 16178 20256
rect 16776 20244 16804 20343
rect 17586 20340 17592 20392
rect 17644 20340 17650 20392
rect 17604 20244 17632 20340
rect 16776 20216 17632 20244
rect 19444 20244 19472 20411
rect 20162 20408 20168 20420
rect 20220 20408 20226 20460
rect 20990 20408 20996 20460
rect 21048 20448 21054 20460
rect 21284 20457 21312 20488
rect 21177 20451 21235 20457
rect 21177 20448 21189 20451
rect 21048 20420 21189 20448
rect 21048 20408 21054 20420
rect 21177 20417 21189 20420
rect 21223 20417 21235 20451
rect 21177 20411 21235 20417
rect 21269 20451 21327 20457
rect 21269 20417 21281 20451
rect 21315 20417 21327 20451
rect 21269 20411 21327 20417
rect 19518 20340 19524 20392
rect 19576 20340 19582 20392
rect 19978 20244 19984 20256
rect 19444 20216 19984 20244
rect 19978 20204 19984 20216
rect 20036 20204 20042 20256
rect 20530 20204 20536 20256
rect 20588 20204 20594 20256
rect 20993 20247 21051 20253
rect 20993 20213 21005 20247
rect 21039 20244 21051 20247
rect 21174 20244 21180 20256
rect 21039 20216 21180 20244
rect 21039 20213 21051 20216
rect 20993 20207 21051 20213
rect 21174 20204 21180 20216
rect 21232 20204 21238 20256
rect 21450 20204 21456 20256
rect 21508 20204 21514 20256
rect 1104 20154 21896 20176
rect 1104 20102 3549 20154
rect 3601 20102 3613 20154
rect 3665 20102 3677 20154
rect 3729 20102 3741 20154
rect 3793 20102 3805 20154
rect 3857 20102 8747 20154
rect 8799 20102 8811 20154
rect 8863 20102 8875 20154
rect 8927 20102 8939 20154
rect 8991 20102 9003 20154
rect 9055 20102 13945 20154
rect 13997 20102 14009 20154
rect 14061 20102 14073 20154
rect 14125 20102 14137 20154
rect 14189 20102 14201 20154
rect 14253 20102 19143 20154
rect 19195 20102 19207 20154
rect 19259 20102 19271 20154
rect 19323 20102 19335 20154
rect 19387 20102 19399 20154
rect 19451 20102 21896 20154
rect 1104 20080 21896 20102
rect 750 20040 756 20052
rect 676 20012 756 20040
rect 676 19576 704 20012
rect 750 20000 756 20012
rect 808 20000 814 20052
rect 1581 20043 1639 20049
rect 1581 20009 1593 20043
rect 1627 20040 1639 20043
rect 1762 20040 1768 20052
rect 1627 20012 1768 20040
rect 1627 20009 1639 20012
rect 1581 20003 1639 20009
rect 1762 20000 1768 20012
rect 1820 20000 1826 20052
rect 2774 20000 2780 20052
rect 2832 20040 2838 20052
rect 3329 20043 3387 20049
rect 2832 20012 3280 20040
rect 2832 20000 2838 20012
rect 2038 19932 2044 19984
rect 2096 19932 2102 19984
rect 3252 19972 3280 20012
rect 3329 20009 3341 20043
rect 3375 20040 3387 20043
rect 4430 20040 4436 20052
rect 3375 20012 4436 20040
rect 3375 20009 3387 20012
rect 3329 20003 3387 20009
rect 4430 20000 4436 20012
rect 4488 20000 4494 20052
rect 5350 20040 5356 20052
rect 4632 20012 5356 20040
rect 3973 19975 4031 19981
rect 3973 19972 3985 19975
rect 3252 19944 3985 19972
rect 3973 19941 3985 19944
rect 4019 19972 4031 19975
rect 4632 19972 4660 20012
rect 5350 20000 5356 20012
rect 5408 20000 5414 20052
rect 5718 20000 5724 20052
rect 5776 20040 5782 20052
rect 6086 20040 6092 20052
rect 5776 20012 6092 20040
rect 5776 20000 5782 20012
rect 6086 20000 6092 20012
rect 6144 20000 6150 20052
rect 8202 20000 8208 20052
rect 8260 20040 8266 20052
rect 8662 20040 8668 20052
rect 8260 20012 8668 20040
rect 8260 20000 8266 20012
rect 8662 20000 8668 20012
rect 8720 20000 8726 20052
rect 11146 20000 11152 20052
rect 11204 20040 11210 20052
rect 11241 20043 11299 20049
rect 11241 20040 11253 20043
rect 11204 20012 11253 20040
rect 11204 20000 11210 20012
rect 11241 20009 11253 20012
rect 11287 20009 11299 20043
rect 11241 20003 11299 20009
rect 11330 20000 11336 20052
rect 11388 20000 11394 20052
rect 11514 20000 11520 20052
rect 11572 20040 11578 20052
rect 13354 20040 13360 20052
rect 11572 20012 13360 20040
rect 11572 20000 11578 20012
rect 4019 19944 4660 19972
rect 5537 19975 5595 19981
rect 4019 19941 4031 19944
rect 3973 19935 4031 19941
rect 5537 19941 5549 19975
rect 5583 19972 5595 19975
rect 5583 19944 5948 19972
rect 5583 19941 5595 19944
rect 5537 19935 5595 19941
rect 1210 19864 1216 19916
rect 1268 19904 1274 19916
rect 2314 19904 2320 19916
rect 1268 19876 2320 19904
rect 1268 19864 1274 19876
rect 2314 19864 2320 19876
rect 2372 19864 2378 19916
rect 3234 19864 3240 19916
rect 3292 19904 3298 19916
rect 4522 19904 4528 19916
rect 3292 19876 4528 19904
rect 3292 19864 3298 19876
rect 4522 19864 4528 19876
rect 4580 19864 4586 19916
rect 5920 19890 5948 19944
rect 10410 19864 10416 19916
rect 10468 19864 10474 19916
rect 11054 19864 11060 19916
rect 11112 19864 11118 19916
rect 750 19796 756 19848
rect 808 19836 814 19848
rect 1489 19839 1547 19845
rect 1489 19836 1501 19839
rect 808 19808 1501 19836
rect 808 19796 814 19808
rect 1489 19805 1501 19808
rect 1535 19805 1547 19839
rect 1489 19799 1547 19805
rect 1762 19796 1768 19848
rect 1820 19836 1826 19848
rect 3789 19839 3847 19845
rect 1820 19808 2360 19836
rect 3789 19832 3801 19839
rect 1820 19796 1826 19808
rect 2332 19780 2360 19808
rect 2575 19809 2633 19815
rect 2575 19806 2587 19809
rect 1854 19728 1860 19780
rect 1912 19728 1918 19780
rect 2314 19728 2320 19780
rect 2372 19768 2378 19780
rect 2574 19775 2587 19806
rect 2621 19775 2633 19809
rect 3786 19805 3801 19832
rect 3835 19805 3847 19839
rect 3786 19799 3847 19805
rect 2574 19769 2633 19775
rect 2574 19768 2602 19769
rect 2372 19740 2602 19768
rect 2372 19728 2378 19740
rect 2774 19728 2780 19780
rect 2832 19768 2838 19780
rect 3786 19768 3814 19799
rect 4430 19796 4436 19848
rect 4488 19836 4494 19848
rect 4767 19839 4825 19845
rect 4767 19836 4779 19839
rect 4488 19808 4779 19836
rect 4488 19796 4494 19808
rect 4767 19805 4779 19808
rect 4813 19805 4825 19839
rect 4767 19799 4825 19805
rect 6365 19839 6423 19845
rect 6365 19805 6377 19839
rect 6411 19836 6423 19839
rect 6638 19836 6644 19848
rect 6411 19808 6644 19836
rect 6411 19805 6423 19808
rect 6365 19799 6423 19805
rect 6638 19796 6644 19808
rect 6696 19796 6702 19848
rect 6914 19796 6920 19848
rect 6972 19796 6978 19848
rect 10134 19796 10140 19848
rect 10192 19836 10198 19848
rect 10229 19839 10287 19845
rect 10229 19836 10241 19839
rect 10192 19808 10241 19836
rect 10192 19796 10198 19808
rect 10229 19805 10241 19808
rect 10275 19805 10287 19839
rect 10229 19799 10287 19805
rect 10321 19839 10379 19845
rect 10321 19805 10333 19839
rect 10367 19836 10379 19839
rect 11072 19836 11100 19864
rect 10367 19808 11100 19836
rect 11348 19836 11376 20000
rect 12636 19913 12664 20012
rect 13354 20000 13360 20012
rect 13412 20000 13418 20052
rect 15378 20000 15384 20052
rect 15436 20040 15442 20052
rect 15933 20043 15991 20049
rect 15436 20012 15700 20040
rect 15436 20000 15442 20012
rect 13633 19975 13691 19981
rect 13633 19941 13645 19975
rect 13679 19972 13691 19975
rect 13722 19972 13728 19984
rect 13679 19944 13728 19972
rect 13679 19941 13691 19944
rect 13633 19935 13691 19941
rect 13722 19932 13728 19944
rect 13780 19972 13786 19984
rect 14737 19975 14795 19981
rect 14737 19972 14749 19975
rect 13780 19944 14749 19972
rect 13780 19932 13786 19944
rect 14737 19941 14749 19944
rect 14783 19941 14795 19975
rect 14737 19935 14795 19941
rect 12621 19907 12679 19913
rect 12621 19873 12633 19907
rect 12667 19873 12679 19907
rect 12621 19867 12679 19873
rect 14093 19907 14151 19913
rect 14093 19873 14105 19907
rect 14139 19904 14151 19907
rect 14458 19904 14464 19916
rect 14139 19876 14464 19904
rect 14139 19873 14151 19876
rect 14093 19867 14151 19873
rect 14458 19864 14464 19876
rect 14516 19864 14522 19916
rect 14642 19864 14648 19916
rect 14700 19904 14706 19916
rect 14826 19904 14832 19916
rect 14700 19876 14832 19904
rect 14700 19864 14706 19876
rect 14826 19864 14832 19876
rect 14884 19904 14890 19916
rect 15013 19907 15071 19913
rect 15013 19904 15025 19907
rect 14884 19876 15025 19904
rect 14884 19864 14890 19876
rect 15013 19873 15025 19876
rect 15059 19873 15071 19907
rect 15013 19867 15071 19873
rect 15102 19864 15108 19916
rect 15160 19913 15166 19916
rect 15160 19907 15188 19913
rect 15176 19873 15188 19907
rect 15160 19867 15188 19873
rect 15289 19907 15347 19913
rect 15289 19873 15301 19907
rect 15335 19904 15347 19907
rect 15672 19904 15700 20012
rect 15933 20009 15945 20043
rect 15979 20040 15991 20043
rect 16022 20040 16028 20052
rect 15979 20012 16028 20040
rect 15979 20009 15991 20012
rect 15933 20003 15991 20009
rect 16022 20000 16028 20012
rect 16080 20000 16086 20052
rect 19978 20000 19984 20052
rect 20036 20040 20042 20052
rect 20625 20043 20683 20049
rect 20625 20040 20637 20043
rect 20036 20012 20637 20040
rect 20036 20000 20042 20012
rect 20625 20009 20637 20012
rect 20671 20009 20683 20043
rect 20625 20003 20683 20009
rect 17497 19975 17555 19981
rect 17497 19972 17509 19975
rect 17328 19944 17509 19972
rect 17328 19916 17356 19944
rect 17497 19941 17509 19944
rect 17543 19941 17555 19975
rect 17497 19935 17555 19941
rect 15335 19876 15700 19904
rect 15335 19873 15347 19876
rect 15289 19867 15347 19873
rect 15160 19864 15166 19867
rect 16942 19864 16948 19916
rect 17000 19864 17006 19916
rect 17310 19864 17316 19916
rect 17368 19864 17374 19916
rect 19245 19907 19303 19913
rect 19245 19904 19257 19907
rect 18984 19876 19257 19904
rect 18984 19848 19012 19876
rect 19245 19873 19257 19876
rect 19291 19873 19303 19907
rect 19245 19867 19303 19873
rect 20346 19864 20352 19916
rect 20404 19904 20410 19916
rect 20404 19876 21312 19904
rect 20404 19864 20410 19876
rect 11517 19839 11575 19845
rect 11517 19836 11529 19839
rect 11348 19808 11529 19836
rect 10367 19805 10379 19808
rect 10321 19799 10379 19805
rect 11517 19805 11529 19808
rect 11563 19805 11575 19839
rect 11517 19799 11575 19805
rect 12066 19796 12072 19848
rect 12124 19836 12130 19848
rect 12124 19815 12922 19836
rect 12124 19809 12937 19815
rect 12124 19808 12891 19809
rect 12124 19796 12130 19808
rect 6043 19771 6101 19777
rect 6043 19768 6055 19771
rect 2832 19740 3814 19768
rect 4080 19740 6055 19768
rect 2832 19728 2838 19740
rect 750 19660 756 19712
rect 808 19700 814 19712
rect 3050 19700 3056 19712
rect 808 19672 3056 19700
rect 808 19660 814 19672
rect 3050 19660 3056 19672
rect 3108 19660 3114 19712
rect 3142 19660 3148 19712
rect 3200 19700 3206 19712
rect 4080 19700 4108 19740
rect 6043 19737 6055 19740
rect 6089 19737 6101 19771
rect 6043 19731 6101 19737
rect 6178 19728 6184 19780
rect 6236 19768 6242 19780
rect 6457 19771 6515 19777
rect 6457 19768 6469 19771
rect 6236 19740 6469 19768
rect 6236 19728 6242 19740
rect 6457 19737 6469 19740
rect 6503 19737 6515 19771
rect 6457 19731 6515 19737
rect 6825 19771 6883 19777
rect 6825 19737 6837 19771
rect 6871 19737 6883 19771
rect 6932 19768 6960 19796
rect 7193 19771 7251 19777
rect 7193 19768 7205 19771
rect 6932 19740 7205 19768
rect 6825 19731 6883 19737
rect 7193 19737 7205 19740
rect 7239 19737 7251 19771
rect 7193 19731 7251 19737
rect 7392 19740 10640 19768
rect 3200 19672 4108 19700
rect 3200 19660 3206 19672
rect 4982 19660 4988 19712
rect 5040 19700 5046 19712
rect 6840 19700 6868 19731
rect 7392 19709 7420 19740
rect 5040 19672 6868 19700
rect 7377 19703 7435 19709
rect 5040 19660 5046 19672
rect 7377 19669 7389 19703
rect 7423 19669 7435 19703
rect 7377 19663 7435 19669
rect 9674 19660 9680 19712
rect 9732 19700 9738 19712
rect 9953 19703 10011 19709
rect 9953 19700 9965 19703
rect 9732 19672 9965 19700
rect 9732 19660 9738 19672
rect 9953 19669 9965 19672
rect 9999 19669 10011 19703
rect 10612 19700 10640 19740
rect 10686 19728 10692 19780
rect 10744 19728 10750 19780
rect 10980 19740 11192 19768
rect 10980 19700 11008 19740
rect 11164 19712 11192 19740
rect 11698 19728 11704 19780
rect 11756 19728 11762 19780
rect 12879 19775 12891 19808
rect 12925 19775 12937 19809
rect 14274 19796 14280 19848
rect 14332 19796 14338 19848
rect 16758 19796 16764 19848
rect 16816 19836 16822 19848
rect 16816 19808 16988 19836
rect 16816 19796 16822 19808
rect 12879 19769 12937 19775
rect 13078 19728 13084 19780
rect 13136 19768 13142 19780
rect 13722 19768 13728 19780
rect 13136 19740 13728 19768
rect 13136 19728 13142 19740
rect 13722 19728 13728 19740
rect 13780 19728 13786 19780
rect 10612 19672 11008 19700
rect 9953 19663 10011 19669
rect 11054 19660 11060 19712
rect 11112 19660 11118 19712
rect 11146 19660 11152 19712
rect 11204 19660 11210 19712
rect 11790 19660 11796 19712
rect 11848 19700 11854 19712
rect 12434 19700 12440 19712
rect 11848 19672 12440 19700
rect 11848 19660 11854 19672
rect 12434 19660 12440 19672
rect 12492 19660 12498 19712
rect 12710 19660 12716 19712
rect 12768 19700 12774 19712
rect 14292 19700 14320 19796
rect 16022 19728 16028 19780
rect 16080 19768 16086 19780
rect 16960 19777 16988 19808
rect 17126 19796 17132 19848
rect 17184 19796 17190 19848
rect 18414 19796 18420 19848
rect 18472 19836 18478 19848
rect 18785 19839 18843 19845
rect 18785 19836 18797 19839
rect 18472 19808 18797 19836
rect 18472 19796 18478 19808
rect 18785 19805 18797 19808
rect 18831 19805 18843 19839
rect 18785 19799 18843 19805
rect 18966 19796 18972 19848
rect 19024 19796 19030 19848
rect 19058 19796 19064 19848
rect 19116 19836 19122 19848
rect 19501 19839 19559 19845
rect 19501 19836 19513 19839
rect 19116 19808 19513 19836
rect 19116 19796 19122 19808
rect 19501 19805 19513 19808
rect 19547 19805 19559 19839
rect 19501 19799 19559 19805
rect 20898 19796 20904 19848
rect 20956 19796 20962 19848
rect 21085 19839 21143 19845
rect 21085 19805 21097 19839
rect 21131 19836 21143 19839
rect 21174 19836 21180 19848
rect 21131 19808 21180 19836
rect 21131 19805 21143 19808
rect 21085 19799 21143 19805
rect 21174 19796 21180 19808
rect 21232 19796 21238 19848
rect 21284 19845 21312 19876
rect 21269 19839 21327 19845
rect 21269 19805 21281 19839
rect 21315 19805 21327 19839
rect 21269 19799 21327 19805
rect 21358 19796 21364 19848
rect 21416 19796 21422 19848
rect 16485 19771 16543 19777
rect 16485 19768 16497 19771
rect 16080 19740 16497 19768
rect 16080 19728 16086 19740
rect 16485 19737 16497 19740
rect 16531 19737 16543 19771
rect 16485 19731 16543 19737
rect 16577 19771 16635 19777
rect 16577 19737 16589 19771
rect 16623 19737 16635 19771
rect 16577 19731 16635 19737
rect 16945 19771 17003 19777
rect 16945 19737 16957 19771
rect 16991 19737 17003 19771
rect 17144 19768 17172 19796
rect 17310 19768 17316 19780
rect 17144 19740 17316 19768
rect 16945 19731 17003 19737
rect 12768 19672 14320 19700
rect 12768 19660 12774 19672
rect 15746 19660 15752 19712
rect 15804 19700 15810 19712
rect 16209 19703 16267 19709
rect 16209 19700 16221 19703
rect 15804 19672 16221 19700
rect 15804 19660 15810 19672
rect 16209 19669 16221 19672
rect 16255 19669 16267 19703
rect 16592 19700 16620 19731
rect 17310 19728 17316 19740
rect 17368 19728 17374 19780
rect 19610 19768 19616 19780
rect 18616 19740 19616 19768
rect 17126 19700 17132 19712
rect 16592 19672 17132 19700
rect 16209 19663 16267 19669
rect 17126 19660 17132 19672
rect 17184 19660 17190 19712
rect 18616 19709 18644 19740
rect 19610 19728 19616 19740
rect 19668 19728 19674 19780
rect 20162 19728 20168 19780
rect 20220 19768 20226 19780
rect 20438 19768 20444 19780
rect 20220 19740 20444 19768
rect 20220 19728 20226 19740
rect 20438 19728 20444 19740
rect 20496 19728 20502 19780
rect 20993 19771 21051 19777
rect 20993 19737 21005 19771
rect 21039 19768 21051 19771
rect 21376 19768 21404 19796
rect 21039 19740 21404 19768
rect 21039 19737 21051 19740
rect 20993 19731 21051 19737
rect 18601 19703 18659 19709
rect 18601 19669 18613 19703
rect 18647 19669 18659 19703
rect 18601 19663 18659 19669
rect 18874 19660 18880 19712
rect 18932 19660 18938 19712
rect 21453 19703 21511 19709
rect 21453 19669 21465 19703
rect 21499 19700 21511 19703
rect 22186 19700 22192 19712
rect 21499 19672 22192 19700
rect 21499 19669 21511 19672
rect 21453 19663 21511 19669
rect 22186 19660 22192 19672
rect 22244 19660 22250 19712
rect 1104 19610 22056 19632
rect 658 19524 664 19576
rect 716 19524 722 19576
rect 1104 19558 6148 19610
rect 6200 19558 6212 19610
rect 6264 19558 6276 19610
rect 6328 19558 6340 19610
rect 6392 19558 6404 19610
rect 6456 19558 11346 19610
rect 11398 19558 11410 19610
rect 11462 19558 11474 19610
rect 11526 19558 11538 19610
rect 11590 19558 11602 19610
rect 11654 19558 16544 19610
rect 16596 19558 16608 19610
rect 16660 19558 16672 19610
rect 16724 19558 16736 19610
rect 16788 19558 16800 19610
rect 16852 19558 21742 19610
rect 21794 19558 21806 19610
rect 21858 19558 21870 19610
rect 21922 19558 21934 19610
rect 21986 19558 21998 19610
rect 22050 19558 22056 19610
rect 1104 19536 22056 19558
rect 2498 19456 2504 19508
rect 2556 19456 2562 19508
rect 3053 19499 3111 19505
rect 3053 19465 3065 19499
rect 3099 19496 3111 19499
rect 3099 19468 5856 19496
rect 3099 19465 3111 19468
rect 3053 19459 3111 19465
rect 1946 19428 1952 19440
rect 1504 19400 1952 19428
rect 1504 19369 1532 19400
rect 1946 19388 1952 19400
rect 2004 19388 2010 19440
rect 2700 19400 3648 19428
rect 2700 19372 2728 19400
rect 1489 19363 1547 19369
rect 1489 19329 1501 19363
rect 1535 19329 1547 19363
rect 1489 19323 1547 19329
rect 1763 19363 1821 19369
rect 1763 19329 1775 19363
rect 1809 19360 1821 19363
rect 2590 19360 2596 19372
rect 1809 19332 2596 19360
rect 1809 19329 1821 19332
rect 1763 19323 1821 19329
rect 2590 19320 2596 19332
rect 2648 19320 2654 19372
rect 2682 19320 2688 19372
rect 2740 19320 2746 19372
rect 2866 19320 2872 19372
rect 2924 19320 2930 19372
rect 3326 19320 3332 19372
rect 3384 19360 3390 19372
rect 3513 19363 3571 19369
rect 3513 19360 3525 19363
rect 3384 19332 3525 19360
rect 3384 19320 3390 19332
rect 3513 19329 3525 19332
rect 3559 19329 3571 19363
rect 3620 19360 3648 19400
rect 4430 19388 4436 19440
rect 4488 19428 4494 19440
rect 4488 19400 5210 19428
rect 4488 19388 4494 19400
rect 3755 19363 3813 19369
rect 3755 19360 3767 19363
rect 3620 19332 3767 19360
rect 3513 19323 3571 19329
rect 3755 19329 3767 19332
rect 3801 19329 3813 19363
rect 3755 19323 3813 19329
rect 4246 19320 4252 19372
rect 4304 19360 4310 19372
rect 5182 19369 5210 19400
rect 5350 19388 5356 19440
rect 5408 19388 5414 19440
rect 5828 19428 5856 19468
rect 5902 19456 5908 19508
rect 5960 19456 5966 19508
rect 6546 19456 6552 19508
rect 6604 19496 6610 19508
rect 7006 19496 7012 19508
rect 6604 19468 7012 19496
rect 6604 19456 6610 19468
rect 7006 19456 7012 19468
rect 7064 19456 7070 19508
rect 7926 19456 7932 19508
rect 7984 19496 7990 19508
rect 8481 19499 8539 19505
rect 8481 19496 8493 19499
rect 7984 19468 8493 19496
rect 7984 19456 7990 19468
rect 8481 19465 8493 19468
rect 8527 19465 8539 19499
rect 8481 19459 8539 19465
rect 9674 19456 9680 19508
rect 9732 19496 9738 19508
rect 9732 19468 10364 19496
rect 9732 19456 9738 19468
rect 9766 19428 9772 19440
rect 5828 19400 9772 19428
rect 9766 19388 9772 19400
rect 9824 19388 9830 19440
rect 4893 19363 4951 19369
rect 4893 19360 4905 19363
rect 4304 19332 4905 19360
rect 4304 19320 4310 19332
rect 4540 19292 4568 19332
rect 4893 19329 4905 19332
rect 4939 19329 4951 19363
rect 4893 19323 4951 19329
rect 5167 19363 5225 19369
rect 5167 19329 5179 19363
rect 5213 19360 5225 19363
rect 5368 19360 5396 19388
rect 10336 19379 10364 19468
rect 11422 19456 11428 19508
rect 11480 19496 11486 19508
rect 11882 19496 11888 19508
rect 11480 19468 11888 19496
rect 11480 19456 11486 19468
rect 11882 19456 11888 19468
rect 11940 19456 11946 19508
rect 12434 19456 12440 19508
rect 12492 19496 12498 19508
rect 12492 19468 15240 19496
rect 12492 19456 12498 19468
rect 11054 19388 11060 19440
rect 11112 19428 11118 19440
rect 11112 19400 12664 19428
rect 11112 19388 11118 19400
rect 10287 19373 10364 19379
rect 5213 19332 5396 19360
rect 5213 19329 5225 19332
rect 5167 19323 5225 19329
rect 5534 19320 5540 19372
rect 5592 19360 5598 19372
rect 7469 19363 7527 19369
rect 7469 19360 7481 19363
rect 5592 19332 7481 19360
rect 5592 19320 5598 19332
rect 7469 19329 7481 19332
rect 7515 19329 7527 19363
rect 7469 19323 7527 19329
rect 7743 19363 7801 19369
rect 7743 19329 7755 19363
rect 7789 19360 7801 19363
rect 8202 19360 8208 19372
rect 7789 19332 8208 19360
rect 7789 19329 7801 19332
rect 7743 19323 7801 19329
rect 8202 19320 8208 19332
rect 8260 19320 8266 19372
rect 9858 19320 9864 19372
rect 9916 19320 9922 19372
rect 10287 19339 10299 19373
rect 10333 19342 10364 19373
rect 10333 19339 10345 19342
rect 10287 19333 10345 19339
rect 10686 19320 10692 19372
rect 10744 19360 10750 19372
rect 10744 19332 11100 19360
rect 10744 19320 10750 19332
rect 9876 19292 9904 19320
rect 10045 19295 10103 19301
rect 10045 19292 10057 19295
rect 4540 19264 4936 19292
rect 9876 19264 10057 19292
rect 4338 19184 4344 19236
rect 4396 19224 4402 19236
rect 4798 19224 4804 19236
rect 4396 19196 4804 19224
rect 4396 19184 4402 19196
rect 4798 19184 4804 19196
rect 4856 19184 4862 19236
rect 4908 19224 4936 19264
rect 10045 19261 10057 19264
rect 10091 19261 10103 19295
rect 11072 19292 11100 19332
rect 11882 19320 11888 19372
rect 11940 19360 11946 19372
rect 12066 19360 12072 19372
rect 11940 19332 12072 19360
rect 11940 19320 11946 19332
rect 12066 19320 12072 19332
rect 12124 19320 12130 19372
rect 12636 19369 12664 19400
rect 13538 19369 13544 19372
rect 12621 19363 12679 19369
rect 12621 19329 12633 19363
rect 12667 19329 12679 19363
rect 12621 19323 12679 19329
rect 13495 19363 13544 19369
rect 13495 19329 13507 19363
rect 13541 19329 13544 19363
rect 13495 19323 13544 19329
rect 13538 19320 13544 19323
rect 13596 19320 13602 19372
rect 14384 19369 14412 19468
rect 15212 19428 15240 19468
rect 15930 19456 15936 19508
rect 15988 19496 15994 19508
rect 16850 19496 16856 19508
rect 15988 19468 16856 19496
rect 15988 19456 15994 19468
rect 16850 19456 16856 19468
rect 16908 19456 16914 19508
rect 17126 19456 17132 19508
rect 17184 19496 17190 19508
rect 17681 19499 17739 19505
rect 17681 19496 17693 19499
rect 17184 19468 17693 19496
rect 17184 19456 17190 19468
rect 17681 19465 17693 19468
rect 17727 19465 17739 19499
rect 17681 19459 17739 19465
rect 15212 19400 16252 19428
rect 14369 19363 14427 19369
rect 14369 19329 14381 19363
rect 14415 19329 14427 19363
rect 14642 19360 14648 19372
rect 14603 19332 14648 19360
rect 14369 19323 14427 19329
rect 14642 19320 14648 19332
rect 14700 19320 14706 19372
rect 15378 19320 15384 19372
rect 15436 19360 15442 19372
rect 15933 19363 15991 19369
rect 15933 19360 15945 19363
rect 15436 19332 15945 19360
rect 15436 19320 15442 19332
rect 15933 19329 15945 19332
rect 15979 19329 15991 19363
rect 15933 19323 15991 19329
rect 16114 19320 16120 19372
rect 16172 19320 16178 19372
rect 16224 19360 16252 19400
rect 16298 19388 16304 19440
rect 16356 19388 16362 19440
rect 17586 19428 17592 19440
rect 16408 19400 17592 19428
rect 16408 19360 16436 19400
rect 17586 19388 17592 19400
rect 17644 19388 17650 19440
rect 18414 19388 18420 19440
rect 18472 19428 18478 19440
rect 19306 19431 19364 19437
rect 19306 19428 19318 19431
rect 18472 19400 19318 19428
rect 18472 19388 18478 19400
rect 19306 19397 19318 19400
rect 19352 19397 19364 19431
rect 19306 19391 19364 19397
rect 16669 19363 16727 19369
rect 16669 19360 16681 19363
rect 16224 19332 16436 19360
rect 16546 19332 16681 19360
rect 12437 19295 12495 19301
rect 12437 19292 12449 19295
rect 11072 19264 12449 19292
rect 10045 19255 10103 19261
rect 12084 19236 12112 19264
rect 12437 19261 12449 19264
rect 12483 19261 12495 19295
rect 12437 19255 12495 19261
rect 13354 19252 13360 19304
rect 13412 19252 13418 19304
rect 13633 19295 13691 19301
rect 13633 19261 13645 19295
rect 13679 19292 13691 19295
rect 13679 19264 14320 19292
rect 13679 19261 13691 19264
rect 13633 19255 13691 19261
rect 4908 19196 5028 19224
rect 4525 19159 4583 19165
rect 4525 19125 4537 19159
rect 4571 19156 4583 19159
rect 4614 19156 4620 19168
rect 4571 19128 4620 19156
rect 4571 19125 4583 19128
rect 4525 19119 4583 19125
rect 4614 19116 4620 19128
rect 4672 19116 4678 19168
rect 5000 19156 5028 19196
rect 8294 19184 8300 19236
rect 8352 19224 8358 19236
rect 9766 19224 9772 19236
rect 8352 19196 9772 19224
rect 8352 19184 8358 19196
rect 9766 19184 9772 19196
rect 9824 19184 9830 19236
rect 11790 19224 11796 19236
rect 10980 19196 11796 19224
rect 5350 19156 5356 19168
rect 5000 19128 5356 19156
rect 5350 19116 5356 19128
rect 5408 19116 5414 19168
rect 6914 19116 6920 19168
rect 6972 19156 6978 19168
rect 7377 19159 7435 19165
rect 7377 19156 7389 19159
rect 6972 19128 7389 19156
rect 6972 19116 6978 19128
rect 7377 19125 7389 19128
rect 7423 19125 7435 19159
rect 7377 19119 7435 19125
rect 7558 19116 7564 19168
rect 7616 19156 7622 19168
rect 8662 19156 8668 19168
rect 7616 19128 8668 19156
rect 7616 19116 7622 19128
rect 8662 19116 8668 19128
rect 8720 19116 8726 19168
rect 9582 19116 9588 19168
rect 9640 19156 9646 19168
rect 10980 19156 11008 19196
rect 11790 19184 11796 19196
rect 11848 19184 11854 19236
rect 12066 19184 12072 19236
rect 12124 19184 12130 19236
rect 13078 19184 13084 19236
rect 13136 19184 13142 19236
rect 14292 19224 14320 19264
rect 15194 19252 15200 19304
rect 15252 19292 15258 19304
rect 16546 19292 16574 19332
rect 16669 19329 16681 19332
rect 16715 19329 16727 19363
rect 16669 19323 16727 19329
rect 16850 19320 16856 19372
rect 16908 19360 16914 19372
rect 16943 19363 17001 19369
rect 16943 19360 16955 19363
rect 16908 19332 16955 19360
rect 16908 19320 16914 19332
rect 16943 19329 16955 19332
rect 16989 19329 17001 19363
rect 18598 19360 18604 19372
rect 16943 19323 17001 19329
rect 17328 19332 18604 19360
rect 15252 19264 16574 19292
rect 15252 19252 15258 19264
rect 14292 19196 14412 19224
rect 9640 19128 11008 19156
rect 11057 19159 11115 19165
rect 9640 19116 9646 19128
rect 11057 19125 11069 19159
rect 11103 19156 11115 19159
rect 12434 19156 12440 19168
rect 11103 19128 12440 19156
rect 11103 19125 11115 19128
rect 11057 19119 11115 19125
rect 12434 19116 12440 19128
rect 12492 19116 12498 19168
rect 14274 19116 14280 19168
rect 14332 19116 14338 19168
rect 14384 19156 14412 19196
rect 15102 19184 15108 19236
rect 15160 19224 15166 19236
rect 15838 19224 15844 19236
rect 15160 19196 15844 19224
rect 15160 19184 15166 19196
rect 15838 19184 15844 19196
rect 15896 19184 15902 19236
rect 15381 19159 15439 19165
rect 15381 19156 15393 19159
rect 14384 19128 15393 19156
rect 15381 19125 15393 19128
rect 15427 19125 15439 19159
rect 15381 19119 15439 19125
rect 16209 19159 16267 19165
rect 16209 19125 16221 19159
rect 16255 19156 16267 19159
rect 16298 19156 16304 19168
rect 16255 19128 16304 19156
rect 16255 19125 16267 19128
rect 16209 19119 16267 19125
rect 16298 19116 16304 19128
rect 16356 19116 16362 19168
rect 16546 19156 16574 19264
rect 17328 19156 17356 19332
rect 18598 19320 18604 19332
rect 18656 19320 18662 19372
rect 18785 19363 18843 19369
rect 18785 19329 18797 19363
rect 18831 19360 18843 19363
rect 18874 19360 18880 19372
rect 18831 19332 18880 19360
rect 18831 19329 18843 19332
rect 18785 19323 18843 19329
rect 18874 19320 18880 19332
rect 18932 19320 18938 19372
rect 20533 19363 20591 19369
rect 20533 19329 20545 19363
rect 20579 19360 20591 19363
rect 20622 19360 20628 19372
rect 20579 19332 20628 19360
rect 20579 19329 20591 19332
rect 20533 19323 20591 19329
rect 20622 19320 20628 19332
rect 20680 19320 20686 19372
rect 21174 19320 21180 19372
rect 21232 19320 21238 19372
rect 18966 19252 18972 19304
rect 19024 19292 19030 19304
rect 19061 19295 19119 19301
rect 19061 19292 19073 19295
rect 19024 19264 19073 19292
rect 19024 19252 19030 19264
rect 19061 19261 19073 19264
rect 19107 19261 19119 19295
rect 19061 19255 19119 19261
rect 20809 19295 20867 19301
rect 20809 19261 20821 19295
rect 20855 19292 20867 19295
rect 20855 19264 21036 19292
rect 20855 19261 20867 19264
rect 20809 19255 20867 19261
rect 20625 19227 20683 19233
rect 20625 19224 20637 19227
rect 19996 19196 20637 19224
rect 16546 19128 17356 19156
rect 18877 19159 18935 19165
rect 18877 19125 18889 19159
rect 18923 19156 18935 19159
rect 19996 19156 20024 19196
rect 20625 19193 20637 19196
rect 20671 19193 20683 19227
rect 20625 19187 20683 19193
rect 21008 19168 21036 19264
rect 18923 19128 20024 19156
rect 18923 19125 18935 19128
rect 18877 19119 18935 19125
rect 20438 19116 20444 19168
rect 20496 19116 20502 19168
rect 20714 19116 20720 19168
rect 20772 19116 20778 19168
rect 20990 19116 20996 19168
rect 21048 19116 21054 19168
rect 21450 19116 21456 19168
rect 21508 19116 21514 19168
rect 1104 19066 21896 19088
rect 1104 19014 3549 19066
rect 3601 19014 3613 19066
rect 3665 19014 3677 19066
rect 3729 19014 3741 19066
rect 3793 19014 3805 19066
rect 3857 19014 8747 19066
rect 8799 19014 8811 19066
rect 8863 19014 8875 19066
rect 8927 19014 8939 19066
rect 8991 19014 9003 19066
rect 9055 19014 13945 19066
rect 13997 19014 14009 19066
rect 14061 19014 14073 19066
rect 14125 19014 14137 19066
rect 14189 19014 14201 19066
rect 14253 19014 19143 19066
rect 19195 19014 19207 19066
rect 19259 19014 19271 19066
rect 19323 19014 19335 19066
rect 19387 19014 19399 19066
rect 19451 19014 21896 19066
rect 1104 18992 21896 19014
rect 1026 18912 1032 18964
rect 1084 18952 1090 18964
rect 4522 18952 4528 18964
rect 1084 18924 4528 18952
rect 1084 18912 1090 18924
rect 4522 18912 4528 18924
rect 4580 18912 4586 18964
rect 5442 18952 5448 18964
rect 4724 18924 5448 18952
rect 1397 18819 1455 18825
rect 1397 18785 1409 18819
rect 1443 18816 1455 18819
rect 1486 18816 1492 18828
rect 1443 18788 1492 18816
rect 1443 18785 1455 18788
rect 1397 18779 1455 18785
rect 1486 18776 1492 18788
rect 1544 18776 1550 18828
rect 1670 18776 1676 18828
rect 1728 18776 1734 18828
rect 2314 18776 2320 18828
rect 2372 18776 2378 18828
rect 3234 18776 3240 18828
rect 3292 18816 3298 18828
rect 3789 18819 3847 18825
rect 3789 18816 3801 18819
rect 3292 18788 3801 18816
rect 3292 18776 3298 18788
rect 3789 18785 3801 18788
rect 3835 18785 3847 18819
rect 3789 18779 3847 18785
rect 4062 18776 4068 18828
rect 4120 18776 4126 18828
rect 4724 18825 4752 18924
rect 5442 18912 5448 18924
rect 5500 18912 5506 18964
rect 5718 18912 5724 18964
rect 5776 18912 5782 18964
rect 7098 18912 7104 18964
rect 7156 18912 7162 18964
rect 9766 18952 9772 18964
rect 7300 18924 9772 18952
rect 7300 18896 7328 18924
rect 9766 18912 9772 18924
rect 9824 18912 9830 18964
rect 10410 18912 10416 18964
rect 10468 18912 10474 18964
rect 12618 18952 12624 18964
rect 11716 18924 12624 18952
rect 7282 18844 7288 18896
rect 7340 18844 7346 18896
rect 11716 18893 11744 18924
rect 12618 18912 12624 18924
rect 12676 18912 12682 18964
rect 12802 18912 12808 18964
rect 12860 18912 12866 18964
rect 13354 18912 13360 18964
rect 13412 18952 13418 18964
rect 13541 18955 13599 18961
rect 13541 18952 13553 18955
rect 13412 18924 13553 18952
rect 13412 18912 13418 18924
rect 13541 18921 13553 18924
rect 13587 18921 13599 18955
rect 13541 18915 13599 18921
rect 15194 18912 15200 18964
rect 15252 18912 15258 18964
rect 15378 18912 15384 18964
rect 15436 18912 15442 18964
rect 16114 18912 16120 18964
rect 16172 18952 16178 18964
rect 16761 18955 16819 18961
rect 16172 18924 16436 18952
rect 16172 18912 16178 18924
rect 11701 18887 11759 18893
rect 10152 18856 11652 18884
rect 10152 18828 10180 18856
rect 11624 18828 11652 18856
rect 11701 18853 11713 18887
rect 11747 18853 11759 18887
rect 12820 18884 12848 18912
rect 14642 18884 14648 18896
rect 12820 18856 14648 18884
rect 11701 18847 11759 18853
rect 14642 18844 14648 18856
rect 14700 18844 14706 18896
rect 15212 18884 15240 18912
rect 16408 18884 16436 18924
rect 16761 18921 16773 18955
rect 16807 18952 16819 18955
rect 16942 18952 16948 18964
rect 16807 18924 16948 18952
rect 16807 18921 16819 18924
rect 16761 18915 16819 18921
rect 16942 18912 16948 18924
rect 17000 18912 17006 18964
rect 19518 18952 19524 18964
rect 19260 18924 19524 18952
rect 15212 18856 15792 18884
rect 16408 18856 17172 18884
rect 4709 18819 4767 18825
rect 4709 18785 4721 18819
rect 4755 18785 4767 18819
rect 4709 18779 4767 18785
rect 5534 18776 5540 18828
rect 5592 18816 5598 18828
rect 6089 18819 6147 18825
rect 6089 18816 6101 18819
rect 5592 18788 6101 18816
rect 5592 18776 5598 18788
rect 6089 18785 6101 18788
rect 6135 18785 6147 18819
rect 6089 18779 6147 18785
rect 8128 18788 9352 18816
rect 2222 18708 2228 18760
rect 2280 18748 2286 18760
rect 2590 18757 2596 18760
rect 2559 18751 2596 18757
rect 2559 18748 2571 18751
rect 2280 18720 2571 18748
rect 2280 18708 2286 18720
rect 2559 18717 2571 18720
rect 2559 18711 2596 18717
rect 2590 18708 2596 18711
rect 2648 18708 2654 18760
rect 4983 18751 5041 18757
rect 4983 18717 4995 18751
rect 5029 18717 5041 18751
rect 7469 18751 7527 18757
rect 4983 18711 5041 18717
rect 6347 18721 6405 18727
rect 4614 18640 4620 18692
rect 4672 18680 4678 18692
rect 4798 18680 4804 18692
rect 4672 18652 4804 18680
rect 4672 18640 4678 18652
rect 4798 18640 4804 18652
rect 4856 18640 4862 18692
rect 4998 18680 5026 18711
rect 5258 18680 5264 18692
rect 4998 18652 5264 18680
rect 5258 18640 5264 18652
rect 5316 18640 5322 18692
rect 6347 18687 6359 18721
rect 6393 18718 6405 18721
rect 6393 18687 6406 18718
rect 7469 18717 7481 18751
rect 7515 18748 7527 18751
rect 7743 18751 7801 18757
rect 7515 18720 7604 18748
rect 7515 18717 7527 18720
rect 7469 18711 7527 18717
rect 7576 18692 7604 18720
rect 7743 18717 7755 18751
rect 7789 18748 7801 18751
rect 7789 18720 7880 18748
rect 7789 18717 7801 18720
rect 7743 18711 7801 18717
rect 7852 18692 7880 18720
rect 6347 18681 6406 18687
rect 6378 18680 6406 18681
rect 7098 18680 7104 18692
rect 6378 18652 7104 18680
rect 7098 18640 7104 18652
rect 7156 18640 7162 18692
rect 7558 18640 7564 18692
rect 7616 18640 7622 18692
rect 7834 18640 7840 18692
rect 7892 18640 7898 18692
rect 3326 18572 3332 18624
rect 3384 18572 3390 18624
rect 4890 18572 4896 18624
rect 4948 18612 4954 18624
rect 5350 18612 5356 18624
rect 4948 18584 5356 18612
rect 4948 18572 4954 18584
rect 5350 18572 5356 18584
rect 5408 18572 5414 18624
rect 5442 18572 5448 18624
rect 5500 18612 5506 18624
rect 8128 18612 8156 18788
rect 8846 18708 8852 18760
rect 8904 18748 8910 18760
rect 9125 18751 9183 18757
rect 9125 18748 9137 18751
rect 8904 18720 9137 18748
rect 8904 18708 8910 18720
rect 9125 18717 9137 18720
rect 9171 18717 9183 18751
rect 9125 18711 9183 18717
rect 8294 18680 8300 18692
rect 8220 18652 8300 18680
rect 8220 18624 8248 18652
rect 8294 18640 8300 18652
rect 8352 18640 8358 18692
rect 5500 18584 8156 18612
rect 5500 18572 5506 18584
rect 8202 18572 8208 18624
rect 8260 18572 8266 18624
rect 8386 18572 8392 18624
rect 8444 18612 8450 18624
rect 8481 18615 8539 18621
rect 8481 18612 8493 18615
rect 8444 18584 8493 18612
rect 8444 18572 8450 18584
rect 8481 18581 8493 18584
rect 8527 18581 8539 18615
rect 9324 18612 9352 18788
rect 9398 18776 9404 18828
rect 9456 18776 9462 18828
rect 10134 18776 10140 18828
rect 10192 18776 10198 18828
rect 11054 18776 11060 18828
rect 11112 18776 11118 18828
rect 11606 18776 11612 18828
rect 11664 18816 11670 18828
rect 11977 18819 12035 18825
rect 11977 18816 11989 18819
rect 11664 18788 11989 18816
rect 11664 18776 11670 18788
rect 11977 18785 11989 18788
rect 12023 18785 12035 18819
rect 11977 18779 12035 18785
rect 12066 18776 12072 18828
rect 12124 18825 12130 18828
rect 12124 18819 12152 18825
rect 12140 18785 12152 18819
rect 12124 18779 12152 18785
rect 12253 18819 12311 18825
rect 12253 18785 12265 18819
rect 12299 18816 12311 18819
rect 12434 18816 12440 18828
rect 12299 18788 12440 18816
rect 12299 18785 12311 18788
rect 12253 18779 12311 18785
rect 12124 18776 12130 18779
rect 12434 18776 12440 18788
rect 12492 18776 12498 18828
rect 15102 18776 15108 18828
rect 15160 18816 15166 18828
rect 15764 18825 15792 18856
rect 15749 18819 15807 18825
rect 15160 18788 15332 18816
rect 15160 18776 15166 18788
rect 9675 18751 9733 18757
rect 9675 18717 9687 18751
rect 9721 18748 9733 18751
rect 11241 18751 11299 18757
rect 11241 18748 11253 18751
rect 9721 18720 9996 18748
rect 9721 18717 9733 18720
rect 9675 18711 9733 18717
rect 9968 18692 9996 18720
rect 11072 18720 11253 18748
rect 9950 18640 9956 18692
rect 10008 18640 10014 18692
rect 11072 18612 11100 18720
rect 11241 18717 11253 18720
rect 11287 18748 11299 18751
rect 11422 18748 11428 18760
rect 11287 18720 11428 18748
rect 11287 18717 11299 18720
rect 11241 18711 11299 18717
rect 11422 18708 11428 18720
rect 11480 18708 11486 18760
rect 12897 18751 12955 18757
rect 12897 18717 12909 18751
rect 12943 18748 12955 18751
rect 15194 18748 15200 18760
rect 12943 18720 15200 18748
rect 12943 18717 12955 18720
rect 12897 18711 12955 18717
rect 15194 18708 15200 18720
rect 15252 18708 15258 18760
rect 15304 18757 15332 18788
rect 15749 18785 15761 18819
rect 15795 18785 15807 18819
rect 15749 18779 15807 18785
rect 15289 18751 15347 18757
rect 15289 18717 15301 18751
rect 15335 18717 15347 18751
rect 15289 18711 15347 18717
rect 16023 18751 16081 18757
rect 16023 18717 16035 18751
rect 16069 18748 16081 18751
rect 16942 18748 16948 18760
rect 16069 18720 16948 18748
rect 16069 18717 16081 18720
rect 16023 18711 16081 18717
rect 16942 18708 16948 18720
rect 17000 18708 17006 18760
rect 17144 18757 17172 18856
rect 17402 18776 17408 18828
rect 17460 18776 17466 18828
rect 19260 18825 19288 18924
rect 19518 18912 19524 18924
rect 19576 18952 19582 18964
rect 19702 18952 19708 18964
rect 19576 18924 19708 18952
rect 19576 18912 19582 18924
rect 19702 18912 19708 18924
rect 19760 18912 19766 18964
rect 20530 18912 20536 18964
rect 20588 18912 20594 18964
rect 21085 18955 21143 18961
rect 21085 18921 21097 18955
rect 21131 18952 21143 18955
rect 21174 18952 21180 18964
rect 21131 18924 21180 18952
rect 21131 18921 21143 18924
rect 21085 18915 21143 18921
rect 21174 18912 21180 18924
rect 21232 18912 21238 18964
rect 20346 18844 20352 18896
rect 20404 18884 20410 18896
rect 20548 18884 20576 18912
rect 20404 18856 21128 18884
rect 20404 18844 20410 18856
rect 19245 18819 19303 18825
rect 19245 18785 19257 18819
rect 19291 18785 19303 18819
rect 19245 18779 19303 18785
rect 20717 18819 20775 18825
rect 20717 18785 20729 18819
rect 20763 18816 20775 18819
rect 20993 18819 21051 18825
rect 20993 18816 21005 18819
rect 20763 18788 21005 18816
rect 20763 18785 20775 18788
rect 20717 18779 20775 18785
rect 20993 18785 21005 18788
rect 21039 18785 21051 18819
rect 20993 18779 21051 18785
rect 17129 18751 17187 18757
rect 17129 18717 17141 18751
rect 17175 18717 17187 18751
rect 17129 18711 17187 18717
rect 17770 18708 17776 18760
rect 17828 18748 17834 18760
rect 19487 18751 19545 18757
rect 19487 18748 19499 18751
rect 17828 18720 18092 18748
rect 17828 18708 17834 18720
rect 17954 18680 17960 18692
rect 12820 18652 17960 18680
rect 9324 18584 11100 18612
rect 8481 18575 8539 18581
rect 11146 18572 11152 18624
rect 11204 18612 11210 18624
rect 12820 18612 12848 18652
rect 17954 18640 17960 18652
rect 18012 18640 18018 18692
rect 18064 18680 18092 18720
rect 19352 18720 19499 18748
rect 19352 18680 19380 18720
rect 19487 18717 19499 18720
rect 19533 18717 19545 18751
rect 19487 18711 19545 18717
rect 19610 18708 19616 18760
rect 19668 18748 19674 18760
rect 20625 18751 20683 18757
rect 20625 18748 20637 18751
rect 19668 18720 20637 18748
rect 19668 18708 19674 18720
rect 20625 18717 20637 18720
rect 20671 18717 20683 18751
rect 20625 18711 20683 18717
rect 20901 18751 20959 18757
rect 20901 18717 20913 18751
rect 20947 18748 20959 18751
rect 21100 18748 21128 18856
rect 21177 18819 21235 18825
rect 21177 18785 21189 18819
rect 21223 18785 21235 18819
rect 21177 18779 21235 18785
rect 20947 18720 21128 18748
rect 20947 18717 20959 18720
rect 20901 18711 20959 18717
rect 18064 18652 19380 18680
rect 20530 18640 20536 18692
rect 20588 18680 20594 18692
rect 21192 18680 21220 18779
rect 21269 18751 21327 18757
rect 21269 18717 21281 18751
rect 21315 18748 21327 18751
rect 22738 18748 22744 18760
rect 21315 18720 22744 18748
rect 21315 18717 21327 18720
rect 21269 18711 21327 18717
rect 22738 18708 22744 18720
rect 22796 18708 22802 18760
rect 20588 18652 21220 18680
rect 20588 18640 20594 18652
rect 22646 18640 22652 18692
rect 22704 18640 22710 18692
rect 11204 18584 12848 18612
rect 11204 18572 11210 18584
rect 14274 18572 14280 18624
rect 14332 18612 14338 18624
rect 19518 18612 19524 18624
rect 14332 18584 19524 18612
rect 14332 18572 14338 18584
rect 19518 18572 19524 18584
rect 19576 18572 19582 18624
rect 20257 18615 20315 18621
rect 20257 18581 20269 18615
rect 20303 18612 20315 18615
rect 20622 18612 20628 18624
rect 20303 18584 20628 18612
rect 20303 18581 20315 18584
rect 20257 18575 20315 18581
rect 20622 18572 20628 18584
rect 20680 18572 20686 18624
rect 21453 18615 21511 18621
rect 21453 18581 21465 18615
rect 21499 18612 21511 18615
rect 22186 18612 22192 18624
rect 21499 18584 22192 18612
rect 21499 18581 21511 18584
rect 21453 18575 21511 18581
rect 22186 18572 22192 18584
rect 22244 18572 22250 18624
rect 1104 18522 22056 18544
rect 1104 18470 6148 18522
rect 6200 18470 6212 18522
rect 6264 18470 6276 18522
rect 6328 18470 6340 18522
rect 6392 18470 6404 18522
rect 6456 18470 11346 18522
rect 11398 18470 11410 18522
rect 11462 18470 11474 18522
rect 11526 18470 11538 18522
rect 11590 18470 11602 18522
rect 11654 18470 16544 18522
rect 16596 18470 16608 18522
rect 16660 18470 16672 18522
rect 16724 18470 16736 18522
rect 16788 18470 16800 18522
rect 16852 18470 21742 18522
rect 21794 18470 21806 18522
rect 21858 18470 21870 18522
rect 21922 18470 21934 18522
rect 21986 18470 21998 18522
rect 22050 18470 22056 18522
rect 22664 18488 22692 18640
rect 1104 18448 22056 18470
rect 22646 18436 22652 18488
rect 22704 18436 22710 18488
rect 3142 18368 3148 18420
rect 3200 18408 3206 18420
rect 5629 18411 5687 18417
rect 5629 18408 5641 18411
rect 3200 18380 5641 18408
rect 3200 18368 3206 18380
rect 5629 18377 5641 18380
rect 5675 18377 5687 18411
rect 5629 18371 5687 18377
rect 6730 18368 6736 18420
rect 6788 18368 6794 18420
rect 6914 18368 6920 18420
rect 6972 18408 6978 18420
rect 7558 18408 7564 18420
rect 6972 18380 7564 18408
rect 6972 18368 6978 18380
rect 7558 18368 7564 18380
rect 7616 18368 7622 18420
rect 7926 18368 7932 18420
rect 7984 18408 7990 18420
rect 8294 18408 8300 18420
rect 7984 18380 8300 18408
rect 7984 18368 7990 18380
rect 8294 18368 8300 18380
rect 8352 18408 8358 18420
rect 8389 18411 8447 18417
rect 8389 18408 8401 18411
rect 8352 18380 8401 18408
rect 8352 18368 8358 18380
rect 8389 18377 8401 18380
rect 8435 18377 8447 18411
rect 8389 18371 8447 18377
rect 8588 18380 9168 18408
rect 934 18300 940 18352
rect 992 18340 998 18352
rect 2041 18343 2099 18349
rect 2041 18340 2053 18343
rect 992 18312 2053 18340
rect 992 18300 998 18312
rect 2041 18309 2053 18312
rect 2087 18309 2099 18343
rect 2041 18303 2099 18309
rect 2225 18343 2283 18349
rect 2225 18309 2237 18343
rect 2271 18340 2283 18343
rect 2958 18340 2964 18352
rect 2271 18312 2964 18340
rect 2271 18309 2283 18312
rect 2225 18303 2283 18309
rect 2958 18300 2964 18312
rect 3016 18300 3022 18352
rect 6748 18340 6776 18368
rect 8110 18340 8116 18352
rect 6748 18312 8116 18340
rect 8110 18300 8116 18312
rect 8168 18340 8174 18352
rect 8588 18340 8616 18380
rect 8168 18312 8616 18340
rect 8665 18343 8723 18349
rect 8168 18300 8174 18312
rect 8665 18309 8677 18343
rect 8711 18340 8723 18343
rect 8846 18340 8852 18352
rect 8711 18312 8852 18340
rect 8711 18309 8723 18312
rect 8665 18303 8723 18309
rect 8846 18300 8852 18312
rect 8904 18300 8910 18352
rect 9140 18349 9168 18380
rect 9214 18368 9220 18420
rect 9272 18408 9278 18420
rect 9493 18411 9551 18417
rect 9493 18408 9505 18411
rect 9272 18380 9505 18408
rect 9272 18368 9278 18380
rect 9493 18377 9505 18380
rect 9539 18377 9551 18411
rect 9493 18371 9551 18377
rect 9677 18411 9735 18417
rect 9677 18377 9689 18411
rect 9723 18377 9735 18411
rect 9677 18371 9735 18377
rect 9125 18343 9183 18349
rect 9125 18309 9137 18343
rect 9171 18309 9183 18343
rect 9692 18340 9720 18371
rect 10594 18368 10600 18420
rect 10652 18408 10658 18420
rect 12710 18408 12716 18420
rect 10652 18380 12716 18408
rect 10652 18368 10658 18380
rect 12710 18368 12716 18380
rect 12768 18368 12774 18420
rect 13078 18368 13084 18420
rect 13136 18368 13142 18420
rect 13722 18368 13728 18420
rect 13780 18408 13786 18420
rect 16117 18411 16175 18417
rect 13780 18380 15792 18408
rect 13780 18368 13786 18380
rect 10686 18340 10692 18352
rect 9692 18312 10692 18340
rect 9125 18303 9183 18309
rect 10686 18300 10692 18312
rect 10744 18300 10750 18352
rect 10870 18300 10876 18352
rect 10928 18340 10934 18352
rect 10928 18312 11928 18340
rect 10928 18300 10934 18312
rect 1489 18275 1547 18281
rect 1489 18241 1501 18275
rect 1535 18272 1547 18275
rect 1946 18272 1952 18284
rect 1535 18244 1952 18272
rect 1535 18241 1547 18244
rect 1489 18235 1547 18241
rect 1946 18232 1952 18244
rect 2004 18232 2010 18284
rect 2682 18281 2688 18284
rect 2651 18275 2688 18281
rect 2651 18272 2663 18275
rect 2240 18244 2663 18272
rect 2240 18080 2268 18244
rect 2651 18241 2663 18244
rect 2651 18235 2688 18241
rect 2682 18232 2688 18235
rect 2740 18232 2746 18284
rect 3789 18275 3847 18281
rect 3789 18241 3801 18275
rect 3835 18272 3847 18275
rect 3835 18244 4108 18272
rect 3835 18241 3847 18244
rect 3789 18235 3847 18241
rect 4080 18216 4108 18244
rect 4982 18232 4988 18284
rect 5040 18232 5046 18284
rect 7098 18272 7104 18284
rect 7059 18244 7104 18272
rect 7098 18232 7104 18244
rect 7156 18232 7162 18284
rect 7466 18232 7472 18284
rect 7524 18272 7530 18284
rect 7926 18272 7932 18284
rect 7524 18244 7932 18272
rect 7524 18232 7530 18244
rect 7926 18232 7932 18244
rect 7984 18232 7990 18284
rect 8757 18275 8815 18281
rect 8757 18241 8769 18275
rect 8803 18272 8815 18275
rect 9950 18272 9956 18284
rect 8803 18244 9956 18272
rect 8803 18241 8815 18244
rect 8757 18235 8815 18241
rect 9950 18232 9956 18244
rect 10008 18232 10014 18284
rect 10226 18232 10232 18284
rect 10284 18272 10290 18284
rect 10319 18275 10377 18281
rect 10319 18272 10331 18275
rect 10284 18244 10331 18272
rect 10284 18232 10290 18244
rect 10319 18241 10331 18244
rect 10365 18241 10377 18275
rect 11900 18272 11928 18312
rect 15654 18300 15660 18352
rect 15712 18300 15718 18352
rect 15764 18340 15792 18380
rect 16117 18377 16129 18411
rect 16163 18408 16175 18411
rect 16206 18408 16212 18420
rect 16163 18380 16212 18408
rect 16163 18377 16175 18380
rect 16117 18371 16175 18377
rect 16206 18368 16212 18380
rect 16264 18368 16270 18420
rect 20070 18408 20076 18420
rect 16314 18380 20076 18408
rect 16314 18340 16342 18380
rect 20070 18368 20076 18380
rect 20128 18368 20134 18420
rect 20346 18368 20352 18420
rect 20404 18368 20410 18420
rect 20438 18368 20444 18420
rect 20496 18368 20502 18420
rect 20530 18368 20536 18420
rect 20588 18368 20594 18420
rect 20714 18368 20720 18420
rect 20772 18408 20778 18420
rect 20772 18380 21220 18408
rect 20772 18368 20778 18380
rect 15764 18312 16342 18340
rect 16927 18305 16985 18311
rect 12311 18275 12369 18281
rect 12311 18272 12323 18275
rect 11900 18244 12323 18272
rect 10319 18235 10377 18241
rect 12311 18241 12323 18244
rect 12357 18241 12369 18275
rect 12311 18235 12369 18241
rect 13814 18232 13820 18284
rect 13872 18272 13878 18284
rect 14151 18275 14209 18281
rect 14151 18272 14163 18275
rect 13872 18244 14163 18272
rect 13872 18232 13878 18244
rect 14151 18241 14163 18244
rect 14197 18241 14209 18275
rect 15672 18272 15700 18300
rect 16301 18275 16359 18281
rect 16301 18272 16313 18275
rect 15672 18244 16313 18272
rect 14151 18235 14209 18241
rect 16301 18241 16313 18244
rect 16347 18241 16359 18275
rect 16301 18235 16359 18241
rect 16390 18232 16396 18284
rect 16448 18272 16454 18284
rect 16927 18272 16939 18305
rect 16448 18271 16939 18272
rect 16973 18271 16985 18305
rect 17954 18300 17960 18352
rect 18012 18340 18018 18352
rect 18938 18343 18996 18349
rect 18938 18340 18950 18343
rect 18012 18312 18950 18340
rect 18012 18300 18018 18312
rect 18938 18309 18950 18312
rect 18984 18340 18996 18343
rect 19058 18340 19064 18352
rect 18984 18312 19064 18340
rect 18984 18309 18996 18312
rect 18938 18303 18996 18309
rect 19058 18300 19064 18312
rect 19116 18300 19122 18352
rect 20364 18281 20392 18368
rect 20456 18340 20484 18368
rect 21192 18349 21220 18380
rect 21177 18343 21235 18349
rect 20456 18312 20852 18340
rect 20824 18281 20852 18312
rect 21177 18309 21189 18343
rect 21223 18309 21235 18343
rect 21177 18303 21235 18309
rect 16448 18265 16985 18271
rect 20349 18275 20407 18281
rect 16448 18244 16970 18265
rect 16448 18232 16454 18244
rect 20349 18241 20361 18275
rect 20395 18241 20407 18275
rect 20349 18235 20407 18241
rect 20533 18275 20591 18281
rect 20533 18241 20545 18275
rect 20579 18272 20591 18275
rect 20809 18275 20867 18281
rect 20579 18244 20668 18272
rect 20579 18241 20591 18244
rect 20533 18235 20591 18241
rect 8392 18216 8444 18222
rect 2314 18164 2320 18216
rect 2372 18204 2378 18216
rect 2409 18207 2467 18213
rect 2409 18204 2421 18207
rect 2372 18176 2421 18204
rect 2372 18164 2378 18176
rect 2409 18173 2421 18176
rect 2455 18173 2467 18207
rect 2409 18167 2467 18173
rect 3418 18164 3424 18216
rect 3476 18204 3482 18216
rect 3973 18207 4031 18213
rect 3973 18204 3985 18207
rect 3476 18176 3985 18204
rect 3476 18164 3482 18176
rect 3973 18173 3985 18176
rect 4019 18173 4031 18207
rect 3973 18167 4031 18173
rect 4062 18164 4068 18216
rect 4120 18164 4126 18216
rect 4154 18164 4160 18216
rect 4212 18204 4218 18216
rect 4709 18207 4767 18213
rect 4709 18204 4721 18207
rect 4212 18176 4721 18204
rect 4212 18164 4218 18176
rect 3878 18096 3884 18148
rect 3936 18136 3942 18148
rect 4433 18139 4491 18145
rect 4433 18136 4445 18139
rect 3936 18108 4445 18136
rect 3936 18096 3942 18108
rect 4433 18105 4445 18108
rect 4479 18105 4491 18139
rect 4433 18099 4491 18105
rect 1578 18028 1584 18080
rect 1636 18028 1642 18080
rect 2222 18028 2228 18080
rect 2280 18028 2286 18080
rect 3421 18071 3479 18077
rect 3421 18037 3433 18071
rect 3467 18068 3479 18071
rect 3970 18068 3976 18080
rect 3467 18040 3976 18068
rect 3467 18037 3479 18040
rect 3421 18031 3479 18037
rect 3970 18028 3976 18040
rect 4028 18028 4034 18080
rect 4540 18068 4568 18176
rect 4709 18173 4721 18176
rect 4755 18173 4767 18207
rect 4709 18167 4767 18173
rect 4798 18164 4804 18216
rect 4856 18213 4862 18216
rect 4856 18207 4884 18213
rect 4872 18173 4884 18207
rect 4856 18167 4884 18173
rect 4856 18164 4862 18167
rect 5350 18164 5356 18216
rect 5408 18164 5414 18216
rect 5534 18164 5540 18216
rect 5592 18204 5598 18216
rect 6825 18207 6883 18213
rect 6825 18204 6837 18207
rect 5592 18176 6837 18204
rect 5592 18164 5598 18176
rect 6825 18173 6837 18176
rect 6871 18173 6883 18207
rect 6825 18167 6883 18173
rect 10042 18164 10048 18216
rect 10100 18164 10106 18216
rect 11790 18164 11796 18216
rect 11848 18204 11854 18216
rect 12069 18207 12127 18213
rect 11848 18176 11928 18204
rect 11848 18164 11854 18176
rect 4798 18068 4804 18080
rect 4540 18040 4804 18068
rect 4798 18028 4804 18040
rect 4856 18028 4862 18080
rect 5368 18068 5396 18164
rect 8392 18158 8444 18164
rect 11900 18136 11928 18176
rect 12069 18173 12081 18207
rect 12115 18173 12127 18207
rect 12069 18167 12127 18173
rect 12084 18136 12112 18167
rect 13078 18164 13084 18216
rect 13136 18204 13142 18216
rect 13909 18207 13967 18213
rect 13909 18204 13921 18207
rect 13136 18176 13921 18204
rect 13136 18164 13142 18176
rect 13909 18173 13921 18176
rect 13955 18173 13967 18207
rect 13909 18167 13967 18173
rect 11900 18108 12112 18136
rect 7282 18068 7288 18080
rect 5368 18040 7288 18068
rect 7282 18028 7288 18040
rect 7340 18028 7346 18080
rect 7834 18028 7840 18080
rect 7892 18028 7898 18080
rect 11054 18028 11060 18080
rect 11112 18028 11118 18080
rect 11146 18028 11152 18080
rect 11204 18068 11210 18080
rect 12802 18068 12808 18080
rect 11204 18040 12808 18068
rect 11204 18028 11210 18040
rect 12802 18028 12808 18040
rect 12860 18028 12866 18080
rect 13924 18068 13952 18167
rect 15378 18164 15384 18216
rect 15436 18204 15442 18216
rect 16666 18204 16672 18216
rect 15436 18176 16672 18204
rect 15436 18164 15442 18176
rect 16666 18164 16672 18176
rect 16724 18164 16730 18216
rect 18693 18207 18751 18213
rect 18693 18173 18705 18207
rect 18739 18173 18751 18207
rect 18693 18167 18751 18173
rect 15194 18096 15200 18148
rect 15252 18136 15258 18148
rect 16390 18136 16396 18148
rect 15252 18108 16396 18136
rect 15252 18096 15258 18108
rect 16390 18096 16396 18108
rect 16448 18096 16454 18148
rect 14734 18068 14740 18080
rect 13924 18040 14740 18068
rect 14734 18028 14740 18040
rect 14792 18028 14798 18080
rect 14921 18071 14979 18077
rect 14921 18037 14933 18071
rect 14967 18068 14979 18071
rect 15286 18068 15292 18080
rect 14967 18040 15292 18068
rect 14967 18037 14979 18040
rect 14921 18031 14979 18037
rect 15286 18028 15292 18040
rect 15344 18028 15350 18080
rect 15746 18028 15752 18080
rect 15804 18068 15810 18080
rect 16206 18068 16212 18080
rect 15804 18040 16212 18068
rect 15804 18028 15810 18040
rect 16206 18028 16212 18040
rect 16264 18028 16270 18080
rect 16574 18028 16580 18080
rect 16632 18068 16638 18080
rect 17681 18071 17739 18077
rect 17681 18068 17693 18071
rect 16632 18040 17693 18068
rect 16632 18028 16638 18040
rect 17681 18037 17693 18040
rect 17727 18037 17739 18071
rect 18708 18068 18736 18167
rect 20640 18145 20668 18244
rect 20809 18241 20821 18275
rect 20855 18241 20867 18275
rect 20809 18235 20867 18241
rect 20073 18139 20131 18145
rect 20073 18105 20085 18139
rect 20119 18136 20131 18139
rect 20625 18139 20683 18145
rect 20119 18108 20576 18136
rect 20119 18105 20131 18108
rect 20073 18099 20131 18105
rect 18966 18068 18972 18080
rect 18708 18040 18972 18068
rect 17681 18031 17739 18037
rect 18966 18028 18972 18040
rect 19024 18028 19030 18080
rect 20548 18068 20576 18108
rect 20625 18105 20637 18139
rect 20671 18105 20683 18139
rect 20625 18099 20683 18105
rect 20714 18068 20720 18080
rect 20548 18040 20720 18068
rect 20714 18028 20720 18040
rect 20772 18028 20778 18080
rect 21450 18028 21456 18080
rect 21508 18028 21514 18080
rect 1104 17978 21896 18000
rect 1104 17926 3549 17978
rect 3601 17926 3613 17978
rect 3665 17926 3677 17978
rect 3729 17926 3741 17978
rect 3793 17926 3805 17978
rect 3857 17926 8747 17978
rect 8799 17926 8811 17978
rect 8863 17926 8875 17978
rect 8927 17926 8939 17978
rect 8991 17926 9003 17978
rect 9055 17926 13945 17978
rect 13997 17926 14009 17978
rect 14061 17926 14073 17978
rect 14125 17926 14137 17978
rect 14189 17926 14201 17978
rect 14253 17926 19143 17978
rect 19195 17926 19207 17978
rect 19259 17926 19271 17978
rect 19323 17926 19335 17978
rect 19387 17926 19399 17978
rect 19451 17926 21896 17978
rect 1104 17904 21896 17926
rect 1762 17824 1768 17876
rect 1820 17864 1826 17876
rect 6086 17864 6092 17876
rect 1820 17836 6092 17864
rect 1820 17824 1826 17836
rect 6086 17824 6092 17836
rect 6144 17824 6150 17876
rect 6178 17824 6184 17876
rect 6236 17864 6242 17876
rect 6236 17836 7144 17864
rect 6236 17824 6242 17836
rect 1581 17799 1639 17805
rect 1581 17765 1593 17799
rect 1627 17796 1639 17799
rect 2498 17796 2504 17808
rect 1627 17768 2504 17796
rect 1627 17765 1639 17768
rect 1581 17759 1639 17765
rect 2498 17756 2504 17768
rect 2556 17756 2562 17808
rect 6730 17756 6736 17808
rect 6788 17756 6794 17808
rect 1765 17731 1823 17737
rect 1765 17697 1777 17731
rect 1811 17728 1823 17731
rect 2038 17728 2044 17740
rect 1811 17700 2044 17728
rect 1811 17697 1823 17700
rect 1765 17691 1823 17697
rect 2038 17688 2044 17700
rect 2096 17688 2102 17740
rect 2406 17688 2412 17740
rect 2464 17688 2470 17740
rect 2682 17688 2688 17740
rect 2740 17688 2746 17740
rect 2823 17731 2881 17737
rect 2823 17697 2835 17731
rect 2869 17728 2881 17731
rect 4062 17728 4068 17740
rect 2869 17700 4068 17728
rect 2869 17697 2881 17700
rect 2823 17691 2881 17697
rect 4062 17688 4068 17700
rect 4120 17688 4126 17740
rect 5718 17728 5724 17740
rect 4172 17700 5724 17728
rect 1397 17663 1455 17669
rect 1397 17629 1409 17663
rect 1443 17660 1455 17663
rect 1670 17660 1676 17672
rect 1443 17632 1676 17660
rect 1443 17629 1455 17632
rect 1397 17623 1455 17629
rect 1670 17620 1676 17632
rect 1728 17620 1734 17672
rect 1949 17663 2007 17669
rect 1949 17629 1961 17663
rect 1995 17660 2007 17663
rect 2130 17660 2136 17672
rect 1995 17632 2136 17660
rect 1995 17629 2007 17632
rect 1949 17623 2007 17629
rect 2130 17620 2136 17632
rect 2188 17620 2194 17672
rect 2958 17620 2964 17672
rect 3016 17620 3022 17672
rect 3694 17620 3700 17672
rect 3752 17660 3758 17672
rect 4172 17660 4200 17700
rect 5718 17688 5724 17700
rect 5776 17688 5782 17740
rect 7006 17688 7012 17740
rect 7064 17688 7070 17740
rect 3752 17632 4200 17660
rect 3752 17620 3758 17632
rect 4246 17620 4252 17672
rect 4304 17660 4310 17672
rect 4706 17660 4712 17672
rect 4304 17632 4712 17660
rect 4304 17620 4310 17632
rect 4706 17620 4712 17632
rect 4764 17620 4770 17672
rect 4801 17663 4859 17669
rect 4801 17629 4813 17663
rect 4847 17629 4859 17663
rect 4801 17623 4859 17629
rect 4816 17592 4844 17623
rect 5902 17620 5908 17672
rect 5960 17660 5966 17672
rect 5995 17663 6053 17669
rect 5995 17660 6007 17663
rect 5960 17632 6007 17660
rect 5960 17620 5966 17632
rect 5995 17629 6007 17632
rect 6041 17660 6053 17663
rect 7024 17660 7052 17688
rect 6041 17632 7052 17660
rect 7116 17650 7144 17836
rect 8570 17824 8576 17876
rect 8628 17864 8634 17876
rect 8628 17836 9674 17864
rect 8628 17824 8634 17836
rect 8665 17799 8723 17805
rect 8665 17765 8677 17799
rect 8711 17765 8723 17799
rect 9646 17796 9674 17836
rect 9950 17824 9956 17876
rect 10008 17824 10014 17876
rect 10042 17824 10048 17876
rect 10100 17864 10106 17876
rect 10100 17836 11376 17864
rect 10100 17824 10106 17836
rect 10060 17796 10088 17824
rect 9646 17768 10088 17796
rect 11348 17796 11376 17836
rect 12066 17824 12072 17876
rect 12124 17864 12130 17876
rect 12894 17864 12900 17876
rect 12124 17836 12900 17864
rect 12124 17824 12130 17836
rect 12894 17824 12900 17836
rect 12952 17864 12958 17876
rect 12952 17836 13308 17864
rect 12952 17824 12958 17836
rect 11348 17768 12664 17796
rect 8665 17759 8723 17765
rect 7196 17740 7248 17746
rect 7196 17682 7248 17688
rect 7466 17660 7472 17672
rect 7282 17650 7472 17660
rect 7116 17632 7472 17650
rect 6041 17629 6053 17632
rect 5995 17623 6053 17629
rect 7116 17622 7310 17632
rect 7466 17620 7472 17632
rect 7524 17620 7530 17672
rect 7558 17620 7564 17672
rect 7616 17660 7622 17672
rect 7653 17663 7711 17669
rect 7653 17660 7665 17663
rect 7616 17632 7665 17660
rect 7616 17620 7622 17632
rect 7653 17629 7665 17632
rect 7699 17629 7711 17663
rect 7653 17623 7711 17629
rect 7745 17663 7803 17669
rect 7745 17629 7757 17663
rect 7791 17660 7803 17663
rect 7834 17660 7840 17672
rect 7791 17632 7840 17660
rect 7791 17629 7803 17632
rect 7745 17623 7803 17629
rect 7834 17620 7840 17632
rect 7892 17620 7898 17672
rect 8110 17620 8116 17672
rect 8168 17620 8174 17672
rect 8294 17620 8300 17672
rect 8352 17660 8358 17672
rect 8680 17660 8708 17759
rect 12636 17740 12664 17768
rect 11790 17688 11796 17740
rect 11848 17728 11854 17740
rect 11974 17728 11980 17740
rect 11848 17700 11980 17728
rect 11848 17688 11854 17700
rect 11974 17688 11980 17700
rect 12032 17688 12038 17740
rect 12618 17688 12624 17740
rect 12676 17688 12682 17740
rect 13280 17728 13308 17836
rect 15930 17824 15936 17876
rect 15988 17864 15994 17876
rect 16114 17864 16120 17876
rect 15988 17836 16120 17864
rect 15988 17824 15994 17836
rect 16114 17824 16120 17836
rect 16172 17824 16178 17876
rect 20898 17824 20904 17876
rect 20956 17824 20962 17876
rect 20990 17824 20996 17876
rect 21048 17824 21054 17876
rect 13633 17799 13691 17805
rect 13633 17765 13645 17799
rect 13679 17796 13691 17799
rect 14737 17799 14795 17805
rect 14737 17796 14749 17799
rect 13679 17768 14749 17796
rect 13679 17765 13691 17768
rect 13633 17759 13691 17765
rect 14737 17765 14749 17768
rect 14783 17765 14795 17799
rect 14737 17759 14795 17765
rect 19705 17799 19763 17805
rect 19705 17765 19717 17799
rect 19751 17796 19763 17799
rect 20806 17796 20812 17808
rect 19751 17768 20812 17796
rect 19751 17765 19763 17768
rect 19705 17759 19763 17765
rect 20806 17756 20812 17768
rect 20864 17756 20870 17808
rect 16212 17740 16264 17746
rect 15013 17731 15071 17737
rect 15013 17728 15025 17731
rect 13280 17700 15025 17728
rect 15013 17697 15025 17700
rect 15059 17697 15071 17731
rect 15013 17691 15071 17697
rect 15286 17688 15292 17740
rect 15344 17688 15350 17740
rect 20073 17731 20131 17737
rect 20073 17697 20085 17731
rect 20119 17728 20131 17731
rect 20441 17731 20499 17737
rect 20441 17728 20453 17731
rect 20119 17700 20453 17728
rect 20119 17697 20131 17700
rect 20073 17691 20131 17697
rect 20441 17697 20453 17700
rect 20487 17697 20499 17731
rect 20441 17691 20499 17697
rect 20622 17688 20628 17740
rect 20680 17688 20686 17740
rect 20916 17728 20944 17824
rect 20916 17700 21128 17728
rect 8352 17632 8708 17660
rect 8352 17620 8358 17632
rect 8938 17620 8944 17672
rect 8996 17620 9002 17672
rect 9214 17660 9220 17672
rect 9175 17632 9220 17660
rect 9214 17620 9220 17632
rect 9272 17620 9278 17672
rect 10594 17660 10600 17672
rect 9876 17632 10600 17660
rect 6822 17592 6828 17604
rect 4816 17564 6828 17592
rect 6822 17552 6828 17564
rect 6880 17552 6886 17604
rect 7006 17552 7012 17604
rect 7064 17592 7070 17604
rect 7377 17595 7435 17601
rect 7377 17592 7389 17595
rect 7064 17564 7389 17592
rect 7064 17552 7070 17564
rect 7377 17561 7389 17564
rect 7423 17561 7435 17595
rect 9876 17592 9904 17632
rect 10594 17620 10600 17632
rect 10652 17620 10658 17672
rect 10686 17620 10692 17672
rect 10744 17620 10750 17672
rect 10963 17663 11021 17669
rect 10963 17629 10975 17663
rect 11009 17660 11021 17663
rect 11808 17660 11836 17688
rect 16212 17682 16264 17688
rect 12863 17663 12921 17669
rect 12863 17660 12875 17663
rect 11009 17632 11836 17660
rect 11900 17632 12875 17660
rect 11009 17629 11021 17632
rect 10963 17623 11021 17629
rect 7377 17555 7435 17561
rect 7484 17564 9904 17592
rect 1670 17484 1676 17536
rect 1728 17524 1734 17536
rect 2590 17524 2596 17536
rect 1728 17496 2596 17524
rect 1728 17484 1734 17496
rect 2590 17484 2596 17496
rect 2648 17484 2654 17536
rect 3050 17484 3056 17536
rect 3108 17524 3114 17536
rect 3605 17527 3663 17533
rect 3605 17524 3617 17527
rect 3108 17496 3617 17524
rect 3108 17484 3114 17496
rect 3605 17493 3617 17496
rect 3651 17493 3663 17527
rect 3605 17487 3663 17493
rect 4614 17484 4620 17536
rect 4672 17484 4678 17536
rect 4982 17484 4988 17536
rect 5040 17524 5046 17536
rect 5353 17527 5411 17533
rect 5353 17524 5365 17527
rect 5040 17496 5365 17524
rect 5040 17484 5046 17496
rect 5353 17493 5365 17496
rect 5399 17524 5411 17527
rect 5902 17524 5908 17536
rect 5399 17496 5908 17524
rect 5399 17493 5411 17496
rect 5353 17487 5411 17493
rect 5902 17484 5908 17496
rect 5960 17484 5966 17536
rect 6086 17484 6092 17536
rect 6144 17524 6150 17536
rect 7484 17524 7512 17564
rect 10410 17552 10416 17604
rect 10468 17552 10474 17604
rect 6144 17496 7512 17524
rect 6144 17484 6150 17496
rect 8110 17484 8116 17536
rect 8168 17524 8174 17536
rect 8481 17527 8539 17533
rect 8481 17524 8493 17527
rect 8168 17496 8493 17524
rect 8168 17484 8174 17496
rect 8481 17493 8493 17496
rect 8527 17493 8539 17527
rect 8481 17487 8539 17493
rect 8754 17484 8760 17536
rect 8812 17524 8818 17536
rect 10428 17524 10456 17552
rect 11900 17536 11928 17632
rect 12863 17629 12875 17632
rect 12909 17660 12921 17663
rect 13354 17660 13360 17672
rect 12909 17632 13360 17660
rect 12909 17629 12921 17632
rect 12863 17623 12921 17629
rect 13354 17620 13360 17632
rect 13412 17620 13418 17672
rect 14093 17663 14151 17669
rect 14093 17629 14105 17663
rect 14139 17629 14151 17663
rect 14093 17623 14151 17629
rect 14277 17663 14335 17669
rect 14277 17629 14289 17663
rect 14323 17660 14335 17663
rect 14458 17660 14464 17672
rect 14323 17632 14464 17660
rect 14323 17629 14335 17632
rect 14277 17623 14335 17629
rect 12618 17552 12624 17604
rect 12676 17592 12682 17604
rect 13078 17592 13084 17604
rect 12676 17564 13084 17592
rect 12676 17552 12682 17564
rect 13078 17552 13084 17564
rect 13136 17552 13142 17604
rect 8812 17496 10456 17524
rect 8812 17484 8818 17496
rect 11698 17484 11704 17536
rect 11756 17484 11762 17536
rect 11882 17484 11888 17536
rect 11940 17484 11946 17536
rect 12066 17484 12072 17536
rect 12124 17524 12130 17536
rect 12434 17524 12440 17536
rect 12124 17496 12440 17524
rect 12124 17484 12130 17496
rect 12434 17484 12440 17496
rect 12492 17484 12498 17536
rect 14108 17524 14136 17623
rect 14458 17620 14464 17632
rect 14516 17620 14522 17672
rect 15102 17620 15108 17672
rect 15160 17669 15166 17672
rect 15160 17663 15188 17669
rect 15176 17629 15188 17663
rect 15160 17623 15188 17629
rect 15160 17620 15166 17623
rect 17034 17620 17040 17672
rect 17092 17660 17098 17672
rect 17681 17663 17739 17669
rect 17681 17660 17693 17663
rect 17092 17632 17693 17660
rect 17092 17620 17098 17632
rect 17681 17629 17693 17632
rect 17727 17629 17739 17663
rect 17681 17623 17739 17629
rect 17954 17620 17960 17672
rect 18012 17620 18018 17672
rect 19058 17620 19064 17672
rect 19116 17660 19122 17672
rect 19429 17663 19487 17669
rect 19429 17660 19441 17663
rect 19116 17632 19441 17660
rect 19116 17620 19122 17632
rect 19429 17629 19441 17632
rect 19475 17629 19487 17663
rect 19429 17623 19487 17629
rect 19518 17620 19524 17672
rect 19576 17660 19582 17672
rect 19889 17663 19947 17669
rect 19889 17660 19901 17663
rect 19576 17632 19901 17660
rect 19576 17620 19582 17632
rect 19889 17629 19901 17632
rect 19935 17629 19947 17663
rect 19889 17623 19947 17629
rect 19981 17663 20039 17669
rect 19981 17629 19993 17663
rect 20027 17629 20039 17663
rect 19981 17623 20039 17629
rect 20349 17663 20407 17669
rect 20349 17629 20361 17663
rect 20395 17629 20407 17663
rect 20349 17623 20407 17629
rect 16022 17552 16028 17604
rect 16080 17592 16086 17604
rect 16485 17595 16543 17601
rect 16485 17592 16497 17595
rect 16080 17564 16497 17592
rect 16080 17552 16086 17564
rect 16485 17561 16497 17564
rect 16531 17561 16543 17595
rect 16485 17555 16543 17561
rect 16574 17552 16580 17604
rect 16632 17552 16638 17604
rect 16945 17595 17003 17601
rect 16945 17561 16957 17595
rect 16991 17592 17003 17595
rect 17770 17592 17776 17604
rect 16991 17564 17776 17592
rect 16991 17561 17003 17564
rect 16945 17555 17003 17561
rect 17770 17552 17776 17564
rect 17828 17552 17834 17604
rect 19996 17592 20024 17623
rect 19260 17564 20024 17592
rect 14826 17524 14832 17536
rect 14108 17496 14832 17524
rect 14826 17484 14832 17496
rect 14884 17484 14890 17536
rect 15286 17484 15292 17536
rect 15344 17524 15350 17536
rect 15933 17527 15991 17533
rect 15933 17524 15945 17527
rect 15344 17496 15945 17524
rect 15344 17484 15350 17496
rect 15933 17493 15945 17496
rect 15979 17493 15991 17527
rect 15933 17487 15991 17493
rect 16114 17484 16120 17536
rect 16172 17524 16178 17536
rect 16209 17527 16267 17533
rect 16209 17524 16221 17527
rect 16172 17496 16221 17524
rect 16172 17484 16178 17496
rect 16209 17493 16221 17496
rect 16255 17493 16267 17527
rect 16209 17487 16267 17493
rect 16666 17484 16672 17536
rect 16724 17524 16730 17536
rect 17218 17524 17224 17536
rect 16724 17496 17224 17524
rect 16724 17484 16730 17496
rect 17218 17484 17224 17496
rect 17276 17484 17282 17536
rect 17310 17484 17316 17536
rect 17368 17484 17374 17536
rect 17494 17484 17500 17536
rect 17552 17484 17558 17536
rect 17862 17484 17868 17536
rect 17920 17524 17926 17536
rect 19260 17533 19288 17564
rect 20364 17536 20392 17623
rect 20530 17620 20536 17672
rect 20588 17660 20594 17672
rect 21100 17669 21128 17700
rect 20901 17663 20959 17669
rect 20901 17660 20913 17663
rect 20588 17632 20913 17660
rect 20588 17620 20594 17632
rect 20901 17629 20913 17632
rect 20947 17629 20959 17663
rect 20901 17623 20959 17629
rect 21085 17663 21143 17669
rect 21085 17629 21097 17663
rect 21131 17629 21143 17663
rect 21085 17623 21143 17629
rect 21266 17620 21272 17672
rect 21324 17620 21330 17672
rect 18693 17527 18751 17533
rect 18693 17524 18705 17527
rect 17920 17496 18705 17524
rect 17920 17484 17926 17496
rect 18693 17493 18705 17496
rect 18739 17493 18751 17527
rect 18693 17487 18751 17493
rect 19245 17527 19303 17533
rect 19245 17493 19257 17527
rect 19291 17493 19303 17527
rect 19245 17487 19303 17493
rect 20346 17484 20352 17536
rect 20404 17484 20410 17536
rect 20625 17527 20683 17533
rect 20625 17493 20637 17527
rect 20671 17524 20683 17527
rect 20898 17524 20904 17536
rect 20671 17496 20904 17524
rect 20671 17493 20683 17496
rect 20625 17487 20683 17493
rect 20898 17484 20904 17496
rect 20956 17484 20962 17536
rect 21453 17527 21511 17533
rect 21453 17493 21465 17527
rect 21499 17524 21511 17527
rect 22186 17524 22192 17536
rect 21499 17496 22192 17524
rect 21499 17493 21511 17496
rect 21453 17487 21511 17493
rect 22186 17484 22192 17496
rect 22244 17484 22250 17536
rect 1104 17434 22056 17456
rect 1104 17382 6148 17434
rect 6200 17382 6212 17434
rect 6264 17382 6276 17434
rect 6328 17382 6340 17434
rect 6392 17382 6404 17434
rect 6456 17382 11346 17434
rect 11398 17382 11410 17434
rect 11462 17382 11474 17434
rect 11526 17382 11538 17434
rect 11590 17382 11602 17434
rect 11654 17382 16544 17434
rect 16596 17382 16608 17434
rect 16660 17382 16672 17434
rect 16724 17382 16736 17434
rect 16788 17382 16800 17434
rect 16852 17382 21742 17434
rect 21794 17382 21806 17434
rect 21858 17382 21870 17434
rect 21922 17382 21934 17434
rect 21986 17382 21998 17434
rect 22050 17382 22056 17434
rect 1104 17360 22056 17382
rect 1673 17323 1731 17329
rect 1673 17289 1685 17323
rect 1719 17320 1731 17323
rect 1762 17320 1768 17332
rect 1719 17292 1768 17320
rect 1719 17289 1731 17292
rect 1673 17283 1731 17289
rect 1762 17280 1768 17292
rect 1820 17280 1826 17332
rect 2682 17320 2688 17332
rect 2332 17292 2688 17320
rect 1578 17212 1584 17264
rect 1636 17212 1642 17264
rect 2332 17116 2360 17292
rect 2682 17280 2688 17292
rect 2740 17320 2746 17332
rect 3421 17323 3479 17329
rect 2740 17292 3372 17320
rect 2740 17280 2746 17292
rect 3344 17252 3372 17292
rect 3421 17289 3433 17323
rect 3467 17320 3479 17323
rect 3878 17320 3884 17332
rect 3467 17292 3884 17320
rect 3467 17289 3479 17292
rect 3421 17283 3479 17289
rect 3878 17280 3884 17292
rect 3936 17280 3942 17332
rect 3970 17280 3976 17332
rect 4028 17320 4034 17332
rect 4982 17320 4988 17332
rect 4028 17292 4988 17320
rect 4028 17280 4034 17292
rect 4982 17280 4988 17292
rect 5040 17280 5046 17332
rect 7466 17280 7472 17332
rect 7524 17320 7530 17332
rect 7524 17292 7742 17320
rect 7524 17280 7530 17292
rect 3694 17252 3700 17264
rect 3344 17224 3700 17252
rect 3694 17212 3700 17224
rect 3752 17212 3758 17264
rect 7006 17212 7012 17264
rect 7064 17252 7070 17264
rect 7193 17255 7251 17261
rect 7193 17252 7205 17255
rect 7064 17224 7205 17252
rect 7064 17212 7070 17224
rect 7193 17221 7205 17224
rect 7239 17221 7251 17255
rect 7193 17215 7251 17221
rect 7558 17212 7564 17264
rect 7616 17212 7622 17264
rect 7714 17252 7742 17292
rect 7834 17280 7840 17332
rect 7892 17320 7898 17332
rect 8481 17323 8539 17329
rect 8481 17320 8493 17323
rect 7892 17292 8493 17320
rect 7892 17280 7898 17292
rect 8481 17289 8493 17292
rect 8527 17289 8539 17323
rect 8481 17283 8539 17289
rect 10226 17280 10232 17332
rect 10284 17320 10290 17332
rect 12986 17320 12992 17332
rect 10284 17292 11008 17320
rect 10284 17280 10290 17292
rect 10980 17264 11008 17292
rect 12176 17292 12992 17320
rect 7929 17255 7987 17261
rect 7929 17252 7941 17255
rect 7714 17224 7941 17252
rect 7929 17221 7941 17224
rect 7975 17221 7987 17255
rect 7929 17215 7987 17221
rect 8110 17212 8116 17264
rect 8168 17252 8174 17264
rect 8297 17255 8355 17261
rect 8297 17252 8309 17255
rect 8168 17224 8309 17252
rect 8168 17212 8174 17224
rect 8297 17221 8309 17224
rect 8343 17221 8355 17255
rect 8297 17215 8355 17221
rect 8570 17212 8576 17264
rect 8628 17212 8634 17264
rect 9766 17212 9772 17264
rect 9824 17252 9830 17264
rect 9824 17224 10180 17252
rect 9824 17212 9830 17224
rect 10152 17214 10180 17224
rect 10211 17217 10269 17223
rect 10211 17214 10223 17217
rect 2651 17197 2709 17203
rect 2651 17196 2663 17197
rect 2590 17144 2596 17196
rect 2648 17163 2663 17196
rect 2697 17163 2709 17197
rect 2648 17157 2709 17163
rect 2648 17156 2694 17157
rect 2648 17144 2654 17156
rect 2774 17144 2780 17196
rect 2832 17184 2838 17196
rect 3789 17187 3847 17193
rect 3789 17184 3801 17187
rect 2832 17156 3801 17184
rect 2832 17144 2838 17156
rect 3789 17153 3801 17156
rect 3835 17153 3847 17187
rect 3789 17147 3847 17153
rect 3896 17156 4108 17184
rect 2409 17119 2467 17125
rect 2409 17116 2421 17119
rect 2332 17088 2421 17116
rect 2409 17085 2421 17088
rect 2455 17085 2467 17119
rect 2409 17079 2467 17085
rect 3326 17076 3332 17128
rect 3384 17116 3390 17128
rect 3896 17116 3924 17156
rect 3384 17088 3924 17116
rect 3973 17119 4031 17125
rect 3384 17076 3390 17088
rect 3973 17085 3985 17119
rect 4019 17085 4031 17119
rect 4080 17116 4108 17156
rect 4982 17144 4988 17196
rect 5040 17144 5046 17196
rect 5905 17187 5963 17193
rect 5905 17153 5917 17187
rect 5951 17153 5963 17187
rect 5905 17147 5963 17153
rect 4433 17119 4491 17125
rect 4433 17116 4445 17119
rect 4080 17088 4445 17116
rect 3973 17079 4031 17085
rect 4433 17085 4445 17088
rect 4479 17085 4491 17119
rect 4706 17116 4712 17128
rect 4433 17079 4491 17085
rect 4538 17088 4712 17116
rect 1854 17008 1860 17060
rect 1912 17048 1918 17060
rect 2314 17048 2320 17060
rect 1912 17020 2320 17048
rect 1912 17008 1918 17020
rect 2314 17008 2320 17020
rect 2372 17008 2378 17060
rect 3786 17048 3792 17060
rect 3344 17020 3792 17048
rect 1210 16940 1216 16992
rect 1268 16980 1274 16992
rect 3344 16980 3372 17020
rect 3786 17008 3792 17020
rect 3844 17008 3850 17060
rect 3988 16992 4016 17079
rect 4338 17008 4344 17060
rect 4396 17048 4402 17060
rect 4538 17048 4566 17088
rect 4706 17076 4712 17088
rect 4764 17076 4770 17128
rect 4826 17119 4884 17125
rect 4826 17085 4838 17119
rect 4872 17116 4884 17119
rect 5534 17116 5540 17128
rect 4872 17088 5540 17116
rect 4872 17085 4884 17088
rect 4826 17079 4884 17085
rect 5534 17076 5540 17088
rect 5592 17076 5598 17128
rect 5920 17116 5948 17147
rect 7466 17144 7472 17196
rect 7524 17184 7530 17196
rect 8588 17184 8616 17212
rect 10152 17186 10223 17214
rect 7524 17156 8616 17184
rect 10211 17183 10223 17186
rect 10257 17183 10269 17217
rect 10962 17212 10968 17264
rect 11020 17212 11026 17264
rect 12176 17252 12204 17292
rect 12986 17280 12992 17292
rect 13044 17280 13050 17332
rect 15010 17280 15016 17332
rect 15068 17280 15074 17332
rect 15286 17280 15292 17332
rect 15344 17280 15350 17332
rect 16206 17280 16212 17332
rect 16264 17280 16270 17332
rect 16850 17280 16856 17332
rect 16908 17320 16914 17332
rect 17310 17320 17316 17332
rect 16908 17292 17316 17320
rect 16908 17280 16914 17292
rect 17310 17280 17316 17292
rect 17368 17280 17374 17332
rect 17678 17280 17684 17332
rect 17736 17320 17742 17332
rect 20625 17323 20683 17329
rect 17736 17292 18828 17320
rect 17736 17280 17742 17292
rect 15304 17252 15332 17280
rect 11072 17224 12204 17252
rect 10211 17177 10269 17183
rect 7524 17144 7530 17156
rect 10594 17144 10600 17196
rect 10652 17184 10658 17196
rect 11072 17184 11100 17224
rect 10652 17156 11100 17184
rect 10652 17144 10658 17156
rect 11238 17144 11244 17196
rect 11296 17184 11302 17196
rect 12176 17193 12204 17224
rect 14844 17224 15332 17252
rect 14844 17193 14872 17224
rect 15654 17212 15660 17264
rect 15712 17212 15718 17264
rect 11517 17187 11575 17193
rect 11517 17184 11529 17187
rect 11296 17156 11529 17184
rect 11296 17144 11302 17156
rect 11517 17153 11529 17156
rect 11563 17153 11575 17187
rect 11517 17147 11575 17153
rect 12161 17187 12219 17193
rect 12161 17153 12173 17187
rect 12207 17153 12219 17187
rect 12161 17147 12219 17153
rect 14829 17187 14887 17193
rect 14829 17153 14841 17187
rect 14875 17153 14887 17187
rect 15439 17187 15497 17193
rect 15439 17184 15451 17187
rect 14829 17147 14887 17153
rect 14934 17156 15451 17184
rect 5994 17116 6000 17128
rect 5920 17088 6000 17116
rect 5994 17076 6000 17088
rect 6052 17076 6058 17128
rect 6546 17076 6552 17128
rect 6604 17116 6610 17128
rect 6604 17088 7038 17116
rect 6604 17076 6610 17088
rect 9858 17076 9864 17128
rect 9916 17116 9922 17128
rect 9953 17119 10011 17125
rect 9953 17116 9965 17119
rect 9916 17088 9965 17116
rect 9916 17076 9922 17088
rect 9953 17085 9965 17088
rect 9999 17085 10011 17119
rect 9953 17079 10011 17085
rect 4396 17020 4566 17048
rect 4396 17008 4402 17020
rect 5442 17008 5448 17060
rect 5500 17048 5506 17060
rect 5721 17051 5779 17057
rect 5721 17048 5733 17051
rect 5500 17020 5733 17048
rect 5500 17008 5506 17020
rect 5721 17017 5733 17020
rect 5767 17017 5779 17051
rect 5721 17011 5779 17017
rect 1268 16952 3372 16980
rect 1268 16940 1274 16952
rect 3418 16940 3424 16992
rect 3476 16980 3482 16992
rect 3970 16980 3976 16992
rect 3476 16952 3976 16980
rect 3476 16940 3482 16952
rect 3970 16940 3976 16952
rect 4028 16940 4034 16992
rect 4062 16940 4068 16992
rect 4120 16980 4126 16992
rect 5629 16983 5687 16989
rect 5629 16980 5641 16983
rect 4120 16952 5641 16980
rect 4120 16940 4126 16952
rect 5629 16949 5641 16952
rect 5675 16949 5687 16983
rect 5629 16943 5687 16949
rect 8938 16940 8944 16992
rect 8996 16980 9002 16992
rect 9490 16980 9496 16992
rect 8996 16952 9496 16980
rect 8996 16940 9002 16952
rect 9490 16940 9496 16952
rect 9548 16940 9554 16992
rect 9968 16980 9996 17079
rect 10870 17076 10876 17128
rect 10928 17116 10934 17128
rect 13262 17125 13268 17128
rect 12345 17119 12403 17125
rect 12345 17116 12357 17119
rect 10928 17088 12357 17116
rect 10928 17076 10934 17088
rect 12345 17085 12357 17088
rect 12391 17085 12403 17119
rect 13081 17119 13139 17125
rect 13081 17116 13093 17119
rect 12345 17079 12403 17085
rect 12912 17088 13093 17116
rect 12802 17008 12808 17060
rect 12860 17008 12866 17060
rect 10410 16980 10416 16992
rect 9968 16952 10416 16980
rect 10410 16940 10416 16952
rect 10468 16980 10474 16992
rect 10686 16980 10692 16992
rect 10468 16952 10692 16980
rect 10468 16940 10474 16952
rect 10686 16940 10692 16952
rect 10744 16940 10750 16992
rect 10962 16940 10968 16992
rect 11020 16940 11026 16992
rect 11146 16940 11152 16992
rect 11204 16980 11210 16992
rect 11701 16983 11759 16989
rect 11701 16980 11713 16983
rect 11204 16952 11713 16980
rect 11204 16940 11210 16952
rect 11701 16949 11713 16952
rect 11747 16949 11759 16983
rect 11701 16943 11759 16949
rect 12434 16940 12440 16992
rect 12492 16980 12498 16992
rect 12618 16980 12624 16992
rect 12492 16952 12624 16980
rect 12492 16940 12498 16952
rect 12618 16940 12624 16952
rect 12676 16940 12682 16992
rect 12912 16980 12940 17088
rect 13081 17085 13093 17088
rect 13127 17085 13139 17119
rect 13081 17079 13139 17085
rect 13219 17119 13268 17125
rect 13219 17085 13231 17119
rect 13265 17085 13268 17119
rect 13219 17079 13268 17085
rect 13262 17076 13268 17079
rect 13320 17076 13326 17128
rect 13354 17076 13360 17128
rect 13412 17076 13418 17128
rect 14734 17076 14740 17128
rect 14792 17116 14798 17128
rect 14934 17116 14962 17156
rect 15439 17153 15451 17156
rect 15485 17153 15497 17187
rect 15672 17184 15700 17212
rect 16669 17187 16727 17193
rect 16669 17184 16681 17187
rect 15672 17156 16681 17184
rect 15439 17147 15497 17153
rect 16669 17153 16681 17156
rect 16715 17153 16727 17187
rect 16669 17147 16727 17153
rect 17586 17144 17592 17196
rect 17644 17144 17650 17196
rect 14792 17088 14962 17116
rect 15197 17119 15255 17125
rect 14792 17076 14798 17088
rect 15197 17085 15209 17119
rect 15243 17085 15255 17119
rect 15197 17079 15255 17085
rect 15212 17048 15240 17079
rect 16850 17076 16856 17128
rect 16908 17076 16914 17128
rect 17678 17076 17684 17128
rect 17736 17125 17742 17128
rect 17736 17119 17764 17125
rect 17752 17085 17764 17119
rect 17736 17079 17764 17085
rect 17736 17076 17742 17079
rect 17860 17076 17866 17128
rect 17918 17076 17924 17128
rect 18800 17125 18828 17292
rect 20625 17289 20637 17323
rect 20671 17289 20683 17323
rect 20625 17283 20683 17289
rect 20717 17323 20775 17329
rect 20717 17289 20729 17323
rect 20763 17289 20775 17323
rect 20717 17283 20775 17289
rect 20640 17252 20668 17283
rect 19168 17224 20668 17252
rect 20732 17252 20760 17283
rect 20898 17280 20904 17332
rect 20956 17320 20962 17332
rect 20956 17292 21312 17320
rect 20956 17280 20962 17292
rect 20732 17224 21220 17252
rect 19168 17193 19196 17224
rect 19518 17193 19524 17196
rect 19153 17187 19211 17193
rect 19153 17153 19165 17187
rect 19199 17153 19211 17187
rect 19512 17184 19524 17193
rect 19479 17156 19524 17184
rect 19153 17147 19211 17153
rect 19512 17147 19524 17156
rect 19518 17144 19524 17147
rect 19576 17144 19582 17196
rect 20714 17144 20720 17196
rect 20772 17184 20778 17196
rect 21192 17193 21220 17224
rect 21284 17193 21312 17292
rect 20901 17187 20959 17193
rect 20901 17184 20913 17187
rect 20772 17156 20913 17184
rect 20772 17144 20778 17156
rect 20901 17153 20913 17156
rect 20947 17153 20959 17187
rect 20901 17147 20959 17153
rect 20993 17187 21051 17193
rect 20993 17153 21005 17187
rect 21039 17153 21051 17187
rect 20993 17147 21051 17153
rect 21177 17187 21235 17193
rect 21177 17153 21189 17187
rect 21223 17153 21235 17187
rect 21177 17147 21235 17153
rect 21269 17187 21327 17193
rect 21269 17153 21281 17187
rect 21315 17153 21327 17187
rect 21269 17147 21327 17153
rect 18785 17119 18843 17125
rect 18785 17085 18797 17119
rect 18831 17085 18843 17119
rect 18785 17079 18843 17085
rect 18966 17076 18972 17128
rect 19024 17116 19030 17128
rect 19245 17119 19303 17125
rect 19245 17116 19257 17119
rect 19024 17088 19257 17116
rect 19024 17076 19030 17088
rect 19245 17085 19257 17088
rect 19291 17085 19303 17119
rect 19245 17079 19303 17085
rect 15212 17020 15332 17048
rect 15304 16992 15332 17020
rect 17310 17008 17316 17060
rect 17368 17008 17374 17060
rect 20346 17008 20352 17060
rect 20404 17048 20410 17060
rect 21008 17048 21036 17147
rect 20404 17020 21036 17048
rect 20404 17008 20410 17020
rect 13538 16980 13544 16992
rect 12912 16952 13544 16980
rect 13538 16940 13544 16952
rect 13596 16940 13602 16992
rect 14001 16983 14059 16989
rect 14001 16949 14013 16983
rect 14047 16980 14059 16983
rect 14274 16980 14280 16992
rect 14047 16952 14280 16980
rect 14047 16949 14059 16952
rect 14001 16943 14059 16949
rect 14274 16940 14280 16952
rect 14332 16940 14338 16992
rect 15286 16940 15292 16992
rect 15344 16940 15350 16992
rect 16206 16940 16212 16992
rect 16264 16980 16270 16992
rect 17034 16980 17040 16992
rect 16264 16952 17040 16980
rect 16264 16940 16270 16952
rect 17034 16940 17040 16952
rect 17092 16940 17098 16992
rect 18506 16940 18512 16992
rect 18564 16940 18570 16992
rect 18969 16983 19027 16989
rect 18969 16949 18981 16983
rect 19015 16980 19027 16983
rect 19518 16980 19524 16992
rect 19015 16952 19524 16980
rect 19015 16949 19027 16952
rect 18969 16943 19027 16949
rect 19518 16940 19524 16952
rect 19576 16940 19582 16992
rect 20162 16940 20168 16992
rect 20220 16980 20226 16992
rect 20530 16980 20536 16992
rect 20220 16952 20536 16980
rect 20220 16940 20226 16952
rect 20530 16940 20536 16952
rect 20588 16940 20594 16992
rect 20622 16940 20628 16992
rect 20680 16980 20686 16992
rect 21085 16983 21143 16989
rect 21085 16980 21097 16983
rect 20680 16952 21097 16980
rect 20680 16940 20686 16952
rect 21085 16949 21097 16952
rect 21131 16949 21143 16983
rect 21085 16943 21143 16949
rect 21450 16940 21456 16992
rect 21508 16940 21514 16992
rect 1104 16890 21896 16912
rect 1104 16838 3549 16890
rect 3601 16838 3613 16890
rect 3665 16838 3677 16890
rect 3729 16838 3741 16890
rect 3793 16838 3805 16890
rect 3857 16838 8747 16890
rect 8799 16838 8811 16890
rect 8863 16838 8875 16890
rect 8927 16838 8939 16890
rect 8991 16838 9003 16890
rect 9055 16838 13945 16890
rect 13997 16838 14009 16890
rect 14061 16838 14073 16890
rect 14125 16838 14137 16890
rect 14189 16838 14201 16890
rect 14253 16838 19143 16890
rect 19195 16838 19207 16890
rect 19259 16838 19271 16890
rect 19323 16838 19335 16890
rect 19387 16838 19399 16890
rect 19451 16838 21896 16890
rect 1104 16816 21896 16838
rect 1946 16736 1952 16788
rect 2004 16736 2010 16788
rect 2869 16779 2927 16785
rect 2869 16745 2881 16779
rect 2915 16776 2927 16779
rect 2958 16776 2964 16788
rect 2915 16748 2964 16776
rect 2915 16745 2927 16748
rect 2869 16739 2927 16745
rect 2958 16736 2964 16748
rect 3016 16736 3022 16788
rect 3602 16736 3608 16788
rect 3660 16776 3666 16788
rect 4525 16779 4583 16785
rect 4525 16776 4537 16779
rect 3660 16748 4537 16776
rect 3660 16736 3666 16748
rect 4525 16745 4537 16748
rect 4571 16745 4583 16779
rect 4525 16739 4583 16745
rect 6730 16736 6736 16788
rect 6788 16736 6794 16788
rect 6822 16736 6828 16788
rect 6880 16736 6886 16788
rect 7558 16736 7564 16788
rect 7616 16776 7622 16788
rect 8481 16779 8539 16785
rect 8481 16776 8493 16779
rect 7616 16748 8493 16776
rect 7616 16736 7622 16748
rect 8481 16745 8493 16748
rect 8527 16745 8539 16779
rect 12158 16776 12164 16788
rect 8481 16739 8539 16745
rect 10336 16748 12164 16776
rect 1964 16708 1992 16736
rect 1872 16680 1992 16708
rect 3988 16680 5212 16708
rect 1872 16649 1900 16680
rect 3988 16652 4016 16680
rect 1857 16643 1915 16649
rect 1857 16609 1869 16643
rect 1903 16609 1915 16643
rect 1857 16603 1915 16609
rect 3970 16600 3976 16652
rect 4028 16600 4034 16652
rect 4890 16600 4896 16652
rect 4948 16640 4954 16652
rect 4985 16643 5043 16649
rect 4985 16640 4997 16643
rect 4948 16612 4997 16640
rect 4948 16600 4954 16612
rect 4985 16609 4997 16612
rect 5031 16609 5043 16643
rect 4985 16603 5043 16609
rect 2131 16575 2189 16581
rect 2131 16541 2143 16575
rect 2177 16572 2189 16575
rect 2222 16572 2228 16584
rect 2177 16544 2228 16572
rect 2177 16541 2189 16544
rect 2131 16535 2189 16541
rect 2222 16532 2228 16544
rect 2280 16532 2286 16584
rect 2590 16532 2596 16584
rect 2648 16572 2654 16584
rect 2774 16572 2780 16584
rect 2648 16544 2780 16572
rect 2648 16532 2654 16544
rect 2774 16532 2780 16544
rect 2832 16532 2838 16584
rect 3605 16575 3663 16581
rect 3605 16541 3617 16575
rect 3651 16572 3663 16575
rect 4338 16572 4344 16584
rect 3651 16544 4344 16572
rect 3651 16541 3663 16544
rect 3605 16535 3663 16541
rect 4338 16532 4344 16544
rect 4396 16532 4402 16584
rect 5184 16581 5212 16680
rect 5626 16600 5632 16652
rect 5684 16600 5690 16652
rect 5902 16600 5908 16652
rect 5960 16600 5966 16652
rect 6181 16643 6239 16649
rect 6181 16609 6193 16643
rect 6227 16640 6239 16643
rect 6748 16640 6776 16736
rect 7006 16708 7012 16720
rect 6227 16612 6776 16640
rect 6840 16680 7012 16708
rect 6227 16609 6239 16612
rect 6181 16603 6239 16609
rect 6086 16581 6092 16584
rect 4433 16575 4491 16581
rect 4433 16541 4445 16575
rect 4479 16541 4491 16575
rect 4433 16535 4491 16541
rect 5169 16575 5227 16581
rect 5169 16541 5181 16575
rect 5215 16541 5227 16575
rect 5169 16535 5227 16541
rect 6043 16575 6092 16581
rect 6043 16541 6055 16575
rect 6089 16541 6092 16575
rect 6043 16535 6092 16541
rect 474 16464 480 16516
rect 532 16504 538 16516
rect 3234 16504 3240 16516
rect 532 16476 3240 16504
rect 532 16464 538 16476
rect 3234 16464 3240 16476
rect 3292 16464 3298 16516
rect 3326 16464 3332 16516
rect 3384 16504 3390 16516
rect 3881 16507 3939 16513
rect 3881 16504 3893 16507
rect 3384 16476 3893 16504
rect 3384 16464 3390 16476
rect 3881 16473 3893 16476
rect 3927 16473 3939 16507
rect 3881 16467 3939 16473
rect 1486 16396 1492 16448
rect 1544 16436 1550 16448
rect 3421 16439 3479 16445
rect 3421 16436 3433 16439
rect 1544 16408 3433 16436
rect 1544 16396 1550 16408
rect 3421 16405 3433 16408
rect 3467 16405 3479 16439
rect 3421 16399 3479 16405
rect 3970 16396 3976 16448
rect 4028 16396 4034 16448
rect 4448 16436 4476 16535
rect 6086 16532 6092 16535
rect 6144 16532 6150 16584
rect 4522 16464 4528 16516
rect 4580 16504 4586 16516
rect 4706 16504 4712 16516
rect 4580 16476 4712 16504
rect 4580 16464 4586 16476
rect 4706 16464 4712 16476
rect 4764 16464 4770 16516
rect 6730 16464 6736 16516
rect 6788 16504 6794 16516
rect 6840 16504 6868 16680
rect 7006 16668 7012 16680
rect 7064 16668 7070 16720
rect 7469 16643 7527 16649
rect 7469 16640 7481 16643
rect 7024 16612 7481 16640
rect 7024 16584 7052 16612
rect 7469 16609 7481 16612
rect 7515 16609 7527 16643
rect 7469 16603 7527 16609
rect 8662 16600 8668 16652
rect 8720 16640 8726 16652
rect 10336 16649 10364 16748
rect 12158 16736 12164 16748
rect 12216 16736 12222 16788
rect 12710 16736 12716 16788
rect 12768 16776 12774 16788
rect 12768 16748 13308 16776
rect 12768 16736 12774 16748
rect 10686 16668 10692 16720
rect 10744 16708 10750 16720
rect 10965 16711 11023 16717
rect 10965 16708 10977 16711
rect 10744 16680 10977 16708
rect 10744 16668 10750 16680
rect 10965 16677 10977 16680
rect 11011 16677 11023 16711
rect 13280 16708 13308 16748
rect 13354 16736 13360 16788
rect 13412 16776 13418 16788
rect 13449 16779 13507 16785
rect 13449 16776 13461 16779
rect 13412 16748 13461 16776
rect 13412 16736 13418 16748
rect 13449 16745 13461 16748
rect 13495 16745 13507 16779
rect 15194 16776 15200 16788
rect 13449 16739 13507 16745
rect 13924 16748 15200 16776
rect 13924 16708 13952 16748
rect 15194 16736 15200 16748
rect 15252 16736 15258 16788
rect 15930 16776 15936 16788
rect 15580 16748 15936 16776
rect 15286 16708 15292 16720
rect 13280 16680 13952 16708
rect 14016 16680 15292 16708
rect 10965 16671 11023 16677
rect 8941 16643 8999 16649
rect 8941 16640 8953 16643
rect 8720 16612 8953 16640
rect 8720 16600 8726 16612
rect 8941 16609 8953 16612
rect 8987 16609 8999 16643
rect 8941 16603 8999 16609
rect 10321 16643 10379 16649
rect 10321 16609 10333 16643
rect 10367 16609 10379 16643
rect 10870 16640 10876 16652
rect 10321 16603 10379 16609
rect 10428 16612 10876 16640
rect 7006 16532 7012 16584
rect 7064 16532 7070 16584
rect 7711 16575 7769 16581
rect 7711 16572 7723 16575
rect 7116 16544 7723 16572
rect 6788 16476 6868 16504
rect 6788 16464 6794 16476
rect 6914 16464 6920 16516
rect 6972 16504 6978 16516
rect 7116 16513 7144 16544
rect 7711 16541 7723 16544
rect 7757 16541 7769 16575
rect 7711 16535 7769 16541
rect 9215 16575 9273 16581
rect 9215 16541 9227 16575
rect 9261 16572 9273 16575
rect 9306 16572 9312 16584
rect 9261 16544 9312 16572
rect 9261 16541 9273 16544
rect 9215 16535 9273 16541
rect 9306 16532 9312 16544
rect 9364 16532 9370 16584
rect 10134 16532 10140 16584
rect 10192 16572 10198 16584
rect 10428 16572 10456 16612
rect 10870 16600 10876 16612
rect 10928 16640 10934 16652
rect 11241 16643 11299 16649
rect 11241 16640 11253 16643
rect 10928 16612 11253 16640
rect 10928 16600 10934 16612
rect 11241 16609 11253 16612
rect 11287 16609 11299 16643
rect 11241 16603 11299 16609
rect 11517 16643 11575 16649
rect 11517 16609 11529 16643
rect 11563 16640 11575 16643
rect 11698 16640 11704 16652
rect 11563 16612 11704 16640
rect 11563 16609 11575 16612
rect 11517 16603 11575 16609
rect 11698 16600 11704 16612
rect 11756 16600 11762 16652
rect 10192 16544 10456 16572
rect 10192 16532 10198 16544
rect 10502 16532 10508 16584
rect 10560 16532 10566 16584
rect 11330 16532 11336 16584
rect 11388 16581 11394 16584
rect 11388 16575 11416 16581
rect 11404 16541 11416 16575
rect 11388 16535 11416 16541
rect 11388 16532 11394 16535
rect 12434 16532 12440 16584
rect 12492 16532 12498 16584
rect 12618 16532 12624 16584
rect 12676 16572 12682 16584
rect 12711 16575 12769 16581
rect 12711 16572 12723 16575
rect 12676 16544 12723 16572
rect 12676 16532 12682 16544
rect 12711 16541 12723 16544
rect 12757 16572 12769 16575
rect 14016 16572 14044 16680
rect 15286 16668 15292 16680
rect 15344 16668 15350 16720
rect 15580 16717 15608 16748
rect 15930 16736 15936 16748
rect 15988 16736 15994 16788
rect 16022 16736 16028 16788
rect 16080 16776 16086 16788
rect 16758 16776 16764 16788
rect 16080 16748 16764 16776
rect 16080 16736 16086 16748
rect 16758 16736 16764 16748
rect 16816 16736 16822 16788
rect 17865 16779 17923 16785
rect 17865 16776 17877 16779
rect 16868 16748 17877 16776
rect 15565 16711 15623 16717
rect 15565 16677 15577 16711
rect 15611 16677 15623 16711
rect 15565 16671 15623 16677
rect 14642 16600 14648 16652
rect 14700 16600 14706 16652
rect 14734 16600 14740 16652
rect 14792 16640 14798 16652
rect 15105 16643 15163 16649
rect 14792 16612 15056 16640
rect 14792 16600 14798 16612
rect 12757 16544 14044 16572
rect 14093 16575 14151 16581
rect 12757 16541 12769 16544
rect 12711 16535 12769 16541
rect 14093 16541 14105 16575
rect 14139 16572 14151 16575
rect 14274 16572 14280 16584
rect 14139 16544 14280 16572
rect 14139 16541 14151 16544
rect 14093 16535 14151 16541
rect 14274 16532 14280 16544
rect 14332 16532 14338 16584
rect 14660 16572 14688 16600
rect 14921 16575 14979 16581
rect 14921 16572 14933 16575
rect 14660 16544 14933 16572
rect 14921 16541 14933 16544
rect 14967 16541 14979 16575
rect 15028 16572 15056 16612
rect 15105 16609 15117 16643
rect 15151 16640 15163 16643
rect 15194 16640 15200 16652
rect 15151 16612 15200 16640
rect 15151 16609 15163 16612
rect 15105 16603 15163 16609
rect 15194 16600 15200 16612
rect 15252 16600 15258 16652
rect 15958 16643 16016 16649
rect 15958 16640 15970 16643
rect 15304 16612 15970 16640
rect 15304 16572 15332 16612
rect 15958 16609 15970 16612
rect 16004 16609 16016 16643
rect 15958 16603 16016 16609
rect 16117 16643 16175 16649
rect 16117 16609 16129 16643
rect 16163 16640 16175 16643
rect 16868 16640 16896 16748
rect 17865 16745 17877 16748
rect 17911 16745 17923 16779
rect 17865 16739 17923 16745
rect 20346 16736 20352 16788
rect 20404 16736 20410 16788
rect 16163 16612 16896 16640
rect 16163 16609 16175 16612
rect 16117 16603 16175 16609
rect 20898 16600 20904 16652
rect 20956 16640 20962 16652
rect 20993 16643 21051 16649
rect 20993 16640 21005 16643
rect 20956 16612 21005 16640
rect 20956 16600 20962 16612
rect 20993 16609 21005 16612
rect 21039 16609 21051 16643
rect 20993 16603 21051 16609
rect 21450 16600 21456 16652
rect 21508 16600 21514 16652
rect 15028 16544 15332 16572
rect 14921 16535 14979 16541
rect 15838 16532 15844 16584
rect 15896 16532 15902 16584
rect 16853 16575 16911 16581
rect 16853 16541 16865 16575
rect 16899 16541 16911 16575
rect 17586 16572 17592 16584
rect 17144 16571 17592 16572
rect 16853 16535 16911 16541
rect 17127 16565 17592 16571
rect 7101 16507 7159 16513
rect 7101 16504 7113 16507
rect 6972 16476 7113 16504
rect 6972 16464 6978 16476
rect 7101 16473 7113 16476
rect 7147 16473 7159 16507
rect 7101 16467 7159 16473
rect 5442 16436 5448 16448
rect 4448 16408 5448 16436
rect 5442 16396 5448 16408
rect 5500 16396 5506 16448
rect 5534 16396 5540 16448
rect 5592 16436 5598 16448
rect 6086 16436 6092 16448
rect 5592 16408 6092 16436
rect 5592 16396 5598 16408
rect 6086 16396 6092 16408
rect 6144 16436 6150 16448
rect 7558 16436 7564 16448
rect 6144 16408 7564 16436
rect 6144 16396 6150 16408
rect 7558 16396 7564 16408
rect 7616 16396 7622 16448
rect 9953 16439 10011 16445
rect 9953 16405 9965 16439
rect 9999 16436 10011 16439
rect 10042 16436 10048 16448
rect 9999 16408 10048 16436
rect 9999 16405 10011 16408
rect 9953 16399 10011 16405
rect 10042 16396 10048 16408
rect 10100 16396 10106 16448
rect 11054 16396 11060 16448
rect 11112 16436 11118 16448
rect 11330 16436 11336 16448
rect 11112 16408 11336 16436
rect 11112 16396 11118 16408
rect 11330 16396 11336 16408
rect 11388 16396 11394 16448
rect 12158 16396 12164 16448
rect 12216 16396 12222 16448
rect 14277 16439 14335 16445
rect 14277 16405 14289 16439
rect 14323 16436 14335 16439
rect 15286 16436 15292 16448
rect 14323 16408 15292 16436
rect 14323 16405 14335 16408
rect 14277 16399 14335 16405
rect 15286 16396 15292 16408
rect 15344 16396 15350 16448
rect 15378 16396 15384 16448
rect 15436 16436 15442 16448
rect 16868 16436 16896 16535
rect 17127 16531 17139 16565
rect 17173 16544 17592 16565
rect 17173 16531 17185 16544
rect 17586 16532 17592 16544
rect 17644 16532 17650 16584
rect 19337 16575 19395 16581
rect 19337 16541 19349 16575
rect 19383 16541 19395 16575
rect 20162 16572 20168 16584
rect 19610 16551 20168 16572
rect 19337 16535 19395 16541
rect 19595 16545 20168 16551
rect 17127 16525 17185 16531
rect 15436 16408 16896 16436
rect 15436 16396 15442 16408
rect 17034 16396 17040 16448
rect 17092 16436 17098 16448
rect 17144 16436 17172 16525
rect 17092 16408 17172 16436
rect 19352 16436 19380 16535
rect 19595 16511 19607 16545
rect 19641 16544 20168 16545
rect 19641 16511 19653 16544
rect 20162 16532 20168 16544
rect 20220 16532 20226 16584
rect 20714 16532 20720 16584
rect 20772 16532 20778 16584
rect 20809 16575 20867 16581
rect 20809 16541 20821 16575
rect 20855 16572 20867 16575
rect 21082 16572 21088 16584
rect 20855 16544 21088 16572
rect 20855 16541 20867 16544
rect 20809 16535 20867 16541
rect 21082 16532 21088 16544
rect 21140 16532 21146 16584
rect 19595 16505 19653 16511
rect 19978 16464 19984 16516
rect 20036 16504 20042 16516
rect 21177 16507 21235 16513
rect 21177 16504 21189 16507
rect 20036 16476 21189 16504
rect 20036 16464 20042 16476
rect 21177 16473 21189 16476
rect 21223 16473 21235 16507
rect 21177 16467 21235 16473
rect 19610 16436 19616 16448
rect 19352 16408 19616 16436
rect 17092 16396 17098 16408
rect 19610 16396 19616 16408
rect 19668 16396 19674 16448
rect 20990 16396 20996 16448
rect 21048 16396 21054 16448
rect 1104 16346 22056 16368
rect 1104 16294 6148 16346
rect 6200 16294 6212 16346
rect 6264 16294 6276 16346
rect 6328 16294 6340 16346
rect 6392 16294 6404 16346
rect 6456 16294 11346 16346
rect 11398 16294 11410 16346
rect 11462 16294 11474 16346
rect 11526 16294 11538 16346
rect 11590 16294 11602 16346
rect 11654 16294 16544 16346
rect 16596 16294 16608 16346
rect 16660 16294 16672 16346
rect 16724 16294 16736 16346
rect 16788 16294 16800 16346
rect 16852 16294 21742 16346
rect 21794 16294 21806 16346
rect 21858 16294 21870 16346
rect 21922 16294 21934 16346
rect 21986 16294 21998 16346
rect 22050 16294 22056 16346
rect 1104 16272 22056 16294
rect 1302 16192 1308 16244
rect 1360 16232 1366 16244
rect 1581 16235 1639 16241
rect 1581 16232 1593 16235
rect 1360 16204 1593 16232
rect 1360 16192 1366 16204
rect 1581 16201 1593 16204
rect 1627 16201 1639 16235
rect 1581 16195 1639 16201
rect 2774 16192 2780 16244
rect 2832 16232 2838 16244
rect 5258 16232 5264 16244
rect 2832 16204 5264 16232
rect 2832 16192 2838 16204
rect 5258 16192 5264 16204
rect 5316 16232 5322 16244
rect 5905 16235 5963 16241
rect 5316 16204 5856 16232
rect 5316 16192 5322 16204
rect 1486 16124 1492 16176
rect 1544 16124 1550 16176
rect 4890 16164 4896 16176
rect 4356 16136 4896 16164
rect 2314 16056 2320 16108
rect 2372 16096 2378 16108
rect 2409 16099 2467 16105
rect 2409 16096 2421 16099
rect 2372 16068 2421 16096
rect 2372 16056 2378 16068
rect 2409 16065 2421 16068
rect 2455 16065 2467 16099
rect 2409 16059 2467 16065
rect 3418 16056 3424 16108
rect 3476 16056 3482 16108
rect 4246 16056 4252 16108
rect 4304 16056 4310 16108
rect 2038 15988 2044 16040
rect 2096 16028 2102 16040
rect 2225 16031 2283 16037
rect 2225 16028 2237 16031
rect 2096 16000 2237 16028
rect 2096 15988 2102 16000
rect 2225 15997 2237 16000
rect 2271 16028 2283 16031
rect 2590 16028 2596 16040
rect 2271 16000 2596 16028
rect 2271 15997 2283 16000
rect 2225 15991 2283 15997
rect 2590 15988 2596 16000
rect 2648 15988 2654 16040
rect 2958 15988 2964 16040
rect 3016 16028 3022 16040
rect 3145 16031 3203 16037
rect 3145 16028 3157 16031
rect 3016 16000 3157 16028
rect 3016 15988 3022 16000
rect 3145 15997 3157 16000
rect 3191 15997 3203 16031
rect 3145 15991 3203 15997
rect 3283 16031 3341 16037
rect 3283 15997 3295 16031
rect 3329 16028 3341 16031
rect 4356 16028 4384 16136
rect 4890 16124 4896 16136
rect 4948 16124 4954 16176
rect 4982 16124 4988 16176
rect 5040 16164 5046 16176
rect 5828 16164 5856 16204
rect 5905 16201 5917 16235
rect 5951 16232 5963 16235
rect 7190 16232 7196 16244
rect 5951 16204 7196 16232
rect 5951 16201 5963 16204
rect 5905 16195 5963 16201
rect 7190 16192 7196 16204
rect 7248 16192 7254 16244
rect 7282 16192 7288 16244
rect 7340 16232 7346 16244
rect 9950 16232 9956 16244
rect 7340 16204 9956 16232
rect 7340 16192 7346 16204
rect 5040 16136 5166 16164
rect 5828 16136 5948 16164
rect 5040 16124 5046 16136
rect 5138 16135 5166 16136
rect 5138 16129 5209 16135
rect 5138 16095 5163 16129
rect 5197 16096 5209 16129
rect 5920 16096 5948 16136
rect 5994 16124 6000 16176
rect 6052 16164 6058 16176
rect 9214 16164 9220 16176
rect 6052 16136 9220 16164
rect 6052 16124 6058 16136
rect 9214 16124 9220 16136
rect 9272 16124 9278 16176
rect 6914 16096 6920 16108
rect 5197 16095 5764 16096
rect 5138 16068 5764 16095
rect 5920 16068 6920 16096
rect 3329 16000 4384 16028
rect 4893 16031 4951 16037
rect 3329 15997 3341 16000
rect 3283 15991 3341 15997
rect 4893 15997 4905 16031
rect 4939 15997 4951 16031
rect 5736 16028 5764 16068
rect 6914 16056 6920 16068
rect 6972 16056 6978 16108
rect 7006 16056 7012 16108
rect 7064 16096 7070 16108
rect 7282 16096 7288 16108
rect 7064 16068 7288 16096
rect 7064 16056 7070 16068
rect 7282 16056 7288 16068
rect 7340 16096 7346 16108
rect 8113 16099 8171 16105
rect 8113 16096 8125 16099
rect 7340 16068 8125 16096
rect 7340 16056 7346 16068
rect 8113 16065 8125 16068
rect 8159 16096 8171 16099
rect 8294 16096 8300 16108
rect 8159 16068 8300 16096
rect 8159 16065 8171 16068
rect 8113 16059 8171 16065
rect 8294 16056 8300 16068
rect 8352 16056 8358 16108
rect 9508 16105 9536 16204
rect 9950 16192 9956 16204
rect 10008 16192 10014 16244
rect 11238 16192 11244 16244
rect 11296 16232 11302 16244
rect 11333 16235 11391 16241
rect 11333 16232 11345 16235
rect 11296 16204 11345 16232
rect 11296 16192 11302 16204
rect 11333 16201 11345 16204
rect 11379 16201 11391 16235
rect 11333 16195 11391 16201
rect 12802 16192 12808 16244
rect 12860 16232 12866 16244
rect 12897 16235 12955 16241
rect 12897 16232 12909 16235
rect 12860 16204 12909 16232
rect 12860 16192 12866 16204
rect 12897 16201 12909 16204
rect 12943 16201 12955 16235
rect 12897 16195 12955 16201
rect 13446 16192 13452 16244
rect 13504 16232 13510 16244
rect 15657 16235 15715 16241
rect 13504 16204 14688 16232
rect 13504 16192 13510 16204
rect 9674 16164 9680 16176
rect 9600 16136 9680 16164
rect 8387 16099 8445 16105
rect 8387 16065 8399 16099
rect 8433 16096 8445 16099
rect 9493 16099 9551 16105
rect 8433 16068 8800 16096
rect 8433 16065 8445 16068
rect 8387 16059 8445 16065
rect 7745 16031 7803 16037
rect 7745 16028 7757 16031
rect 5736 16000 7757 16028
rect 4893 15991 4951 15997
rect 7745 15997 7757 16000
rect 7791 15997 7803 16031
rect 7745 15991 7803 15997
rect 8772 16028 8800 16068
rect 9493 16065 9505 16099
rect 9539 16065 9551 16099
rect 9493 16059 9551 16065
rect 9600 16028 9628 16136
rect 9674 16124 9680 16136
rect 9732 16124 9738 16176
rect 12434 16164 12440 16176
rect 11900 16136 12440 16164
rect 10594 16105 10600 16108
rect 10551 16099 10600 16105
rect 10551 16065 10563 16099
rect 10597 16065 10600 16099
rect 10551 16059 10600 16065
rect 10594 16056 10600 16059
rect 10652 16056 10658 16108
rect 11900 16105 11928 16136
rect 12434 16124 12440 16136
rect 12492 16124 12498 16176
rect 13630 16124 13636 16176
rect 13688 16124 13694 16176
rect 14660 16164 14688 16204
rect 15657 16201 15669 16235
rect 15703 16232 15715 16235
rect 15930 16232 15936 16244
rect 15703 16204 15936 16232
rect 15703 16201 15715 16204
rect 15657 16195 15715 16201
rect 15930 16192 15936 16204
rect 15988 16192 15994 16244
rect 16038 16204 17080 16232
rect 15378 16164 15384 16176
rect 14660 16136 15384 16164
rect 11885 16099 11943 16105
rect 11885 16065 11897 16099
rect 11931 16065 11943 16099
rect 11885 16059 11943 16065
rect 12066 16056 12072 16108
rect 12124 16096 12130 16108
rect 12159 16099 12217 16105
rect 12159 16096 12171 16099
rect 12124 16068 12171 16096
rect 12124 16056 12130 16068
rect 12159 16065 12171 16068
rect 12205 16096 12217 16099
rect 12205 16068 12572 16096
rect 12205 16065 12217 16068
rect 12159 16059 12217 16065
rect 8772 16000 9628 16028
rect 2498 15920 2504 15972
rect 2556 15960 2562 15972
rect 2869 15963 2927 15969
rect 2869 15960 2881 15963
rect 2556 15932 2881 15960
rect 2556 15920 2562 15932
rect 2869 15929 2881 15932
rect 2915 15929 2927 15963
rect 4908 15960 4936 15991
rect 2869 15923 2927 15929
rect 3804 15932 4384 15960
rect 4908 15932 5028 15960
rect 3804 15904 3832 15932
rect 3786 15852 3792 15904
rect 3844 15852 3850 15904
rect 3878 15852 3884 15904
rect 3936 15892 3942 15904
rect 4356 15901 4384 15932
rect 5000 15904 5028 15932
rect 4065 15895 4123 15901
rect 4065 15892 4077 15895
rect 3936 15864 4077 15892
rect 3936 15852 3942 15864
rect 4065 15861 4077 15864
rect 4111 15861 4123 15895
rect 4065 15855 4123 15861
rect 4341 15895 4399 15901
rect 4341 15861 4353 15895
rect 4387 15861 4399 15895
rect 4341 15855 4399 15861
rect 4982 15852 4988 15904
rect 5040 15892 5046 15904
rect 5350 15892 5356 15904
rect 5040 15864 5356 15892
rect 5040 15852 5046 15864
rect 5350 15852 5356 15864
rect 5408 15852 5414 15904
rect 7760 15892 7788 15991
rect 8772 15892 8800 16000
rect 9674 15988 9680 16040
rect 9732 15988 9738 16040
rect 10042 15988 10048 16040
rect 10100 16028 10106 16040
rect 10137 16031 10195 16037
rect 10137 16028 10149 16031
rect 10100 16000 10149 16028
rect 10100 15988 10106 16000
rect 10137 15997 10149 16000
rect 10183 15997 10195 16031
rect 10137 15991 10195 15997
rect 10226 15988 10232 16040
rect 10284 16028 10290 16040
rect 10410 16028 10416 16040
rect 10284 16000 10416 16028
rect 10284 15988 10290 16000
rect 10410 15988 10416 16000
rect 10468 15988 10474 16040
rect 10689 16031 10747 16037
rect 10689 15997 10701 16031
rect 10735 16028 10747 16031
rect 10870 16028 10876 16040
rect 10735 16000 10876 16028
rect 10735 15997 10747 16000
rect 10689 15991 10747 15997
rect 10870 15988 10876 16000
rect 10928 15988 10934 16040
rect 7760 15864 8800 15892
rect 9122 15852 9128 15904
rect 9180 15852 9186 15904
rect 10686 15852 10692 15904
rect 10744 15892 10750 15904
rect 12544 15892 12572 16068
rect 13078 16056 13084 16108
rect 13136 16096 13142 16108
rect 13539 16099 13597 16105
rect 13539 16096 13551 16099
rect 13136 16068 13551 16096
rect 13136 16056 13142 16068
rect 13539 16065 13551 16068
rect 13585 16096 13597 16099
rect 13648 16096 13676 16124
rect 13585 16068 13676 16096
rect 13585 16065 13597 16068
rect 13539 16059 13597 16065
rect 14660 16040 14688 16136
rect 15378 16124 15384 16136
rect 15436 16124 15442 16176
rect 16038 16164 16066 16204
rect 15470 16136 16066 16164
rect 14919 16099 14977 16105
rect 14919 16065 14931 16099
rect 14965 16096 14977 16099
rect 15470 16096 15498 16136
rect 16114 16124 16120 16176
rect 16172 16164 16178 16176
rect 17052 16164 17080 16204
rect 17310 16192 17316 16244
rect 17368 16232 17374 16244
rect 17681 16235 17739 16241
rect 17681 16232 17693 16235
rect 17368 16204 17693 16232
rect 17368 16192 17374 16204
rect 17681 16201 17693 16204
rect 17727 16201 17739 16235
rect 17681 16195 17739 16201
rect 17954 16192 17960 16244
rect 18012 16232 18018 16244
rect 18322 16232 18328 16244
rect 18012 16204 18328 16232
rect 18012 16192 18018 16204
rect 18322 16192 18328 16204
rect 18380 16192 18386 16244
rect 18785 16235 18843 16241
rect 18785 16201 18797 16235
rect 18831 16201 18843 16235
rect 18785 16195 18843 16201
rect 20625 16235 20683 16241
rect 20625 16201 20637 16235
rect 20671 16232 20683 16235
rect 20714 16232 20720 16244
rect 20671 16204 20720 16232
rect 20671 16201 20683 16204
rect 20625 16195 20683 16201
rect 18800 16164 18828 16195
rect 20714 16192 20720 16204
rect 20772 16192 20778 16244
rect 20806 16192 20812 16244
rect 20864 16192 20870 16244
rect 20990 16192 20996 16244
rect 21048 16192 21054 16244
rect 21082 16192 21088 16244
rect 21140 16192 21146 16244
rect 16172 16136 16342 16164
rect 17052 16136 17356 16164
rect 18800 16136 19288 16164
rect 16172 16124 16178 16136
rect 14965 16068 15498 16096
rect 14965 16065 14977 16068
rect 14919 16059 14977 16065
rect 15838 16056 15844 16108
rect 15896 16096 15902 16108
rect 16209 16099 16267 16105
rect 16209 16096 16221 16099
rect 15896 16068 16221 16096
rect 15896 16056 15902 16068
rect 16209 16065 16221 16068
rect 16255 16065 16267 16099
rect 16314 16096 16342 16136
rect 16850 16096 16856 16108
rect 16314 16068 16856 16096
rect 16209 16059 16267 16065
rect 16850 16056 16856 16068
rect 16908 16105 16914 16108
rect 16908 16099 16969 16105
rect 16908 16065 16923 16099
rect 16957 16065 16969 16099
rect 16908 16059 16969 16065
rect 16908 16056 16914 16059
rect 13262 15988 13268 16040
rect 13320 15988 13326 16040
rect 14642 15988 14648 16040
rect 14700 15988 14706 16040
rect 15746 15988 15752 16040
rect 15804 16028 15810 16040
rect 16669 16031 16727 16037
rect 16669 16028 16681 16031
rect 15804 16000 16681 16028
rect 15804 15988 15810 16000
rect 16224 15972 16252 16000
rect 16669 15997 16681 16000
rect 16715 15997 16727 16031
rect 16669 15991 16727 15997
rect 14200 15932 14780 15960
rect 14200 15892 14228 15932
rect 10744 15864 14228 15892
rect 10744 15852 10750 15864
rect 14274 15852 14280 15904
rect 14332 15852 14338 15904
rect 14752 15892 14780 15932
rect 16206 15920 16212 15972
rect 16264 15920 16270 15972
rect 17328 15960 17356 16136
rect 18322 16056 18328 16108
rect 18380 16056 18386 16108
rect 18690 16056 18696 16108
rect 18748 16096 18754 16108
rect 19260 16105 19288 16136
rect 18969 16099 19027 16105
rect 18969 16096 18981 16099
rect 18748 16068 18981 16096
rect 18748 16056 18754 16068
rect 18969 16065 18981 16068
rect 19015 16065 19027 16099
rect 18969 16059 19027 16065
rect 19061 16099 19119 16105
rect 19061 16065 19073 16099
rect 19107 16065 19119 16099
rect 19061 16059 19119 16065
rect 19245 16099 19303 16105
rect 19245 16065 19257 16099
rect 19291 16065 19303 16099
rect 19855 16099 19913 16105
rect 19855 16096 19867 16099
rect 19245 16059 19303 16065
rect 19352 16068 19867 16096
rect 17402 15988 17408 16040
rect 17460 16028 17466 16040
rect 17862 16028 17868 16040
rect 17460 16000 17868 16028
rect 17460 15988 17466 16000
rect 17862 15988 17868 16000
rect 17920 15988 17926 16040
rect 18874 15988 18880 16040
rect 18932 16028 18938 16040
rect 19076 16028 19104 16059
rect 18932 16000 19104 16028
rect 18932 15988 18938 16000
rect 19242 15960 19248 15972
rect 17328 15932 19248 15960
rect 19242 15920 19248 15932
rect 19300 15960 19306 15972
rect 19352 15960 19380 16068
rect 19855 16065 19867 16068
rect 19901 16065 19913 16099
rect 20824 16096 20852 16192
rect 21008 16164 21036 16192
rect 21008 16136 21312 16164
rect 21284 16105 21312 16136
rect 20993 16099 21051 16105
rect 20993 16096 21005 16099
rect 20824 16068 21005 16096
rect 19855 16059 19913 16065
rect 20993 16065 21005 16068
rect 21039 16065 21051 16099
rect 20993 16059 21051 16065
rect 21269 16099 21327 16105
rect 21269 16065 21281 16099
rect 21315 16065 21327 16099
rect 21269 16059 21327 16065
rect 19610 15988 19616 16040
rect 19668 15988 19674 16040
rect 19300 15932 19380 15960
rect 19300 15920 19306 15932
rect 16114 15892 16120 15904
rect 14752 15864 16120 15892
rect 16114 15852 16120 15864
rect 16172 15852 16178 15904
rect 16298 15852 16304 15904
rect 16356 15892 16362 15904
rect 17402 15892 17408 15904
rect 16356 15864 17408 15892
rect 16356 15852 16362 15864
rect 17402 15852 17408 15864
rect 17460 15852 17466 15904
rect 18414 15852 18420 15904
rect 18472 15852 18478 15904
rect 19058 15852 19064 15904
rect 19116 15892 19122 15904
rect 19153 15895 19211 15901
rect 19153 15892 19165 15895
rect 19116 15864 19165 15892
rect 19116 15852 19122 15864
rect 19153 15861 19165 15864
rect 19199 15861 19211 15895
rect 19153 15855 19211 15861
rect 21450 15852 21456 15904
rect 21508 15852 21514 15904
rect 1104 15802 21896 15824
rect 1104 15750 3549 15802
rect 3601 15750 3613 15802
rect 3665 15750 3677 15802
rect 3729 15750 3741 15802
rect 3793 15750 3805 15802
rect 3857 15750 8747 15802
rect 8799 15750 8811 15802
rect 8863 15750 8875 15802
rect 8927 15750 8939 15802
rect 8991 15750 9003 15802
rect 9055 15750 13945 15802
rect 13997 15750 14009 15802
rect 14061 15750 14073 15802
rect 14125 15750 14137 15802
rect 14189 15750 14201 15802
rect 14253 15750 19143 15802
rect 19195 15750 19207 15802
rect 19259 15750 19271 15802
rect 19323 15750 19335 15802
rect 19387 15750 19399 15802
rect 19451 15750 21896 15802
rect 1104 15728 21896 15750
rect 2406 15648 2412 15700
rect 2464 15648 2470 15700
rect 2869 15691 2927 15697
rect 2869 15657 2881 15691
rect 2915 15688 2927 15691
rect 4246 15688 4252 15700
rect 2915 15660 4252 15688
rect 2915 15657 2927 15660
rect 2869 15651 2927 15657
rect 4246 15648 4252 15660
rect 4304 15648 4310 15700
rect 4338 15648 4344 15700
rect 4396 15688 4402 15700
rect 5905 15691 5963 15697
rect 5905 15688 5917 15691
rect 4396 15660 5917 15688
rect 4396 15648 4402 15660
rect 5905 15657 5917 15660
rect 5951 15657 5963 15691
rect 5905 15651 5963 15657
rect 9122 15648 9128 15700
rect 9180 15648 9186 15700
rect 9214 15648 9220 15700
rect 9272 15688 9278 15700
rect 13909 15691 13967 15697
rect 13909 15688 13921 15691
rect 9272 15660 13921 15688
rect 9272 15648 9278 15660
rect 13909 15657 13921 15660
rect 13955 15657 13967 15691
rect 13909 15651 13967 15657
rect 14274 15648 14280 15700
rect 14332 15648 14338 15700
rect 17037 15691 17095 15697
rect 17037 15657 17049 15691
rect 17083 15688 17095 15691
rect 18322 15688 18328 15700
rect 17083 15660 18328 15688
rect 17083 15657 17095 15660
rect 17037 15651 17095 15657
rect 18322 15648 18328 15660
rect 18380 15648 18386 15700
rect 18414 15648 18420 15700
rect 18472 15688 18478 15700
rect 18877 15691 18935 15697
rect 18877 15688 18889 15691
rect 18472 15660 18889 15688
rect 18472 15648 18478 15660
rect 18877 15657 18889 15660
rect 18923 15657 18935 15691
rect 18877 15651 18935 15657
rect 19058 15648 19064 15700
rect 19116 15648 19122 15700
rect 19518 15648 19524 15700
rect 19576 15688 19582 15700
rect 19576 15660 20668 15688
rect 19576 15648 19582 15660
rect 3142 15580 3148 15632
rect 3200 15580 3206 15632
rect 3970 15580 3976 15632
rect 4028 15580 4034 15632
rect 4522 15580 4528 15632
rect 4580 15620 4586 15632
rect 4580 15592 4844 15620
rect 4580 15580 4586 15592
rect 1397 15487 1455 15493
rect 1397 15453 1409 15487
rect 1443 15453 1455 15487
rect 1397 15447 1455 15453
rect 1412 15416 1440 15447
rect 1670 15444 1676 15496
rect 1728 15444 1734 15496
rect 2038 15444 2044 15496
rect 2096 15444 2102 15496
rect 3053 15487 3111 15493
rect 3053 15453 3065 15487
rect 3099 15484 3111 15487
rect 3160 15484 3188 15580
rect 3988 15493 4016 15580
rect 4065 15555 4123 15561
rect 4065 15521 4077 15555
rect 4111 15552 4123 15555
rect 4154 15552 4160 15564
rect 4111 15524 4160 15552
rect 4111 15521 4123 15524
rect 4065 15515 4123 15521
rect 4154 15512 4160 15524
rect 4212 15512 4218 15564
rect 4338 15512 4344 15564
rect 4396 15552 4402 15564
rect 4709 15555 4767 15561
rect 4709 15552 4721 15555
rect 4396 15524 4721 15552
rect 4396 15512 4402 15524
rect 4709 15521 4721 15524
rect 4755 15521 4767 15555
rect 4816 15552 4844 15592
rect 4985 15555 5043 15561
rect 4985 15552 4997 15555
rect 4816 15524 4997 15552
rect 4709 15515 4767 15521
rect 4985 15521 4997 15524
rect 5031 15521 5043 15555
rect 4985 15515 5043 15521
rect 5074 15512 5080 15564
rect 5132 15561 5138 15564
rect 5132 15555 5160 15561
rect 5148 15552 5160 15555
rect 5442 15552 5448 15564
rect 5148 15524 5448 15552
rect 5148 15521 5160 15524
rect 5132 15515 5160 15521
rect 5132 15512 5138 15515
rect 5442 15512 5448 15524
rect 5500 15512 5506 15564
rect 9140 15552 9168 15648
rect 10778 15580 10784 15632
rect 10836 15620 10842 15632
rect 10836 15592 12848 15620
rect 10836 15580 10842 15592
rect 7682 15524 9168 15552
rect 12069 15555 12127 15561
rect 12069 15521 12081 15555
rect 12115 15552 12127 15555
rect 12618 15552 12624 15564
rect 12115 15524 12624 15552
rect 12115 15521 12127 15524
rect 12069 15515 12127 15521
rect 12618 15512 12624 15524
rect 12676 15512 12682 15564
rect 12710 15512 12716 15564
rect 12768 15512 12774 15564
rect 12820 15552 12848 15592
rect 12989 15555 13047 15561
rect 12989 15552 13001 15555
rect 12820 15524 13001 15552
rect 12989 15521 13001 15524
rect 13035 15521 13047 15555
rect 12989 15515 13047 15521
rect 13265 15555 13323 15561
rect 13265 15521 13277 15555
rect 13311 15552 13323 15555
rect 14292 15552 14320 15648
rect 18690 15580 18696 15632
rect 18748 15580 18754 15632
rect 13311 15524 14320 15552
rect 13311 15521 13323 15524
rect 13265 15515 13323 15521
rect 14550 15512 14556 15564
rect 14608 15512 14614 15564
rect 15378 15512 15384 15564
rect 15436 15552 15442 15564
rect 15562 15552 15568 15564
rect 15436 15524 15568 15552
rect 15436 15512 15442 15524
rect 15562 15512 15568 15524
rect 15620 15512 15626 15564
rect 18874 15512 18880 15564
rect 18932 15512 18938 15564
rect 19076 15561 19104 15648
rect 19061 15555 19119 15561
rect 19061 15521 19073 15555
rect 19107 15521 19119 15555
rect 20640 15552 20668 15660
rect 20898 15648 20904 15700
rect 20956 15648 20962 15700
rect 20640 15524 21036 15552
rect 19061 15515 19119 15521
rect 3099 15456 3188 15484
rect 3973 15487 4031 15493
rect 3099 15453 3111 15456
rect 3053 15447 3111 15453
rect 3973 15453 3985 15487
rect 4019 15453 4031 15487
rect 3973 15447 4031 15453
rect 4246 15444 4252 15496
rect 4304 15444 4310 15496
rect 5258 15444 5264 15496
rect 5316 15444 5322 15496
rect 5902 15444 5908 15496
rect 5960 15484 5966 15496
rect 6181 15487 6239 15493
rect 6181 15484 6193 15487
rect 5960 15456 6193 15484
rect 5960 15444 5966 15456
rect 6181 15453 6193 15456
rect 6227 15453 6239 15487
rect 6181 15447 6239 15453
rect 7009 15487 7067 15493
rect 7009 15453 7021 15487
rect 7055 15484 7067 15487
rect 8018 15484 8024 15496
rect 7055 15456 8024 15484
rect 7055 15453 7067 15456
rect 7009 15447 7067 15453
rect 8018 15444 8024 15456
rect 8076 15444 8082 15496
rect 8662 15444 8668 15496
rect 8720 15484 8726 15496
rect 9214 15484 9220 15496
rect 8720 15456 9220 15484
rect 8720 15444 8726 15456
rect 9214 15444 9220 15456
rect 9272 15444 9278 15496
rect 9459 15487 9517 15493
rect 9459 15484 9471 15487
rect 9324 15456 9471 15484
rect 2056 15416 2084 15444
rect 9324 15428 9352 15456
rect 9459 15453 9471 15456
rect 9505 15453 9517 15487
rect 9459 15447 9517 15453
rect 11882 15444 11888 15496
rect 11940 15484 11946 15496
rect 13170 15493 13176 15496
rect 12253 15487 12311 15493
rect 12253 15484 12265 15487
rect 11940 15456 12265 15484
rect 11940 15444 11946 15456
rect 12253 15453 12265 15456
rect 12299 15453 12311 15487
rect 12253 15447 12311 15453
rect 13127 15487 13176 15493
rect 13127 15453 13139 15487
rect 13173 15453 13176 15487
rect 13127 15447 13176 15453
rect 13142 15446 13176 15447
rect 13170 15444 13176 15446
rect 13228 15444 13234 15496
rect 14093 15487 14151 15493
rect 14093 15453 14105 15487
rect 14139 15484 14151 15487
rect 14366 15484 14372 15496
rect 14139 15456 14372 15484
rect 14139 15453 14151 15456
rect 14093 15447 14151 15453
rect 14366 15444 14372 15456
rect 14424 15444 14430 15496
rect 14795 15487 14853 15493
rect 14795 15453 14807 15487
rect 14841 15453 14853 15487
rect 14795 15447 14853 15453
rect 1412 15388 2084 15416
rect 3237 15419 3295 15425
rect 3237 15385 3249 15419
rect 3283 15416 3295 15419
rect 6641 15419 6699 15425
rect 3283 15388 4292 15416
rect 3283 15385 3295 15388
rect 3237 15379 3295 15385
rect 3050 15308 3056 15360
rect 3108 15348 3114 15360
rect 3329 15351 3387 15357
rect 3329 15348 3341 15351
rect 3108 15320 3341 15348
rect 3108 15308 3114 15320
rect 3329 15317 3341 15320
rect 3375 15317 3387 15351
rect 3329 15311 3387 15317
rect 3789 15351 3847 15357
rect 3789 15317 3801 15351
rect 3835 15348 3847 15351
rect 4062 15348 4068 15360
rect 3835 15320 4068 15348
rect 3835 15317 3847 15320
rect 3789 15311 3847 15317
rect 4062 15308 4068 15320
rect 4120 15308 4126 15360
rect 4264 15348 4292 15388
rect 6641 15385 6653 15419
rect 6687 15416 6699 15419
rect 6730 15416 6736 15428
rect 6687 15388 6736 15416
rect 6687 15385 6699 15388
rect 6641 15379 6699 15385
rect 6730 15376 6736 15388
rect 6788 15376 6794 15428
rect 6917 15419 6975 15425
rect 6917 15385 6929 15419
rect 6963 15385 6975 15419
rect 6917 15379 6975 15385
rect 5534 15348 5540 15360
rect 4264 15320 5540 15348
rect 5534 15308 5540 15320
rect 5592 15308 5598 15360
rect 5994 15308 6000 15360
rect 6052 15308 6058 15360
rect 6932 15348 6960 15379
rect 7374 15376 7380 15428
rect 7432 15376 7438 15428
rect 7466 15376 7472 15428
rect 7524 15376 7530 15428
rect 7745 15419 7803 15425
rect 7745 15385 7757 15419
rect 7791 15416 7803 15419
rect 7834 15416 7840 15428
rect 7791 15388 7840 15416
rect 7791 15385 7803 15388
rect 7745 15379 7803 15385
rect 7834 15376 7840 15388
rect 7892 15376 7898 15428
rect 9306 15376 9312 15428
rect 9364 15376 9370 15428
rect 14810 15416 14838 15447
rect 15194 15444 15200 15496
rect 15252 15484 15258 15496
rect 16206 15484 16212 15496
rect 15252 15456 16212 15484
rect 15252 15444 15258 15456
rect 16206 15444 16212 15456
rect 16264 15444 16270 15496
rect 17126 15444 17132 15496
rect 17184 15484 17190 15496
rect 17221 15487 17279 15493
rect 17221 15484 17233 15487
rect 17184 15456 17233 15484
rect 17184 15444 17190 15456
rect 17221 15453 17233 15456
rect 17267 15453 17279 15487
rect 17221 15447 17279 15453
rect 17313 15487 17371 15493
rect 17313 15453 17325 15487
rect 17359 15484 17371 15487
rect 18785 15487 18843 15493
rect 17359 15456 18552 15484
rect 17359 15453 17371 15456
rect 17313 15447 17371 15453
rect 13738 15388 14838 15416
rect 17236 15416 17264 15447
rect 17558 15419 17616 15425
rect 17558 15416 17570 15419
rect 17236 15388 17570 15416
rect 7006 15348 7012 15360
rect 6932 15320 7012 15348
rect 7006 15308 7012 15320
rect 7064 15348 7070 15360
rect 7484 15348 7512 15376
rect 7064 15320 7512 15348
rect 7064 15308 7070 15320
rect 7558 15308 7564 15360
rect 7616 15348 7622 15360
rect 7929 15351 7987 15357
rect 7929 15348 7941 15351
rect 7616 15320 7941 15348
rect 7616 15308 7622 15320
rect 7929 15317 7941 15320
rect 7975 15317 7987 15351
rect 7929 15311 7987 15317
rect 10226 15308 10232 15360
rect 10284 15308 10290 15360
rect 11698 15308 11704 15360
rect 11756 15348 11762 15360
rect 12066 15348 12072 15360
rect 11756 15320 12072 15348
rect 11756 15308 11762 15320
rect 12066 15308 12072 15320
rect 12124 15348 12130 15360
rect 13738 15348 13766 15388
rect 17558 15385 17570 15388
rect 17604 15385 17616 15419
rect 18524 15416 18552 15456
rect 18785 15453 18797 15487
rect 18831 15484 18843 15487
rect 18892 15484 18920 15512
rect 18831 15456 18920 15484
rect 18831 15453 18843 15456
rect 18785 15447 18843 15453
rect 19150 15444 19156 15496
rect 19208 15484 19214 15496
rect 19245 15487 19303 15493
rect 19245 15484 19257 15487
rect 19208 15456 19257 15484
rect 19208 15444 19214 15456
rect 19245 15453 19257 15456
rect 19291 15453 19303 15487
rect 19245 15447 19303 15453
rect 19512 15487 19570 15493
rect 19512 15453 19524 15487
rect 19558 15484 19570 15487
rect 19794 15484 19800 15496
rect 19558 15456 19800 15484
rect 19558 15453 19570 15456
rect 19512 15447 19570 15453
rect 19794 15444 19800 15456
rect 19852 15444 19858 15496
rect 20714 15444 20720 15496
rect 20772 15484 20778 15496
rect 21008 15493 21036 15524
rect 20809 15487 20867 15493
rect 20809 15484 20821 15487
rect 20772 15456 20821 15484
rect 20772 15444 20778 15456
rect 20809 15453 20821 15456
rect 20855 15453 20867 15487
rect 20809 15447 20867 15453
rect 20993 15487 21051 15493
rect 20993 15453 21005 15487
rect 21039 15453 21051 15487
rect 20993 15447 21051 15453
rect 21174 15444 21180 15496
rect 21232 15444 21238 15496
rect 18966 15416 18972 15428
rect 18524 15388 18972 15416
rect 17558 15379 17616 15385
rect 18966 15376 18972 15388
rect 19024 15416 19030 15428
rect 19168 15416 19196 15444
rect 21082 15416 21088 15428
rect 19024 15388 19196 15416
rect 20548 15388 21088 15416
rect 19024 15376 19030 15388
rect 12124 15320 13766 15348
rect 12124 15308 12130 15320
rect 13814 15308 13820 15360
rect 13872 15348 13878 15360
rect 14277 15351 14335 15357
rect 14277 15348 14289 15351
rect 13872 15320 14289 15348
rect 13872 15308 13878 15320
rect 14277 15317 14289 15320
rect 14323 15317 14335 15351
rect 14277 15311 14335 15317
rect 15562 15308 15568 15360
rect 15620 15308 15626 15360
rect 16850 15308 16856 15360
rect 16908 15348 16914 15360
rect 18414 15348 18420 15360
rect 16908 15320 18420 15348
rect 16908 15308 16914 15320
rect 18414 15308 18420 15320
rect 18472 15308 18478 15360
rect 19061 15351 19119 15357
rect 19061 15317 19073 15351
rect 19107 15348 19119 15351
rect 20548 15348 20576 15388
rect 21082 15376 21088 15388
rect 21140 15376 21146 15428
rect 21545 15419 21603 15425
rect 21545 15385 21557 15419
rect 21591 15416 21603 15419
rect 22554 15416 22560 15428
rect 21591 15388 22560 15416
rect 21591 15385 21603 15388
rect 21545 15379 21603 15385
rect 22554 15376 22560 15388
rect 22612 15376 22618 15428
rect 19107 15320 20576 15348
rect 20625 15351 20683 15357
rect 19107 15317 19119 15320
rect 19061 15311 19119 15317
rect 20625 15317 20637 15351
rect 20671 15348 20683 15351
rect 20714 15348 20720 15360
rect 20671 15320 20720 15348
rect 20671 15317 20683 15320
rect 20625 15311 20683 15317
rect 20714 15308 20720 15320
rect 20772 15308 20778 15360
rect 1104 15258 22056 15280
rect 1104 15206 6148 15258
rect 6200 15206 6212 15258
rect 6264 15206 6276 15258
rect 6328 15206 6340 15258
rect 6392 15206 6404 15258
rect 6456 15206 11346 15258
rect 11398 15206 11410 15258
rect 11462 15206 11474 15258
rect 11526 15206 11538 15258
rect 11590 15206 11602 15258
rect 11654 15206 16544 15258
rect 16596 15206 16608 15258
rect 16660 15206 16672 15258
rect 16724 15206 16736 15258
rect 16788 15206 16800 15258
rect 16852 15206 21742 15258
rect 21794 15206 21806 15258
rect 21858 15206 21870 15258
rect 21922 15206 21934 15258
rect 21986 15206 21998 15258
rect 22050 15206 22056 15258
rect 1104 15184 22056 15206
rect 22186 15172 22192 15224
rect 22244 15212 22250 15224
rect 22554 15212 22560 15224
rect 22244 15184 22560 15212
rect 22244 15172 22250 15184
rect 22554 15172 22560 15184
rect 22612 15172 22618 15224
rect 3142 15144 3148 15156
rect 1854 15116 3148 15144
rect 1854 15047 1882 15116
rect 3142 15104 3148 15116
rect 3200 15144 3206 15156
rect 4801 15147 4859 15153
rect 3200 15116 4660 15144
rect 3200 15104 3206 15116
rect 4632 15076 4660 15116
rect 4801 15113 4813 15147
rect 4847 15144 4859 15147
rect 5902 15144 5908 15156
rect 4847 15116 5908 15144
rect 4847 15113 4859 15116
rect 4801 15107 4859 15113
rect 5902 15104 5908 15116
rect 5960 15104 5966 15156
rect 7374 15144 7380 15156
rect 6564 15116 7380 15144
rect 5074 15076 5080 15088
rect 4632 15048 5080 15076
rect 1839 15041 1897 15047
rect 1839 15007 1851 15041
rect 1885 15007 1897 15041
rect 5074 15036 5080 15048
rect 5132 15036 5138 15088
rect 1839 15001 1897 15007
rect 3970 14968 3976 15020
rect 4028 15017 4034 15020
rect 4028 15011 4056 15017
rect 4044 14977 4056 15011
rect 4028 14971 4056 14977
rect 4028 14968 4034 14971
rect 4154 14968 4160 15020
rect 4212 14968 4218 15020
rect 5092 15008 5120 15036
rect 5167 15011 5225 15017
rect 5167 15008 5179 15011
rect 5092 14980 5179 15008
rect 5167 14977 5179 14980
rect 5213 14977 5225 15011
rect 5167 14971 5225 14977
rect 5718 14968 5724 15020
rect 5776 15008 5782 15020
rect 6564 15017 6592 15116
rect 7374 15104 7380 15116
rect 7432 15104 7438 15156
rect 8294 15104 8300 15156
rect 8352 15144 8358 15156
rect 9490 15144 9496 15156
rect 8352 15116 9496 15144
rect 8352 15104 8358 15116
rect 9490 15104 9496 15116
rect 9548 15144 9554 15156
rect 9548 15116 12664 15144
rect 9548 15104 9554 15116
rect 8923 15041 8981 15047
rect 6549 15011 6607 15017
rect 5776 14980 6482 15008
rect 5776 14968 5782 14980
rect 6104 14952 6132 14980
rect 1581 14943 1639 14949
rect 1581 14909 1593 14943
rect 1627 14909 1639 14943
rect 1581 14903 1639 14909
rect 1596 14804 1624 14903
rect 2958 14900 2964 14952
rect 3016 14900 3022 14952
rect 3145 14943 3203 14949
rect 3145 14909 3157 14943
rect 3191 14940 3203 14943
rect 3881 14943 3939 14949
rect 3191 14912 3740 14940
rect 3191 14909 3203 14912
rect 3145 14903 3203 14909
rect 2593 14875 2651 14881
rect 2593 14841 2605 14875
rect 2639 14872 2651 14875
rect 3585 14875 3643 14881
rect 3585 14872 3597 14875
rect 2639 14844 3597 14872
rect 2639 14841 2651 14844
rect 2593 14835 2651 14841
rect 3585 14841 3597 14844
rect 3631 14841 3643 14875
rect 3585 14835 3643 14841
rect 1854 14804 1860 14816
rect 1596 14776 1860 14804
rect 1854 14764 1860 14776
rect 1912 14764 1918 14816
rect 3712 14804 3740 14912
rect 3881 14909 3893 14943
rect 3927 14940 3939 14943
rect 4893 14943 4951 14949
rect 4893 14940 4905 14943
rect 3927 14912 4566 14940
rect 3927 14909 3939 14912
rect 3881 14903 3939 14909
rect 3970 14804 3976 14816
rect 3712 14776 3976 14804
rect 3970 14764 3976 14776
rect 4028 14804 4034 14816
rect 4246 14804 4252 14816
rect 4028 14776 4252 14804
rect 4028 14764 4034 14776
rect 4246 14764 4252 14776
rect 4304 14764 4310 14816
rect 4538 14804 4566 14912
rect 4632 14912 4905 14940
rect 4632 14884 4660 14912
rect 4893 14909 4905 14912
rect 4939 14909 4951 14943
rect 4893 14903 4951 14909
rect 6086 14900 6092 14952
rect 6144 14900 6150 14952
rect 6362 14900 6368 14952
rect 6420 14900 6426 14952
rect 6454 14940 6482 14980
rect 6549 14977 6561 15011
rect 6595 14977 6607 15011
rect 6549 14971 6607 14977
rect 8202 14968 8208 15020
rect 8260 15008 8266 15020
rect 8923 15008 8935 15041
rect 8260 15007 8935 15008
rect 8969 15007 8981 15041
rect 9214 15036 9220 15088
rect 9272 15076 9278 15088
rect 9272 15048 9674 15076
rect 9272 15036 9278 15048
rect 8260 15001 8981 15007
rect 9646 15008 9674 15048
rect 10318 15047 10324 15088
rect 10303 15041 10324 15047
rect 10045 15011 10103 15017
rect 10045 15008 10057 15011
rect 8260 14980 8966 15001
rect 9646 14980 10057 15008
rect 8260 14968 8266 14980
rect 10045 14977 10057 14980
rect 10091 14977 10103 15011
rect 10303 15007 10315 15041
rect 10376 15036 10382 15088
rect 12434 15076 12440 15088
rect 12084 15048 12440 15076
rect 10349 15010 10364 15036
rect 12084 15017 12112 15048
rect 12434 15036 12440 15048
rect 12492 15036 12498 15088
rect 12636 15076 12664 15116
rect 12710 15104 12716 15156
rect 12768 15144 12774 15156
rect 13081 15147 13139 15153
rect 13081 15144 13093 15147
rect 12768 15116 13093 15144
rect 12768 15104 12774 15116
rect 13081 15113 13093 15116
rect 13127 15113 13139 15147
rect 15746 15144 15752 15156
rect 13081 15107 13139 15113
rect 13924 15116 15752 15144
rect 13924 15076 13952 15116
rect 15746 15104 15752 15116
rect 15804 15144 15810 15156
rect 16114 15144 16120 15156
rect 15804 15116 16120 15144
rect 15804 15104 15810 15116
rect 16114 15104 16120 15116
rect 16172 15104 16178 15156
rect 16390 15104 16396 15156
rect 16448 15144 16454 15156
rect 17126 15144 17132 15156
rect 16448 15116 17132 15144
rect 16448 15104 16454 15116
rect 17126 15104 17132 15116
rect 17184 15104 17190 15156
rect 18785 15147 18843 15153
rect 18785 15113 18797 15147
rect 18831 15144 18843 15147
rect 18874 15144 18880 15156
rect 18831 15116 18880 15144
rect 18831 15113 18843 15116
rect 18785 15107 18843 15113
rect 18874 15104 18880 15116
rect 18932 15104 18938 15156
rect 19794 15104 19800 15156
rect 19852 15104 19858 15156
rect 20714 15104 20720 15156
rect 20772 15104 20778 15156
rect 12636 15048 13952 15076
rect 12069 15011 12127 15017
rect 10349 15007 10361 15010
rect 10303 15001 10361 15007
rect 10045 14971 10103 14977
rect 12069 14977 12081 15011
rect 12115 14977 12127 15011
rect 12069 14971 12127 14977
rect 12343 15011 12401 15017
rect 12343 14977 12355 15011
rect 12389 15008 12401 15011
rect 12389 14980 12848 15008
rect 12389 14977 12401 14980
rect 12343 14971 12401 14977
rect 7466 14949 7472 14952
rect 7285 14943 7343 14949
rect 7285 14940 7297 14943
rect 6454 14912 7297 14940
rect 7285 14909 7297 14912
rect 7331 14909 7343 14943
rect 7285 14903 7343 14909
rect 7423 14943 7472 14949
rect 7423 14909 7435 14943
rect 7469 14909 7472 14943
rect 7423 14903 7472 14909
rect 7466 14900 7472 14903
rect 7524 14900 7530 14952
rect 7558 14900 7564 14952
rect 7616 14900 7622 14952
rect 7926 14900 7932 14952
rect 7984 14940 7990 14952
rect 8662 14940 8668 14952
rect 7984 14912 8668 14940
rect 7984 14900 7990 14912
rect 8662 14900 8668 14912
rect 8720 14900 8726 14952
rect 12820 14884 12848 14980
rect 15562 14968 15568 15020
rect 15620 14968 15626 15020
rect 18046 15008 18052 15020
rect 18007 14980 18052 15008
rect 18046 14968 18052 14980
rect 18104 14968 18110 15020
rect 19812 15017 19840 15104
rect 19797 15011 19855 15017
rect 19797 14977 19809 15011
rect 19843 14977 19855 15011
rect 19797 14971 19855 14977
rect 20257 15011 20315 15017
rect 20257 14977 20269 15011
rect 20303 14977 20315 15011
rect 20732 15008 20760 15104
rect 20809 15011 20867 15017
rect 20809 15008 20821 15011
rect 20732 14980 20821 15008
rect 20257 14971 20315 14977
rect 20809 14977 20821 14980
rect 20855 14977 20867 15011
rect 20809 14971 20867 14977
rect 12894 14900 12900 14952
rect 12952 14940 12958 14952
rect 13725 14943 13783 14949
rect 13725 14940 13737 14943
rect 12952 14912 13737 14940
rect 12952 14900 12958 14912
rect 13725 14909 13737 14912
rect 13771 14909 13783 14943
rect 13725 14903 13783 14909
rect 13909 14943 13967 14949
rect 13909 14909 13921 14943
rect 13955 14940 13967 14943
rect 14274 14940 14280 14952
rect 13955 14912 14280 14940
rect 13955 14909 13967 14912
rect 13909 14903 13967 14909
rect 14274 14900 14280 14912
rect 14332 14900 14338 14952
rect 14826 14949 14832 14952
rect 14645 14943 14703 14949
rect 14645 14940 14657 14943
rect 14476 14912 14657 14940
rect 4614 14832 4620 14884
rect 4672 14832 4678 14884
rect 5828 14844 6868 14872
rect 4890 14804 4896 14816
rect 4538 14776 4896 14804
rect 4890 14764 4896 14776
rect 4948 14764 4954 14816
rect 5166 14764 5172 14816
rect 5224 14804 5230 14816
rect 5828 14804 5856 14844
rect 5224 14776 5856 14804
rect 5905 14807 5963 14813
rect 5224 14764 5230 14776
rect 5905 14773 5917 14807
rect 5951 14804 5963 14807
rect 6546 14804 6552 14816
rect 5951 14776 6552 14804
rect 5951 14773 5963 14776
rect 5905 14767 5963 14773
rect 6546 14764 6552 14776
rect 6604 14764 6610 14816
rect 6840 14804 6868 14844
rect 6914 14832 6920 14884
rect 6972 14872 6978 14884
rect 7009 14875 7067 14881
rect 7009 14872 7021 14875
rect 6972 14844 7021 14872
rect 6972 14832 6978 14844
rect 7009 14841 7021 14844
rect 7055 14841 7067 14875
rect 7009 14835 7067 14841
rect 9324 14844 10180 14872
rect 7466 14804 7472 14816
rect 6840 14776 7472 14804
rect 7466 14764 7472 14776
rect 7524 14764 7530 14816
rect 8202 14764 8208 14816
rect 8260 14764 8266 14816
rect 8386 14764 8392 14816
rect 8444 14804 8450 14816
rect 9324 14804 9352 14844
rect 8444 14776 9352 14804
rect 9677 14807 9735 14813
rect 8444 14764 8450 14776
rect 9677 14773 9689 14807
rect 9723 14804 9735 14807
rect 10042 14804 10048 14816
rect 9723 14776 10048 14804
rect 9723 14773 9735 14776
rect 9677 14767 9735 14773
rect 10042 14764 10048 14776
rect 10100 14764 10106 14816
rect 10152 14804 10180 14844
rect 10704 14844 11192 14872
rect 10704 14804 10732 14844
rect 10152 14776 10732 14804
rect 11054 14764 11060 14816
rect 11112 14764 11118 14816
rect 11164 14804 11192 14844
rect 12802 14832 12808 14884
rect 12860 14832 12866 14884
rect 13538 14832 13544 14884
rect 13596 14872 13602 14884
rect 13596 14844 14320 14872
rect 13596 14832 13602 14844
rect 13630 14804 13636 14816
rect 11164 14776 13636 14804
rect 13630 14764 13636 14776
rect 13688 14764 13694 14816
rect 14292 14804 14320 14844
rect 14366 14832 14372 14884
rect 14424 14832 14430 14884
rect 14476 14804 14504 14912
rect 14645 14909 14657 14912
rect 14691 14909 14703 14943
rect 14645 14903 14703 14909
rect 14783 14943 14832 14949
rect 14783 14909 14795 14943
rect 14829 14909 14832 14943
rect 14783 14903 14832 14909
rect 14826 14900 14832 14903
rect 14884 14900 14890 14952
rect 14921 14943 14979 14949
rect 14921 14909 14933 14943
rect 14967 14940 14979 14943
rect 15580 14940 15608 14968
rect 14967 14912 15608 14940
rect 14967 14909 14979 14912
rect 14921 14903 14979 14909
rect 17678 14900 17684 14952
rect 17736 14940 17742 14952
rect 17773 14943 17831 14949
rect 17773 14940 17785 14943
rect 17736 14912 17785 14940
rect 17736 14900 17742 14912
rect 17773 14909 17785 14912
rect 17819 14909 17831 14943
rect 20272 14940 20300 14971
rect 20898 14968 20904 15020
rect 20956 14968 20962 15020
rect 21085 15011 21143 15017
rect 21085 14977 21097 15011
rect 21131 14977 21143 15011
rect 21085 14971 21143 14977
rect 21269 15011 21327 15017
rect 21269 14977 21281 15011
rect 21315 15008 21327 15011
rect 22738 15008 22744 15020
rect 21315 14980 22744 15008
rect 21315 14977 21327 14980
rect 21269 14971 21327 14977
rect 21100 14940 21128 14971
rect 22738 14968 22744 14980
rect 22796 14968 22802 15020
rect 17773 14903 17831 14909
rect 19628 14912 20300 14940
rect 20640 14912 21128 14940
rect 19628 14881 19656 14912
rect 20640 14881 20668 14912
rect 19613 14875 19671 14881
rect 15304 14844 16436 14872
rect 14292 14776 14504 14804
rect 14826 14764 14832 14816
rect 14884 14804 14890 14816
rect 15304 14804 15332 14844
rect 16408 14816 16436 14844
rect 19613 14841 19625 14875
rect 19659 14841 19671 14875
rect 20625 14875 20683 14881
rect 19613 14835 19671 14841
rect 19720 14844 20484 14872
rect 14884 14776 15332 14804
rect 14884 14764 14890 14776
rect 15562 14764 15568 14816
rect 15620 14764 15626 14816
rect 16390 14764 16396 14816
rect 16448 14764 16454 14816
rect 17310 14764 17316 14816
rect 17368 14804 17374 14816
rect 19720 14804 19748 14844
rect 17368 14776 19748 14804
rect 17368 14764 17374 14776
rect 20346 14764 20352 14816
rect 20404 14764 20410 14816
rect 20456 14804 20484 14844
rect 20625 14841 20637 14875
rect 20671 14841 20683 14875
rect 22738 14872 22744 14884
rect 20625 14835 20683 14841
rect 20732 14844 22744 14872
rect 20732 14804 20760 14844
rect 22738 14832 22744 14844
rect 22796 14832 22802 14884
rect 20456 14776 20760 14804
rect 20990 14764 20996 14816
rect 21048 14764 21054 14816
rect 21450 14764 21456 14816
rect 21508 14764 21514 14816
rect 1104 14714 21896 14736
rect 1104 14662 3549 14714
rect 3601 14662 3613 14714
rect 3665 14662 3677 14714
rect 3729 14662 3741 14714
rect 3793 14662 3805 14714
rect 3857 14662 8747 14714
rect 8799 14662 8811 14714
rect 8863 14662 8875 14714
rect 8927 14662 8939 14714
rect 8991 14662 9003 14714
rect 9055 14662 13945 14714
rect 13997 14662 14009 14714
rect 14061 14662 14073 14714
rect 14125 14662 14137 14714
rect 14189 14662 14201 14714
rect 14253 14662 19143 14714
rect 19195 14662 19207 14714
rect 19259 14662 19271 14714
rect 19323 14662 19335 14714
rect 19387 14662 19399 14714
rect 19451 14662 21896 14714
rect 1104 14640 21896 14662
rect 1762 14560 1768 14612
rect 1820 14560 1826 14612
rect 3329 14603 3387 14609
rect 3329 14569 3341 14603
rect 3375 14600 3387 14603
rect 4338 14600 4344 14612
rect 3375 14572 4344 14600
rect 3375 14569 3387 14572
rect 3329 14563 3387 14569
rect 4338 14560 4344 14572
rect 4396 14560 4402 14612
rect 5258 14560 5264 14612
rect 5316 14560 5322 14612
rect 6454 14600 6460 14612
rect 5552 14572 6460 14600
rect 4246 14492 4252 14544
rect 4304 14492 4310 14544
rect 3418 14424 3424 14476
rect 3476 14464 3482 14476
rect 3602 14464 3608 14476
rect 3476 14436 3608 14464
rect 3476 14424 3482 14436
rect 3602 14424 3608 14436
rect 3660 14424 3666 14476
rect 4264 14464 4292 14492
rect 4080 14436 4292 14464
rect 1210 14356 1216 14408
rect 1268 14396 1274 14408
rect 1673 14399 1731 14405
rect 1673 14396 1685 14399
rect 1268 14368 1685 14396
rect 1268 14356 1274 14368
rect 1673 14365 1685 14368
rect 1719 14365 1731 14399
rect 1673 14359 1731 14365
rect 2317 14399 2375 14405
rect 2317 14365 2329 14399
rect 2363 14365 2375 14399
rect 2317 14359 2375 14365
rect 2591 14399 2649 14405
rect 2591 14365 2603 14399
rect 2637 14396 2649 14399
rect 4080 14396 4108 14436
rect 2637 14368 4108 14396
rect 4249 14399 4307 14405
rect 2637 14365 2649 14368
rect 2591 14359 2649 14365
rect 4249 14365 4261 14399
rect 4295 14396 4307 14399
rect 4295 14368 4384 14396
rect 4295 14365 4307 14368
rect 4249 14359 4307 14365
rect 2332 14328 2360 14359
rect 4356 14340 4384 14368
rect 4507 14369 4565 14375
rect 2682 14328 2688 14340
rect 2332 14300 2688 14328
rect 2682 14288 2688 14300
rect 2740 14328 2746 14340
rect 4338 14328 4344 14340
rect 2740 14300 4344 14328
rect 2740 14288 2746 14300
rect 4338 14288 4344 14300
rect 4396 14288 4402 14340
rect 4507 14335 4519 14369
rect 4553 14366 4565 14369
rect 4553 14335 4566 14366
rect 4614 14356 4620 14408
rect 4672 14396 4678 14408
rect 5552 14396 5580 14572
rect 4672 14368 5580 14396
rect 5629 14399 5687 14405
rect 4672 14356 4678 14368
rect 5629 14365 5641 14399
rect 5675 14365 5687 14399
rect 5902 14396 5908 14408
rect 5863 14368 5908 14396
rect 5629 14359 5687 14365
rect 4507 14329 4566 14335
rect 4538 14328 4566 14329
rect 4706 14328 4712 14340
rect 4538 14300 4712 14328
rect 4706 14288 4712 14300
rect 4764 14328 4770 14340
rect 5350 14328 5356 14340
rect 4764 14300 5356 14328
rect 4764 14288 4770 14300
rect 5350 14288 5356 14300
rect 5408 14288 5414 14340
rect 1210 14220 1216 14272
rect 1268 14260 1274 14272
rect 2406 14260 2412 14272
rect 1268 14232 2412 14260
rect 1268 14220 1274 14232
rect 2406 14220 2412 14232
rect 2464 14220 2470 14272
rect 3234 14220 3240 14272
rect 3292 14260 3298 14272
rect 5644 14260 5672 14359
rect 5902 14356 5908 14368
rect 5960 14396 5966 14408
rect 6288 14396 6316 14572
rect 6454 14560 6460 14572
rect 6512 14560 6518 14612
rect 6641 14603 6699 14609
rect 6641 14569 6653 14603
rect 6687 14600 6699 14603
rect 7466 14600 7472 14612
rect 6687 14572 7472 14600
rect 6687 14569 6699 14572
rect 6641 14563 6699 14569
rect 7466 14560 7472 14572
rect 7524 14560 7530 14612
rect 8018 14560 8024 14612
rect 8076 14560 8082 14612
rect 9766 14560 9772 14612
rect 9824 14600 9830 14612
rect 10962 14600 10968 14612
rect 9824 14572 10968 14600
rect 9824 14560 9830 14572
rect 10962 14560 10968 14572
rect 11020 14560 11026 14612
rect 11606 14560 11612 14612
rect 11664 14600 11670 14612
rect 12894 14600 12900 14612
rect 11664 14572 12900 14600
rect 11664 14560 11670 14572
rect 12894 14560 12900 14572
rect 12952 14560 12958 14612
rect 13630 14560 13636 14612
rect 13688 14560 13694 14612
rect 14366 14560 14372 14612
rect 14424 14600 14430 14612
rect 15105 14603 15163 14609
rect 15105 14600 15117 14603
rect 14424 14572 15117 14600
rect 14424 14560 14430 14572
rect 15105 14569 15117 14572
rect 15151 14569 15163 14603
rect 15105 14563 15163 14569
rect 15562 14560 15568 14612
rect 15620 14560 15626 14612
rect 19610 14600 19616 14612
rect 19536 14572 19616 14600
rect 6362 14492 6368 14544
rect 6420 14532 6426 14544
rect 7006 14532 7012 14544
rect 6420 14504 7012 14532
rect 6420 14492 6426 14504
rect 7006 14492 7012 14504
rect 7064 14492 7070 14544
rect 10226 14492 10232 14544
rect 10284 14532 10290 14544
rect 10505 14535 10563 14541
rect 10505 14532 10517 14535
rect 10284 14504 10517 14532
rect 10284 14492 10290 14504
rect 10505 14501 10517 14504
rect 10551 14501 10563 14535
rect 10505 14495 10563 14501
rect 6546 14424 6552 14476
rect 6604 14464 6610 14476
rect 6730 14464 6736 14476
rect 6604 14436 6736 14464
rect 6604 14424 6610 14436
rect 6730 14424 6736 14436
rect 6788 14424 6794 14476
rect 10045 14467 10103 14473
rect 10045 14433 10057 14467
rect 10091 14464 10103 14467
rect 10134 14464 10140 14476
rect 10091 14436 10140 14464
rect 10091 14433 10103 14436
rect 10045 14427 10103 14433
rect 10134 14424 10140 14436
rect 10192 14424 10198 14476
rect 10594 14424 10600 14476
rect 10652 14464 10658 14476
rect 10898 14467 10956 14473
rect 10898 14464 10910 14467
rect 10652 14436 10910 14464
rect 10652 14424 10658 14436
rect 10898 14433 10910 14436
rect 10944 14433 10956 14467
rect 10898 14427 10956 14433
rect 11606 14424 11612 14476
rect 11664 14424 11670 14476
rect 12434 14424 12440 14476
rect 12492 14424 12498 14476
rect 12710 14424 12716 14476
rect 12768 14424 12774 14476
rect 12851 14467 12909 14473
rect 12851 14433 12863 14467
rect 12897 14464 12909 14467
rect 13354 14464 13360 14476
rect 12897 14436 13360 14464
rect 12897 14433 12909 14436
rect 12851 14427 12909 14433
rect 13354 14424 13360 14436
rect 13412 14464 13418 14476
rect 13538 14464 13544 14476
rect 13412 14436 13544 14464
rect 13412 14424 13418 14436
rect 13538 14424 13544 14436
rect 13596 14424 13602 14476
rect 7009 14399 7067 14405
rect 7009 14396 7021 14399
rect 5960 14368 6224 14396
rect 6288 14368 7021 14396
rect 5960 14356 5966 14368
rect 6196 14328 6224 14368
rect 7009 14365 7021 14368
rect 7055 14365 7067 14399
rect 7251 14399 7309 14405
rect 7251 14396 7263 14399
rect 7009 14359 7067 14365
rect 7114 14368 7263 14396
rect 7114 14340 7142 14368
rect 7251 14365 7263 14368
rect 7297 14365 7309 14399
rect 7251 14359 7309 14365
rect 9858 14356 9864 14408
rect 9916 14356 9922 14408
rect 10778 14356 10784 14408
rect 10836 14356 10842 14408
rect 11054 14356 11060 14408
rect 11112 14356 11118 14408
rect 11624 14396 11652 14424
rect 11793 14399 11851 14405
rect 11793 14396 11805 14399
rect 11624 14368 11805 14396
rect 11793 14365 11805 14368
rect 11839 14365 11851 14399
rect 11793 14359 11851 14365
rect 11882 14356 11888 14408
rect 11940 14396 11946 14408
rect 11977 14399 12035 14405
rect 11977 14396 11989 14399
rect 11940 14368 11989 14396
rect 11940 14356 11946 14368
rect 11977 14365 11989 14368
rect 12023 14365 12035 14399
rect 11977 14359 12035 14365
rect 12986 14356 12992 14408
rect 13044 14356 13050 14408
rect 14090 14356 14096 14408
rect 14148 14356 14154 14408
rect 14335 14399 14393 14405
rect 14335 14396 14347 14399
rect 14200 14368 14347 14396
rect 7098 14328 7104 14340
rect 6196 14300 7104 14328
rect 7098 14288 7104 14300
rect 7156 14288 7162 14340
rect 14200 14328 14228 14368
rect 14335 14365 14347 14368
rect 14381 14365 14393 14399
rect 14335 14359 14393 14365
rect 15473 14399 15531 14405
rect 15473 14365 15485 14399
rect 15519 14396 15531 14399
rect 15580 14396 15608 14560
rect 15657 14535 15715 14541
rect 15657 14501 15669 14535
rect 15703 14501 15715 14535
rect 15657 14495 15715 14501
rect 15672 14408 15700 14495
rect 17678 14424 17684 14476
rect 17736 14464 17742 14476
rect 19536 14473 19564 14572
rect 19610 14560 19616 14572
rect 19668 14560 19674 14612
rect 20346 14560 20352 14612
rect 20404 14560 20410 14612
rect 20898 14560 20904 14612
rect 20956 14560 20962 14612
rect 20990 14560 20996 14612
rect 21048 14560 21054 14612
rect 19521 14467 19579 14473
rect 19521 14464 19533 14467
rect 17736 14436 19533 14464
rect 17736 14424 17742 14436
rect 19521 14433 19533 14436
rect 19567 14433 19579 14467
rect 19521 14427 19579 14433
rect 15519 14368 15608 14396
rect 15519 14365 15531 14368
rect 15473 14359 15531 14365
rect 15654 14356 15660 14408
rect 15712 14356 15718 14408
rect 15746 14356 15752 14408
rect 15804 14356 15810 14408
rect 16298 14356 16304 14408
rect 16356 14396 16362 14408
rect 19763 14399 19821 14405
rect 19763 14396 19775 14399
rect 16356 14368 19775 14396
rect 16356 14356 16362 14368
rect 19763 14365 19775 14368
rect 19809 14365 19821 14399
rect 19763 14359 19821 14365
rect 11624 14300 12020 14328
rect 7282 14260 7288 14272
rect 3292 14232 7288 14260
rect 3292 14220 3298 14232
rect 7282 14220 7288 14232
rect 7340 14260 7346 14272
rect 7926 14260 7932 14272
rect 7340 14232 7932 14260
rect 7340 14220 7346 14232
rect 7926 14220 7932 14232
rect 7984 14220 7990 14272
rect 10962 14220 10968 14272
rect 11020 14260 11026 14272
rect 11624 14260 11652 14300
rect 11020 14232 11652 14260
rect 11020 14220 11026 14232
rect 11698 14220 11704 14272
rect 11756 14220 11762 14272
rect 11992 14260 12020 14300
rect 14016 14300 14228 14328
rect 14016 14260 14044 14300
rect 14550 14288 14556 14340
rect 14608 14288 14614 14340
rect 15194 14288 15200 14340
rect 15252 14328 15258 14340
rect 20364 14328 20392 14560
rect 20533 14535 20591 14541
rect 20533 14501 20545 14535
rect 20579 14532 20591 14535
rect 20916 14532 20944 14560
rect 20579 14504 20944 14532
rect 20579 14501 20591 14504
rect 20533 14495 20591 14501
rect 20916 14405 20944 14504
rect 21008 14464 21036 14560
rect 21177 14467 21235 14473
rect 21177 14464 21189 14467
rect 21008 14436 21189 14464
rect 21177 14433 21189 14436
rect 21223 14433 21235 14467
rect 21177 14427 21235 14433
rect 20901 14399 20959 14405
rect 20901 14365 20913 14399
rect 20947 14365 20959 14399
rect 20901 14359 20959 14365
rect 20993 14399 21051 14405
rect 20993 14365 21005 14399
rect 21039 14365 21051 14399
rect 20993 14359 21051 14365
rect 21008 14328 21036 14359
rect 21082 14356 21088 14408
rect 21140 14396 21146 14408
rect 21269 14399 21327 14405
rect 21269 14396 21281 14399
rect 21140 14368 21281 14396
rect 21140 14356 21146 14368
rect 21269 14365 21281 14368
rect 21315 14365 21327 14399
rect 21269 14359 21327 14365
rect 15252 14300 18000 14328
rect 20364 14300 21036 14328
rect 15252 14288 15258 14300
rect 11992 14232 14044 14260
rect 14090 14220 14096 14272
rect 14148 14260 14154 14272
rect 14568 14260 14596 14288
rect 17972 14272 18000 14300
rect 14148 14232 14596 14260
rect 14148 14220 14154 14232
rect 15930 14220 15936 14272
rect 15988 14220 15994 14272
rect 17954 14220 17960 14272
rect 18012 14220 18018 14272
rect 21174 14220 21180 14272
rect 21232 14220 21238 14272
rect 21453 14263 21511 14269
rect 21453 14229 21465 14263
rect 21499 14260 21511 14263
rect 22186 14260 22192 14272
rect 21499 14232 22192 14260
rect 21499 14229 21511 14232
rect 21453 14223 21511 14229
rect 22186 14220 22192 14232
rect 22244 14220 22250 14272
rect 1104 14170 22056 14192
rect 1104 14118 6148 14170
rect 6200 14118 6212 14170
rect 6264 14118 6276 14170
rect 6328 14118 6340 14170
rect 6392 14118 6404 14170
rect 6456 14118 11346 14170
rect 11398 14118 11410 14170
rect 11462 14118 11474 14170
rect 11526 14118 11538 14170
rect 11590 14118 11602 14170
rect 11654 14118 16544 14170
rect 16596 14118 16608 14170
rect 16660 14118 16672 14170
rect 16724 14118 16736 14170
rect 16788 14118 16800 14170
rect 16852 14118 21742 14170
rect 21794 14118 21806 14170
rect 21858 14118 21870 14170
rect 21922 14118 21934 14170
rect 21986 14118 21998 14170
rect 22050 14118 22056 14170
rect 1104 14096 22056 14118
rect 1857 14059 1915 14065
rect 1857 14056 1869 14059
rect 1504 14028 1869 14056
rect 934 13948 940 14000
rect 992 13988 998 14000
rect 1504 13988 1532 14028
rect 1857 14025 1869 14028
rect 1903 14025 1915 14059
rect 1857 14019 1915 14025
rect 4154 14016 4160 14068
rect 4212 14056 4218 14068
rect 4249 14059 4307 14065
rect 4249 14056 4261 14059
rect 4212 14028 4261 14056
rect 4212 14016 4218 14028
rect 4249 14025 4261 14028
rect 4295 14025 4307 14059
rect 4249 14019 4307 14025
rect 4430 14016 4436 14068
rect 4488 14016 4494 14068
rect 5258 14016 5264 14068
rect 5316 14016 5322 14068
rect 5350 14016 5356 14068
rect 5408 14016 5414 14068
rect 5626 14016 5632 14068
rect 5684 14056 5690 14068
rect 5905 14059 5963 14065
rect 5905 14056 5917 14059
rect 5684 14028 5917 14056
rect 5684 14016 5690 14028
rect 5905 14025 5917 14028
rect 5951 14025 5963 14059
rect 8021 14059 8079 14065
rect 8021 14056 8033 14059
rect 5905 14019 5963 14025
rect 6378 14028 8033 14056
rect 4448 13988 4476 14016
rect 992 13960 1532 13988
rect 1596 13960 4476 13988
rect 992 13948 998 13960
rect 1596 13929 1624 13960
rect 1581 13923 1639 13929
rect 1581 13889 1593 13923
rect 1627 13889 1639 13923
rect 1581 13883 1639 13889
rect 1762 13880 1768 13932
rect 1820 13880 1826 13932
rect 3234 13920 3240 13932
rect 1964 13892 3240 13920
rect 1964 13864 1992 13892
rect 3234 13880 3240 13892
rect 3292 13880 3298 13932
rect 3418 13880 3424 13932
rect 3476 13920 3482 13932
rect 3511 13923 3569 13929
rect 3511 13920 3523 13923
rect 3476 13892 3523 13920
rect 3476 13880 3482 13892
rect 3511 13889 3523 13892
rect 3557 13889 3569 13923
rect 3511 13883 3569 13889
rect 4430 13880 4436 13932
rect 4488 13920 4494 13932
rect 5074 13920 5080 13932
rect 4488 13892 5080 13920
rect 4488 13880 4494 13892
rect 5074 13880 5080 13892
rect 5132 13920 5138 13932
rect 5167 13923 5225 13929
rect 5167 13920 5179 13923
rect 5132 13892 5179 13920
rect 5132 13880 5138 13892
rect 5167 13889 5179 13892
rect 5213 13889 5225 13923
rect 5276 13920 5304 14016
rect 5368 13988 5396 14016
rect 6270 13988 6276 14000
rect 5368 13960 6276 13988
rect 6270 13948 6276 13960
rect 6328 13948 6334 14000
rect 6378 13920 6406 14028
rect 8021 14025 8033 14028
rect 8067 14025 8079 14059
rect 8021 14019 8079 14025
rect 8864 14028 11008 14056
rect 6546 13948 6552 14000
rect 6604 13988 6610 14000
rect 6733 13991 6791 13997
rect 6733 13988 6745 13991
rect 6604 13960 6745 13988
rect 6604 13948 6610 13960
rect 6733 13957 6745 13960
rect 6779 13957 6791 13991
rect 6733 13951 6791 13957
rect 7006 13948 7012 14000
rect 7064 13948 7070 14000
rect 5276 13892 6406 13920
rect 5167 13883 5225 13889
rect 7098 13880 7104 13932
rect 7156 13880 7162 13932
rect 7374 13880 7380 13932
rect 7432 13920 7438 13932
rect 7469 13923 7527 13929
rect 7469 13920 7481 13923
rect 7432 13892 7481 13920
rect 7432 13880 7438 13892
rect 7469 13889 7481 13892
rect 7515 13889 7527 13923
rect 7469 13883 7527 13889
rect 7558 13880 7564 13932
rect 7616 13920 7622 13932
rect 7834 13920 7840 13932
rect 7892 13929 7898 13932
rect 7892 13923 7909 13929
rect 7616 13892 7840 13920
rect 7616 13880 7622 13892
rect 7834 13880 7840 13892
rect 7897 13889 7909 13923
rect 7892 13883 7909 13889
rect 7892 13880 7898 13883
rect 6552 13864 6604 13870
rect 1946 13812 1952 13864
rect 2004 13812 2010 13864
rect 2866 13812 2872 13864
rect 2924 13852 2930 13864
rect 3050 13852 3056 13864
rect 2924 13824 3056 13852
rect 2924 13812 2930 13824
rect 3050 13812 3056 13824
rect 3108 13812 3114 13864
rect 4338 13812 4344 13864
rect 4396 13852 4402 13864
rect 4893 13855 4951 13861
rect 4893 13852 4905 13855
rect 4396 13824 4905 13852
rect 4396 13812 4402 13824
rect 4893 13821 4905 13824
rect 4939 13821 4951 13855
rect 4893 13815 4951 13821
rect 8864 13861 8892 14028
rect 9950 13929 9956 13932
rect 9907 13923 9956 13929
rect 9907 13889 9919 13923
rect 9953 13889 9956 13923
rect 9907 13883 9956 13889
rect 9950 13880 9956 13883
rect 10008 13880 10014 13932
rect 10042 13880 10048 13932
rect 10100 13880 10106 13932
rect 10689 13923 10747 13929
rect 10689 13889 10701 13923
rect 10735 13920 10747 13923
rect 10781 13923 10839 13929
rect 10781 13920 10793 13923
rect 10735 13892 10793 13920
rect 10735 13889 10747 13892
rect 10689 13883 10747 13889
rect 10781 13889 10793 13892
rect 10827 13889 10839 13923
rect 10781 13883 10839 13889
rect 10870 13880 10876 13932
rect 10928 13880 10934 13932
rect 8849 13855 8907 13861
rect 8849 13821 8861 13855
rect 8895 13821 8907 13855
rect 8849 13815 8907 13821
rect 9033 13855 9091 13861
rect 9033 13821 9045 13855
rect 9079 13852 9091 13855
rect 9214 13852 9220 13864
rect 9079 13824 9220 13852
rect 9079 13821 9091 13824
rect 9033 13815 9091 13821
rect 9214 13812 9220 13824
rect 9272 13812 9278 13864
rect 9769 13855 9827 13861
rect 9769 13821 9781 13855
rect 9815 13852 9827 13855
rect 10226 13852 10232 13864
rect 9815 13824 10232 13852
rect 9815 13821 9827 13824
rect 9769 13815 9827 13821
rect 10226 13812 10232 13824
rect 10284 13852 10290 13864
rect 10888 13852 10916 13880
rect 10284 13824 10916 13852
rect 10980 13852 11008 14028
rect 11054 14016 11060 14068
rect 11112 14056 11118 14068
rect 11241 14059 11299 14065
rect 11241 14056 11253 14059
rect 11112 14028 11253 14056
rect 11112 14016 11118 14028
rect 11241 14025 11253 14028
rect 11287 14025 11299 14059
rect 11241 14019 11299 14025
rect 11698 14016 11704 14068
rect 11756 14016 11762 14068
rect 12066 14016 12072 14068
rect 12124 14056 12130 14068
rect 12897 14059 12955 14065
rect 12124 14028 12204 14056
rect 12124 14016 12130 14028
rect 11057 13923 11115 13929
rect 11057 13889 11069 13923
rect 11103 13920 11115 13923
rect 11716 13920 11744 14016
rect 11974 13948 11980 14000
rect 12032 13948 12038 14000
rect 12176 13959 12204 14028
rect 12897 14025 12909 14059
rect 12943 14056 12955 14059
rect 12986 14056 12992 14068
rect 12943 14028 12992 14056
rect 12943 14025 12955 14028
rect 12897 14019 12955 14025
rect 12986 14016 12992 14028
rect 13044 14016 13050 14068
rect 13170 14016 13176 14068
rect 13228 14056 13234 14068
rect 13538 14056 13544 14068
rect 13228 14028 13544 14056
rect 13228 14016 13234 14028
rect 13538 14016 13544 14028
rect 13596 14016 13602 14068
rect 14458 14016 14464 14068
rect 14516 14056 14522 14068
rect 14734 14056 14740 14068
rect 14516 14028 14740 14056
rect 14516 14016 14522 14028
rect 14734 14016 14740 14028
rect 14792 14056 14798 14068
rect 15105 14059 15163 14065
rect 15105 14056 15117 14059
rect 14792 14028 15117 14056
rect 14792 14016 14798 14028
rect 15105 14025 15117 14028
rect 15151 14025 15163 14059
rect 16574 14056 16580 14068
rect 15105 14019 15163 14025
rect 15488 14028 16580 14056
rect 12143 13953 12204 13959
rect 11103 13892 11744 13920
rect 11885 13923 11943 13929
rect 11103 13889 11115 13892
rect 11057 13883 11115 13889
rect 11885 13889 11897 13923
rect 11931 13920 11943 13923
rect 11992 13920 12020 13948
rect 11931 13892 12020 13920
rect 12143 13919 12155 13953
rect 12189 13922 12204 13953
rect 14274 13948 14280 14000
rect 14332 13988 14338 14000
rect 15194 13988 15200 14000
rect 14332 13960 15200 13988
rect 14332 13948 14338 13960
rect 15194 13948 15200 13960
rect 15252 13988 15258 14000
rect 15488 13997 15516 14028
rect 16574 14016 16580 14028
rect 16632 14016 16638 14068
rect 20809 14059 20867 14065
rect 20809 14025 20821 14059
rect 20855 14056 20867 14059
rect 21082 14056 21088 14068
rect 20855 14028 21088 14056
rect 20855 14025 20867 14028
rect 20809 14019 20867 14025
rect 21082 14016 21088 14028
rect 21140 14016 21146 14068
rect 21174 14016 21180 14068
rect 21232 14016 21238 14068
rect 15381 13991 15439 13997
rect 15381 13988 15393 13991
rect 15252 13960 15393 13988
rect 15252 13948 15258 13960
rect 15381 13957 15393 13960
rect 15427 13957 15439 13991
rect 15381 13951 15439 13957
rect 15473 13991 15531 13997
rect 15473 13957 15485 13991
rect 15519 13957 15531 13991
rect 15473 13951 15531 13957
rect 16114 13948 16120 14000
rect 16172 13948 16178 14000
rect 16206 13948 16212 14000
rect 16264 13948 16270 14000
rect 19061 13991 19119 13997
rect 19061 13957 19073 13991
rect 19107 13988 19119 13991
rect 19794 13988 19800 14000
rect 19107 13960 19800 13988
rect 19107 13957 19119 13960
rect 19061 13951 19119 13957
rect 19794 13948 19800 13960
rect 19852 13948 19858 14000
rect 20070 13948 20076 14000
rect 20128 13948 20134 14000
rect 12189 13919 12201 13922
rect 12143 13913 12201 13919
rect 11931 13889 11943 13892
rect 11885 13883 11943 13889
rect 12894 13880 12900 13932
rect 12952 13920 12958 13932
rect 13170 13920 13176 13932
rect 12952 13892 13176 13920
rect 12952 13880 12958 13892
rect 13170 13880 13176 13892
rect 13228 13880 13234 13932
rect 15838 13880 15844 13932
rect 15896 13880 15902 13932
rect 16132 13920 16160 13948
rect 16669 13923 16727 13929
rect 16669 13920 16681 13923
rect 16132 13892 16681 13920
rect 16669 13889 16681 13892
rect 16715 13889 16727 13923
rect 16669 13883 16727 13889
rect 16942 13880 16948 13932
rect 17000 13880 17006 13932
rect 18966 13880 18972 13932
rect 19024 13880 19030 13932
rect 19429 13923 19487 13929
rect 19429 13889 19441 13923
rect 19475 13920 19487 13923
rect 19518 13920 19524 13932
rect 19475 13892 19524 13920
rect 19475 13889 19487 13892
rect 19429 13883 19487 13889
rect 19518 13880 19524 13892
rect 19576 13880 19582 13932
rect 19696 13923 19754 13929
rect 19696 13889 19708 13923
rect 19742 13920 19754 13923
rect 20088 13920 20116 13948
rect 20714 13920 20720 13932
rect 19742 13892 20720 13920
rect 19742 13889 19754 13892
rect 19696 13883 19754 13889
rect 20714 13880 20720 13892
rect 20772 13880 20778 13932
rect 21192 13929 21220 14016
rect 21177 13923 21235 13929
rect 21177 13889 21189 13923
rect 21223 13889 21235 13923
rect 21177 13883 21235 13889
rect 11146 13852 11152 13864
rect 10980 13824 11152 13852
rect 10284 13812 10290 13824
rect 11146 13812 11152 13824
rect 11204 13812 11210 13864
rect 16146 13824 16344 13852
rect 6552 13806 6604 13812
rect 566 13744 572 13796
rect 624 13744 630 13796
rect 1394 13744 1400 13796
rect 1452 13744 1458 13796
rect 2424 13756 3372 13784
rect 584 13592 612 13744
rect 2424 13728 2452 13756
rect 2406 13676 2412 13728
rect 2464 13676 2470 13728
rect 2866 13676 2872 13728
rect 2924 13716 2930 13728
rect 3234 13716 3240 13728
rect 2924 13688 3240 13716
rect 2924 13676 2930 13688
rect 3234 13676 3240 13688
rect 3292 13676 3298 13728
rect 3344 13716 3372 13756
rect 4246 13744 4252 13796
rect 4304 13784 4310 13796
rect 4614 13784 4620 13796
rect 4304 13756 4620 13784
rect 4304 13744 4310 13756
rect 4614 13744 4620 13756
rect 4672 13744 4678 13796
rect 9490 13744 9496 13796
rect 9548 13744 9554 13796
rect 5902 13716 5908 13728
rect 3344 13688 5908 13716
rect 5902 13676 5908 13688
rect 5960 13676 5966 13728
rect 9766 13676 9772 13728
rect 9824 13716 9830 13728
rect 10965 13719 11023 13725
rect 10965 13716 10977 13719
rect 9824 13688 10977 13716
rect 9824 13676 9830 13688
rect 10965 13685 10977 13688
rect 11011 13685 11023 13719
rect 10965 13679 11023 13685
rect 11330 13676 11336 13728
rect 11388 13716 11394 13728
rect 13354 13716 13360 13728
rect 11388 13688 13360 13716
rect 11388 13676 11394 13688
rect 13354 13676 13360 13688
rect 13412 13676 13418 13728
rect 16316 13716 16344 13824
rect 16390 13744 16396 13796
rect 16448 13744 16454 13796
rect 17681 13787 17739 13793
rect 17681 13753 17693 13787
rect 17727 13753 17739 13787
rect 17681 13747 17739 13753
rect 17696 13716 17724 13747
rect 16316 13688 17724 13716
rect 18874 13676 18880 13728
rect 18932 13716 18938 13728
rect 21266 13716 21272 13728
rect 18932 13688 21272 13716
rect 18932 13676 18938 13688
rect 21266 13676 21272 13688
rect 21324 13676 21330 13728
rect 21450 13676 21456 13728
rect 21508 13676 21514 13728
rect 1104 13626 21896 13648
rect 566 13540 572 13592
rect 624 13540 630 13592
rect 1104 13574 3549 13626
rect 3601 13574 3613 13626
rect 3665 13574 3677 13626
rect 3729 13574 3741 13626
rect 3793 13574 3805 13626
rect 3857 13574 8747 13626
rect 8799 13574 8811 13626
rect 8863 13574 8875 13626
rect 8927 13574 8939 13626
rect 8991 13574 9003 13626
rect 9055 13574 13945 13626
rect 13997 13574 14009 13626
rect 14061 13574 14073 13626
rect 14125 13574 14137 13626
rect 14189 13574 14201 13626
rect 14253 13574 19143 13626
rect 19195 13574 19207 13626
rect 19259 13574 19271 13626
rect 19323 13574 19335 13626
rect 19387 13574 19399 13626
rect 19451 13574 21896 13626
rect 1104 13552 21896 13574
rect 934 13472 940 13524
rect 992 13512 998 13524
rect 1765 13515 1823 13521
rect 1765 13512 1777 13515
rect 992 13484 1777 13512
rect 992 13472 998 13484
rect 1765 13481 1777 13484
rect 1811 13481 1823 13515
rect 1765 13475 1823 13481
rect 3237 13515 3295 13521
rect 3237 13481 3249 13515
rect 3283 13512 3295 13515
rect 3418 13512 3424 13524
rect 3283 13484 3424 13512
rect 3283 13481 3295 13484
rect 3237 13475 3295 13481
rect 3418 13472 3424 13484
rect 3476 13472 3482 13524
rect 4154 13472 4160 13524
rect 4212 13512 4218 13524
rect 4212 13484 5394 13512
rect 4212 13472 4218 13484
rect 1394 13336 1400 13388
rect 1452 13376 1458 13388
rect 1946 13376 1952 13388
rect 1452 13348 1952 13376
rect 1452 13336 1458 13348
rect 1946 13336 1952 13348
rect 2004 13376 2010 13388
rect 2225 13379 2283 13385
rect 2225 13376 2237 13379
rect 2004 13348 2237 13376
rect 2004 13336 2010 13348
rect 2225 13345 2237 13348
rect 2271 13345 2283 13379
rect 2225 13339 2283 13345
rect 3878 13336 3884 13388
rect 3936 13376 3942 13388
rect 4433 13379 4491 13385
rect 4433 13376 4445 13379
rect 3936 13348 4445 13376
rect 3936 13336 3942 13348
rect 4433 13345 4445 13348
rect 4479 13345 4491 13379
rect 4433 13339 4491 13345
rect 4706 13336 4712 13388
rect 4764 13336 4770 13388
rect 4890 13385 4896 13388
rect 4847 13379 4896 13385
rect 4847 13345 4859 13379
rect 4893 13345 4896 13379
rect 4847 13339 4896 13345
rect 4890 13336 4896 13339
rect 4948 13336 4954 13388
rect 4995 13379 5053 13385
rect 4995 13345 5007 13379
rect 5041 13376 5053 13379
rect 5366 13376 5394 13484
rect 5534 13472 5540 13524
rect 5592 13512 5598 13524
rect 5813 13515 5871 13521
rect 5813 13512 5825 13515
rect 5592 13484 5825 13512
rect 5592 13472 5598 13484
rect 5813 13481 5825 13484
rect 5859 13481 5871 13515
rect 5813 13475 5871 13481
rect 7098 13472 7104 13524
rect 7156 13472 7162 13524
rect 8481 13515 8539 13521
rect 8481 13481 8493 13515
rect 8527 13512 8539 13515
rect 9490 13512 9496 13524
rect 8527 13484 9496 13512
rect 8527 13481 8539 13484
rect 8481 13475 8539 13481
rect 9490 13472 9496 13484
rect 9548 13472 9554 13524
rect 10042 13472 10048 13524
rect 10100 13512 10106 13524
rect 10410 13512 10416 13524
rect 10100 13484 10416 13512
rect 10100 13472 10106 13484
rect 10410 13472 10416 13484
rect 10468 13472 10474 13524
rect 10962 13472 10968 13524
rect 11020 13512 11026 13524
rect 11974 13512 11980 13524
rect 11020 13484 11560 13512
rect 11020 13472 11026 13484
rect 7282 13404 7288 13456
rect 7340 13444 7346 13456
rect 7340 13416 7512 13444
rect 7340 13404 7346 13416
rect 7484 13388 7512 13416
rect 6089 13379 6147 13385
rect 6089 13376 6101 13379
rect 5041 13348 5394 13376
rect 5736 13348 6101 13376
rect 5041 13345 5053 13348
rect 4995 13339 5053 13345
rect 5736 13320 5764 13348
rect 6089 13345 6101 13348
rect 6135 13345 6147 13379
rect 6089 13339 6147 13345
rect 7466 13336 7472 13388
rect 7524 13336 7530 13388
rect 8294 13336 8300 13388
rect 8352 13336 8358 13388
rect 9769 13379 9827 13385
rect 9769 13345 9781 13379
rect 9815 13376 9827 13379
rect 9858 13376 9864 13388
rect 9815 13348 9864 13376
rect 9815 13345 9827 13348
rect 9769 13339 9827 13345
rect 9858 13336 9864 13348
rect 9916 13336 9922 13388
rect 10410 13336 10416 13388
rect 10468 13336 10474 13388
rect 10686 13336 10692 13388
rect 10744 13336 10750 13388
rect 10870 13385 10876 13388
rect 10827 13379 10876 13385
rect 10827 13345 10839 13379
rect 10873 13345 10876 13379
rect 10827 13339 10876 13345
rect 10842 13336 10876 13339
rect 10928 13376 10934 13388
rect 11330 13376 11336 13388
rect 10928 13348 11336 13376
rect 10928 13336 10934 13348
rect 11330 13336 11336 13348
rect 11388 13336 11394 13388
rect 1673 13311 1731 13317
rect 1673 13277 1685 13311
rect 1719 13308 1731 13311
rect 2130 13308 2136 13320
rect 1719 13280 2136 13308
rect 1719 13277 1731 13280
rect 1673 13271 1731 13277
rect 2130 13268 2136 13280
rect 2188 13268 2194 13320
rect 2499 13311 2557 13317
rect 2499 13277 2511 13311
rect 2545 13308 2557 13311
rect 2590 13308 2596 13320
rect 2545 13280 2596 13308
rect 2545 13277 2557 13280
rect 2499 13271 2557 13277
rect 2590 13268 2596 13280
rect 2648 13268 2654 13320
rect 2958 13268 2964 13320
rect 3016 13308 3022 13320
rect 3786 13308 3792 13320
rect 3016 13280 3792 13308
rect 3016 13268 3022 13280
rect 3786 13268 3792 13280
rect 3844 13268 3850 13320
rect 3970 13268 3976 13320
rect 4028 13268 4034 13320
rect 5718 13268 5724 13320
rect 5776 13268 5782 13320
rect 5810 13268 5816 13320
rect 5868 13308 5874 13320
rect 5997 13311 6055 13317
rect 5997 13308 6009 13311
rect 5868 13280 6009 13308
rect 5868 13268 5874 13280
rect 5997 13277 6009 13280
rect 6043 13277 6055 13311
rect 5997 13271 6055 13277
rect 6270 13268 6276 13320
rect 6328 13308 6334 13320
rect 6363 13311 6421 13317
rect 6363 13308 6375 13311
rect 6328 13280 6375 13308
rect 6328 13268 6334 13280
rect 6363 13277 6375 13280
rect 6409 13277 6421 13311
rect 6363 13271 6421 13277
rect 7743 13311 7801 13317
rect 7743 13277 7755 13311
rect 7789 13308 7801 13311
rect 7834 13308 7840 13320
rect 7789 13280 7840 13308
rect 7789 13277 7801 13280
rect 7743 13271 7801 13277
rect 7834 13268 7840 13280
rect 7892 13268 7898 13320
rect 8312 13308 8340 13336
rect 9125 13311 9183 13317
rect 9125 13308 9137 13311
rect 8312 13280 9137 13308
rect 9125 13277 9137 13280
rect 9171 13277 9183 13311
rect 9125 13271 9183 13277
rect 9214 13268 9220 13320
rect 9272 13308 9278 13320
rect 9674 13308 9680 13320
rect 9272 13280 9680 13308
rect 9272 13268 9278 13280
rect 9674 13268 9680 13280
rect 9732 13308 9738 13320
rect 9950 13308 9956 13320
rect 9732 13280 9956 13308
rect 9732 13268 9738 13280
rect 9950 13268 9956 13280
rect 10008 13268 10014 13320
rect 10842 13314 10914 13336
rect 10962 13268 10968 13320
rect 11020 13268 11026 13320
rect 11532 13308 11560 13484
rect 11716 13484 11980 13512
rect 11716 13385 11744 13484
rect 11974 13472 11980 13484
rect 12032 13472 12038 13524
rect 12434 13472 12440 13524
rect 12492 13512 12498 13524
rect 12713 13515 12771 13521
rect 12713 13512 12725 13515
rect 12492 13484 12725 13512
rect 12492 13472 12498 13484
rect 12713 13481 12725 13484
rect 12759 13481 12771 13515
rect 12713 13475 12771 13481
rect 14292 13484 15700 13512
rect 11701 13379 11759 13385
rect 11701 13345 11713 13379
rect 11747 13345 11759 13379
rect 11701 13339 11759 13345
rect 14093 13379 14151 13385
rect 14093 13345 14105 13379
rect 14139 13376 14151 13379
rect 14182 13376 14188 13388
rect 14139 13348 14188 13376
rect 14139 13345 14151 13348
rect 14093 13339 14151 13345
rect 14182 13336 14188 13348
rect 14240 13336 14246 13388
rect 14292 13385 14320 13484
rect 14734 13404 14740 13456
rect 14792 13404 14798 13456
rect 14277 13379 14335 13385
rect 14277 13345 14289 13379
rect 14323 13345 14335 13379
rect 15130 13379 15188 13385
rect 15130 13376 15142 13379
rect 14277 13339 14335 13345
rect 14366 13348 15142 13376
rect 11943 13311 12001 13317
rect 11943 13308 11955 13311
rect 11532 13280 11955 13308
rect 11943 13277 11955 13280
rect 11989 13277 12001 13311
rect 13262 13308 13268 13320
rect 11943 13271 12001 13277
rect 12360 13280 13268 13308
rect 7852 13240 7880 13268
rect 8570 13240 8576 13252
rect 5460 13212 6592 13240
rect 7852 13212 8576 13240
rect 1302 13132 1308 13184
rect 1360 13172 1366 13184
rect 5460 13172 5488 13212
rect 1360 13144 5488 13172
rect 1360 13132 1366 13144
rect 5626 13132 5632 13184
rect 5684 13132 5690 13184
rect 5718 13132 5724 13184
rect 5776 13172 5782 13184
rect 6454 13172 6460 13184
rect 5776 13144 6460 13172
rect 5776 13132 5782 13144
rect 6454 13132 6460 13144
rect 6512 13132 6518 13184
rect 6564 13172 6592 13212
rect 8570 13200 8576 13212
rect 8628 13200 8634 13252
rect 11698 13200 11704 13252
rect 11756 13240 11762 13252
rect 12360 13240 12388 13280
rect 13262 13268 13268 13280
rect 13320 13308 13326 13320
rect 14366 13308 14394 13348
rect 15130 13345 15142 13348
rect 15176 13345 15188 13379
rect 15672 13376 15700 13484
rect 15746 13472 15752 13524
rect 15804 13512 15810 13524
rect 15933 13515 15991 13521
rect 15933 13512 15945 13515
rect 15804 13484 15945 13512
rect 15804 13472 15810 13484
rect 15933 13481 15945 13484
rect 15979 13481 15991 13515
rect 15933 13475 15991 13481
rect 16574 13472 16580 13524
rect 16632 13512 16638 13524
rect 17129 13515 17187 13521
rect 17129 13512 17141 13515
rect 16632 13484 17141 13512
rect 16632 13472 16638 13484
rect 17129 13481 17141 13484
rect 17175 13481 17187 13515
rect 17129 13475 17187 13481
rect 17696 13484 18920 13512
rect 15838 13376 15844 13388
rect 15672 13348 15844 13376
rect 15130 13339 15188 13345
rect 15838 13336 15844 13348
rect 15896 13336 15902 13388
rect 16114 13336 16120 13388
rect 16172 13336 16178 13388
rect 13320 13280 14394 13308
rect 13320 13268 13326 13280
rect 15010 13268 15016 13320
rect 15068 13268 15074 13320
rect 15286 13268 15292 13320
rect 15344 13268 15350 13320
rect 16375 13281 16433 13287
rect 13814 13240 13820 13252
rect 11756 13212 12388 13240
rect 12452 13212 13820 13240
rect 11756 13200 11762 13212
rect 12452 13184 12480 13212
rect 13814 13200 13820 13212
rect 13872 13200 13878 13252
rect 16375 13247 16387 13281
rect 16421 13278 16433 13281
rect 16421 13252 16436 13278
rect 17034 13268 17040 13320
rect 17092 13308 17098 13320
rect 17696 13317 17724 13484
rect 18892 13444 18920 13484
rect 18966 13472 18972 13524
rect 19024 13512 19030 13524
rect 19245 13515 19303 13521
rect 19245 13512 19257 13515
rect 19024 13484 19257 13512
rect 19024 13472 19030 13484
rect 19245 13481 19257 13484
rect 19291 13481 19303 13515
rect 19245 13475 19303 13481
rect 20806 13472 20812 13524
rect 20864 13512 20870 13524
rect 21177 13515 21235 13521
rect 21177 13512 21189 13515
rect 20864 13484 21189 13512
rect 20864 13472 20870 13484
rect 21177 13481 21189 13484
rect 21223 13481 21235 13515
rect 21177 13475 21235 13481
rect 19058 13444 19064 13456
rect 18892 13416 19064 13444
rect 19058 13404 19064 13416
rect 19116 13404 19122 13456
rect 20824 13376 20852 13472
rect 20272 13348 20852 13376
rect 17681 13311 17739 13317
rect 17681 13308 17693 13311
rect 17092 13280 17693 13308
rect 17092 13268 17098 13280
rect 17681 13277 17693 13280
rect 17727 13277 17739 13311
rect 17681 13271 17739 13277
rect 17948 13311 18006 13317
rect 17948 13277 17960 13311
rect 17994 13308 18006 13311
rect 18506 13308 18512 13320
rect 17994 13280 18512 13308
rect 17994 13277 18006 13280
rect 17948 13271 18006 13277
rect 18506 13268 18512 13280
rect 18564 13308 18570 13320
rect 19429 13311 19487 13317
rect 19429 13308 19441 13311
rect 18564 13280 19441 13308
rect 18564 13268 18570 13280
rect 19429 13277 19441 13280
rect 19475 13277 19487 13311
rect 19429 13271 19487 13277
rect 19610 13268 19616 13320
rect 19668 13268 19674 13320
rect 19887 13311 19945 13317
rect 19887 13277 19899 13311
rect 19933 13308 19945 13311
rect 19978 13308 19984 13320
rect 19933 13280 19984 13308
rect 19933 13277 19945 13280
rect 19887 13271 19945 13277
rect 19978 13268 19984 13280
rect 20036 13308 20042 13320
rect 20272 13308 20300 13348
rect 20036 13280 20300 13308
rect 20036 13268 20042 13280
rect 20714 13268 20720 13320
rect 20772 13308 20778 13320
rect 21545 13311 21603 13317
rect 21545 13308 21557 13311
rect 20772 13280 21557 13308
rect 20772 13268 20778 13280
rect 21545 13277 21557 13280
rect 21591 13277 21603 13311
rect 21545 13271 21603 13277
rect 16375 13241 16396 13247
rect 16390 13200 16396 13241
rect 16448 13200 16454 13252
rect 18598 13200 18604 13252
rect 18656 13240 18662 13252
rect 19628 13240 19656 13268
rect 18656 13212 19656 13240
rect 18656 13200 18662 13212
rect 8941 13175 8999 13181
rect 8941 13172 8953 13175
rect 6564 13144 8953 13172
rect 8941 13141 8953 13144
rect 8987 13141 8999 13175
rect 8941 13135 8999 13141
rect 9214 13132 9220 13184
rect 9272 13172 9278 13184
rect 11609 13175 11667 13181
rect 11609 13172 11621 13175
rect 9272 13144 11621 13172
rect 9272 13132 9278 13144
rect 11609 13141 11621 13144
rect 11655 13141 11667 13175
rect 11609 13135 11667 13141
rect 12434 13132 12440 13184
rect 12492 13132 12498 13184
rect 19058 13132 19064 13184
rect 19116 13132 19122 13184
rect 20622 13132 20628 13184
rect 20680 13132 20686 13184
rect 21358 13132 21364 13184
rect 21416 13132 21422 13184
rect 1104 13082 22056 13104
rect 1104 13030 6148 13082
rect 6200 13030 6212 13082
rect 6264 13030 6276 13082
rect 6328 13030 6340 13082
rect 6392 13030 6404 13082
rect 6456 13030 11346 13082
rect 11398 13030 11410 13082
rect 11462 13030 11474 13082
rect 11526 13030 11538 13082
rect 11590 13030 11602 13082
rect 11654 13030 16544 13082
rect 16596 13030 16608 13082
rect 16660 13030 16672 13082
rect 16724 13030 16736 13082
rect 16788 13030 16800 13082
rect 16852 13030 21742 13082
rect 21794 13030 21806 13082
rect 21858 13030 21870 13082
rect 21922 13030 21934 13082
rect 21986 13030 21998 13082
rect 22050 13030 22056 13082
rect 1104 13008 22056 13030
rect 13722 12968 13728 12980
rect 1688 12940 13728 12968
rect 1688 12909 1716 12940
rect 13722 12928 13728 12940
rect 13780 12928 13786 12980
rect 14461 12971 14519 12977
rect 14461 12937 14473 12971
rect 14507 12968 14519 12971
rect 14734 12968 14740 12980
rect 14507 12940 14740 12968
rect 14507 12937 14519 12940
rect 14461 12931 14519 12937
rect 14734 12928 14740 12940
rect 14792 12928 14798 12980
rect 15286 12928 15292 12980
rect 15344 12968 15350 12980
rect 15841 12971 15899 12977
rect 15841 12968 15853 12971
rect 15344 12940 15853 12968
rect 15344 12928 15350 12940
rect 15841 12937 15853 12940
rect 15887 12937 15899 12971
rect 15841 12931 15899 12937
rect 16390 12928 16396 12980
rect 16448 12928 16454 12980
rect 18598 12928 18604 12980
rect 18656 12928 18662 12980
rect 19058 12928 19064 12980
rect 19116 12928 19122 12980
rect 21358 12968 21364 12980
rect 20456 12940 21364 12968
rect 1673 12903 1731 12909
rect 1673 12869 1685 12903
rect 1719 12869 1731 12903
rect 1673 12863 1731 12869
rect 4157 12903 4215 12909
rect 4157 12869 4169 12903
rect 4203 12900 4215 12903
rect 5810 12900 5816 12912
rect 4203 12872 5816 12900
rect 4203 12869 4215 12872
rect 4157 12863 4215 12869
rect 5810 12860 5816 12872
rect 5868 12860 5874 12912
rect 6641 12903 6699 12909
rect 6641 12900 6653 12903
rect 6288 12872 6653 12900
rect 6288 12844 6316 12872
rect 6641 12869 6653 12872
rect 6687 12869 6699 12903
rect 6641 12863 6699 12869
rect 6917 12903 6975 12909
rect 6917 12869 6929 12903
rect 6963 12900 6975 12903
rect 7098 12900 7104 12912
rect 6963 12872 7104 12900
rect 6963 12869 6975 12872
rect 6917 12863 6975 12869
rect 7098 12860 7104 12872
rect 7156 12860 7162 12912
rect 7374 12860 7380 12912
rect 7432 12860 7438 12912
rect 7558 12860 7564 12912
rect 7616 12900 7622 12912
rect 7745 12903 7803 12909
rect 7745 12900 7757 12903
rect 7616 12872 7757 12900
rect 7616 12860 7622 12872
rect 7745 12869 7757 12872
rect 7791 12869 7803 12903
rect 9306 12900 9312 12912
rect 7745 12863 7803 12869
rect 8954 12872 9312 12900
rect 2222 12792 2228 12844
rect 2280 12832 2286 12844
rect 2498 12832 2504 12844
rect 2280 12804 2504 12832
rect 2280 12792 2286 12804
rect 2498 12792 2504 12804
rect 2556 12792 2562 12844
rect 3234 12792 3240 12844
rect 3292 12792 3298 12844
rect 3510 12792 3516 12844
rect 3568 12792 3574 12844
rect 4614 12792 4620 12844
rect 4672 12832 4678 12844
rect 4951 12835 5009 12841
rect 4951 12832 4963 12835
rect 4672 12804 4963 12832
rect 4672 12792 4678 12804
rect 4951 12801 4963 12804
rect 4997 12801 5009 12835
rect 4951 12795 5009 12801
rect 5350 12792 5356 12844
rect 5408 12792 5414 12844
rect 5718 12792 5724 12844
rect 5776 12832 5782 12844
rect 6270 12832 6276 12844
rect 5776 12804 6276 12832
rect 5776 12792 5782 12804
rect 6270 12792 6276 12804
rect 6328 12792 6334 12844
rect 7006 12792 7012 12844
rect 7064 12792 7070 12844
rect 7282 12792 7288 12844
rect 7340 12832 7346 12844
rect 8846 12832 8852 12844
rect 7340 12804 8852 12832
rect 7340 12792 7346 12804
rect 8846 12792 8852 12804
rect 8904 12792 8910 12844
rect 8954 12841 8982 12872
rect 9306 12860 9312 12872
rect 9364 12860 9370 12912
rect 10410 12900 10416 12912
rect 9692 12872 10416 12900
rect 8939 12835 8997 12841
rect 8939 12801 8951 12835
rect 8985 12801 8997 12835
rect 8939 12795 8997 12801
rect 1394 12724 1400 12776
rect 1452 12724 1458 12776
rect 2314 12724 2320 12776
rect 2372 12724 2378 12776
rect 3375 12767 3433 12773
rect 3375 12733 3387 12767
rect 3421 12764 3433 12767
rect 3694 12764 3700 12776
rect 3421 12736 3700 12764
rect 3421 12733 3433 12736
rect 3375 12727 3433 12733
rect 3694 12724 3700 12736
rect 3752 12724 3758 12776
rect 4709 12767 4767 12773
rect 4709 12733 4721 12767
rect 4755 12733 4767 12767
rect 4709 12727 4767 12733
rect 1412 12696 1440 12724
rect 1412 12668 2912 12696
rect 1486 12588 1492 12640
rect 1544 12628 1550 12640
rect 1765 12631 1823 12637
rect 1765 12628 1777 12631
rect 1544 12600 1777 12628
rect 1544 12588 1550 12600
rect 1765 12597 1777 12600
rect 1811 12597 1823 12631
rect 2884 12628 2912 12668
rect 2958 12656 2964 12708
rect 3016 12656 3022 12708
rect 4724 12628 4752 12727
rect 2884 12600 4752 12628
rect 1765 12591 1823 12597
rect 4798 12588 4804 12640
rect 4856 12628 4862 12640
rect 5368 12628 5396 12792
rect 6546 12724 6552 12776
rect 6604 12724 6610 12776
rect 7742 12724 7748 12776
rect 7800 12764 7806 12776
rect 8665 12767 8723 12773
rect 7800 12736 7972 12764
rect 7800 12724 7806 12736
rect 5718 12656 5724 12708
rect 5776 12656 5782 12708
rect 7944 12705 7972 12736
rect 8665 12733 8677 12767
rect 8711 12733 8723 12767
rect 8665 12727 8723 12733
rect 7929 12699 7987 12705
rect 7929 12665 7941 12699
rect 7975 12665 7987 12699
rect 8680 12696 8708 12727
rect 9692 12705 9720 12872
rect 10410 12860 10416 12872
rect 10468 12860 10474 12912
rect 11146 12860 11152 12912
rect 11204 12900 11210 12912
rect 12526 12900 12532 12912
rect 11204 12872 12532 12900
rect 11204 12860 11210 12872
rect 10318 12832 10324 12844
rect 10279 12804 10324 12832
rect 10318 12792 10324 12804
rect 10376 12832 10382 12844
rect 12084 12841 12112 12872
rect 12526 12860 12532 12872
rect 12584 12860 12590 12912
rect 16408 12900 16436 12928
rect 18616 12900 18644 12928
rect 13004 12872 16436 12900
rect 18340 12872 18644 12900
rect 19076 12900 19104 12928
rect 19076 12872 20300 12900
rect 12069 12835 12127 12841
rect 10376 12804 10916 12832
rect 10376 12792 10382 12804
rect 10045 12767 10103 12773
rect 10045 12733 10057 12767
rect 10091 12733 10103 12767
rect 10045 12727 10103 12733
rect 9677 12699 9735 12705
rect 8680 12668 8800 12696
rect 7929 12659 7987 12665
rect 4856 12600 5396 12628
rect 4856 12588 4862 12600
rect 5626 12588 5632 12640
rect 5684 12628 5690 12640
rect 6362 12628 6368 12640
rect 5684 12600 6368 12628
rect 5684 12588 5690 12600
rect 6362 12588 6368 12600
rect 6420 12588 6426 12640
rect 8772 12628 8800 12668
rect 9677 12665 9689 12699
rect 9723 12665 9735 12699
rect 9677 12659 9735 12665
rect 10060 12640 10088 12727
rect 10042 12628 10048 12640
rect 8772 12600 10048 12628
rect 10042 12588 10048 12600
rect 10100 12628 10106 12640
rect 10318 12628 10324 12640
rect 10100 12600 10324 12628
rect 10100 12588 10106 12600
rect 10318 12588 10324 12600
rect 10376 12588 10382 12640
rect 10888 12628 10916 12804
rect 12069 12801 12081 12835
rect 12115 12801 12127 12835
rect 12069 12795 12127 12801
rect 12343 12835 12401 12841
rect 12343 12801 12355 12835
rect 12389 12832 12401 12835
rect 12802 12832 12808 12844
rect 12389 12804 12808 12832
rect 12389 12801 12401 12804
rect 12343 12795 12401 12801
rect 12802 12792 12808 12804
rect 12860 12832 12866 12844
rect 12860 12804 12940 12832
rect 12860 12792 12866 12804
rect 10962 12724 10968 12776
rect 11020 12724 11026 12776
rect 11146 12724 11152 12776
rect 11204 12764 11210 12776
rect 11698 12764 11704 12776
rect 11204 12736 11704 12764
rect 11204 12724 11210 12736
rect 11698 12724 11704 12736
rect 11756 12724 11762 12776
rect 10980 12696 11008 12724
rect 12912 12708 12940 12804
rect 11057 12699 11115 12705
rect 11057 12696 11069 12699
rect 10980 12668 11069 12696
rect 11057 12665 11069 12668
rect 11103 12665 11115 12699
rect 11057 12659 11115 12665
rect 12894 12656 12900 12708
rect 12952 12656 12958 12708
rect 13004 12628 13032 12872
rect 13723 12835 13781 12841
rect 13723 12801 13735 12835
rect 13769 12832 13781 12835
rect 13814 12832 13820 12844
rect 13769 12804 13820 12832
rect 13769 12801 13781 12804
rect 13723 12795 13781 12801
rect 13814 12792 13820 12804
rect 13872 12792 13878 12844
rect 14550 12792 14556 12844
rect 14608 12832 14614 12844
rect 14829 12835 14887 12841
rect 14829 12832 14841 12835
rect 14608 12804 14841 12832
rect 14608 12792 14614 12804
rect 14829 12801 14841 12804
rect 14875 12801 14887 12835
rect 14829 12795 14887 12801
rect 15010 12792 15016 12844
rect 15068 12832 15074 12844
rect 15103 12835 15161 12841
rect 15103 12832 15115 12835
rect 15068 12804 15115 12832
rect 15068 12792 15074 12804
rect 15103 12801 15115 12804
rect 15149 12801 15161 12835
rect 15103 12795 15161 12801
rect 16850 12792 16856 12844
rect 16908 12832 16914 12844
rect 17770 12832 17776 12844
rect 16908 12804 17776 12832
rect 16908 12792 16914 12804
rect 17770 12792 17776 12804
rect 17828 12792 17834 12844
rect 18340 12841 18368 12872
rect 18325 12835 18383 12841
rect 18325 12801 18337 12835
rect 18371 12801 18383 12835
rect 18325 12795 18383 12801
rect 18506 12792 18512 12844
rect 18564 12832 18570 12844
rect 18599 12835 18657 12841
rect 18599 12832 18611 12835
rect 18564 12804 18611 12832
rect 18564 12792 18570 12804
rect 18599 12801 18611 12804
rect 18645 12801 18657 12835
rect 19518 12832 19524 12844
rect 18599 12795 18657 12801
rect 19352 12804 19524 12832
rect 13449 12767 13507 12773
rect 13449 12733 13461 12767
rect 13495 12733 13507 12767
rect 14568 12764 14596 12792
rect 13449 12727 13507 12733
rect 14108 12736 14596 12764
rect 13464 12640 13492 12727
rect 10888 12600 13032 12628
rect 13078 12588 13084 12640
rect 13136 12588 13142 12640
rect 13446 12588 13452 12640
rect 13504 12628 13510 12640
rect 14108 12628 14136 12736
rect 17954 12724 17960 12776
rect 18012 12724 18018 12776
rect 19352 12705 19380 12804
rect 19518 12792 19524 12804
rect 19576 12832 19582 12844
rect 19705 12835 19763 12841
rect 19705 12832 19717 12835
rect 19576 12804 19717 12832
rect 19576 12792 19582 12804
rect 19705 12801 19717 12804
rect 19751 12801 19763 12835
rect 19705 12795 19763 12801
rect 19794 12792 19800 12844
rect 19852 12792 19858 12844
rect 20272 12841 20300 12872
rect 20456 12841 20484 12940
rect 21358 12928 21364 12940
rect 21416 12928 21422 12980
rect 20622 12860 20628 12912
rect 20680 12860 20686 12912
rect 20809 12903 20867 12909
rect 20809 12869 20821 12903
rect 20855 12900 20867 12903
rect 21545 12903 21603 12909
rect 21545 12900 21557 12903
rect 20855 12872 21557 12900
rect 20855 12869 20867 12872
rect 20809 12863 20867 12869
rect 21545 12869 21557 12872
rect 21591 12869 21603 12903
rect 21545 12863 21603 12869
rect 20257 12835 20315 12841
rect 20257 12801 20269 12835
rect 20303 12801 20315 12835
rect 20257 12795 20315 12801
rect 20441 12835 20499 12841
rect 20441 12801 20453 12835
rect 20487 12801 20499 12835
rect 20640 12832 20668 12860
rect 21269 12835 21327 12841
rect 21269 12832 21281 12835
rect 20640 12804 21281 12832
rect 20441 12795 20499 12801
rect 21269 12801 21281 12804
rect 21315 12801 21327 12835
rect 21269 12795 21327 12801
rect 19886 12764 19892 12776
rect 19444 12736 19892 12764
rect 19337 12699 19395 12705
rect 19337 12665 19349 12699
rect 19383 12665 19395 12699
rect 19337 12659 19395 12665
rect 13504 12600 14136 12628
rect 13504 12588 13510 12600
rect 19058 12588 19064 12640
rect 19116 12628 19122 12640
rect 19444 12628 19472 12736
rect 19886 12724 19892 12736
rect 19944 12724 19950 12776
rect 19978 12724 19984 12776
rect 20036 12724 20042 12776
rect 20898 12724 20904 12776
rect 20956 12764 20962 12776
rect 21545 12767 21603 12773
rect 21545 12764 21557 12767
rect 20956 12736 21557 12764
rect 20956 12724 20962 12736
rect 21545 12733 21557 12736
rect 21591 12733 21603 12767
rect 21545 12727 21603 12733
rect 20533 12699 20591 12705
rect 19904 12668 20484 12696
rect 19116 12600 19472 12628
rect 19116 12588 19122 12600
rect 19610 12588 19616 12640
rect 19668 12628 19674 12640
rect 19794 12628 19800 12640
rect 19668 12600 19800 12628
rect 19668 12588 19674 12600
rect 19794 12588 19800 12600
rect 19852 12588 19858 12640
rect 19904 12637 19932 12668
rect 19889 12631 19947 12637
rect 19889 12597 19901 12631
rect 19935 12597 19947 12631
rect 19889 12591 19947 12597
rect 20070 12588 20076 12640
rect 20128 12588 20134 12640
rect 20456 12628 20484 12668
rect 20533 12665 20545 12699
rect 20579 12696 20591 12699
rect 21361 12699 21419 12705
rect 21361 12696 21373 12699
rect 20579 12668 21373 12696
rect 20579 12665 20591 12668
rect 20533 12659 20591 12665
rect 21361 12665 21373 12668
rect 21407 12665 21419 12699
rect 21361 12659 21419 12665
rect 20714 12628 20720 12640
rect 20456 12600 20720 12628
rect 20714 12588 20720 12600
rect 20772 12588 20778 12640
rect 21082 12588 21088 12640
rect 21140 12588 21146 12640
rect 1104 12538 21896 12560
rect 1104 12486 3549 12538
rect 3601 12486 3613 12538
rect 3665 12486 3677 12538
rect 3729 12486 3741 12538
rect 3793 12486 3805 12538
rect 3857 12486 8747 12538
rect 8799 12486 8811 12538
rect 8863 12486 8875 12538
rect 8927 12486 8939 12538
rect 8991 12486 9003 12538
rect 9055 12486 13945 12538
rect 13997 12486 14009 12538
rect 14061 12486 14073 12538
rect 14125 12486 14137 12538
rect 14189 12486 14201 12538
rect 14253 12486 19143 12538
rect 19195 12486 19207 12538
rect 19259 12486 19271 12538
rect 19323 12486 19335 12538
rect 19387 12486 19399 12538
rect 19451 12486 21896 12538
rect 1104 12464 21896 12486
rect 22186 12452 22192 12504
rect 22244 12452 22250 12504
rect 1578 12384 1584 12436
rect 1636 12384 1642 12436
rect 3329 12427 3387 12433
rect 2148 12396 3280 12424
rect 2148 12368 2176 12396
rect 2130 12316 2136 12368
rect 2188 12316 2194 12368
rect 2222 12316 2228 12368
rect 2280 12356 2286 12368
rect 3252 12356 3280 12396
rect 3329 12393 3341 12427
rect 3375 12424 3387 12427
rect 3878 12424 3884 12436
rect 3375 12396 3884 12424
rect 3375 12393 3387 12396
rect 3329 12387 3387 12393
rect 3878 12384 3884 12396
rect 3936 12384 3942 12436
rect 3970 12384 3976 12436
rect 4028 12424 4034 12436
rect 4341 12427 4399 12433
rect 4341 12424 4353 12427
rect 4028 12396 4353 12424
rect 4028 12384 4034 12396
rect 4341 12393 4353 12396
rect 4387 12393 4399 12427
rect 4341 12387 4399 12393
rect 4706 12384 4712 12436
rect 4764 12424 4770 12436
rect 5166 12424 5172 12436
rect 4764 12396 5172 12424
rect 4764 12384 4770 12396
rect 5166 12384 5172 12396
rect 5224 12384 5230 12436
rect 5721 12427 5779 12433
rect 5721 12393 5733 12427
rect 5767 12424 5779 12427
rect 6454 12424 6460 12436
rect 5767 12396 6460 12424
rect 5767 12393 5779 12396
rect 5721 12387 5779 12393
rect 6454 12384 6460 12396
rect 6512 12384 6518 12436
rect 7006 12384 7012 12436
rect 7064 12424 7070 12436
rect 7101 12427 7159 12433
rect 7101 12424 7113 12427
rect 7064 12396 7113 12424
rect 7064 12384 7070 12396
rect 7101 12393 7113 12396
rect 7147 12393 7159 12427
rect 7101 12387 7159 12393
rect 7466 12384 7472 12436
rect 7524 12384 7530 12436
rect 7742 12384 7748 12436
rect 7800 12424 7806 12436
rect 10226 12424 10232 12436
rect 7800 12396 10232 12424
rect 7800 12384 7806 12396
rect 10226 12384 10232 12396
rect 10284 12384 10290 12436
rect 10336 12396 11468 12424
rect 4062 12356 4068 12368
rect 2280 12328 2360 12356
rect 3252 12328 4068 12356
rect 2280 12316 2286 12328
rect 2332 12297 2360 12328
rect 4062 12316 4068 12328
rect 4120 12316 4126 12368
rect 4246 12316 4252 12368
rect 4304 12356 4310 12368
rect 4304 12328 4752 12356
rect 4304 12316 4310 12328
rect 4724 12300 4752 12328
rect 6822 12316 6828 12368
rect 6880 12356 6886 12368
rect 7484 12356 7512 12384
rect 6880 12328 7512 12356
rect 8481 12359 8539 12365
rect 6880 12316 6886 12328
rect 8481 12325 8493 12359
rect 8527 12356 8539 12359
rect 10336 12356 10364 12396
rect 8527 12328 10364 12356
rect 8527 12325 8539 12328
rect 8481 12319 8539 12325
rect 2317 12291 2375 12297
rect 2317 12257 2329 12291
rect 2363 12257 2375 12291
rect 4614 12288 4620 12300
rect 2317 12251 2375 12257
rect 3896 12260 4620 12288
rect 2225 12223 2283 12229
rect 2225 12189 2237 12223
rect 2271 12189 2283 12223
rect 2225 12183 2283 12189
rect 2591 12223 2649 12229
rect 2591 12189 2603 12223
rect 2637 12220 2649 12223
rect 3896 12220 3924 12260
rect 4614 12248 4620 12260
rect 4672 12248 4678 12300
rect 4706 12248 4712 12300
rect 4764 12248 4770 12300
rect 7282 12248 7288 12300
rect 7340 12288 7346 12300
rect 7469 12291 7527 12297
rect 7469 12288 7481 12291
rect 7340 12260 7481 12288
rect 7340 12248 7346 12260
rect 7469 12257 7481 12260
rect 7515 12257 7527 12291
rect 7469 12251 7527 12257
rect 10045 12291 10103 12297
rect 10045 12257 10057 12291
rect 10091 12288 10103 12291
rect 10134 12288 10140 12300
rect 10091 12260 10140 12288
rect 10091 12257 10103 12260
rect 10045 12251 10103 12257
rect 10134 12248 10140 12260
rect 10192 12248 10198 12300
rect 10502 12248 10508 12300
rect 10560 12248 10566 12300
rect 10594 12248 10600 12300
rect 10652 12288 10658 12300
rect 10781 12291 10839 12297
rect 10781 12288 10793 12291
rect 10652 12260 10793 12288
rect 10652 12248 10658 12260
rect 10781 12257 10793 12260
rect 10827 12257 10839 12291
rect 10781 12251 10839 12257
rect 11057 12291 11115 12297
rect 11057 12257 11069 12291
rect 11103 12288 11115 12291
rect 11440 12288 11468 12396
rect 12526 12384 12532 12436
rect 12584 12424 12590 12436
rect 12894 12424 12900 12436
rect 12584 12396 12900 12424
rect 12584 12384 12590 12396
rect 12636 12297 12664 12396
rect 12894 12384 12900 12396
rect 12952 12424 12958 12436
rect 13446 12424 13452 12436
rect 12952 12396 13452 12424
rect 12952 12384 12958 12396
rect 13446 12384 13452 12396
rect 13504 12384 13510 12436
rect 13722 12384 13728 12436
rect 13780 12424 13786 12436
rect 14918 12424 14924 12436
rect 13780 12396 14924 12424
rect 13780 12384 13786 12396
rect 14918 12384 14924 12396
rect 14976 12384 14982 12436
rect 16114 12424 16120 12436
rect 15028 12396 16120 12424
rect 13630 12316 13636 12368
rect 13688 12316 13694 12368
rect 11103 12260 11468 12288
rect 12621 12291 12679 12297
rect 11103 12257 11115 12260
rect 11057 12251 11115 12257
rect 12621 12257 12633 12291
rect 12667 12257 12679 12291
rect 14734 12288 14740 12300
rect 12621 12251 12679 12257
rect 13740 12260 14740 12288
rect 2637 12192 3924 12220
rect 3973 12223 4031 12229
rect 2637 12189 2649 12192
rect 2591 12183 2649 12189
rect 3973 12189 3985 12223
rect 4019 12220 4031 12223
rect 4983 12223 5041 12229
rect 4019 12192 4936 12220
rect 4019 12189 4031 12192
rect 3973 12183 4031 12189
rect 1486 12112 1492 12164
rect 1544 12112 1550 12164
rect 2240 12152 2268 12183
rect 3878 12152 3884 12164
rect 2240 12124 3884 12152
rect 3878 12112 3884 12124
rect 3936 12112 3942 12164
rect 4249 12155 4307 12161
rect 4249 12121 4261 12155
rect 4295 12121 4307 12155
rect 4908 12152 4936 12192
rect 4983 12189 4995 12223
rect 5029 12220 5041 12223
rect 5074 12220 5080 12232
rect 5029 12192 5080 12220
rect 5029 12189 5041 12192
rect 4983 12183 5041 12189
rect 5074 12180 5080 12192
rect 5132 12180 5138 12232
rect 5626 12180 5632 12232
rect 5684 12220 5690 12232
rect 6089 12223 6147 12229
rect 6089 12220 6101 12223
rect 5684 12192 6101 12220
rect 5684 12180 5690 12192
rect 6089 12189 6101 12192
rect 6135 12189 6147 12223
rect 6089 12183 6147 12189
rect 6363 12223 6421 12229
rect 6363 12189 6375 12223
rect 6409 12220 6421 12223
rect 7190 12220 7196 12232
rect 6409 12192 7196 12220
rect 6409 12189 6421 12192
rect 6363 12183 6421 12189
rect 7190 12180 7196 12192
rect 7248 12180 7254 12232
rect 7650 12180 7656 12232
rect 7708 12220 7714 12232
rect 7743 12223 7801 12229
rect 7743 12220 7755 12223
rect 7708 12192 7755 12220
rect 7708 12180 7714 12192
rect 7743 12189 7755 12192
rect 7789 12220 7801 12223
rect 9306 12220 9312 12232
rect 7789 12192 9312 12220
rect 7789 12189 7801 12192
rect 7743 12183 7801 12189
rect 9306 12180 9312 12192
rect 9364 12180 9370 12232
rect 9674 12180 9680 12232
rect 9732 12220 9738 12232
rect 9858 12220 9864 12232
rect 9732 12192 9864 12220
rect 9732 12180 9738 12192
rect 9858 12180 9864 12192
rect 9916 12180 9922 12232
rect 10962 12229 10968 12232
rect 10919 12223 10968 12229
rect 10919 12189 10931 12223
rect 10965 12189 10968 12223
rect 10919 12183 10968 12189
rect 10962 12180 10968 12183
rect 11020 12180 11026 12232
rect 12895 12223 12953 12229
rect 12895 12189 12907 12223
rect 12941 12220 12953 12223
rect 12986 12220 12992 12232
rect 12941 12192 12992 12220
rect 12941 12189 12953 12192
rect 12895 12183 12953 12189
rect 12986 12180 12992 12192
rect 13044 12220 13050 12232
rect 13740 12220 13768 12260
rect 14734 12248 14740 12260
rect 14792 12248 14798 12300
rect 15028 12297 15056 12396
rect 16114 12384 16120 12396
rect 16172 12384 16178 12436
rect 16942 12384 16948 12436
rect 17000 12424 17006 12436
rect 17586 12424 17592 12436
rect 17000 12396 17592 12424
rect 17000 12384 17006 12396
rect 17586 12384 17592 12396
rect 17644 12384 17650 12436
rect 18782 12384 18788 12436
rect 18840 12384 18846 12436
rect 19521 12427 19579 12433
rect 19521 12393 19533 12427
rect 19567 12424 19579 12427
rect 19978 12424 19984 12436
rect 19567 12396 19984 12424
rect 19567 12393 19579 12396
rect 19521 12387 19579 12393
rect 19978 12384 19984 12396
rect 20036 12384 20042 12436
rect 20070 12384 20076 12436
rect 20128 12384 20134 12436
rect 20349 12427 20407 12433
rect 20349 12393 20361 12427
rect 20395 12424 20407 12427
rect 20898 12424 20904 12436
rect 20395 12396 20904 12424
rect 20395 12393 20407 12396
rect 20349 12387 20407 12393
rect 20898 12384 20904 12396
rect 20956 12384 20962 12436
rect 21453 12427 21511 12433
rect 21453 12393 21465 12427
rect 21499 12424 21511 12427
rect 22204 12424 22232 12452
rect 21499 12396 22232 12424
rect 21499 12393 21511 12396
rect 21453 12387 21511 12393
rect 16025 12359 16083 12365
rect 16025 12325 16037 12359
rect 16071 12356 16083 12359
rect 16390 12356 16396 12368
rect 16071 12328 16396 12356
rect 16071 12325 16083 12328
rect 16025 12319 16083 12325
rect 16390 12316 16396 12328
rect 16448 12316 16454 12368
rect 17770 12316 17776 12368
rect 17828 12356 17834 12368
rect 18598 12356 18604 12368
rect 17828 12328 18604 12356
rect 17828 12316 17834 12328
rect 18598 12316 18604 12328
rect 18656 12316 18662 12368
rect 18800 12356 18828 12384
rect 18966 12356 18972 12368
rect 18800 12328 18972 12356
rect 18966 12316 18972 12328
rect 19024 12316 19030 12368
rect 15013 12291 15071 12297
rect 15013 12257 15025 12291
rect 15059 12257 15071 12291
rect 15013 12251 15071 12257
rect 16850 12248 16856 12300
rect 16908 12248 16914 12300
rect 20088 12288 20116 12384
rect 20990 12356 20996 12368
rect 17503 12260 19104 12288
rect 13044 12192 13768 12220
rect 13044 12180 13050 12192
rect 13814 12180 13820 12232
rect 13872 12220 13878 12232
rect 13872 12193 15330 12220
rect 13872 12192 15283 12193
rect 13872 12180 13878 12192
rect 8202 12152 8208 12164
rect 4908 12124 8208 12152
rect 4249 12115 4307 12121
rect 2038 12044 2044 12096
rect 2096 12044 2102 12096
rect 3234 12044 3240 12096
rect 3292 12084 3298 12096
rect 3418 12084 3424 12096
rect 3292 12056 3424 12084
rect 3292 12044 3298 12056
rect 3418 12044 3424 12056
rect 3476 12044 3482 12096
rect 3789 12087 3847 12093
rect 3789 12053 3801 12087
rect 3835 12084 3847 12087
rect 4264 12084 4292 12115
rect 8202 12112 8208 12124
rect 8260 12112 8266 12164
rect 11624 12124 11836 12152
rect 3835 12056 4292 12084
rect 3835 12053 3847 12056
rect 3789 12047 3847 12053
rect 6362 12044 6368 12096
rect 6420 12084 6426 12096
rect 6822 12084 6828 12096
rect 6420 12056 6828 12084
rect 6420 12044 6426 12056
rect 6822 12044 6828 12056
rect 6880 12044 6886 12096
rect 7282 12044 7288 12096
rect 7340 12084 7346 12096
rect 8110 12084 8116 12096
rect 7340 12056 8116 12084
rect 7340 12044 7346 12056
rect 8110 12044 8116 12056
rect 8168 12044 8174 12096
rect 9490 12044 9496 12096
rect 9548 12084 9554 12096
rect 11624 12084 11652 12124
rect 9548 12056 11652 12084
rect 9548 12044 9554 12056
rect 11698 12044 11704 12096
rect 11756 12044 11762 12096
rect 11808 12084 11836 12124
rect 11974 12112 11980 12164
rect 12032 12152 12038 12164
rect 13446 12152 13452 12164
rect 12032 12124 13452 12152
rect 12032 12112 12038 12124
rect 13446 12112 13452 12124
rect 13504 12112 13510 12164
rect 15271 12159 15283 12192
rect 15317 12190 15330 12193
rect 15317 12159 15332 12190
rect 15930 12180 15936 12232
rect 15988 12220 15994 12232
rect 17095 12223 17153 12229
rect 17095 12220 17107 12223
rect 15988 12192 17107 12220
rect 15988 12180 15994 12192
rect 17095 12189 17107 12192
rect 17141 12220 17153 12223
rect 17218 12220 17224 12232
rect 17141 12192 17224 12220
rect 17141 12189 17153 12192
rect 17095 12183 17153 12189
rect 17218 12180 17224 12192
rect 17276 12180 17282 12232
rect 15271 12153 15332 12159
rect 15304 12152 15332 12153
rect 17503 12152 17531 12260
rect 19076 12232 19104 12260
rect 19628 12260 20116 12288
rect 20180 12328 20996 12356
rect 18233 12223 18291 12229
rect 18233 12220 18245 12223
rect 15304 12124 17531 12152
rect 17880 12192 18245 12220
rect 14642 12084 14648 12096
rect 11808 12056 14648 12084
rect 14642 12044 14648 12056
rect 14700 12044 14706 12096
rect 15654 12044 15660 12096
rect 15712 12084 15718 12096
rect 16114 12084 16120 12096
rect 15712 12056 16120 12084
rect 15712 12044 15718 12056
rect 16114 12044 16120 12056
rect 16172 12044 16178 12096
rect 17218 12044 17224 12096
rect 17276 12084 17282 12096
rect 17586 12084 17592 12096
rect 17276 12056 17592 12084
rect 17276 12044 17282 12056
rect 17586 12044 17592 12056
rect 17644 12044 17650 12096
rect 17678 12044 17684 12096
rect 17736 12084 17742 12096
rect 17880 12093 17908 12192
rect 18233 12189 18245 12192
rect 18279 12189 18291 12223
rect 18233 12183 18291 12189
rect 18414 12180 18420 12232
rect 18472 12180 18478 12232
rect 18693 12223 18751 12229
rect 18693 12189 18705 12223
rect 18739 12189 18751 12223
rect 18693 12183 18751 12189
rect 18708 12096 18736 12183
rect 19058 12180 19064 12232
rect 19116 12180 19122 12232
rect 19426 12180 19432 12232
rect 19484 12180 19490 12232
rect 19628 12229 19656 12260
rect 19613 12223 19671 12229
rect 19613 12189 19625 12223
rect 19659 12189 19671 12223
rect 19613 12183 19671 12189
rect 19886 12180 19892 12232
rect 19944 12180 19950 12232
rect 19978 12180 19984 12232
rect 20036 12180 20042 12232
rect 20180 12229 20208 12328
rect 20990 12316 20996 12328
rect 21048 12316 21054 12368
rect 20622 12288 20628 12300
rect 20272 12260 20628 12288
rect 20272 12229 20300 12260
rect 20622 12248 20628 12260
rect 20680 12248 20686 12300
rect 20165 12223 20223 12229
rect 20165 12189 20177 12223
rect 20211 12189 20223 12223
rect 20165 12183 20223 12189
rect 20257 12223 20315 12229
rect 20257 12189 20269 12223
rect 20303 12189 20315 12223
rect 20257 12183 20315 12189
rect 20438 12180 20444 12232
rect 20496 12180 20502 12232
rect 20530 12180 20536 12232
rect 20588 12180 20594 12232
rect 20714 12180 20720 12232
rect 20772 12220 20778 12232
rect 20901 12223 20959 12229
rect 20901 12220 20913 12223
rect 20772 12192 20913 12220
rect 20772 12180 20778 12192
rect 20901 12189 20913 12192
rect 20947 12189 20959 12223
rect 20901 12183 20959 12189
rect 21269 12223 21327 12229
rect 21269 12189 21281 12223
rect 21315 12220 21327 12223
rect 22830 12220 22836 12232
rect 21315 12192 22836 12220
rect 21315 12189 21327 12192
rect 21269 12183 21327 12189
rect 22830 12180 22836 12192
rect 22888 12180 22894 12232
rect 20622 12152 20628 12164
rect 19720 12124 20628 12152
rect 17865 12087 17923 12093
rect 17865 12084 17877 12087
rect 17736 12056 17877 12084
rect 17736 12044 17742 12056
rect 17865 12053 17877 12056
rect 17911 12053 17923 12087
rect 17865 12047 17923 12053
rect 18322 12044 18328 12096
rect 18380 12044 18386 12096
rect 18506 12044 18512 12096
rect 18564 12044 18570 12096
rect 18690 12044 18696 12096
rect 18748 12044 18754 12096
rect 19720 12093 19748 12124
rect 20622 12112 20628 12124
rect 20680 12112 20686 12164
rect 22186 12152 22192 12164
rect 21008 12124 22192 12152
rect 19705 12087 19763 12093
rect 19705 12053 19717 12087
rect 19751 12053 19763 12087
rect 19705 12047 19763 12053
rect 20165 12087 20223 12093
rect 20165 12053 20177 12087
rect 20211 12084 20223 12087
rect 20346 12084 20352 12096
rect 20211 12056 20352 12084
rect 20211 12053 20223 12056
rect 20165 12047 20223 12053
rect 20346 12044 20352 12056
rect 20404 12044 20410 12096
rect 20717 12087 20775 12093
rect 20717 12053 20729 12087
rect 20763 12084 20775 12087
rect 21008 12084 21036 12124
rect 22186 12112 22192 12124
rect 22244 12112 22250 12164
rect 20763 12056 21036 12084
rect 20763 12053 20775 12056
rect 20717 12047 20775 12053
rect 21082 12044 21088 12096
rect 21140 12044 21146 12096
rect 1104 11994 22056 12016
rect 1104 11942 6148 11994
rect 6200 11942 6212 11994
rect 6264 11942 6276 11994
rect 6328 11942 6340 11994
rect 6392 11942 6404 11994
rect 6456 11942 11346 11994
rect 11398 11942 11410 11994
rect 11462 11942 11474 11994
rect 11526 11942 11538 11994
rect 11590 11942 11602 11994
rect 11654 11942 16544 11994
rect 16596 11942 16608 11994
rect 16660 11942 16672 11994
rect 16724 11942 16736 11994
rect 16788 11942 16800 11994
rect 16852 11942 21742 11994
rect 21794 11942 21806 11994
rect 21858 11942 21870 11994
rect 21922 11942 21934 11994
rect 21986 11942 21998 11994
rect 22050 11942 22056 11994
rect 1104 11920 22056 11942
rect 1397 11883 1455 11889
rect 1397 11849 1409 11883
rect 1443 11880 1455 11883
rect 1578 11880 1584 11892
rect 1443 11852 1584 11880
rect 1443 11849 1455 11852
rect 1397 11843 1455 11849
rect 1578 11840 1584 11852
rect 1636 11840 1642 11892
rect 2682 11840 2688 11892
rect 2740 11840 2746 11892
rect 4522 11880 4528 11892
rect 3326 11852 4528 11880
rect 1412 11784 1716 11812
rect 1412 11756 1440 11784
rect 1394 11704 1400 11756
rect 1452 11704 1458 11756
rect 1688 11753 1716 11784
rect 1762 11772 1768 11824
rect 1820 11772 1826 11824
rect 3326 11812 3354 11852
rect 4522 11840 4528 11852
rect 4580 11840 4586 11892
rect 4706 11840 4712 11892
rect 4764 11880 4770 11892
rect 4982 11880 4988 11892
rect 4764 11852 4988 11880
rect 4764 11840 4770 11852
rect 4982 11840 4988 11852
rect 5040 11880 5046 11892
rect 5626 11880 5632 11892
rect 5040 11852 5632 11880
rect 5040 11840 5046 11852
rect 5626 11840 5632 11852
rect 5684 11840 5690 11892
rect 5721 11883 5779 11889
rect 5721 11849 5733 11883
rect 5767 11880 5779 11883
rect 6546 11880 6552 11892
rect 5767 11852 6552 11880
rect 5767 11849 5779 11852
rect 5721 11843 5779 11849
rect 6546 11840 6552 11852
rect 6604 11840 6610 11892
rect 6730 11840 6736 11892
rect 6788 11880 6794 11892
rect 6917 11883 6975 11889
rect 6917 11880 6929 11883
rect 6788 11852 6929 11880
rect 6788 11840 6794 11852
rect 6917 11849 6929 11852
rect 6963 11849 6975 11883
rect 6917 11843 6975 11849
rect 8202 11840 8208 11892
rect 8260 11880 8266 11892
rect 14277 11883 14335 11889
rect 14277 11880 14289 11883
rect 8260 11852 14289 11880
rect 8260 11840 8266 11852
rect 14277 11849 14289 11852
rect 14323 11849 14335 11883
rect 14277 11843 14335 11849
rect 16040 11852 16342 11880
rect 2240 11784 3354 11812
rect 3436 11784 5212 11812
rect 1581 11747 1639 11753
rect 1581 11713 1593 11747
rect 1627 11713 1639 11747
rect 1581 11707 1639 11713
rect 1673 11747 1731 11753
rect 1673 11713 1685 11747
rect 1719 11713 1731 11747
rect 1780 11744 1808 11772
rect 1947 11747 2005 11753
rect 1947 11744 1959 11747
rect 1780 11716 1959 11744
rect 1673 11707 1731 11713
rect 1947 11713 1959 11716
rect 1993 11744 2005 11747
rect 2240 11744 2268 11784
rect 1993 11716 2268 11744
rect 1993 11713 2005 11716
rect 1947 11707 2005 11713
rect 1596 11540 1624 11707
rect 2314 11704 2320 11756
rect 2372 11744 2378 11756
rect 2866 11744 2872 11756
rect 2372 11716 2872 11744
rect 2372 11704 2378 11716
rect 2866 11704 2872 11716
rect 2924 11704 2930 11756
rect 3329 11747 3387 11753
rect 3329 11713 3341 11747
rect 3375 11744 3387 11747
rect 3436 11744 3464 11784
rect 3375 11716 3464 11744
rect 3375 11713 3387 11716
rect 3329 11707 3387 11713
rect 3510 11704 3516 11756
rect 3568 11744 3574 11756
rect 3603 11747 3661 11753
rect 3603 11744 3615 11747
rect 3568 11716 3615 11744
rect 3568 11704 3574 11716
rect 3603 11713 3615 11716
rect 3649 11744 3661 11747
rect 3970 11744 3976 11756
rect 3649 11716 3976 11744
rect 3649 11713 3661 11716
rect 3603 11707 3661 11713
rect 3970 11704 3976 11716
rect 4028 11704 4034 11756
rect 4706 11704 4712 11756
rect 4764 11704 4770 11756
rect 4982 11744 4988 11756
rect 4943 11716 4988 11744
rect 4982 11704 4988 11716
rect 5040 11704 5046 11756
rect 5184 11744 5212 11784
rect 5258 11772 5264 11824
rect 5316 11812 5322 11824
rect 5902 11812 5908 11824
rect 5316 11784 5908 11812
rect 5316 11772 5322 11784
rect 5902 11772 5908 11784
rect 5960 11772 5966 11824
rect 5994 11772 6000 11824
rect 6052 11812 6058 11824
rect 6052 11784 6408 11812
rect 6052 11772 6058 11784
rect 6270 11744 6276 11756
rect 5184 11716 6276 11744
rect 6270 11704 6276 11716
rect 6328 11704 6334 11756
rect 6380 11728 6408 11784
rect 9600 11784 10272 11812
rect 9600 11756 9628 11784
rect 6439 11747 6497 11753
rect 6439 11728 6451 11747
rect 6380 11713 6451 11728
rect 6485 11744 6497 11747
rect 6485 11713 6500 11744
rect 6380 11700 6500 11713
rect 7098 11704 7104 11756
rect 7156 11704 7162 11756
rect 7374 11704 7380 11756
rect 7432 11704 7438 11756
rect 8570 11704 8576 11756
rect 8628 11704 8634 11756
rect 9582 11704 9588 11756
rect 9640 11704 9646 11756
rect 10042 11704 10048 11756
rect 10100 11704 10106 11756
rect 10244 11744 10272 11784
rect 14458 11772 14464 11824
rect 14516 11812 14522 11824
rect 14826 11812 14832 11824
rect 14516 11784 14832 11812
rect 14516 11772 14522 11784
rect 14826 11772 14832 11784
rect 14884 11812 14890 11824
rect 15013 11815 15071 11821
rect 15013 11812 15025 11815
rect 14884 11784 15025 11812
rect 14884 11772 14890 11784
rect 15013 11781 15025 11784
rect 15059 11781 15071 11815
rect 15013 11775 15071 11781
rect 15381 11815 15439 11821
rect 15381 11781 15393 11815
rect 15427 11812 15439 11815
rect 16040 11812 16068 11852
rect 15427 11784 16068 11812
rect 16117 11815 16175 11821
rect 15427 11781 15439 11784
rect 15381 11775 15439 11781
rect 16117 11781 16129 11815
rect 16163 11812 16175 11815
rect 16314 11812 16342 11852
rect 18506 11840 18512 11892
rect 18564 11840 18570 11892
rect 19058 11840 19064 11892
rect 19116 11840 19122 11892
rect 19518 11840 19524 11892
rect 19576 11880 19582 11892
rect 19794 11880 19800 11892
rect 19576 11852 19800 11880
rect 19576 11840 19582 11852
rect 19794 11840 19800 11852
rect 19852 11840 19858 11892
rect 20346 11840 20352 11892
rect 20404 11840 20410 11892
rect 20438 11840 20444 11892
rect 20496 11880 20502 11892
rect 21361 11883 21419 11889
rect 21361 11880 21373 11883
rect 20496 11852 21373 11880
rect 20496 11840 20502 11852
rect 21361 11849 21373 11852
rect 21407 11849 21419 11883
rect 21361 11843 21419 11849
rect 16574 11812 16580 11824
rect 16163 11784 16252 11812
rect 16314 11784 16580 11812
rect 16163 11781 16175 11784
rect 16117 11775 16175 11781
rect 16224 11756 16252 11784
rect 16574 11772 16580 11784
rect 16632 11772 16638 11824
rect 18524 11812 18552 11840
rect 16960 11784 18552 11812
rect 10303 11747 10361 11753
rect 10303 11744 10315 11747
rect 10244 11716 10315 11744
rect 10303 11713 10315 11716
rect 10349 11744 10361 11747
rect 10349 11716 11560 11744
rect 10349 11713 10361 11716
rect 10303 11707 10361 11713
rect 3050 11636 3056 11688
rect 3108 11676 3114 11688
rect 3234 11676 3240 11688
rect 3108 11648 3240 11676
rect 3108 11636 3114 11648
rect 3234 11636 3240 11648
rect 3292 11636 3298 11688
rect 5552 11648 6224 11676
rect 3050 11540 3056 11552
rect 1596 11512 3056 11540
rect 3050 11500 3056 11512
rect 3108 11500 3114 11552
rect 4341 11543 4399 11549
rect 4341 11509 4353 11543
rect 4387 11540 4399 11543
rect 5552 11540 5580 11648
rect 6196 11608 6224 11648
rect 7006 11636 7012 11688
rect 7064 11676 7070 11688
rect 7558 11676 7564 11688
rect 7064 11648 7564 11676
rect 7064 11636 7070 11648
rect 7558 11636 7564 11648
rect 7616 11636 7622 11688
rect 8294 11636 8300 11688
rect 8352 11636 8358 11688
rect 8435 11679 8493 11685
rect 8435 11645 8447 11679
rect 8481 11676 8493 11679
rect 9766 11676 9772 11688
rect 8481 11648 9772 11676
rect 8481 11645 8493 11648
rect 8435 11639 8493 11645
rect 9766 11636 9772 11648
rect 9824 11636 9830 11688
rect 8021 11611 8079 11617
rect 8021 11608 8033 11611
rect 6196 11580 8033 11608
rect 8021 11577 8033 11580
rect 8067 11577 8079 11611
rect 11532 11608 11560 11716
rect 11882 11704 11888 11756
rect 11940 11744 11946 11756
rect 11940 11716 12572 11744
rect 11940 11704 11946 11716
rect 12544 11688 12572 11716
rect 13354 11704 13360 11756
rect 13412 11704 13418 11756
rect 13538 11753 13544 11756
rect 13495 11747 13544 11753
rect 13495 11713 13507 11747
rect 13541 11713 13544 11747
rect 13495 11707 13544 11713
rect 13538 11704 13544 11707
rect 13596 11704 13602 11756
rect 13630 11704 13636 11756
rect 13688 11704 13694 11756
rect 14274 11704 14280 11756
rect 14332 11744 14338 11756
rect 15102 11744 15108 11756
rect 14332 11716 15108 11744
rect 14332 11704 14338 11716
rect 15102 11704 15108 11716
rect 15160 11744 15166 11756
rect 15289 11747 15347 11753
rect 15289 11744 15301 11747
rect 15160 11716 15301 11744
rect 15160 11704 15166 11716
rect 15289 11713 15301 11716
rect 15335 11713 15347 11747
rect 15289 11707 15347 11713
rect 15746 11704 15752 11756
rect 15804 11704 15810 11756
rect 11606 11636 11612 11688
rect 11664 11676 11670 11688
rect 12437 11679 12495 11685
rect 12437 11676 12449 11679
rect 11664 11648 12449 11676
rect 11664 11636 11670 11648
rect 12437 11645 12449 11648
rect 12483 11645 12495 11679
rect 12437 11639 12495 11645
rect 12526 11636 12532 11688
rect 12584 11676 12590 11688
rect 12621 11679 12679 11685
rect 12621 11676 12633 11679
rect 12584 11648 12633 11676
rect 12584 11636 12590 11648
rect 12621 11645 12633 11648
rect 12667 11645 12679 11679
rect 12621 11639 12679 11645
rect 16038 11662 16068 11710
rect 16206 11704 16212 11756
rect 16264 11704 16270 11756
rect 16960 11753 16988 11784
rect 19076 11763 19104 11840
rect 20364 11812 20392 11840
rect 20364 11784 21036 11812
rect 19059 11757 19117 11763
rect 16945 11747 17003 11753
rect 16945 11713 16957 11747
rect 16991 11713 17003 11747
rect 16945 11707 17003 11713
rect 17034 11704 17040 11756
rect 17092 11744 17098 11756
rect 17221 11747 17279 11753
rect 17221 11744 17233 11747
rect 17092 11716 17233 11744
rect 17092 11704 17098 11716
rect 17221 11713 17233 11716
rect 17267 11744 17279 11747
rect 17310 11744 17316 11756
rect 17267 11716 17316 11744
rect 17267 11713 17279 11716
rect 17221 11707 17279 11713
rect 17310 11704 17316 11716
rect 17368 11704 17374 11756
rect 17488 11747 17546 11753
rect 17488 11713 17500 11747
rect 17534 11744 17546 11747
rect 18690 11744 18696 11756
rect 17534 11716 18696 11744
rect 17534 11713 17546 11716
rect 17488 11707 17546 11713
rect 18690 11704 18696 11716
rect 18748 11704 18754 11756
rect 19059 11723 19071 11757
rect 19105 11723 19117 11757
rect 19059 11717 19117 11723
rect 19794 11704 19800 11756
rect 19852 11744 19858 11756
rect 21008 11753 21036 11784
rect 20533 11747 20591 11753
rect 20533 11744 20545 11747
rect 19852 11716 20545 11744
rect 19852 11704 19858 11716
rect 20533 11713 20545 11716
rect 20579 11713 20591 11747
rect 20533 11707 20591 11713
rect 20993 11747 21051 11753
rect 20993 11713 21005 11747
rect 21039 11713 21051 11747
rect 20993 11707 21051 11713
rect 21174 11704 21180 11756
rect 21232 11744 21238 11756
rect 21545 11747 21603 11753
rect 21545 11744 21557 11747
rect 21232 11716 21557 11744
rect 21232 11704 21238 11716
rect 21545 11713 21557 11716
rect 21591 11713 21603 11747
rect 21545 11707 21603 11713
rect 12986 11608 12992 11620
rect 11532 11580 12992 11608
rect 8021 11571 8079 11577
rect 12986 11568 12992 11580
rect 13044 11568 13050 11620
rect 13078 11568 13084 11620
rect 13136 11568 13142 11620
rect 16038 11608 16066 11662
rect 18506 11636 18512 11688
rect 18564 11676 18570 11688
rect 18785 11679 18843 11685
rect 18785 11676 18797 11679
rect 18564 11648 18797 11676
rect 18564 11636 18570 11648
rect 18785 11645 18797 11648
rect 18831 11645 18843 11679
rect 18785 11639 18843 11645
rect 19978 11636 19984 11688
rect 20036 11636 20042 11688
rect 20257 11679 20315 11685
rect 20257 11645 20269 11679
rect 20303 11645 20315 11679
rect 20257 11639 20315 11645
rect 16390 11608 16396 11620
rect 16038 11580 16396 11608
rect 16390 11568 16396 11580
rect 16448 11568 16454 11620
rect 19797 11611 19855 11617
rect 19797 11577 19809 11611
rect 19843 11608 19855 11611
rect 19996 11608 20024 11636
rect 20272 11608 20300 11639
rect 19843 11580 20300 11608
rect 19843 11577 19855 11580
rect 19797 11571 19855 11577
rect 20990 11568 20996 11620
rect 21048 11568 21054 11620
rect 4387 11512 5580 11540
rect 4387 11509 4399 11512
rect 4341 11503 4399 11509
rect 5718 11500 5724 11552
rect 5776 11540 5782 11552
rect 6549 11543 6607 11549
rect 6549 11540 6561 11543
rect 5776 11512 6561 11540
rect 5776 11500 5782 11512
rect 6549 11509 6561 11512
rect 6595 11509 6607 11543
rect 6549 11503 6607 11509
rect 6638 11500 6644 11552
rect 6696 11540 6702 11552
rect 7282 11540 7288 11552
rect 6696 11512 7288 11540
rect 6696 11500 6702 11512
rect 7282 11500 7288 11512
rect 7340 11540 7346 11552
rect 7926 11540 7932 11552
rect 7340 11512 7932 11540
rect 7340 11500 7346 11512
rect 7926 11500 7932 11512
rect 7984 11500 7990 11552
rect 8110 11500 8116 11552
rect 8168 11540 8174 11552
rect 9217 11543 9275 11549
rect 9217 11540 9229 11543
rect 8168 11512 9229 11540
rect 8168 11500 8174 11512
rect 9217 11509 9229 11512
rect 9263 11509 9275 11543
rect 9217 11503 9275 11509
rect 11057 11543 11115 11549
rect 11057 11509 11069 11543
rect 11103 11540 11115 11543
rect 12342 11540 12348 11552
rect 11103 11512 12348 11540
rect 11103 11509 11115 11512
rect 11057 11503 11115 11509
rect 12342 11500 12348 11512
rect 12400 11500 12406 11552
rect 13354 11500 13360 11552
rect 13412 11540 13418 11552
rect 13630 11540 13636 11552
rect 13412 11512 13636 11540
rect 13412 11500 13418 11512
rect 13630 11500 13636 11512
rect 13688 11500 13694 11552
rect 16301 11543 16359 11549
rect 16301 11509 16313 11543
rect 16347 11540 16359 11543
rect 16482 11540 16488 11552
rect 16347 11512 16488 11540
rect 16347 11509 16359 11512
rect 16301 11503 16359 11509
rect 16482 11500 16488 11512
rect 16540 11500 16546 11552
rect 17037 11543 17095 11549
rect 17037 11509 17049 11543
rect 17083 11540 17095 11543
rect 17862 11540 17868 11552
rect 17083 11512 17868 11540
rect 17083 11509 17095 11512
rect 17037 11503 17095 11509
rect 17862 11500 17868 11512
rect 17920 11500 17926 11552
rect 18601 11543 18659 11549
rect 18601 11509 18613 11543
rect 18647 11540 18659 11543
rect 18782 11540 18788 11552
rect 18647 11512 18788 11540
rect 18647 11509 18659 11512
rect 18601 11503 18659 11509
rect 18782 11500 18788 11512
rect 18840 11500 18846 11552
rect 1104 11450 21896 11472
rect 1104 11398 3549 11450
rect 3601 11398 3613 11450
rect 3665 11398 3677 11450
rect 3729 11398 3741 11450
rect 3793 11398 3805 11450
rect 3857 11398 8747 11450
rect 8799 11398 8811 11450
rect 8863 11398 8875 11450
rect 8927 11398 8939 11450
rect 8991 11398 9003 11450
rect 9055 11398 13945 11450
rect 13997 11398 14009 11450
rect 14061 11398 14073 11450
rect 14125 11398 14137 11450
rect 14189 11398 14201 11450
rect 14253 11398 19143 11450
rect 19195 11398 19207 11450
rect 19259 11398 19271 11450
rect 19323 11398 19335 11450
rect 19387 11398 19399 11450
rect 19451 11398 21896 11450
rect 1104 11376 21896 11398
rect 2222 11296 2228 11348
rect 2280 11336 2286 11348
rect 3329 11339 3387 11345
rect 2280 11308 3004 11336
rect 2280 11296 2286 11308
rect 934 11228 940 11280
rect 992 11268 998 11280
rect 1857 11271 1915 11277
rect 1857 11268 1869 11271
rect 992 11240 1869 11268
rect 992 11228 998 11240
rect 1857 11237 1869 11240
rect 1903 11237 1915 11271
rect 1857 11231 1915 11237
rect 2332 11209 2360 11308
rect 2317 11203 2375 11209
rect 2317 11169 2329 11203
rect 2363 11169 2375 11203
rect 2317 11163 2375 11169
rect 1578 11092 1584 11144
rect 1636 11132 1642 11144
rect 1673 11135 1731 11141
rect 1673 11132 1685 11135
rect 1636 11104 1685 11132
rect 1636 11092 1642 11104
rect 1673 11101 1685 11104
rect 1719 11101 1731 11135
rect 2976 11132 3004 11308
rect 3329 11305 3341 11339
rect 3375 11305 3387 11339
rect 3329 11299 3387 11305
rect 3344 11200 3372 11299
rect 3418 11296 3424 11348
rect 3476 11296 3482 11348
rect 3602 11296 3608 11348
rect 3660 11336 3666 11348
rect 3970 11336 3976 11348
rect 3660 11308 3976 11336
rect 3660 11296 3666 11308
rect 3970 11296 3976 11308
rect 4028 11296 4034 11348
rect 4062 11296 4068 11348
rect 4120 11336 4126 11348
rect 6733 11339 6791 11345
rect 4120 11308 6500 11336
rect 4120 11296 4126 11308
rect 3436 11268 3464 11296
rect 4982 11268 4988 11280
rect 3436 11240 4988 11268
rect 4982 11228 4988 11240
rect 5040 11268 5046 11280
rect 6472 11268 6500 11308
rect 6733 11305 6745 11339
rect 6779 11336 6791 11339
rect 7098 11336 7104 11348
rect 6779 11308 7104 11336
rect 6779 11305 6791 11308
rect 6733 11299 6791 11305
rect 7098 11296 7104 11308
rect 7156 11296 7162 11348
rect 7193 11339 7251 11345
rect 7193 11305 7205 11339
rect 7239 11305 7251 11339
rect 7193 11299 7251 11305
rect 7208 11268 7236 11299
rect 8202 11296 8208 11348
rect 8260 11336 8266 11348
rect 8941 11339 8999 11345
rect 8941 11336 8953 11339
rect 8260 11308 8953 11336
rect 8260 11296 8266 11308
rect 8941 11305 8953 11308
rect 8987 11305 8999 11339
rect 8941 11299 8999 11305
rect 9030 11296 9036 11348
rect 9088 11336 9094 11348
rect 9674 11336 9680 11348
rect 9088 11308 9680 11336
rect 9088 11296 9094 11308
rect 9674 11296 9680 11308
rect 9732 11296 9738 11348
rect 10778 11336 10784 11348
rect 9968 11308 10784 11336
rect 5040 11240 5672 11268
rect 6472 11240 7236 11268
rect 8481 11271 8539 11277
rect 5040 11228 5046 11240
rect 4246 11200 4252 11212
rect 3344 11172 4252 11200
rect 4246 11160 4252 11172
rect 4304 11160 4310 11212
rect 4893 11203 4951 11209
rect 4893 11169 4905 11203
rect 4939 11200 4951 11203
rect 5442 11200 5448 11212
rect 4939 11172 5448 11200
rect 4939 11169 4951 11172
rect 4893 11163 4951 11169
rect 5442 11160 5448 11172
rect 5500 11160 5506 11212
rect 5534 11160 5540 11212
rect 5592 11160 5598 11212
rect 5644 11200 5672 11240
rect 8481 11237 8493 11271
rect 8527 11268 8539 11271
rect 9861 11271 9919 11277
rect 9861 11268 9873 11271
rect 8527 11240 9873 11268
rect 8527 11237 8539 11240
rect 8481 11231 8539 11237
rect 9861 11237 9873 11240
rect 9907 11237 9919 11271
rect 9861 11231 9919 11237
rect 5994 11209 6000 11212
rect 5813 11203 5871 11209
rect 5813 11200 5825 11203
rect 5644 11172 5825 11200
rect 5813 11169 5825 11172
rect 5859 11169 5871 11203
rect 5813 11163 5871 11169
rect 5951 11203 6000 11209
rect 5951 11169 5963 11203
rect 5997 11169 6000 11203
rect 5951 11163 6000 11169
rect 5994 11160 6000 11163
rect 6052 11160 6058 11212
rect 6454 11160 6460 11212
rect 6512 11200 6518 11212
rect 6512 11172 6960 11200
rect 6512 11160 6518 11172
rect 2575 11105 2633 11111
rect 2575 11102 2587 11105
rect 1673 11095 1731 11101
rect 934 11024 940 11076
rect 992 11064 998 11076
rect 2406 11064 2412 11076
rect 992 11036 2412 11064
rect 992 11024 998 11036
rect 2406 11024 2412 11036
rect 2464 11064 2470 11076
rect 2574 11071 2587 11102
rect 2621 11071 2633 11105
rect 2976 11104 4200 11132
rect 4172 11076 4200 11104
rect 4430 11092 4436 11144
rect 4488 11132 4494 11144
rect 4617 11135 4675 11141
rect 4617 11132 4629 11135
rect 4488 11104 4629 11132
rect 4488 11092 4494 11104
rect 4617 11101 4629 11104
rect 4663 11101 4675 11135
rect 4617 11095 4675 11101
rect 5077 11135 5135 11141
rect 5077 11101 5089 11135
rect 5123 11101 5135 11135
rect 5077 11095 5135 11101
rect 2574 11065 2633 11071
rect 2574 11064 2602 11065
rect 2464 11036 2602 11064
rect 2464 11024 2470 11036
rect 3050 11024 3056 11076
rect 3108 11064 3114 11076
rect 3786 11064 3792 11076
rect 3108 11036 3792 11064
rect 3108 11024 3114 11036
rect 3786 11024 3792 11036
rect 3844 11024 3850 11076
rect 4154 11024 4160 11076
rect 4212 11024 4218 11076
rect 4246 11024 4252 11076
rect 4304 11024 4310 11076
rect 4798 11024 4804 11076
rect 4856 11064 4862 11076
rect 5092 11064 5120 11095
rect 6086 11092 6092 11144
rect 6144 11092 6150 11144
rect 6822 11092 6828 11144
rect 6880 11092 6886 11144
rect 6932 11141 6960 11172
rect 7282 11160 7288 11212
rect 7340 11200 7346 11212
rect 7469 11203 7527 11209
rect 7469 11200 7481 11203
rect 7340 11172 7481 11200
rect 7340 11160 7346 11172
rect 7469 11169 7481 11172
rect 7515 11169 7527 11203
rect 9766 11200 9772 11212
rect 7469 11163 7527 11169
rect 8266 11172 9168 11200
rect 6917 11135 6975 11141
rect 6917 11101 6929 11135
rect 6963 11101 6975 11135
rect 7742 11132 7748 11144
rect 7703 11104 7748 11132
rect 6917 11095 6975 11101
rect 7742 11092 7748 11104
rect 7800 11092 7806 11144
rect 4856 11036 5120 11064
rect 6840 11064 6868 11092
rect 8266 11064 8294 11172
rect 9030 11092 9036 11144
rect 9088 11092 9094 11144
rect 9140 11141 9168 11172
rect 9416 11172 9772 11200
rect 9416 11141 9444 11172
rect 9766 11160 9772 11172
rect 9824 11160 9830 11212
rect 9968 11200 9996 11308
rect 10778 11296 10784 11308
rect 10836 11336 10842 11348
rect 10836 11308 11928 11336
rect 10836 11296 10842 11308
rect 10870 11228 10876 11280
rect 10928 11228 10934 11280
rect 11790 11228 11796 11280
rect 11848 11228 11854 11280
rect 10137 11203 10195 11209
rect 10137 11200 10149 11203
rect 9968 11172 10149 11200
rect 10137 11169 10149 11172
rect 10183 11169 10195 11203
rect 10137 11163 10195 11169
rect 10275 11203 10333 11209
rect 10275 11169 10287 11203
rect 10321 11200 10333 11203
rect 10888 11200 10916 11228
rect 10321 11172 10916 11200
rect 10321 11169 10333 11172
rect 10275 11163 10333 11169
rect 11330 11160 11336 11212
rect 11388 11160 11394 11212
rect 11900 11200 11928 11308
rect 12066 11296 12072 11348
rect 12124 11336 12130 11348
rect 12989 11339 13047 11345
rect 12989 11336 13001 11339
rect 12124 11308 13001 11336
rect 12124 11296 12130 11308
rect 12989 11305 13001 11308
rect 13035 11305 13047 11339
rect 12989 11299 13047 11305
rect 13354 11296 13360 11348
rect 13412 11336 13418 11348
rect 15105 11339 15163 11345
rect 15105 11336 15117 11339
rect 13412 11308 15117 11336
rect 13412 11296 13418 11308
rect 15105 11305 15117 11308
rect 15151 11305 15163 11339
rect 15286 11336 15292 11348
rect 15105 11299 15163 11305
rect 15212 11308 15292 11336
rect 13538 11268 13544 11280
rect 13372 11240 13544 11268
rect 12066 11200 12072 11212
rect 11900 11172 12072 11200
rect 12066 11160 12072 11172
rect 12124 11160 12130 11212
rect 13372 11200 13400 11240
rect 13538 11228 13544 11240
rect 13596 11228 13602 11280
rect 12222 11172 13400 11200
rect 9125 11135 9183 11141
rect 9125 11101 9137 11135
rect 9171 11101 9183 11135
rect 9125 11095 9183 11101
rect 9217 11135 9275 11141
rect 9217 11101 9229 11135
rect 9263 11101 9275 11135
rect 9217 11095 9275 11101
rect 9401 11135 9459 11141
rect 9401 11101 9413 11135
rect 9447 11101 9459 11135
rect 9401 11095 9459 11101
rect 6840 11036 8294 11064
rect 9048 11064 9076 11092
rect 9232 11064 9260 11095
rect 10410 11092 10416 11144
rect 10468 11092 10474 11144
rect 11149 11135 11207 11141
rect 11149 11101 11161 11135
rect 11195 11132 11207 11135
rect 11238 11132 11244 11144
rect 11195 11104 11244 11132
rect 11195 11101 11207 11104
rect 11149 11095 11207 11101
rect 11238 11092 11244 11104
rect 11296 11092 11302 11144
rect 12222 11141 12250 11172
rect 13446 11160 13452 11212
rect 13504 11200 13510 11212
rect 14090 11200 14096 11212
rect 13504 11172 14096 11200
rect 13504 11160 13510 11172
rect 14090 11160 14096 11172
rect 14148 11160 14154 11212
rect 12207 11135 12265 11141
rect 12207 11101 12219 11135
rect 12253 11101 12265 11135
rect 12207 11095 12265 11101
rect 12342 11092 12348 11144
rect 12400 11092 12406 11144
rect 12986 11092 12992 11144
rect 13044 11132 13050 11144
rect 14367 11135 14425 11141
rect 13044 11104 14320 11132
rect 13044 11092 13050 11104
rect 9048 11036 9260 11064
rect 4856 11024 4862 11036
rect 11054 11024 11060 11076
rect 11112 11024 11118 11076
rect 13538 11064 13544 11076
rect 13372 11036 13544 11064
rect 2866 10956 2872 11008
rect 2924 10996 2930 11008
rect 6638 10996 6644 11008
rect 2924 10968 6644 10996
rect 2924 10956 2930 10968
rect 6638 10956 6644 10968
rect 6696 10956 6702 11008
rect 7006 10956 7012 11008
rect 7064 10996 7070 11008
rect 10962 10996 10968 11008
rect 7064 10968 10968 10996
rect 7064 10956 7070 10968
rect 10962 10956 10968 10968
rect 11020 10956 11026 11008
rect 12066 10956 12072 11008
rect 12124 10996 12130 11008
rect 13372 10996 13400 11036
rect 13538 11024 13544 11036
rect 13596 11024 13602 11076
rect 14292 11064 14320 11104
rect 14367 11101 14379 11135
rect 14413 11132 14425 11135
rect 15212 11132 15240 11308
rect 15286 11296 15292 11308
rect 15344 11336 15350 11348
rect 15344 11308 16252 11336
rect 15344 11296 15350 11308
rect 15562 11160 15568 11212
rect 15620 11160 15626 11212
rect 15807 11135 15865 11141
rect 15807 11132 15819 11135
rect 14413 11104 15240 11132
rect 15286 11104 15819 11132
rect 14413 11101 14425 11104
rect 14367 11095 14425 11101
rect 14918 11064 14924 11076
rect 14292 11036 14924 11064
rect 14918 11024 14924 11036
rect 14976 11064 14982 11076
rect 15286 11064 15314 11104
rect 15807 11101 15819 11104
rect 15853 11132 15865 11135
rect 15930 11132 15936 11144
rect 15853 11104 15936 11132
rect 15853 11101 15865 11104
rect 15807 11095 15865 11101
rect 15930 11092 15936 11104
rect 15988 11092 15994 11144
rect 16224 11132 16252 11308
rect 16574 11296 16580 11348
rect 16632 11296 16638 11348
rect 17678 11336 17684 11348
rect 17604 11308 17684 11336
rect 17604 11209 17632 11308
rect 17678 11296 17684 11308
rect 17736 11296 17742 11348
rect 18414 11296 18420 11348
rect 18472 11336 18478 11348
rect 18693 11339 18751 11345
rect 18693 11336 18705 11339
rect 18472 11308 18705 11336
rect 18472 11296 18478 11308
rect 18693 11305 18705 11308
rect 18739 11305 18751 11339
rect 18693 11299 18751 11305
rect 19794 11296 19800 11348
rect 19852 11296 19858 11348
rect 19334 11268 19340 11280
rect 17696 11240 19340 11268
rect 17589 11203 17647 11209
rect 17589 11169 17601 11203
rect 17635 11169 17647 11203
rect 17589 11163 17647 11169
rect 17696 11132 17724 11240
rect 19334 11228 19340 11240
rect 19392 11228 19398 11280
rect 19429 11271 19487 11277
rect 19429 11237 19441 11271
rect 19475 11268 19487 11271
rect 19702 11268 19708 11280
rect 19475 11240 19708 11268
rect 19475 11237 19487 11240
rect 19429 11231 19487 11237
rect 19702 11228 19708 11240
rect 19760 11228 19766 11280
rect 19981 11203 20039 11209
rect 19981 11200 19993 11203
rect 17788 11172 19993 11200
rect 17788 11144 17816 11172
rect 19981 11169 19993 11172
rect 20027 11169 20039 11203
rect 19981 11163 20039 11169
rect 16224 11104 17724 11132
rect 17770 11092 17776 11144
rect 17828 11092 17834 11144
rect 17862 11092 17868 11144
rect 17920 11092 17926 11144
rect 18322 11092 18328 11144
rect 18380 11092 18386 11144
rect 18782 11092 18788 11144
rect 18840 11132 18846 11144
rect 18877 11135 18935 11141
rect 18877 11132 18889 11135
rect 18840 11104 18889 11132
rect 18840 11092 18846 11104
rect 18877 11101 18889 11104
rect 18923 11101 18935 11135
rect 18877 11095 18935 11101
rect 19613 11135 19671 11141
rect 19613 11101 19625 11135
rect 19659 11101 19671 11135
rect 19613 11095 19671 11101
rect 14976 11036 15314 11064
rect 14976 11024 14982 11036
rect 16298 11024 16304 11076
rect 16356 11064 16362 11076
rect 18601 11067 18659 11073
rect 18601 11064 18613 11067
rect 16356 11036 18613 11064
rect 16356 11024 16362 11036
rect 18601 11033 18613 11036
rect 18647 11033 18659 11067
rect 18601 11027 18659 11033
rect 12124 10968 13400 10996
rect 12124 10956 12130 10968
rect 13446 10956 13452 11008
rect 13504 10996 13510 11008
rect 18138 10996 18144 11008
rect 13504 10968 18144 10996
rect 13504 10956 13510 10968
rect 18138 10956 18144 10968
rect 18196 10956 18202 11008
rect 19628 10996 19656 11095
rect 19702 11092 19708 11144
rect 19760 11092 19766 11144
rect 20226 11067 20284 11073
rect 20226 11064 20238 11067
rect 19870 11036 20238 11064
rect 19702 10996 19708 11008
rect 19628 10968 19708 10996
rect 19702 10956 19708 10968
rect 19760 10996 19766 11008
rect 19870 10996 19898 11036
rect 20226 11033 20238 11036
rect 20272 11033 20284 11067
rect 20226 11027 20284 11033
rect 19760 10968 19898 10996
rect 19760 10956 19766 10968
rect 21358 10956 21364 11008
rect 21416 10956 21422 11008
rect 1104 10906 22056 10928
rect 1104 10854 6148 10906
rect 6200 10854 6212 10906
rect 6264 10854 6276 10906
rect 6328 10854 6340 10906
rect 6392 10854 6404 10906
rect 6456 10854 11346 10906
rect 11398 10854 11410 10906
rect 11462 10854 11474 10906
rect 11526 10854 11538 10906
rect 11590 10854 11602 10906
rect 11654 10854 16544 10906
rect 16596 10854 16608 10906
rect 16660 10854 16672 10906
rect 16724 10854 16736 10906
rect 16788 10854 16800 10906
rect 16852 10854 21742 10906
rect 21794 10854 21806 10906
rect 21858 10854 21870 10906
rect 21922 10854 21934 10906
rect 21986 10854 21998 10906
rect 22050 10854 22056 10906
rect 1104 10832 22056 10854
rect 3786 10752 3792 10804
rect 3844 10792 3850 10804
rect 6181 10795 6239 10801
rect 6181 10792 6193 10795
rect 3844 10764 6193 10792
rect 3844 10752 3850 10764
rect 6181 10761 6193 10764
rect 6227 10761 6239 10795
rect 6181 10755 6239 10761
rect 6362 10752 6368 10804
rect 6420 10792 6426 10804
rect 7650 10792 7656 10804
rect 6420 10764 7656 10792
rect 6420 10752 6426 10764
rect 7650 10752 7656 10764
rect 7708 10752 7714 10804
rect 8297 10795 8355 10801
rect 8297 10761 8309 10795
rect 8343 10792 8355 10795
rect 8570 10792 8576 10804
rect 8343 10764 8576 10792
rect 8343 10761 8355 10764
rect 8297 10755 8355 10761
rect 8570 10752 8576 10764
rect 8628 10752 8634 10804
rect 9677 10795 9735 10801
rect 9677 10761 9689 10795
rect 9723 10792 9735 10795
rect 10410 10792 10416 10804
rect 9723 10764 10416 10792
rect 9723 10761 9735 10764
rect 9677 10755 9735 10761
rect 10410 10752 10416 10764
rect 10468 10752 10474 10804
rect 11057 10795 11115 10801
rect 11057 10761 11069 10795
rect 11103 10792 11115 10795
rect 11882 10792 11888 10804
rect 11103 10764 11888 10792
rect 11103 10761 11115 10764
rect 11057 10755 11115 10761
rect 11882 10752 11888 10764
rect 11940 10752 11946 10804
rect 13262 10792 13268 10804
rect 12636 10764 13268 10792
rect 1210 10684 1216 10736
rect 1268 10724 1274 10736
rect 1673 10727 1731 10733
rect 1673 10724 1685 10727
rect 1268 10696 1685 10724
rect 1268 10684 1274 10696
rect 1673 10693 1685 10696
rect 1719 10693 1731 10727
rect 4430 10724 4436 10736
rect 1673 10687 1731 10693
rect 4080 10696 4436 10724
rect 2317 10659 2375 10665
rect 2317 10625 2329 10659
rect 2363 10656 2375 10659
rect 2363 10628 2728 10656
rect 2363 10625 2375 10628
rect 2317 10619 2375 10625
rect 2700 10600 2728 10628
rect 3510 10616 3516 10668
rect 3568 10616 3574 10668
rect 2406 10548 2412 10600
rect 2464 10588 2470 10600
rect 2501 10591 2559 10597
rect 2501 10588 2513 10591
rect 2464 10560 2513 10588
rect 2464 10548 2470 10560
rect 2501 10557 2513 10560
rect 2547 10557 2559 10591
rect 2501 10551 2559 10557
rect 2682 10548 2688 10600
rect 2740 10548 2746 10600
rect 2866 10548 2872 10600
rect 2924 10588 2930 10600
rect 3237 10591 3295 10597
rect 3237 10588 3249 10591
rect 2924 10560 3249 10588
rect 2924 10548 2930 10560
rect 3237 10557 3249 10560
rect 3283 10557 3295 10591
rect 3237 10551 3295 10557
rect 3375 10591 3433 10597
rect 3375 10557 3387 10591
rect 3421 10588 3433 10591
rect 3878 10588 3884 10600
rect 3421 10560 3884 10588
rect 3421 10557 3433 10560
rect 3375 10551 3433 10557
rect 3878 10548 3884 10560
rect 3936 10548 3942 10600
rect 4080 10588 4108 10696
rect 4430 10684 4436 10696
rect 4488 10684 4494 10736
rect 9122 10684 9128 10736
rect 9180 10724 9186 10736
rect 9180 10696 10272 10724
rect 9180 10684 9186 10696
rect 10244 10668 10272 10696
rect 4525 10659 4583 10665
rect 4525 10625 4537 10659
rect 4571 10656 4583 10659
rect 4706 10656 4712 10668
rect 4571 10628 4712 10656
rect 4571 10625 4583 10628
rect 4525 10619 4583 10625
rect 4706 10616 4712 10628
rect 4764 10616 4770 10668
rect 5350 10616 5356 10668
rect 5408 10665 5414 10668
rect 5408 10659 5436 10665
rect 5424 10625 5436 10659
rect 5408 10619 5436 10625
rect 5408 10616 5414 10619
rect 5534 10616 5540 10668
rect 5592 10616 5598 10668
rect 6641 10659 6699 10665
rect 6641 10625 6653 10659
rect 6687 10656 6699 10659
rect 6822 10656 6828 10668
rect 6687 10628 6828 10656
rect 6687 10625 6699 10628
rect 6641 10619 6699 10625
rect 6822 10616 6828 10628
rect 6880 10616 6886 10668
rect 7527 10659 7585 10665
rect 7527 10656 7539 10659
rect 6932 10628 7539 10656
rect 4341 10591 4399 10597
rect 4341 10588 4353 10591
rect 4080 10560 4353 10588
rect 4341 10557 4353 10560
rect 4387 10557 4399 10591
rect 5261 10591 5319 10597
rect 5261 10588 5273 10591
rect 4341 10551 4399 10557
rect 4448 10560 5273 10588
rect 1210 10480 1216 10532
rect 1268 10520 1274 10532
rect 2961 10523 3019 10529
rect 1268 10492 1882 10520
rect 1268 10480 1274 10492
rect 1762 10412 1768 10464
rect 1820 10412 1826 10464
rect 1854 10452 1882 10492
rect 2961 10489 2973 10523
rect 3007 10520 3019 10523
rect 3050 10520 3056 10532
rect 3007 10492 3056 10520
rect 3007 10489 3019 10492
rect 2961 10483 3019 10489
rect 3050 10480 3056 10492
rect 3108 10480 3114 10532
rect 3896 10520 3924 10548
rect 4448 10520 4476 10560
rect 5261 10557 5273 10560
rect 5307 10557 5319 10591
rect 5261 10551 5319 10557
rect 3896 10492 4476 10520
rect 4982 10480 4988 10532
rect 5040 10480 5046 10532
rect 6932 10464 6960 10628
rect 7527 10625 7539 10628
rect 7573 10625 7585 10659
rect 7527 10619 7585 10625
rect 8939 10659 8997 10665
rect 8939 10625 8951 10659
rect 8985 10656 8997 10659
rect 9582 10656 9588 10668
rect 8985 10628 9588 10656
rect 8985 10625 8997 10628
rect 8939 10619 8997 10625
rect 9582 10616 9588 10628
rect 9640 10616 9646 10668
rect 9674 10616 9680 10668
rect 9732 10656 9738 10668
rect 10042 10656 10048 10668
rect 9732 10628 10048 10656
rect 9732 10616 9738 10628
rect 10042 10616 10048 10628
rect 10100 10616 10106 10668
rect 10226 10616 10232 10668
rect 10284 10616 10290 10668
rect 10318 10616 10324 10668
rect 10376 10656 10382 10668
rect 12636 10665 12664 10764
rect 13262 10752 13268 10764
rect 13320 10792 13326 10804
rect 13446 10792 13452 10804
rect 13320 10764 13452 10792
rect 13320 10752 13326 10764
rect 13446 10752 13452 10764
rect 13504 10752 13510 10804
rect 14090 10752 14096 10804
rect 14148 10792 14154 10804
rect 14148 10764 14596 10792
rect 14148 10752 14154 10764
rect 12621 10659 12679 10665
rect 10376 10628 10419 10656
rect 10376 10616 10382 10628
rect 12621 10625 12633 10659
rect 12667 10625 12679 10659
rect 12621 10619 12679 10625
rect 13538 10616 13544 10668
rect 13596 10616 13602 10668
rect 13630 10616 13636 10668
rect 13688 10665 13694 10668
rect 14568 10665 14596 10764
rect 14642 10752 14648 10804
rect 14700 10792 14706 10804
rect 17034 10792 17040 10804
rect 14700 10764 17040 10792
rect 14700 10752 14706 10764
rect 17034 10752 17040 10764
rect 17092 10752 17098 10804
rect 17310 10752 17316 10804
rect 17368 10792 17374 10804
rect 17770 10792 17776 10804
rect 17368 10764 17776 10792
rect 17368 10752 17374 10764
rect 17770 10752 17776 10764
rect 17828 10752 17834 10804
rect 19334 10752 19340 10804
rect 19392 10792 19398 10804
rect 19794 10792 19800 10804
rect 19392 10764 19800 10792
rect 19392 10752 19398 10764
rect 19794 10752 19800 10764
rect 19852 10752 19858 10804
rect 19886 10752 19892 10804
rect 19944 10792 19950 10804
rect 20533 10795 20591 10801
rect 20533 10792 20545 10795
rect 19944 10764 20545 10792
rect 19944 10752 19950 10764
rect 20533 10761 20545 10764
rect 20579 10761 20591 10795
rect 20533 10755 20591 10761
rect 21453 10795 21511 10801
rect 21453 10761 21465 10795
rect 21499 10792 21511 10795
rect 22186 10792 22192 10804
rect 21499 10764 22192 10792
rect 21499 10761 21511 10764
rect 21453 10755 21511 10761
rect 22186 10752 22192 10764
rect 22244 10752 22250 10804
rect 19306 10696 19564 10724
rect 13688 10659 13716 10665
rect 13704 10625 13716 10659
rect 13688 10619 13716 10625
rect 14553 10659 14611 10665
rect 14553 10625 14565 10659
rect 14599 10625 14611 10659
rect 14553 10619 14611 10625
rect 13688 10616 13694 10619
rect 14734 10616 14740 10668
rect 14792 10656 14798 10668
rect 14827 10659 14885 10665
rect 14827 10656 14839 10659
rect 14792 10628 14839 10656
rect 14792 10616 14798 10628
rect 14827 10625 14839 10628
rect 14873 10656 14885 10659
rect 17555 10659 17613 10665
rect 17555 10656 17567 10659
rect 14873 10628 17567 10656
rect 14873 10625 14885 10628
rect 14827 10619 14885 10625
rect 17555 10625 17567 10628
rect 17601 10656 17613 10659
rect 19306 10656 19334 10696
rect 17601 10628 19334 10656
rect 17601 10625 17613 10628
rect 17555 10619 17613 10625
rect 19426 10616 19432 10668
rect 19484 10616 19490 10668
rect 19536 10656 19564 10696
rect 20714 10684 20720 10736
rect 20772 10724 20778 10736
rect 21177 10727 21235 10733
rect 21177 10724 21189 10727
rect 20772 10696 21189 10724
rect 20772 10684 20778 10696
rect 21177 10693 21189 10696
rect 21223 10693 21235 10727
rect 21177 10687 21235 10693
rect 19763 10659 19821 10665
rect 19763 10656 19775 10659
rect 19536 10628 19775 10656
rect 19763 10625 19775 10628
rect 19809 10625 19821 10659
rect 19763 10619 19821 10625
rect 7282 10548 7288 10600
rect 7340 10548 7346 10600
rect 8665 10591 8723 10597
rect 8665 10557 8677 10591
rect 8711 10557 8723 10591
rect 8665 10551 8723 10557
rect 3602 10452 3608 10464
rect 1854 10424 3608 10452
rect 3602 10412 3608 10424
rect 3660 10412 3666 10464
rect 4154 10412 4160 10464
rect 4212 10412 4218 10464
rect 5718 10412 5724 10464
rect 5776 10452 5782 10464
rect 5902 10452 5908 10464
rect 5776 10424 5908 10452
rect 5776 10412 5782 10424
rect 5902 10412 5908 10424
rect 5960 10412 5966 10464
rect 6454 10412 6460 10464
rect 6512 10412 6518 10464
rect 6914 10412 6920 10464
rect 6972 10412 6978 10464
rect 7300 10452 7328 10548
rect 7558 10452 7564 10464
rect 7300 10424 7564 10452
rect 7558 10412 7564 10424
rect 7616 10452 7622 10464
rect 8680 10452 8708 10551
rect 11882 10548 11888 10600
rect 11940 10588 11946 10600
rect 12526 10588 12532 10600
rect 11940 10560 12532 10588
rect 11940 10548 11946 10560
rect 12526 10548 12532 10560
rect 12584 10588 12590 10600
rect 12805 10591 12863 10597
rect 12805 10588 12817 10591
rect 12584 10560 12817 10588
rect 12584 10548 12590 10560
rect 12805 10557 12817 10560
rect 12851 10588 12863 10591
rect 13265 10591 13323 10597
rect 12851 10560 13124 10588
rect 12851 10557 12863 10560
rect 12805 10551 12863 10557
rect 13096 10464 13124 10560
rect 13265 10557 13277 10591
rect 13311 10588 13323 10591
rect 13354 10588 13360 10600
rect 13311 10560 13360 10588
rect 13311 10557 13323 10560
rect 13265 10551 13323 10557
rect 13354 10548 13360 10560
rect 13412 10548 13418 10600
rect 13817 10591 13875 10597
rect 13817 10557 13829 10591
rect 13863 10588 13875 10591
rect 13863 10560 14504 10588
rect 13863 10557 13875 10560
rect 13817 10551 13875 10557
rect 14476 10520 14504 10560
rect 17218 10548 17224 10600
rect 17276 10588 17282 10600
rect 17313 10591 17371 10597
rect 17313 10588 17325 10591
rect 17276 10560 17325 10588
rect 17276 10548 17282 10560
rect 17313 10557 17325 10560
rect 17359 10557 17371 10591
rect 17313 10551 17371 10557
rect 14476 10492 14596 10520
rect 7616 10424 8708 10452
rect 7616 10412 7622 10424
rect 9030 10412 9036 10464
rect 9088 10452 9094 10464
rect 10318 10452 10324 10464
rect 9088 10424 10324 10452
rect 9088 10412 9094 10424
rect 10318 10412 10324 10424
rect 10376 10412 10382 10464
rect 13078 10412 13084 10464
rect 13136 10412 13142 10464
rect 13722 10412 13728 10464
rect 13780 10452 13786 10464
rect 14461 10455 14519 10461
rect 14461 10452 14473 10455
rect 13780 10424 14473 10452
rect 13780 10412 13786 10424
rect 14461 10421 14473 10424
rect 14507 10421 14519 10455
rect 14568 10452 14596 10492
rect 15286 10480 15292 10532
rect 15344 10520 15350 10532
rect 15746 10520 15752 10532
rect 15344 10492 15752 10520
rect 15344 10480 15350 10492
rect 15746 10480 15752 10492
rect 15804 10480 15810 10532
rect 15565 10455 15623 10461
rect 15565 10452 15577 10455
rect 14568 10424 15577 10452
rect 14461 10415 14519 10421
rect 15565 10421 15577 10424
rect 15611 10421 15623 10455
rect 17328 10452 17356 10551
rect 18414 10548 18420 10600
rect 18472 10548 18478 10600
rect 19518 10548 19524 10600
rect 19576 10548 19582 10600
rect 18432 10520 18460 10548
rect 17972 10492 18460 10520
rect 17972 10452 18000 10492
rect 17328 10424 18000 10452
rect 15565 10415 15623 10421
rect 18322 10412 18328 10464
rect 18380 10412 18386 10464
rect 19245 10455 19303 10461
rect 19245 10421 19257 10455
rect 19291 10452 19303 10455
rect 20346 10452 20352 10464
rect 19291 10424 20352 10452
rect 19291 10421 19303 10424
rect 19245 10415 19303 10421
rect 20346 10412 20352 10424
rect 20404 10412 20410 10464
rect 1104 10362 21896 10384
rect 1104 10310 3549 10362
rect 3601 10310 3613 10362
rect 3665 10310 3677 10362
rect 3729 10310 3741 10362
rect 3793 10310 3805 10362
rect 3857 10310 8747 10362
rect 8799 10310 8811 10362
rect 8863 10310 8875 10362
rect 8927 10310 8939 10362
rect 8991 10310 9003 10362
rect 9055 10310 13945 10362
rect 13997 10310 14009 10362
rect 14061 10310 14073 10362
rect 14125 10310 14137 10362
rect 14189 10310 14201 10362
rect 14253 10310 19143 10362
rect 19195 10310 19207 10362
rect 19259 10310 19271 10362
rect 19323 10310 19335 10362
rect 19387 10310 19399 10362
rect 19451 10310 21896 10362
rect 1104 10288 21896 10310
rect 1486 10208 1492 10260
rect 1544 10248 1550 10260
rect 1670 10248 1676 10260
rect 1544 10220 1676 10248
rect 1544 10208 1550 10220
rect 1670 10208 1676 10220
rect 1728 10208 1734 10260
rect 2133 10251 2191 10257
rect 2133 10217 2145 10251
rect 2179 10248 2191 10251
rect 2774 10248 2780 10260
rect 2179 10220 2780 10248
rect 2179 10217 2191 10220
rect 2133 10211 2191 10217
rect 2774 10208 2780 10220
rect 2832 10208 2838 10260
rect 3326 10208 3332 10260
rect 3384 10208 3390 10260
rect 3970 10208 3976 10260
rect 4028 10208 4034 10260
rect 4525 10251 4583 10257
rect 4525 10217 4537 10251
rect 4571 10217 4583 10251
rect 4525 10211 4583 10217
rect 3050 10140 3056 10192
rect 3108 10180 3114 10192
rect 4540 10180 4568 10211
rect 5994 10208 6000 10260
rect 6052 10248 6058 10260
rect 6089 10251 6147 10257
rect 6089 10248 6101 10251
rect 6052 10220 6101 10248
rect 6052 10208 6058 10220
rect 6089 10217 6101 10220
rect 6135 10217 6147 10251
rect 10413 10251 10471 10257
rect 6089 10211 6147 10217
rect 6656 10220 10088 10248
rect 3108 10152 4568 10180
rect 3108 10140 3114 10152
rect 6656 10124 6684 10220
rect 6748 10152 7420 10180
rect 1394 10072 1400 10124
rect 1452 10112 1458 10124
rect 2317 10115 2375 10121
rect 2317 10112 2329 10115
rect 1452 10084 2329 10112
rect 1452 10072 1458 10084
rect 2317 10081 2329 10084
rect 2363 10081 2375 10115
rect 4062 10112 4068 10124
rect 2317 10075 2375 10081
rect 3804 10084 4068 10112
rect 1857 10047 1915 10053
rect 1857 10013 1869 10047
rect 1903 10044 1915 10047
rect 2130 10044 2136 10056
rect 1903 10016 2136 10044
rect 1903 10013 1915 10016
rect 1857 10007 1915 10013
rect 2130 10004 2136 10016
rect 2188 10004 2194 10056
rect 2591 10047 2649 10053
rect 2591 10013 2603 10047
rect 2637 10044 2649 10047
rect 3050 10044 3056 10056
rect 2637 10016 3056 10044
rect 2637 10013 2649 10016
rect 2591 10007 2649 10013
rect 3050 10004 3056 10016
rect 3108 10004 3114 10056
rect 3804 9976 3832 10084
rect 4062 10072 4068 10084
rect 4120 10112 4126 10124
rect 5077 10115 5135 10121
rect 5077 10112 5089 10115
rect 4120 10084 5089 10112
rect 4120 10072 4126 10084
rect 5077 10081 5089 10084
rect 5123 10081 5135 10115
rect 5077 10075 5135 10081
rect 6638 10072 6644 10124
rect 6696 10072 6702 10124
rect 4522 10004 4528 10056
rect 4580 10044 4586 10056
rect 5351 10047 5409 10053
rect 5351 10044 5363 10047
rect 4580 10016 5363 10044
rect 4580 10004 4586 10016
rect 5351 10013 5363 10016
rect 5397 10044 5409 10047
rect 6362 10044 6368 10056
rect 5397 10016 6368 10044
rect 5397 10013 5409 10016
rect 5351 10007 5409 10013
rect 6362 10004 6368 10016
rect 6420 10004 6426 10056
rect 6454 10004 6460 10056
rect 6512 10004 6518 10056
rect 2148 9948 3832 9976
rect 2148 9920 2176 9948
rect 3878 9936 3884 9988
rect 3936 9936 3942 9988
rect 4433 9979 4491 9985
rect 4433 9945 4445 9979
rect 4479 9976 4491 9979
rect 6472 9976 6500 10004
rect 4479 9948 6500 9976
rect 4479 9945 4491 9948
rect 4433 9939 4491 9945
rect 2130 9868 2136 9920
rect 2188 9868 2194 9920
rect 2866 9868 2872 9920
rect 2924 9908 2930 9920
rect 4614 9908 4620 9920
rect 2924 9880 4620 9908
rect 2924 9868 2930 9880
rect 4614 9868 4620 9880
rect 4672 9908 4678 9920
rect 6748 9908 6776 10152
rect 6825 10115 6883 10121
rect 6825 10081 6837 10115
rect 6871 10112 6883 10115
rect 7006 10112 7012 10124
rect 6871 10084 7012 10112
rect 6871 10081 6883 10084
rect 6825 10075 6883 10081
rect 7006 10072 7012 10084
rect 7064 10072 7070 10124
rect 7282 10072 7288 10124
rect 7340 10072 7346 10124
rect 7392 10112 7420 10152
rect 8294 10140 8300 10192
rect 8352 10180 8358 10192
rect 8573 10183 8631 10189
rect 8573 10180 8585 10183
rect 8352 10152 8585 10180
rect 8352 10140 8358 10152
rect 8573 10149 8585 10152
rect 8619 10149 8631 10183
rect 10060 10180 10088 10220
rect 10413 10217 10425 10251
rect 10459 10248 10471 10251
rect 10502 10248 10508 10260
rect 10459 10220 10508 10248
rect 10459 10217 10471 10220
rect 10413 10211 10471 10217
rect 10502 10208 10508 10220
rect 10560 10208 10566 10260
rect 14550 10248 14556 10260
rect 10612 10220 14556 10248
rect 10612 10180 10640 10220
rect 14550 10208 14556 10220
rect 14608 10208 14614 10260
rect 15930 10208 15936 10260
rect 15988 10248 15994 10260
rect 18046 10248 18052 10260
rect 15988 10220 18052 10248
rect 15988 10208 15994 10220
rect 18046 10208 18052 10220
rect 18104 10208 18110 10260
rect 18598 10208 18604 10260
rect 18656 10248 18662 10260
rect 20254 10248 20260 10260
rect 18656 10220 20260 10248
rect 18656 10208 18662 10220
rect 20254 10208 20260 10220
rect 20312 10208 20318 10260
rect 20346 10208 20352 10260
rect 20404 10208 20410 10260
rect 20898 10208 20904 10260
rect 20956 10208 20962 10260
rect 12066 10180 12072 10192
rect 10060 10152 10640 10180
rect 11808 10152 12072 10180
rect 8573 10143 8631 10149
rect 7561 10115 7619 10121
rect 7561 10112 7573 10115
rect 7392 10084 7573 10112
rect 7561 10081 7573 10084
rect 7607 10081 7619 10115
rect 7561 10075 7619 10081
rect 7650 10072 7656 10124
rect 7708 10121 7714 10124
rect 7708 10115 7736 10121
rect 7724 10081 7736 10115
rect 7708 10075 7736 10081
rect 7708 10072 7714 10075
rect 10410 10072 10416 10124
rect 10468 10112 10474 10124
rect 11808 10112 11836 10152
rect 12066 10140 12072 10152
rect 12124 10180 12130 10192
rect 12124 10152 12480 10180
rect 12124 10140 12130 10152
rect 10468 10084 11836 10112
rect 10468 10072 10474 10084
rect 11882 10072 11888 10124
rect 11940 10072 11946 10124
rect 12342 10072 12348 10124
rect 12400 10072 12406 10124
rect 12452 10112 12480 10152
rect 18138 10140 18144 10192
rect 18196 10140 18202 10192
rect 18414 10140 18420 10192
rect 18472 10180 18478 10192
rect 18472 10152 19288 10180
rect 18472 10140 18478 10152
rect 12621 10115 12679 10121
rect 12621 10112 12633 10115
rect 12452 10084 12633 10112
rect 12621 10081 12633 10084
rect 12667 10081 12679 10115
rect 12621 10075 12679 10081
rect 12710 10072 12716 10124
rect 12768 10121 12774 10124
rect 12768 10115 12817 10121
rect 12768 10081 12771 10115
rect 12805 10112 12817 10115
rect 12805 10084 13492 10112
rect 12805 10081 12817 10084
rect 12768 10075 12817 10081
rect 12768 10072 12774 10075
rect 7834 10004 7840 10056
rect 7892 10004 7898 10056
rect 8754 10004 8760 10056
rect 8812 10004 8818 10056
rect 9401 10047 9459 10053
rect 9401 10013 9413 10047
rect 9447 10013 9459 10047
rect 9674 10044 9680 10056
rect 9635 10016 9680 10044
rect 9401 10007 9459 10013
rect 9416 9976 9444 10007
rect 9674 10004 9680 10016
rect 9732 10044 9738 10056
rect 10686 10044 10692 10056
rect 9732 10016 10692 10044
rect 9732 10004 9738 10016
rect 10686 10004 10692 10016
rect 10744 10004 10750 10056
rect 11698 10004 11704 10056
rect 11756 10044 11762 10056
rect 11756 10016 11928 10044
rect 11756 10004 11762 10016
rect 11790 9976 11796 9988
rect 9416 9948 11796 9976
rect 11790 9936 11796 9948
rect 11848 9936 11854 9988
rect 4672 9880 6776 9908
rect 4672 9868 4678 9880
rect 8478 9868 8484 9920
rect 8536 9868 8542 9920
rect 9122 9868 9128 9920
rect 9180 9908 9186 9920
rect 11900 9908 11928 10016
rect 12894 10004 12900 10056
rect 12952 10004 12958 10056
rect 13464 10044 13492 10084
rect 13538 10072 13544 10124
rect 13596 10072 13602 10124
rect 15102 10072 15108 10124
rect 15160 10072 15166 10124
rect 16758 10072 16764 10124
rect 16816 10112 16822 10124
rect 16816 10084 19012 10112
rect 16816 10072 16822 10084
rect 14921 10047 14979 10053
rect 13464 10016 14688 10044
rect 14366 9976 14372 9988
rect 13372 9948 14372 9976
rect 13372 9908 13400 9948
rect 14366 9936 14372 9948
rect 14424 9936 14430 9988
rect 9180 9880 13400 9908
rect 9180 9868 9186 9880
rect 14274 9868 14280 9920
rect 14332 9908 14338 9920
rect 14553 9911 14611 9917
rect 14553 9908 14565 9911
rect 14332 9880 14565 9908
rect 14332 9868 14338 9880
rect 14553 9877 14565 9880
rect 14599 9877 14611 9911
rect 14660 9908 14688 10016
rect 14921 10013 14933 10047
rect 14967 10044 14979 10047
rect 14967 10016 15976 10044
rect 14967 10013 14979 10016
rect 14921 10007 14979 10013
rect 14829 9979 14887 9985
rect 14829 9945 14841 9979
rect 14875 9976 14887 9979
rect 15010 9976 15016 9988
rect 14875 9948 15016 9976
rect 14875 9945 14887 9948
rect 14829 9939 14887 9945
rect 15010 9936 15016 9948
rect 15068 9936 15074 9988
rect 15286 9936 15292 9988
rect 15344 9936 15350 9988
rect 15948 9976 15976 10016
rect 16022 10004 16028 10056
rect 16080 10004 16086 10056
rect 16299 10047 16357 10053
rect 16299 10013 16311 10047
rect 16345 10044 16357 10047
rect 16390 10044 16396 10056
rect 16345 10016 16396 10044
rect 16345 10013 16357 10016
rect 16299 10007 16357 10013
rect 16390 10004 16396 10016
rect 16448 10004 16454 10056
rect 17957 10047 18015 10053
rect 17957 10013 17969 10047
rect 18003 10013 18015 10047
rect 17957 10007 18015 10013
rect 17972 9976 18000 10007
rect 18138 10004 18144 10056
rect 18196 10004 18202 10056
rect 18322 10004 18328 10056
rect 18380 10044 18386 10056
rect 18601 10047 18659 10053
rect 18601 10044 18613 10047
rect 18380 10016 18613 10044
rect 18380 10004 18386 10016
rect 18601 10013 18613 10016
rect 18647 10013 18659 10047
rect 18601 10007 18659 10013
rect 18782 10004 18788 10056
rect 18840 10004 18846 10056
rect 18340 9976 18368 10004
rect 15396 9948 15884 9976
rect 15948 9948 17080 9976
rect 17972 9948 18368 9976
rect 18509 9979 18567 9985
rect 15396 9908 15424 9948
rect 14660 9880 15424 9908
rect 15657 9911 15715 9917
rect 14553 9871 14611 9877
rect 15657 9877 15669 9911
rect 15703 9908 15715 9911
rect 15746 9908 15752 9920
rect 15703 9880 15752 9908
rect 15703 9877 15715 9880
rect 15657 9871 15715 9877
rect 15746 9868 15752 9880
rect 15804 9868 15810 9920
rect 15856 9917 15884 9948
rect 17052 9917 17080 9948
rect 18509 9945 18521 9979
rect 18555 9976 18567 9979
rect 18693 9979 18751 9985
rect 18693 9976 18705 9979
rect 18555 9948 18705 9976
rect 18555 9945 18567 9948
rect 18509 9939 18567 9945
rect 18693 9945 18705 9948
rect 18739 9945 18751 9979
rect 18693 9939 18751 9945
rect 15841 9911 15899 9917
rect 15841 9877 15853 9911
rect 15887 9877 15899 9911
rect 15841 9871 15899 9877
rect 17037 9911 17095 9917
rect 17037 9877 17049 9911
rect 17083 9877 17095 9911
rect 17037 9871 17095 9877
rect 17678 9868 17684 9920
rect 17736 9908 17742 9920
rect 18877 9911 18935 9917
rect 18877 9908 18889 9911
rect 17736 9880 18889 9908
rect 17736 9868 17742 9880
rect 18877 9877 18889 9880
rect 18923 9877 18935 9911
rect 18984 9908 19012 10084
rect 19260 10056 19288 10152
rect 19058 10004 19064 10056
rect 19116 10004 19122 10056
rect 19242 10004 19248 10056
rect 19300 10004 19306 10056
rect 20364 10044 20392 10208
rect 20717 10047 20775 10053
rect 20717 10044 20729 10047
rect 19503 10017 19561 10023
rect 19503 9983 19515 10017
rect 19549 10014 19561 10017
rect 20364 10016 20729 10044
rect 19549 9983 19564 10014
rect 20717 10013 20729 10016
rect 20763 10013 20775 10047
rect 20717 10007 20775 10013
rect 19503 9977 19564 9983
rect 19536 9976 19564 9977
rect 19794 9976 19800 9988
rect 19536 9948 19800 9976
rect 19794 9936 19800 9948
rect 19852 9936 19858 9988
rect 19904 9948 20576 9976
rect 19904 9908 19932 9948
rect 20548 9920 20576 9948
rect 21174 9936 21180 9988
rect 21232 9936 21238 9988
rect 21545 9979 21603 9985
rect 21545 9945 21557 9979
rect 21591 9976 21603 9979
rect 22278 9976 22284 9988
rect 21591 9948 22284 9976
rect 21591 9945 21603 9948
rect 21545 9939 21603 9945
rect 22278 9936 22284 9948
rect 22336 9936 22342 9988
rect 18984 9880 19932 9908
rect 18877 9871 18935 9877
rect 20254 9868 20260 9920
rect 20312 9868 20318 9920
rect 20530 9868 20536 9920
rect 20588 9868 20594 9920
rect 1104 9818 22056 9840
rect 1104 9766 6148 9818
rect 6200 9766 6212 9818
rect 6264 9766 6276 9818
rect 6328 9766 6340 9818
rect 6392 9766 6404 9818
rect 6456 9766 11346 9818
rect 11398 9766 11410 9818
rect 11462 9766 11474 9818
rect 11526 9766 11538 9818
rect 11590 9766 11602 9818
rect 11654 9766 16544 9818
rect 16596 9766 16608 9818
rect 16660 9766 16672 9818
rect 16724 9766 16736 9818
rect 16788 9766 16800 9818
rect 16852 9766 21742 9818
rect 21794 9766 21806 9818
rect 21858 9766 21870 9818
rect 21922 9766 21934 9818
rect 21986 9766 21998 9818
rect 22050 9766 22056 9818
rect 1104 9744 22056 9766
rect 3050 9664 3056 9716
rect 3108 9704 3114 9716
rect 5074 9704 5080 9716
rect 3108 9676 5080 9704
rect 3108 9664 3114 9676
rect 5074 9664 5080 9676
rect 5132 9664 5138 9716
rect 6638 9664 6644 9716
rect 6696 9704 6702 9716
rect 7558 9704 7564 9716
rect 6696 9676 7564 9704
rect 6696 9664 6702 9676
rect 7558 9664 7564 9676
rect 7616 9664 7622 9716
rect 8478 9704 8484 9716
rect 8220 9676 8484 9704
rect 1486 9596 1492 9648
rect 1544 9596 1550 9648
rect 1857 9639 1915 9645
rect 1857 9605 1869 9639
rect 1903 9636 1915 9639
rect 1946 9636 1952 9648
rect 1903 9608 1952 9636
rect 1903 9605 1915 9608
rect 1857 9599 1915 9605
rect 1946 9596 1952 9608
rect 2004 9596 2010 9648
rect 8220 9636 8248 9676
rect 8478 9664 8484 9676
rect 8536 9664 8542 9716
rect 8956 9676 10456 9704
rect 7116 9608 8248 9636
rect 2222 9528 2228 9580
rect 2280 9528 2286 9580
rect 2498 9528 2504 9580
rect 2556 9568 2562 9580
rect 3510 9577 3516 9580
rect 2593 9571 2651 9577
rect 2593 9568 2605 9571
rect 2556 9540 2605 9568
rect 2556 9528 2562 9540
rect 2593 9537 2605 9540
rect 2639 9537 2651 9571
rect 2593 9531 2651 9537
rect 3467 9571 3516 9577
rect 3467 9537 3479 9571
rect 3513 9537 3516 9571
rect 3467 9531 3516 9537
rect 3510 9528 3516 9531
rect 3568 9528 3574 9580
rect 4249 9571 4307 9577
rect 4249 9537 4261 9571
rect 4295 9568 4307 9571
rect 4706 9568 4712 9580
rect 4295 9540 4712 9568
rect 4295 9537 4307 9540
rect 4249 9531 4307 9537
rect 4706 9528 4712 9540
rect 4764 9528 4770 9580
rect 5258 9528 5264 9580
rect 5316 9528 5322 9580
rect 5442 9577 5448 9580
rect 5399 9571 5448 9577
rect 5399 9537 5411 9571
rect 5445 9537 5448 9571
rect 5399 9531 5448 9537
rect 5442 9528 5448 9531
rect 5500 9528 5506 9580
rect 6457 9571 6515 9577
rect 6457 9537 6469 9571
rect 6503 9568 6515 9571
rect 6546 9568 6552 9580
rect 6503 9540 6552 9568
rect 6503 9537 6515 9540
rect 6457 9531 6515 9537
rect 6546 9528 6552 9540
rect 6604 9528 6610 9580
rect 6914 9528 6920 9580
rect 6972 9568 6978 9580
rect 7116 9577 7144 9608
rect 7101 9571 7159 9577
rect 6972 9540 7052 9568
rect 6972 9528 6978 9540
rect 1578 9460 1584 9512
rect 1636 9500 1642 9512
rect 1854 9500 1860 9512
rect 1636 9472 1860 9500
rect 1636 9460 1642 9472
rect 1854 9460 1860 9472
rect 1912 9460 1918 9512
rect 2409 9503 2467 9509
rect 2409 9469 2421 9503
rect 2455 9500 2467 9503
rect 3329 9503 3387 9509
rect 3329 9500 3341 9503
rect 2455 9472 2544 9500
rect 2455 9469 2467 9472
rect 2409 9463 2467 9469
rect 2516 9444 2544 9472
rect 2884 9472 3341 9500
rect 2884 9444 2912 9472
rect 3329 9469 3341 9472
rect 3375 9469 3387 9503
rect 3329 9463 3387 9469
rect 3605 9503 3663 9509
rect 3605 9469 3617 9503
rect 3651 9500 3663 9503
rect 3970 9500 3976 9512
rect 3651 9472 3976 9500
rect 3651 9469 3663 9472
rect 3605 9463 3663 9469
rect 3970 9460 3976 9472
rect 4028 9460 4034 9512
rect 4341 9503 4399 9509
rect 4341 9469 4353 9503
rect 4387 9500 4399 9503
rect 4430 9500 4436 9512
rect 4387 9472 4436 9500
rect 4387 9469 4399 9472
rect 4341 9463 4399 9469
rect 4430 9460 4436 9472
rect 4488 9460 4494 9512
rect 4525 9503 4583 9509
rect 4525 9469 4537 9503
rect 4571 9500 4583 9503
rect 4614 9500 4620 9512
rect 4571 9472 4620 9500
rect 4571 9469 4583 9472
rect 4525 9463 4583 9469
rect 4614 9460 4620 9472
rect 4672 9460 4678 9512
rect 5276 9500 5304 9528
rect 4816 9472 5304 9500
rect 4816 9444 4844 9472
rect 5534 9460 5540 9512
rect 5592 9460 5598 9512
rect 5718 9460 5724 9512
rect 5776 9500 5782 9512
rect 7024 9500 7052 9540
rect 7101 9537 7113 9571
rect 7147 9537 7159 9571
rect 7650 9568 7656 9580
rect 7611 9540 7656 9568
rect 7101 9531 7159 9537
rect 7650 9528 7656 9540
rect 7708 9528 7714 9580
rect 7742 9528 7748 9580
rect 7800 9568 7806 9580
rect 8956 9577 8984 9676
rect 10428 9636 10456 9676
rect 10502 9664 10508 9716
rect 10560 9704 10566 9716
rect 10597 9707 10655 9713
rect 10597 9704 10609 9707
rect 10560 9676 10609 9704
rect 10560 9664 10566 9676
rect 10597 9673 10609 9676
rect 10643 9673 10655 9707
rect 13262 9704 13268 9716
rect 10597 9667 10655 9673
rect 12268 9676 13268 9704
rect 10428 9608 11928 9636
rect 8941 9571 8999 9577
rect 8941 9568 8953 9571
rect 7800 9540 8953 9568
rect 7800 9528 7806 9540
rect 8941 9537 8953 9540
rect 8987 9537 8999 9571
rect 8941 9531 8999 9537
rect 9122 9528 9128 9580
rect 9180 9528 9186 9580
rect 9950 9528 9956 9580
rect 10008 9528 10014 9580
rect 10594 9528 10600 9580
rect 10652 9528 10658 9580
rect 10873 9571 10931 9577
rect 10873 9537 10885 9571
rect 10919 9568 10931 9571
rect 11698 9568 11704 9580
rect 10919 9540 11704 9568
rect 10919 9537 10931 9540
rect 10873 9531 10931 9537
rect 11698 9528 11704 9540
rect 11756 9528 11762 9580
rect 7377 9503 7435 9509
rect 7377 9500 7389 9503
rect 5776 9472 6960 9500
rect 7024 9472 7389 9500
rect 5776 9460 5782 9472
rect 2498 9392 2504 9444
rect 2556 9392 2562 9444
rect 2866 9392 2872 9444
rect 2924 9392 2930 9444
rect 3050 9392 3056 9444
rect 3108 9392 3114 9444
rect 4062 9392 4068 9444
rect 4120 9432 4126 9444
rect 4120 9404 4384 9432
rect 4120 9392 4126 9404
rect 2041 9367 2099 9373
rect 2041 9333 2053 9367
rect 2087 9364 2099 9367
rect 4246 9364 4252 9376
rect 2087 9336 4252 9364
rect 2087 9333 2099 9336
rect 2041 9327 2099 9333
rect 4246 9324 4252 9336
rect 4304 9324 4310 9376
rect 4356 9364 4384 9404
rect 4798 9392 4804 9444
rect 4856 9392 4862 9444
rect 4985 9435 5043 9441
rect 4985 9401 4997 9435
rect 5031 9432 5043 9435
rect 5074 9432 5080 9444
rect 5031 9404 5080 9432
rect 5031 9401 5043 9404
rect 4985 9395 5043 9401
rect 5074 9392 5080 9404
rect 5132 9392 5138 9444
rect 6932 9441 6960 9472
rect 7377 9469 7389 9472
rect 7423 9469 7435 9503
rect 7377 9463 7435 9469
rect 8757 9503 8815 9509
rect 8757 9469 8769 9503
rect 8803 9500 8815 9503
rect 9140 9500 9168 9528
rect 9677 9503 9735 9509
rect 9677 9500 9689 9503
rect 8803 9472 9168 9500
rect 9508 9472 9689 9500
rect 8803 9469 8815 9472
rect 8757 9463 8815 9469
rect 6181 9435 6239 9441
rect 6181 9401 6193 9435
rect 6227 9432 6239 9435
rect 6917 9435 6975 9441
rect 6227 9404 6868 9432
rect 6227 9401 6239 9404
rect 6181 9395 6239 9401
rect 6549 9367 6607 9373
rect 6549 9364 6561 9367
rect 4356 9336 6561 9364
rect 6549 9333 6561 9336
rect 6595 9333 6607 9367
rect 6840 9364 6868 9404
rect 6917 9401 6929 9435
rect 6963 9401 6975 9435
rect 6917 9395 6975 9401
rect 8389 9435 8447 9441
rect 8389 9401 8401 9435
rect 8435 9432 8447 9435
rect 9401 9435 9459 9441
rect 9401 9432 9413 9435
rect 8435 9404 9413 9432
rect 8435 9401 8447 9404
rect 8389 9395 8447 9401
rect 9401 9401 9413 9404
rect 9447 9401 9459 9435
rect 9401 9395 9459 9401
rect 8294 9364 8300 9376
rect 6840 9336 8300 9364
rect 6549 9327 6607 9333
rect 8294 9324 8300 9336
rect 8352 9324 8358 9376
rect 9508 9364 9536 9472
rect 9677 9469 9689 9472
rect 9723 9469 9735 9503
rect 9677 9463 9735 9469
rect 9815 9503 9873 9509
rect 9815 9469 9827 9503
rect 9861 9500 9873 9503
rect 10612 9500 10640 9528
rect 11900 9512 11928 9608
rect 12069 9571 12127 9577
rect 12069 9537 12081 9571
rect 12115 9568 12127 9571
rect 12268 9568 12296 9676
rect 13262 9664 13268 9676
rect 13320 9664 13326 9716
rect 14936 9676 15424 9704
rect 13814 9596 13820 9648
rect 13872 9636 13878 9648
rect 13909 9639 13967 9645
rect 13909 9636 13921 9639
rect 13872 9608 13921 9636
rect 13872 9596 13878 9608
rect 13909 9605 13921 9608
rect 13955 9605 13967 9639
rect 13909 9599 13967 9605
rect 14274 9596 14280 9648
rect 14332 9636 14338 9648
rect 14826 9636 14832 9648
rect 14332 9608 14832 9636
rect 14332 9596 14338 9608
rect 14826 9596 14832 9608
rect 14884 9596 14890 9648
rect 12115 9552 12130 9568
rect 12176 9552 12296 9568
rect 12115 9540 12296 9552
rect 12115 9537 12204 9540
rect 12069 9531 12204 9537
rect 12102 9524 12204 9531
rect 13262 9528 13268 9580
rect 13320 9528 13326 9580
rect 14936 9568 14964 9676
rect 15010 9596 15016 9648
rect 15068 9636 15074 9648
rect 15105 9639 15163 9645
rect 15105 9636 15117 9639
rect 15068 9608 15117 9636
rect 15068 9596 15074 9608
rect 15105 9605 15117 9608
rect 15151 9605 15163 9639
rect 15105 9599 15163 9605
rect 15286 9596 15292 9648
rect 15344 9596 15350 9648
rect 15396 9636 15424 9676
rect 15562 9664 15568 9716
rect 15620 9704 15626 9716
rect 16022 9704 16028 9716
rect 15620 9676 16028 9704
rect 15620 9664 15626 9676
rect 16022 9664 16028 9676
rect 16080 9664 16086 9716
rect 18598 9704 18604 9716
rect 17512 9676 18604 9704
rect 15396 9608 15700 9636
rect 14568 9540 14964 9568
rect 9861 9472 10640 9500
rect 9861 9469 9873 9472
rect 9815 9463 9873 9469
rect 11882 9460 11888 9512
rect 11940 9460 11946 9512
rect 12253 9503 12311 9509
rect 12253 9469 12265 9503
rect 12299 9500 12311 9503
rect 12342 9500 12348 9512
rect 12299 9472 12348 9500
rect 12299 9469 12311 9472
rect 12253 9463 12311 9469
rect 12342 9460 12348 9472
rect 12400 9460 12406 9512
rect 12989 9503 13047 9509
rect 12989 9500 13001 9503
rect 12452 9472 13001 9500
rect 12066 9392 12072 9444
rect 12124 9432 12130 9444
rect 12452 9432 12480 9472
rect 12989 9469 13001 9472
rect 13035 9469 13047 9503
rect 12989 9463 13047 9469
rect 13127 9503 13185 9509
rect 13127 9469 13139 9503
rect 13173 9500 13185 9503
rect 14568 9500 14596 9540
rect 15194 9528 15200 9580
rect 15252 9528 15258 9580
rect 15304 9568 15332 9596
rect 15565 9571 15623 9577
rect 15565 9568 15577 9571
rect 15304 9540 15577 9568
rect 15565 9537 15577 9540
rect 15611 9537 15623 9571
rect 15672 9568 15700 9608
rect 15746 9596 15752 9648
rect 15804 9636 15810 9648
rect 15933 9639 15991 9645
rect 15933 9636 15945 9639
rect 15804 9608 15945 9636
rect 15804 9596 15810 9608
rect 15933 9605 15945 9608
rect 15979 9636 15991 9639
rect 16206 9636 16212 9648
rect 15979 9608 16212 9636
rect 15979 9605 15991 9608
rect 15933 9599 15991 9605
rect 16206 9596 16212 9608
rect 16264 9596 16270 9648
rect 16114 9568 16120 9580
rect 15672 9540 16120 9568
rect 15565 9531 15623 9537
rect 16114 9528 16120 9540
rect 16172 9528 16178 9580
rect 16298 9528 16304 9580
rect 16356 9568 16362 9580
rect 17512 9568 17540 9676
rect 18598 9664 18604 9676
rect 18656 9664 18662 9716
rect 19153 9707 19211 9713
rect 19153 9673 19165 9707
rect 19199 9704 19211 9707
rect 19199 9676 19288 9704
rect 19199 9673 19211 9676
rect 19153 9667 19211 9673
rect 17696 9608 18083 9636
rect 17696 9577 17724 9608
rect 18055 9580 18083 9608
rect 18046 9577 18052 9580
rect 16356 9540 17540 9568
rect 17681 9571 17739 9577
rect 16356 9528 16362 9540
rect 17681 9537 17693 9571
rect 17727 9537 17739 9571
rect 18040 9568 18052 9577
rect 18007 9540 18052 9568
rect 17681 9531 17739 9537
rect 18040 9531 18052 9540
rect 18046 9528 18052 9531
rect 18104 9528 18110 9580
rect 18598 9528 18604 9580
rect 18656 9568 18662 9580
rect 19150 9568 19156 9580
rect 18656 9540 19156 9568
rect 18656 9528 18662 9540
rect 19150 9528 19156 9540
rect 19208 9528 19214 9580
rect 19260 9568 19288 9676
rect 19518 9664 19524 9716
rect 19576 9704 19582 9716
rect 20533 9707 20591 9713
rect 20533 9704 20545 9707
rect 19576 9676 20545 9704
rect 19576 9664 19582 9676
rect 20533 9673 20545 9676
rect 20579 9673 20591 9707
rect 20533 9667 20591 9673
rect 19610 9636 19616 9648
rect 19536 9608 19616 9636
rect 19536 9577 19564 9608
rect 19610 9596 19616 9608
rect 19668 9636 19674 9648
rect 19978 9636 19984 9648
rect 19668 9608 19984 9636
rect 19668 9596 19674 9608
rect 19978 9596 19984 9608
rect 20036 9596 20042 9648
rect 19429 9571 19487 9577
rect 19429 9568 19441 9571
rect 19260 9540 19441 9568
rect 19429 9537 19441 9540
rect 19475 9537 19487 9571
rect 19429 9531 19487 9537
rect 19521 9571 19579 9577
rect 19521 9537 19533 9571
rect 19567 9537 19579 9571
rect 19521 9531 19579 9537
rect 19794 9528 19800 9580
rect 19852 9528 19858 9580
rect 19886 9528 19892 9580
rect 19944 9568 19950 9580
rect 20162 9568 20168 9580
rect 19944 9540 20168 9568
rect 19944 9528 19950 9540
rect 20162 9528 20168 9540
rect 20220 9528 20226 9580
rect 20254 9528 20260 9580
rect 20312 9568 20318 9580
rect 20901 9571 20959 9577
rect 20901 9568 20913 9571
rect 20312 9540 20913 9568
rect 20312 9528 20318 9540
rect 20901 9537 20913 9540
rect 20947 9537 20959 9571
rect 20901 9531 20959 9537
rect 21082 9528 21088 9580
rect 21140 9528 21146 9580
rect 21266 9528 21272 9580
rect 21324 9568 21330 9580
rect 21453 9571 21511 9577
rect 21453 9568 21465 9571
rect 21324 9540 21465 9568
rect 21324 9528 21330 9540
rect 21453 9537 21465 9540
rect 21499 9537 21511 9571
rect 21453 9531 21511 9537
rect 13173 9472 14596 9500
rect 13173 9469 13185 9472
rect 13127 9463 13185 9469
rect 15286 9460 15292 9512
rect 15344 9460 15350 9512
rect 12124 9404 12480 9432
rect 12124 9392 12130 9404
rect 12710 9392 12716 9444
rect 12768 9392 12774 9444
rect 14550 9392 14556 9444
rect 14608 9392 14614 9444
rect 16132 9441 16160 9528
rect 17770 9460 17776 9512
rect 17828 9460 17834 9512
rect 16117 9435 16175 9441
rect 16117 9401 16129 9435
rect 16163 9401 16175 9435
rect 16117 9395 16175 9401
rect 16206 9392 16212 9444
rect 16264 9432 16270 9444
rect 16264 9404 17816 9432
rect 16264 9392 16270 9404
rect 9674 9364 9680 9376
rect 9508 9336 9680 9364
rect 9674 9324 9680 9336
rect 9732 9324 9738 9376
rect 9858 9324 9864 9376
rect 9916 9364 9922 9376
rect 10318 9364 10324 9376
rect 9916 9336 10324 9364
rect 9916 9324 9922 9336
rect 10318 9324 10324 9336
rect 10376 9324 10382 9376
rect 10686 9324 10692 9376
rect 10744 9324 10750 9376
rect 11330 9324 11336 9376
rect 11388 9364 11394 9376
rect 12250 9364 12256 9376
rect 11388 9336 12256 9364
rect 11388 9324 11394 9336
rect 12250 9324 12256 9336
rect 12308 9324 12314 9376
rect 13446 9324 13452 9376
rect 13504 9364 13510 9376
rect 14568 9364 14596 9392
rect 13504 9336 14596 9364
rect 13504 9324 13510 9336
rect 17218 9324 17224 9376
rect 17276 9364 17282 9376
rect 17497 9367 17555 9373
rect 17497 9364 17509 9367
rect 17276 9336 17509 9364
rect 17276 9324 17282 9336
rect 17497 9333 17509 9336
rect 17543 9333 17555 9367
rect 17788 9364 17816 9404
rect 18708 9404 19380 9432
rect 18708 9364 18736 9404
rect 17788 9336 18736 9364
rect 17497 9327 17555 9333
rect 18782 9324 18788 9376
rect 18840 9364 18846 9376
rect 19245 9367 19303 9373
rect 19245 9364 19257 9367
rect 18840 9336 19257 9364
rect 18840 9324 18846 9336
rect 19245 9333 19257 9336
rect 19291 9333 19303 9367
rect 19352 9364 19380 9404
rect 20346 9392 20352 9444
rect 20404 9432 20410 9444
rect 21085 9435 21143 9441
rect 21085 9432 21097 9435
rect 20404 9404 21097 9432
rect 20404 9392 20410 9404
rect 21085 9401 21097 9404
rect 21131 9401 21143 9435
rect 21085 9395 21143 9401
rect 22278 9364 22284 9376
rect 19352 9336 22284 9364
rect 19245 9327 19303 9333
rect 22278 9324 22284 9336
rect 22336 9324 22342 9376
rect 1104 9274 21896 9296
rect 1104 9222 3549 9274
rect 3601 9222 3613 9274
rect 3665 9222 3677 9274
rect 3729 9222 3741 9274
rect 3793 9222 3805 9274
rect 3857 9222 8747 9274
rect 8799 9222 8811 9274
rect 8863 9222 8875 9274
rect 8927 9222 8939 9274
rect 8991 9222 9003 9274
rect 9055 9222 13945 9274
rect 13997 9222 14009 9274
rect 14061 9222 14073 9274
rect 14125 9222 14137 9274
rect 14189 9222 14201 9274
rect 14253 9222 19143 9274
rect 19195 9222 19207 9274
rect 19259 9222 19271 9274
rect 19323 9222 19335 9274
rect 19387 9222 19399 9274
rect 19451 9222 21896 9274
rect 1104 9200 21896 9222
rect 1762 9120 1768 9172
rect 1820 9120 1826 9172
rect 2240 9132 3832 9160
rect 2240 9092 2268 9132
rect 1412 9064 2268 9092
rect 1412 9036 1440 9064
rect 3804 9036 3832 9132
rect 4062 9120 4068 9172
rect 4120 9160 4126 9172
rect 4522 9160 4528 9172
rect 4120 9132 4528 9160
rect 4120 9120 4126 9132
rect 4522 9120 4528 9132
rect 4580 9120 4586 9172
rect 4801 9163 4859 9169
rect 4801 9129 4813 9163
rect 4847 9160 4859 9163
rect 5626 9160 5632 9172
rect 4847 9132 5632 9160
rect 4847 9129 4859 9132
rect 4801 9123 4859 9129
rect 5626 9120 5632 9132
rect 5684 9120 5690 9172
rect 6638 9160 6644 9172
rect 5736 9132 6644 9160
rect 5169 9095 5227 9101
rect 5169 9061 5181 9095
rect 5215 9061 5227 9095
rect 5736 9092 5764 9132
rect 6638 9120 6644 9132
rect 6696 9120 6702 9172
rect 7834 9120 7840 9172
rect 7892 9160 7898 9172
rect 8021 9163 8079 9169
rect 8021 9160 8033 9163
rect 7892 9132 8033 9160
rect 7892 9120 7898 9132
rect 8021 9129 8033 9132
rect 8067 9129 8079 9163
rect 9490 9160 9496 9172
rect 8021 9123 8079 9129
rect 9048 9132 9496 9160
rect 5169 9055 5227 9061
rect 5644 9064 5764 9092
rect 1394 8984 1400 9036
rect 1452 8984 1458 9036
rect 2130 8984 2136 9036
rect 2188 8984 2194 9036
rect 3786 8984 3792 9036
rect 3844 8984 3850 9036
rect 4522 8984 4528 9036
rect 4580 9024 4586 9036
rect 5184 9024 5212 9055
rect 4580 8996 5212 9024
rect 4580 8984 4586 8996
rect 5442 8984 5448 9036
rect 5500 9024 5506 9036
rect 5644 9033 5672 9064
rect 5629 9027 5687 9033
rect 5629 9024 5641 9027
rect 5500 8996 5641 9024
rect 5500 8984 5506 8996
rect 5629 8993 5641 8996
rect 5675 8993 5687 9027
rect 5629 8987 5687 8993
rect 6914 8984 6920 9036
rect 6972 9024 6978 9036
rect 7009 9027 7067 9033
rect 7009 9024 7021 9027
rect 6972 8996 7021 9024
rect 6972 8984 6978 8996
rect 7009 8993 7021 8996
rect 7055 8993 7067 9027
rect 7009 8987 7067 8993
rect 8478 8984 8484 9036
rect 8536 9024 8542 9036
rect 9048 9033 9076 9132
rect 9490 9120 9496 9132
rect 9548 9160 9554 9172
rect 9548 9132 9996 9160
rect 9548 9120 9554 9132
rect 9033 9027 9091 9033
rect 9033 9024 9045 9027
rect 8536 8996 9045 9024
rect 8536 8984 8542 8996
rect 9033 8993 9045 8996
rect 9079 8993 9091 9027
rect 9968 9024 9996 9132
rect 10042 9120 10048 9172
rect 10100 9120 10106 9172
rect 11609 9163 11667 9169
rect 10612 9132 11560 9160
rect 10612 9033 10640 9132
rect 10597 9027 10655 9033
rect 10597 9024 10609 9027
rect 9968 8996 10609 9024
rect 9033 8987 9091 8993
rect 10597 8993 10609 8996
rect 10643 8993 10655 9027
rect 10597 8987 10655 8993
rect 2375 8959 2433 8965
rect 2375 8956 2387 8959
rect 492 8928 2387 8956
rect 492 8832 520 8928
rect 2375 8925 2387 8928
rect 2421 8956 2433 8959
rect 2498 8956 2504 8968
rect 2421 8928 2504 8956
rect 2421 8925 2433 8928
rect 2375 8919 2433 8925
rect 2498 8916 2504 8928
rect 2556 8916 2562 8968
rect 3418 8916 3424 8968
rect 3476 8956 3482 8968
rect 3602 8956 3608 8968
rect 3476 8928 3608 8956
rect 3476 8916 3482 8928
rect 3602 8916 3608 8928
rect 3660 8916 3666 8968
rect 4062 8956 4068 8968
rect 4023 8928 4068 8956
rect 4062 8916 4068 8928
rect 4120 8916 4126 8968
rect 4154 8916 4160 8968
rect 4212 8956 4218 8968
rect 5353 8959 5411 8965
rect 5353 8956 5365 8959
rect 4212 8928 5365 8956
rect 4212 8916 4218 8928
rect 5353 8925 5365 8928
rect 5399 8925 5411 8959
rect 5353 8919 5411 8925
rect 5903 8959 5961 8965
rect 5903 8925 5915 8959
rect 5949 8956 5961 8959
rect 6822 8956 6828 8968
rect 5949 8928 6828 8956
rect 5949 8925 5961 8928
rect 5903 8919 5961 8925
rect 6822 8916 6828 8928
rect 6880 8916 6886 8968
rect 7283 8959 7341 8965
rect 7283 8925 7295 8959
rect 7329 8956 7341 8959
rect 7650 8956 7656 8968
rect 7329 8928 7656 8956
rect 7329 8925 7341 8928
rect 7283 8919 7341 8925
rect 7650 8916 7656 8928
rect 7708 8916 7714 8968
rect 8386 8916 8392 8968
rect 8444 8956 8450 8968
rect 8573 8959 8631 8965
rect 8573 8956 8585 8959
rect 8444 8928 8585 8956
rect 8444 8916 8450 8928
rect 8573 8925 8585 8928
rect 8619 8925 8631 8959
rect 8573 8919 8631 8925
rect 9307 8959 9365 8965
rect 9307 8925 9319 8959
rect 9353 8956 9365 8959
rect 9353 8928 10732 8956
rect 9353 8925 9365 8928
rect 9307 8919 9365 8925
rect 1486 8848 1492 8900
rect 1544 8848 1550 8900
rect 2682 8848 2688 8900
rect 2740 8888 2746 8900
rect 10318 8888 10324 8900
rect 2740 8860 10324 8888
rect 2740 8848 2746 8860
rect 10318 8848 10324 8860
rect 10376 8848 10382 8900
rect 474 8780 480 8832
rect 532 8780 538 8832
rect 3145 8823 3203 8829
rect 3145 8789 3157 8823
rect 3191 8820 3203 8823
rect 5902 8820 5908 8832
rect 3191 8792 5908 8820
rect 3191 8789 3203 8792
rect 3145 8783 3203 8789
rect 5902 8780 5908 8792
rect 5960 8780 5966 8832
rect 6638 8780 6644 8832
rect 6696 8780 6702 8832
rect 6914 8780 6920 8832
rect 6972 8820 6978 8832
rect 7098 8820 7104 8832
rect 6972 8792 7104 8820
rect 6972 8780 6978 8792
rect 7098 8780 7104 8792
rect 7156 8780 7162 8832
rect 8389 8823 8447 8829
rect 8389 8789 8401 8823
rect 8435 8820 8447 8823
rect 9214 8820 9220 8832
rect 8435 8792 9220 8820
rect 8435 8789 8447 8792
rect 8389 8783 8447 8789
rect 9214 8780 9220 8792
rect 9272 8780 9278 8832
rect 9674 8780 9680 8832
rect 9732 8820 9738 8832
rect 10410 8820 10416 8832
rect 9732 8792 10416 8820
rect 9732 8780 9738 8792
rect 10410 8780 10416 8792
rect 10468 8780 10474 8832
rect 10704 8820 10732 8928
rect 10778 8916 10784 8968
rect 10836 8956 10842 8968
rect 10836 8955 10870 8956
rect 10836 8949 10897 8955
rect 10836 8916 10851 8949
rect 10839 8915 10851 8916
rect 10885 8915 10897 8949
rect 10839 8909 10897 8915
rect 11330 8820 11336 8832
rect 10704 8792 11336 8820
rect 11330 8780 11336 8792
rect 11388 8780 11394 8832
rect 11532 8820 11560 9132
rect 11609 9129 11621 9163
rect 11655 9160 11667 9163
rect 12710 9160 12716 9172
rect 11655 9132 12716 9160
rect 11655 9129 11667 9132
rect 11609 9123 11667 9129
rect 12710 9120 12716 9132
rect 12768 9120 12774 9172
rect 12894 9120 12900 9172
rect 12952 9160 12958 9172
rect 12989 9163 13047 9169
rect 12989 9160 13001 9163
rect 12952 9132 13001 9160
rect 12952 9120 12958 9132
rect 12989 9129 13001 9132
rect 13035 9129 13047 9163
rect 12989 9123 13047 9129
rect 14108 9132 14780 9160
rect 11790 8984 11796 9036
rect 11848 9024 11854 9036
rect 14108 9033 14136 9132
rect 11977 9027 12035 9033
rect 11977 9024 11989 9027
rect 11848 8996 11989 9024
rect 11848 8984 11854 8996
rect 11977 8993 11989 8996
rect 12023 8993 12035 9027
rect 11977 8987 12035 8993
rect 14093 9027 14151 9033
rect 14093 8993 14105 9027
rect 14139 8993 14151 9027
rect 14752 9024 14780 9132
rect 15102 9120 15108 9172
rect 15160 9120 15166 9172
rect 15194 9120 15200 9172
rect 15252 9160 15258 9172
rect 16485 9163 16543 9169
rect 16485 9160 16497 9163
rect 15252 9132 16497 9160
rect 15252 9120 15258 9132
rect 16485 9129 16497 9132
rect 16531 9129 16543 9163
rect 17126 9160 17132 9172
rect 16485 9123 16543 9129
rect 16776 9132 17132 9160
rect 14826 9052 14832 9104
rect 14884 9092 14890 9104
rect 14884 9064 15516 9092
rect 14884 9052 14890 9064
rect 15488 9033 15516 9064
rect 15473 9027 15531 9033
rect 14752 8996 15424 9024
rect 14093 8987 14151 8993
rect 12250 8916 12256 8968
rect 12308 8956 12314 8968
rect 14335 8959 14393 8965
rect 14335 8956 14347 8959
rect 12308 8928 12351 8956
rect 12406 8928 14347 8956
rect 12308 8916 12314 8928
rect 12406 8900 12434 8928
rect 14335 8925 14347 8928
rect 14381 8925 14393 8959
rect 14335 8919 14393 8925
rect 12342 8848 12348 8900
rect 12400 8860 12434 8900
rect 12400 8848 12406 8860
rect 13078 8848 13084 8900
rect 13136 8888 13142 8900
rect 15102 8888 15108 8900
rect 13136 8860 15108 8888
rect 13136 8848 13142 8860
rect 15102 8848 15108 8860
rect 15160 8848 15166 8900
rect 15396 8888 15424 8996
rect 15473 8993 15485 9027
rect 15519 8993 15531 9027
rect 15473 8987 15531 8993
rect 15488 8956 15516 8987
rect 15747 8959 15805 8965
rect 15488 8928 15700 8956
rect 15562 8888 15568 8900
rect 15396 8860 15568 8888
rect 15562 8848 15568 8860
rect 15620 8848 15626 8900
rect 15672 8888 15700 8928
rect 15747 8925 15759 8959
rect 15793 8956 15805 8959
rect 15838 8956 15844 8968
rect 15793 8928 15844 8956
rect 15793 8925 15805 8928
rect 15747 8919 15805 8925
rect 15838 8916 15844 8928
rect 15896 8916 15902 8968
rect 16206 8888 16212 8900
rect 15672 8860 16212 8888
rect 16206 8848 16212 8860
rect 16264 8848 16270 8900
rect 12250 8820 12256 8832
rect 11532 8792 12256 8820
rect 12250 8780 12256 8792
rect 12308 8780 12314 8832
rect 13446 8780 13452 8832
rect 13504 8820 13510 8832
rect 16776 8820 16804 9132
rect 17126 9120 17132 9132
rect 17184 9120 17190 9172
rect 17218 9120 17224 9172
rect 17276 9160 17282 9172
rect 17954 9160 17960 9172
rect 17276 9132 17960 9160
rect 17276 9120 17282 9132
rect 17954 9120 17960 9132
rect 18012 9120 18018 9172
rect 18138 9120 18144 9172
rect 18196 9160 18202 9172
rect 18325 9163 18383 9169
rect 18325 9160 18337 9163
rect 18196 9132 18337 9160
rect 18196 9120 18202 9132
rect 18325 9129 18337 9132
rect 18371 9129 18383 9163
rect 19334 9160 19340 9172
rect 18325 9123 18383 9129
rect 18708 9132 19340 9160
rect 18708 9024 18736 9132
rect 19334 9120 19340 9132
rect 19392 9120 19398 9172
rect 19429 9163 19487 9169
rect 19429 9129 19441 9163
rect 19475 9160 19487 9163
rect 21266 9160 21272 9172
rect 19475 9132 21272 9160
rect 19475 9129 19487 9132
rect 19429 9123 19487 9129
rect 21266 9120 21272 9132
rect 21324 9120 21330 9172
rect 21358 9120 21364 9172
rect 21416 9120 21422 9172
rect 21450 9120 21456 9172
rect 21508 9120 21514 9172
rect 18785 9095 18843 9101
rect 18785 9061 18797 9095
rect 18831 9061 18843 9095
rect 18785 9055 18843 9061
rect 17880 8996 18736 9024
rect 16853 8959 16911 8965
rect 16853 8925 16865 8959
rect 16899 8956 16911 8959
rect 16899 8928 16988 8956
rect 17126 8935 17132 8968
rect 16899 8925 16911 8928
rect 16853 8919 16911 8925
rect 16960 8832 16988 8928
rect 17111 8929 17132 8935
rect 17111 8895 17123 8929
rect 17184 8916 17190 8968
rect 17218 8916 17224 8968
rect 17276 8956 17282 8968
rect 17880 8956 17908 8996
rect 17276 8928 17908 8956
rect 17276 8916 17282 8928
rect 17954 8916 17960 8968
rect 18012 8956 18018 8968
rect 18233 8959 18291 8965
rect 18233 8956 18245 8959
rect 18012 8928 18245 8956
rect 18012 8916 18018 8928
rect 18233 8925 18245 8928
rect 18279 8925 18291 8959
rect 18233 8919 18291 8925
rect 18509 8959 18567 8965
rect 18509 8925 18521 8959
rect 18555 8925 18567 8959
rect 18509 8919 18567 8925
rect 18693 8959 18751 8965
rect 18693 8925 18705 8959
rect 18739 8956 18751 8959
rect 18800 8956 18828 9055
rect 20990 9052 20996 9104
rect 21048 9052 21054 9104
rect 21376 9024 21404 9120
rect 21192 8996 21404 9024
rect 18739 8928 18828 8956
rect 18739 8925 18751 8928
rect 18693 8919 18751 8925
rect 17157 8898 17172 8916
rect 17157 8895 17169 8898
rect 17111 8889 17169 8895
rect 18524 8888 18552 8919
rect 18966 8916 18972 8968
rect 19024 8916 19030 8968
rect 19426 8956 19432 8968
rect 19352 8955 19432 8956
rect 19337 8949 19432 8955
rect 19337 8915 19349 8949
rect 19383 8928 19432 8949
rect 19383 8915 19395 8928
rect 19426 8916 19432 8928
rect 19484 8916 19490 8968
rect 19518 8916 19524 8968
rect 19576 8916 19582 8968
rect 21192 8965 21220 8996
rect 19613 8959 19671 8965
rect 19613 8925 19625 8959
rect 19659 8926 19671 8959
rect 19887 8959 19945 8965
rect 19659 8925 19748 8926
rect 19613 8919 19748 8925
rect 19887 8925 19899 8959
rect 19933 8956 19945 8959
rect 21177 8959 21235 8965
rect 19933 8928 20300 8956
rect 19933 8925 19945 8928
rect 19887 8919 19945 8925
rect 19337 8909 19395 8915
rect 19628 8898 19748 8919
rect 17880 8860 18552 8888
rect 19720 8888 19748 8898
rect 19978 8888 19984 8900
rect 19720 8860 19984 8888
rect 13504 8792 16804 8820
rect 13504 8780 13510 8792
rect 16942 8780 16948 8832
rect 17000 8780 17006 8832
rect 17126 8780 17132 8832
rect 17184 8820 17190 8832
rect 17880 8829 17908 8860
rect 19978 8848 19984 8860
rect 20036 8848 20042 8900
rect 20162 8848 20168 8900
rect 20220 8848 20226 8900
rect 17865 8823 17923 8829
rect 17865 8820 17877 8823
rect 17184 8792 17877 8820
rect 17184 8780 17190 8792
rect 17865 8789 17877 8792
rect 17911 8789 17923 8823
rect 17865 8783 17923 8789
rect 18598 8780 18604 8832
rect 18656 8780 18662 8832
rect 19426 8780 19432 8832
rect 19484 8820 19490 8832
rect 20180 8820 20208 8848
rect 20272 8832 20300 8928
rect 21177 8925 21189 8959
rect 21223 8925 21235 8959
rect 21177 8919 21235 8925
rect 21266 8916 21272 8968
rect 21324 8916 21330 8968
rect 19484 8792 20208 8820
rect 19484 8780 19490 8792
rect 20254 8780 20260 8832
rect 20312 8780 20318 8832
rect 20622 8780 20628 8832
rect 20680 8780 20686 8832
rect 1104 8730 22056 8752
rect 1104 8678 6148 8730
rect 6200 8678 6212 8730
rect 6264 8678 6276 8730
rect 6328 8678 6340 8730
rect 6392 8678 6404 8730
rect 6456 8678 11346 8730
rect 11398 8678 11410 8730
rect 11462 8678 11474 8730
rect 11526 8678 11538 8730
rect 11590 8678 11602 8730
rect 11654 8678 16544 8730
rect 16596 8678 16608 8730
rect 16660 8678 16672 8730
rect 16724 8678 16736 8730
rect 16788 8678 16800 8730
rect 16852 8678 21742 8730
rect 21794 8678 21806 8730
rect 21858 8678 21870 8730
rect 21922 8678 21934 8730
rect 21986 8678 21998 8730
rect 22050 8678 22056 8730
rect 1104 8656 22056 8678
rect 1765 8619 1823 8625
rect 1765 8585 1777 8619
rect 1811 8616 1823 8619
rect 2958 8616 2964 8628
rect 1811 8588 2964 8616
rect 1811 8585 1823 8588
rect 1765 8579 1823 8585
rect 2958 8576 2964 8588
rect 3016 8576 3022 8628
rect 3326 8576 3332 8628
rect 3384 8616 3390 8628
rect 4433 8619 4491 8625
rect 4433 8616 4445 8619
rect 3384 8588 4445 8616
rect 3384 8576 3390 8588
rect 4433 8585 4445 8588
rect 4479 8585 4491 8619
rect 4614 8616 4620 8628
rect 4433 8579 4491 8585
rect 4540 8588 4620 8616
rect 4246 8508 4252 8560
rect 4304 8548 4310 8560
rect 4540 8548 4568 8588
rect 4614 8576 4620 8588
rect 4672 8616 4678 8628
rect 7098 8616 7104 8628
rect 4672 8588 7104 8616
rect 4672 8576 4678 8588
rect 7098 8576 7104 8588
rect 7156 8576 7162 8628
rect 7282 8576 7288 8628
rect 7340 8616 7346 8628
rect 7469 8619 7527 8625
rect 7469 8616 7481 8619
rect 7340 8588 7481 8616
rect 7340 8576 7346 8588
rect 7469 8585 7481 8588
rect 7515 8585 7527 8619
rect 7469 8579 7527 8585
rect 8036 8588 8524 8616
rect 4304 8520 4568 8548
rect 4304 8508 4310 8520
rect 4890 8508 4896 8560
rect 4948 8508 4954 8560
rect 7558 8548 7564 8560
rect 6196 8520 7564 8548
rect 1486 8440 1492 8492
rect 1544 8440 1550 8492
rect 2406 8480 2412 8492
rect 2240 8452 2412 8480
rect 2240 8276 2268 8452
rect 2406 8440 2412 8452
rect 2464 8480 2470 8492
rect 2501 8483 2559 8489
rect 2501 8480 2513 8483
rect 2464 8452 2513 8480
rect 2464 8440 2470 8452
rect 2501 8449 2513 8452
rect 2547 8449 2559 8483
rect 2501 8443 2559 8449
rect 2682 8440 2688 8492
rect 2740 8440 2746 8492
rect 3418 8489 3424 8492
rect 3375 8483 3424 8489
rect 3375 8449 3387 8483
rect 3421 8449 3424 8483
rect 3375 8443 3424 8449
rect 3418 8440 3424 8443
rect 3476 8440 3482 8492
rect 3510 8440 3516 8492
rect 3568 8440 3574 8492
rect 4154 8440 4160 8492
rect 4212 8480 4218 8492
rect 4341 8483 4399 8489
rect 4341 8480 4353 8483
rect 4212 8452 4353 8480
rect 4212 8440 4218 8452
rect 4341 8449 4353 8452
rect 4387 8449 4399 8483
rect 4908 8480 4936 8508
rect 5043 8483 5101 8489
rect 5043 8480 5055 8483
rect 4908 8452 5055 8480
rect 4341 8443 4399 8449
rect 5043 8449 5055 8452
rect 5089 8449 5101 8483
rect 5043 8443 5101 8449
rect 5534 8440 5540 8492
rect 5592 8440 5598 8492
rect 2317 8415 2375 8421
rect 2317 8381 2329 8415
rect 2363 8412 2375 8415
rect 2700 8412 2728 8440
rect 2363 8384 2728 8412
rect 2363 8381 2375 8384
rect 2317 8375 2375 8381
rect 2866 8372 2872 8424
rect 2924 8412 2930 8424
rect 3237 8415 3295 8421
rect 3237 8412 3249 8415
rect 2924 8384 3249 8412
rect 2924 8372 2930 8384
rect 3237 8381 3249 8384
rect 3283 8381 3295 8415
rect 3237 8375 3295 8381
rect 3878 8372 3884 8424
rect 3936 8412 3942 8424
rect 4801 8415 4859 8421
rect 4801 8412 4813 8415
rect 3936 8384 4813 8412
rect 3936 8372 3942 8384
rect 4801 8381 4813 8384
rect 4847 8381 4859 8415
rect 4801 8375 4859 8381
rect 2958 8304 2964 8356
rect 3016 8304 3022 8356
rect 4246 8344 4252 8356
rect 3896 8316 4252 8344
rect 3896 8276 3924 8316
rect 4246 8304 4252 8316
rect 4304 8304 4310 8356
rect 5552 8344 5580 8440
rect 6196 8412 6224 8520
rect 7558 8508 7564 8520
rect 7616 8548 7622 8560
rect 8036 8548 8064 8588
rect 8496 8560 8524 8588
rect 8570 8576 8576 8628
rect 8628 8576 8634 8628
rect 9306 8576 9312 8628
rect 9364 8616 9370 8628
rect 9950 8616 9956 8628
rect 9364 8588 9956 8616
rect 9364 8576 9370 8588
rect 9950 8576 9956 8588
rect 10008 8576 10014 8628
rect 10318 8576 10324 8628
rect 10376 8616 10382 8628
rect 11241 8619 11299 8625
rect 10376 8588 11100 8616
rect 10376 8576 10382 8588
rect 7616 8520 8064 8548
rect 7616 8508 7622 8520
rect 6270 8440 6276 8492
rect 6328 8480 6334 8492
rect 8036 8489 8064 8520
rect 8478 8508 8484 8560
rect 8536 8508 8542 8560
rect 6699 8483 6757 8489
rect 6699 8480 6711 8483
rect 6328 8452 6711 8480
rect 6328 8440 6334 8452
rect 6699 8449 6711 8452
rect 6745 8449 6757 8483
rect 6699 8443 6757 8449
rect 8021 8483 8079 8489
rect 8021 8449 8033 8483
rect 8067 8449 8079 8483
rect 8021 8443 8079 8449
rect 8295 8483 8353 8489
rect 8295 8449 8307 8483
rect 8341 8480 8353 8483
rect 8588 8480 8616 8576
rect 11072 8548 11100 8588
rect 11241 8585 11253 8619
rect 11287 8616 11299 8619
rect 11698 8616 11704 8628
rect 11287 8588 11704 8616
rect 11287 8585 11299 8588
rect 11241 8579 11299 8585
rect 11698 8576 11704 8588
rect 11756 8576 11762 8628
rect 12434 8576 12440 8628
rect 12492 8616 12498 8628
rect 12529 8619 12587 8625
rect 12529 8616 12541 8619
rect 12492 8588 12541 8616
rect 12492 8576 12498 8588
rect 12529 8585 12541 8588
rect 12575 8585 12587 8619
rect 12529 8579 12587 8585
rect 13262 8576 13268 8628
rect 13320 8616 13326 8628
rect 13909 8619 13967 8625
rect 13909 8616 13921 8619
rect 13320 8588 13921 8616
rect 13320 8576 13326 8588
rect 13909 8585 13921 8588
rect 13955 8585 13967 8619
rect 13909 8579 13967 8585
rect 14016 8588 14688 8616
rect 14016 8548 14044 8588
rect 11072 8520 14044 8548
rect 14660 8548 14688 8588
rect 15286 8576 15292 8628
rect 15344 8576 15350 8628
rect 18325 8619 18383 8625
rect 16546 8588 17954 8616
rect 16546 8548 16574 8588
rect 17678 8548 17684 8560
rect 14660 8520 16574 8548
rect 17227 8520 17684 8548
rect 14519 8493 14577 8499
rect 14519 8492 14531 8493
rect 8341 8452 8616 8480
rect 9401 8483 9459 8489
rect 8341 8449 8353 8452
rect 8295 8443 8353 8449
rect 9401 8449 9413 8483
rect 9447 8480 9459 8483
rect 9490 8480 9496 8492
rect 9447 8452 9496 8480
rect 9447 8449 9459 8452
rect 9401 8443 9459 8449
rect 9490 8440 9496 8452
rect 9548 8440 9554 8492
rect 10318 8440 10324 8492
rect 10376 8440 10382 8492
rect 11517 8483 11575 8489
rect 11517 8449 11529 8483
rect 11563 8480 11575 8483
rect 11698 8480 11704 8492
rect 11563 8452 11704 8480
rect 11563 8449 11575 8452
rect 10474 8424 10548 8446
rect 11517 8443 11575 8449
rect 11698 8440 11704 8452
rect 11756 8440 11762 8492
rect 11791 8483 11849 8489
rect 11791 8449 11803 8483
rect 11837 8480 11849 8483
rect 11882 8480 11888 8492
rect 11837 8452 11888 8480
rect 11837 8449 11849 8452
rect 11791 8443 11849 8449
rect 11882 8440 11888 8452
rect 11940 8440 11946 8492
rect 12084 8440 12090 8492
rect 12142 8480 12148 8492
rect 13078 8480 13084 8492
rect 12142 8452 13084 8480
rect 12142 8440 12148 8452
rect 13078 8440 13084 8452
rect 13136 8440 13142 8492
rect 13171 8483 13229 8489
rect 13171 8449 13183 8483
rect 13217 8480 13229 8483
rect 13262 8480 13268 8492
rect 13217 8452 13268 8480
rect 13217 8449 13229 8452
rect 13171 8443 13229 8449
rect 13262 8440 13268 8452
rect 13320 8440 13326 8492
rect 14182 8440 14188 8492
rect 14240 8480 14246 8492
rect 14277 8483 14335 8489
rect 14277 8480 14289 8483
rect 14240 8452 14289 8480
rect 14240 8440 14246 8452
rect 14277 8449 14289 8452
rect 14323 8449 14335 8483
rect 14277 8443 14335 8449
rect 14458 8440 14464 8492
rect 14516 8459 14531 8492
rect 14565 8459 14577 8493
rect 17227 8489 17255 8520
rect 17678 8508 17684 8520
rect 17736 8508 17742 8560
rect 17926 8548 17954 8588
rect 18325 8585 18337 8619
rect 18371 8616 18383 8619
rect 18966 8616 18972 8628
rect 18371 8588 18972 8616
rect 18371 8585 18383 8588
rect 18325 8579 18383 8585
rect 18966 8576 18972 8588
rect 19024 8576 19030 8628
rect 19306 8588 20392 8616
rect 19306 8548 19334 8588
rect 20364 8560 20392 8588
rect 20622 8576 20628 8628
rect 20680 8576 20686 8628
rect 21174 8576 21180 8628
rect 21232 8616 21238 8628
rect 21361 8619 21419 8625
rect 21361 8616 21373 8619
rect 21232 8588 21373 8616
rect 21232 8576 21238 8588
rect 21361 8585 21373 8588
rect 21407 8585 21419 8619
rect 21361 8579 21419 8585
rect 19886 8548 19892 8560
rect 17926 8520 19334 8548
rect 19720 8520 19892 8548
rect 14516 8453 14577 8459
rect 16853 8483 16911 8489
rect 14516 8440 14522 8453
rect 16853 8449 16865 8483
rect 16899 8480 16911 8483
rect 16960 8480 17154 8484
rect 17212 8483 17270 8489
rect 17212 8480 17224 8483
rect 16899 8456 17224 8480
rect 16899 8452 16988 8456
rect 17126 8452 17224 8456
rect 16899 8449 16911 8452
rect 16853 8443 16911 8449
rect 17212 8449 17224 8452
rect 17258 8449 17270 8483
rect 17212 8443 17270 8449
rect 17954 8440 17960 8492
rect 18012 8480 18018 8492
rect 18843 8483 18901 8489
rect 18843 8480 18855 8483
rect 18012 8452 18855 8480
rect 18012 8440 18018 8452
rect 18843 8449 18855 8452
rect 18889 8480 18901 8483
rect 19720 8480 19748 8520
rect 19886 8508 19892 8520
rect 19944 8508 19950 8560
rect 20346 8508 20352 8560
rect 20404 8508 20410 8560
rect 18889 8452 19748 8480
rect 18889 8449 18901 8452
rect 18843 8443 18901 8449
rect 19794 8440 19800 8492
rect 19852 8480 19858 8492
rect 20223 8483 20281 8489
rect 20223 8480 20235 8483
rect 19852 8452 20235 8480
rect 19852 8440 19858 8452
rect 20223 8449 20235 8452
rect 20269 8449 20281 8483
rect 20640 8480 20668 8576
rect 21545 8483 21603 8489
rect 21545 8480 21557 8483
rect 20640 8452 21557 8480
rect 20223 8443 20281 8449
rect 21545 8449 21557 8452
rect 21591 8449 21603 8483
rect 21545 8443 21603 8449
rect 6457 8415 6515 8421
rect 6457 8412 6469 8415
rect 6196 8384 6469 8412
rect 6457 8381 6469 8384
rect 6503 8381 6515 8415
rect 6457 8375 6515 8381
rect 9585 8415 9643 8421
rect 9585 8381 9597 8415
rect 9631 8412 9643 8415
rect 9674 8412 9680 8424
rect 9631 8384 9680 8412
rect 9631 8381 9643 8384
rect 9585 8375 9643 8381
rect 9674 8372 9680 8384
rect 9732 8412 9738 8424
rect 10134 8412 10140 8424
rect 9732 8384 10140 8412
rect 9732 8372 9738 8384
rect 10134 8372 10140 8384
rect 10192 8372 10198 8424
rect 10474 8421 10508 8424
rect 10459 8415 10508 8421
rect 10459 8381 10471 8415
rect 10505 8381 10508 8415
rect 10459 8375 10508 8381
rect 10502 8372 10508 8375
rect 10560 8372 10566 8424
rect 10594 8372 10600 8424
rect 10652 8372 10658 8424
rect 12250 8372 12256 8424
rect 12308 8412 12314 8424
rect 12894 8412 12900 8424
rect 12308 8384 12900 8412
rect 12308 8372 12314 8384
rect 12894 8372 12900 8384
rect 12952 8372 12958 8424
rect 15378 8372 15384 8424
rect 15436 8412 15442 8424
rect 16298 8412 16304 8424
rect 15436 8384 16304 8412
rect 15436 8372 15442 8384
rect 16298 8372 16304 8384
rect 16356 8372 16362 8424
rect 16758 8372 16764 8424
rect 16816 8412 16822 8424
rect 16945 8415 17003 8421
rect 16945 8412 16957 8415
rect 16816 8384 16957 8412
rect 16816 8372 16822 8384
rect 16945 8381 16957 8384
rect 16991 8381 17003 8415
rect 16945 8375 17003 8381
rect 18322 8372 18328 8424
rect 18380 8412 18386 8424
rect 18506 8412 18512 8424
rect 18380 8384 18512 8412
rect 18380 8372 18386 8384
rect 18506 8372 18512 8384
rect 18564 8412 18570 8424
rect 18601 8415 18659 8421
rect 18601 8412 18613 8415
rect 18564 8384 18613 8412
rect 18564 8372 18570 8384
rect 18601 8381 18613 8384
rect 18647 8381 18659 8415
rect 18601 8375 18659 8381
rect 19978 8372 19984 8424
rect 20036 8372 20042 8424
rect 5813 8347 5871 8353
rect 5813 8344 5825 8347
rect 5552 8316 5825 8344
rect 5813 8313 5825 8316
rect 5859 8313 5871 8347
rect 5813 8307 5871 8313
rect 9033 8347 9091 8353
rect 9033 8313 9045 8347
rect 9079 8344 9091 8347
rect 10045 8347 10103 8353
rect 10045 8344 10057 8347
rect 9079 8316 10057 8344
rect 9079 8313 9091 8316
rect 9033 8307 9091 8313
rect 10045 8313 10057 8316
rect 10091 8313 10103 8347
rect 10045 8307 10103 8313
rect 16558 8316 16988 8344
rect 2240 8248 3924 8276
rect 4157 8279 4215 8285
rect 4157 8245 4169 8279
rect 4203 8276 4215 8279
rect 4614 8276 4620 8288
rect 4203 8248 4620 8276
rect 4203 8245 4215 8248
rect 4157 8239 4215 8245
rect 4614 8236 4620 8248
rect 4672 8236 4678 8288
rect 5258 8236 5264 8288
rect 5316 8276 5322 8288
rect 6730 8276 6736 8288
rect 5316 8248 6736 8276
rect 5316 8236 5322 8248
rect 6730 8236 6736 8248
rect 6788 8236 6794 8288
rect 6914 8236 6920 8288
rect 6972 8276 6978 8288
rect 7834 8276 7840 8288
rect 6972 8248 7840 8276
rect 6972 8236 6978 8248
rect 7834 8236 7840 8248
rect 7892 8236 7898 8288
rect 8018 8236 8024 8288
rect 8076 8276 8082 8288
rect 8938 8276 8944 8288
rect 8076 8248 8944 8276
rect 8076 8236 8082 8248
rect 8938 8236 8944 8248
rect 8996 8236 9002 8288
rect 9306 8236 9312 8288
rect 9364 8276 9370 8288
rect 9490 8276 9496 8288
rect 9364 8248 9496 8276
rect 9364 8236 9370 8248
rect 9490 8236 9496 8248
rect 9548 8276 9554 8288
rect 11146 8276 11152 8288
rect 9548 8248 11152 8276
rect 9548 8236 9554 8248
rect 11146 8236 11152 8248
rect 11204 8276 11210 8288
rect 11606 8276 11612 8288
rect 11204 8248 11612 8276
rect 11204 8236 11210 8248
rect 11606 8236 11612 8248
rect 11664 8236 11670 8288
rect 11790 8236 11796 8288
rect 11848 8276 11854 8288
rect 14274 8276 14280 8288
rect 11848 8248 14280 8276
rect 11848 8236 11854 8248
rect 14274 8236 14280 8248
rect 14332 8236 14338 8288
rect 14366 8236 14372 8288
rect 14424 8276 14430 8288
rect 15470 8276 15476 8288
rect 14424 8248 15476 8276
rect 14424 8236 14430 8248
rect 15470 8236 15476 8248
rect 15528 8236 15534 8288
rect 16298 8236 16304 8288
rect 16356 8276 16362 8288
rect 16558 8276 16586 8316
rect 16960 8288 16988 8316
rect 16356 8248 16586 8276
rect 16356 8236 16362 8248
rect 16666 8236 16672 8288
rect 16724 8236 16730 8288
rect 16942 8236 16948 8288
rect 17000 8276 17006 8288
rect 18340 8276 18368 8372
rect 19610 8304 19616 8356
rect 19668 8304 19674 8356
rect 17000 8248 18368 8276
rect 19996 8276 20024 8372
rect 20993 8347 21051 8353
rect 20993 8313 21005 8347
rect 21039 8344 21051 8347
rect 21174 8344 21180 8356
rect 21039 8316 21180 8344
rect 21039 8313 21051 8316
rect 20993 8307 21051 8313
rect 21174 8304 21180 8316
rect 21232 8304 21238 8356
rect 20346 8276 20352 8288
rect 19996 8248 20352 8276
rect 17000 8236 17006 8248
rect 20346 8236 20352 8248
rect 20404 8236 20410 8288
rect 1104 8186 21896 8208
rect 1104 8134 3549 8186
rect 3601 8134 3613 8186
rect 3665 8134 3677 8186
rect 3729 8134 3741 8186
rect 3793 8134 3805 8186
rect 3857 8134 8747 8186
rect 8799 8134 8811 8186
rect 8863 8134 8875 8186
rect 8927 8134 8939 8186
rect 8991 8134 9003 8186
rect 9055 8134 13945 8186
rect 13997 8134 14009 8186
rect 14061 8134 14073 8186
rect 14125 8134 14137 8186
rect 14189 8134 14201 8186
rect 14253 8134 19143 8186
rect 19195 8134 19207 8186
rect 19259 8134 19271 8186
rect 19323 8134 19335 8186
rect 19387 8134 19399 8186
rect 19451 8134 21896 8186
rect 1104 8112 21896 8134
rect 2332 8044 3004 8072
rect 2332 7945 2360 8044
rect 2976 8004 3004 8044
rect 3234 8032 3240 8084
rect 3292 8072 3298 8084
rect 3329 8075 3387 8081
rect 3329 8072 3341 8075
rect 3292 8044 3341 8072
rect 3292 8032 3298 8044
rect 3329 8041 3341 8044
rect 3375 8041 3387 8075
rect 3329 8035 3387 8041
rect 3881 8075 3939 8081
rect 3881 8041 3893 8075
rect 3927 8072 3939 8075
rect 4154 8072 4160 8084
rect 3927 8044 4160 8072
rect 3927 8041 3939 8044
rect 3881 8035 3939 8041
rect 4154 8032 4160 8044
rect 4212 8032 4218 8084
rect 4614 8032 4620 8084
rect 4672 8072 4678 8084
rect 4672 8044 4936 8072
rect 4672 8032 4678 8044
rect 4062 8004 4068 8016
rect 2976 7976 4068 8004
rect 4062 7964 4068 7976
rect 4120 7964 4126 8016
rect 4908 8004 4936 8044
rect 4982 8032 4988 8084
rect 5040 8072 5046 8084
rect 5169 8075 5227 8081
rect 5169 8072 5181 8075
rect 5040 8044 5181 8072
rect 5040 8032 5046 8044
rect 5169 8041 5181 8044
rect 5215 8041 5227 8075
rect 5169 8035 5227 8041
rect 5626 8032 5632 8084
rect 5684 8072 5690 8084
rect 6362 8072 6368 8084
rect 5684 8044 6368 8072
rect 5684 8032 5690 8044
rect 6362 8032 6368 8044
rect 6420 8072 6426 8084
rect 6914 8072 6920 8084
rect 6420 8044 6920 8072
rect 6420 8032 6426 8044
rect 6914 8032 6920 8044
rect 6972 8032 6978 8084
rect 7282 8032 7288 8084
rect 7340 8072 7346 8084
rect 7742 8072 7748 8084
rect 7340 8044 7748 8072
rect 7340 8032 7346 8044
rect 7742 8032 7748 8044
rect 7800 8032 7806 8084
rect 8570 8032 8576 8084
rect 8628 8032 8634 8084
rect 8846 8032 8852 8084
rect 8904 8072 8910 8084
rect 8904 8044 10548 8072
rect 8904 8032 8910 8044
rect 4908 7976 6592 8004
rect 2317 7939 2375 7945
rect 2317 7905 2329 7939
rect 2363 7905 2375 7939
rect 4080 7936 4108 7964
rect 4157 7939 4215 7945
rect 4157 7936 4169 7939
rect 4080 7908 4169 7936
rect 2317 7899 2375 7905
rect 4157 7905 4169 7908
rect 4203 7905 4215 7939
rect 4157 7899 4215 7905
rect 5810 7896 5816 7948
rect 5868 7936 5874 7948
rect 6181 7939 6239 7945
rect 6181 7936 6193 7939
rect 5868 7908 6193 7936
rect 5868 7896 5874 7908
rect 6181 7905 6193 7908
rect 6227 7905 6239 7939
rect 6564 7936 6592 7976
rect 6638 7964 6644 8016
rect 6696 8004 6702 8016
rect 6825 8007 6883 8013
rect 6825 8004 6837 8007
rect 6696 7976 6837 8004
rect 6696 7964 6702 7976
rect 6825 7973 6837 7976
rect 6871 7973 6883 8007
rect 6825 7967 6883 7973
rect 7834 7964 7840 8016
rect 7892 8004 7898 8016
rect 8110 8004 8116 8016
rect 7892 7976 8116 8004
rect 7892 7964 7898 7976
rect 8110 7964 8116 7976
rect 8168 7964 8174 8016
rect 8386 7964 8392 8016
rect 8444 7964 8450 8016
rect 8588 8004 8616 8032
rect 10520 8004 10548 8044
rect 10594 8032 10600 8084
rect 10652 8032 10658 8084
rect 15286 8072 15292 8084
rect 11072 8044 15292 8072
rect 11072 8004 11100 8044
rect 15286 8032 15292 8044
rect 15344 8032 15350 8084
rect 17954 8072 17960 8084
rect 16224 8044 17960 8072
rect 11698 8004 11704 8016
rect 8588 7976 9628 8004
rect 10520 7976 11100 8004
rect 11164 7976 11704 8004
rect 9600 7945 9628 7976
rect 11164 7945 11192 7976
rect 11698 7964 11704 7976
rect 11756 7964 11762 8016
rect 11790 7964 11796 8016
rect 11848 7964 11854 8016
rect 12894 7964 12900 8016
rect 12952 8004 12958 8016
rect 13538 8004 13544 8016
rect 12952 7976 13544 8004
rect 12952 7964 12958 7976
rect 13538 7964 13544 7976
rect 13596 7964 13602 8016
rect 15102 7964 15108 8016
rect 15160 8004 15166 8016
rect 15841 8007 15899 8013
rect 15841 8004 15853 8007
rect 15160 7976 15853 8004
rect 15160 7964 15166 7976
rect 15841 7973 15853 7976
rect 15887 7973 15899 8007
rect 15841 7967 15899 7973
rect 9585 7939 9643 7945
rect 6564 7908 9168 7936
rect 6181 7899 6239 7905
rect 2498 7828 2504 7880
rect 2556 7828 2562 7880
rect 2591 7871 2649 7877
rect 2591 7837 2603 7871
rect 2637 7868 2649 7871
rect 2682 7868 2688 7880
rect 2637 7840 2688 7868
rect 2637 7837 2649 7840
rect 2591 7831 2649 7837
rect 2682 7828 2688 7840
rect 2740 7868 2746 7880
rect 3786 7868 3792 7880
rect 2740 7840 3792 7868
rect 2740 7828 2746 7840
rect 3786 7828 3792 7840
rect 3844 7828 3850 7880
rect 4062 7828 4068 7880
rect 4120 7828 4126 7880
rect 4399 7871 4457 7877
rect 4399 7868 4411 7871
rect 4264 7840 4411 7868
rect 1489 7803 1547 7809
rect 1489 7769 1501 7803
rect 1535 7800 1547 7803
rect 2133 7803 2191 7809
rect 2133 7800 2145 7803
rect 1535 7772 2145 7800
rect 1535 7769 1547 7772
rect 1489 7763 1547 7769
rect 2133 7769 2145 7772
rect 2179 7769 2191 7803
rect 2516 7800 2544 7828
rect 4264 7800 4292 7840
rect 4399 7837 4411 7840
rect 4445 7868 4457 7871
rect 4522 7868 4528 7880
rect 4445 7840 4528 7868
rect 4445 7837 4457 7840
rect 4399 7831 4457 7837
rect 4522 7828 4528 7840
rect 4580 7828 4586 7880
rect 6362 7828 6368 7880
rect 6420 7828 6426 7880
rect 7098 7828 7104 7880
rect 7156 7828 7162 7880
rect 7280 7877 7286 7880
rect 7239 7871 7286 7877
rect 7239 7837 7251 7871
rect 7285 7837 7286 7871
rect 7239 7831 7286 7837
rect 7280 7828 7286 7831
rect 7338 7828 7344 7880
rect 7374 7828 7380 7880
rect 7432 7828 7438 7880
rect 8202 7828 8208 7880
rect 8260 7828 8266 7880
rect 8294 7828 8300 7880
rect 8352 7828 8358 7880
rect 8386 7828 8392 7880
rect 8444 7868 8450 7880
rect 9140 7877 9168 7908
rect 9585 7905 9597 7939
rect 9631 7905 9643 7939
rect 9585 7899 9643 7905
rect 11149 7939 11207 7945
rect 11149 7905 11161 7939
rect 11195 7905 11207 7939
rect 11149 7899 11207 7905
rect 12066 7896 12072 7948
rect 12124 7896 12130 7948
rect 12342 7896 12348 7948
rect 12400 7896 12406 7948
rect 16224 7936 16252 8044
rect 17954 8032 17960 8044
rect 18012 8032 18018 8084
rect 18506 8032 18512 8084
rect 18564 8072 18570 8084
rect 18564 8044 20392 8072
rect 18564 8032 18570 8044
rect 17678 7964 17684 8016
rect 17736 8004 17742 8016
rect 17862 8004 17868 8016
rect 17736 7976 17868 8004
rect 17736 7964 17742 7976
rect 17862 7964 17868 7976
rect 17920 7964 17926 8016
rect 18046 7964 18052 8016
rect 18104 8004 18110 8016
rect 18785 8007 18843 8013
rect 18785 8004 18797 8007
rect 18104 7976 18797 8004
rect 18104 7964 18110 7976
rect 18785 7973 18797 7976
rect 18831 7973 18843 8007
rect 20364 8004 20392 8044
rect 21082 8032 21088 8084
rect 21140 8072 21146 8084
rect 21453 8075 21511 8081
rect 21453 8072 21465 8075
rect 21140 8044 21465 8072
rect 21140 8032 21146 8044
rect 21453 8041 21465 8044
rect 21499 8041 21511 8075
rect 21453 8035 21511 8041
rect 22094 8004 22100 8016
rect 20364 7976 22100 8004
rect 18785 7967 18843 7973
rect 22094 7964 22100 7976
rect 22152 7964 22158 8016
rect 15856 7908 16252 7936
rect 8573 7871 8631 7877
rect 8444 7858 8524 7868
rect 8573 7858 8585 7871
rect 8444 7840 8585 7858
rect 8444 7828 8450 7840
rect 8496 7837 8585 7840
rect 8619 7837 8631 7871
rect 8496 7831 8631 7837
rect 9125 7871 9183 7877
rect 9125 7837 9137 7871
rect 9171 7837 9183 7871
rect 9125 7831 9183 7837
rect 9859 7871 9917 7877
rect 9859 7837 9871 7871
rect 9905 7868 9917 7871
rect 11333 7871 11391 7877
rect 9905 7840 11192 7868
rect 9905 7837 9917 7840
rect 9859 7831 9917 7837
rect 8496 7830 8616 7831
rect 5534 7800 5540 7812
rect 2516 7772 4292 7800
rect 4632 7772 5540 7800
rect 2133 7763 2191 7769
rect 1765 7735 1823 7741
rect 1765 7701 1777 7735
rect 1811 7732 1823 7735
rect 2038 7732 2044 7744
rect 1811 7704 2044 7732
rect 1811 7701 1823 7704
rect 1765 7695 1823 7701
rect 2038 7692 2044 7704
rect 2096 7692 2102 7744
rect 2148 7732 2176 7763
rect 2866 7732 2872 7744
rect 2148 7704 2872 7732
rect 2866 7692 2872 7704
rect 2924 7692 2930 7744
rect 3878 7692 3884 7744
rect 3936 7732 3942 7744
rect 4632 7732 4660 7772
rect 5534 7760 5540 7772
rect 5592 7760 5598 7812
rect 5721 7803 5779 7809
rect 5721 7769 5733 7803
rect 5767 7800 5779 7803
rect 8220 7800 8248 7828
rect 5767 7772 6408 7800
rect 5767 7769 5779 7772
rect 5721 7763 5779 7769
rect 3936 7704 4660 7732
rect 3936 7692 3942 7704
rect 4706 7692 4712 7744
rect 4764 7732 4770 7744
rect 5813 7735 5871 7741
rect 5813 7732 5825 7735
rect 4764 7704 5825 7732
rect 4764 7692 4770 7704
rect 5813 7701 5825 7704
rect 5859 7701 5871 7735
rect 6380 7732 6408 7772
rect 7852 7772 8248 7800
rect 7852 7732 7880 7772
rect 8754 7760 8760 7812
rect 8812 7800 8818 7812
rect 10778 7800 10784 7812
rect 8812 7772 10784 7800
rect 8812 7760 8818 7772
rect 10778 7760 10784 7772
rect 10836 7760 10842 7812
rect 11164 7800 11192 7840
rect 11333 7837 11345 7871
rect 11379 7837 11391 7871
rect 11333 7831 11391 7837
rect 11238 7800 11244 7812
rect 11164 7772 11244 7800
rect 11238 7760 11244 7772
rect 11296 7760 11302 7812
rect 6380 7704 7880 7732
rect 5813 7695 5871 7701
rect 8018 7692 8024 7744
rect 8076 7692 8082 7744
rect 8110 7692 8116 7744
rect 8168 7692 8174 7744
rect 8386 7692 8392 7744
rect 8444 7732 8450 7744
rect 8941 7735 8999 7741
rect 8941 7732 8953 7735
rect 8444 7704 8953 7732
rect 8444 7692 8450 7704
rect 8941 7701 8953 7704
rect 8987 7701 8999 7735
rect 8941 7695 8999 7701
rect 10042 7692 10048 7744
rect 10100 7732 10106 7744
rect 10962 7732 10968 7744
rect 10100 7704 10968 7732
rect 10100 7692 10106 7704
rect 10962 7692 10968 7704
rect 11020 7692 11026 7744
rect 11348 7732 11376 7831
rect 12158 7828 12164 7880
rect 12216 7877 12222 7880
rect 12216 7871 12244 7877
rect 12232 7837 12244 7871
rect 12216 7831 12244 7837
rect 12216 7828 12222 7831
rect 13722 7828 13728 7880
rect 13780 7828 13786 7880
rect 13998 7828 14004 7880
rect 14056 7828 14062 7880
rect 14090 7828 14096 7880
rect 14148 7828 14154 7880
rect 15856 7877 15884 7908
rect 16298 7896 16304 7948
rect 16356 7896 16362 7948
rect 19426 7936 19432 7948
rect 17788 7908 19432 7936
rect 17788 7880 17816 7908
rect 19426 7896 19432 7908
rect 19484 7896 19490 7948
rect 14335 7871 14393 7877
rect 14335 7837 14347 7871
rect 14381 7837 14393 7871
rect 14335 7831 14393 7837
rect 15657 7871 15715 7877
rect 15657 7837 15669 7871
rect 15703 7837 15715 7871
rect 15657 7831 15715 7837
rect 15841 7871 15899 7877
rect 15841 7837 15853 7871
rect 15887 7837 15899 7871
rect 16543 7871 16601 7877
rect 15841 7831 15899 7837
rect 15948 7868 16160 7870
rect 16543 7868 16555 7871
rect 15948 7842 16555 7868
rect 14016 7800 14044 7828
rect 14350 7800 14378 7831
rect 14016 7772 14378 7800
rect 11974 7732 11980 7744
rect 11348 7704 11980 7732
rect 11974 7692 11980 7704
rect 12032 7732 12038 7744
rect 12894 7732 12900 7744
rect 12032 7704 12900 7732
rect 12032 7692 12038 7704
rect 12894 7692 12900 7704
rect 12952 7692 12958 7744
rect 12986 7692 12992 7744
rect 13044 7692 13050 7744
rect 13814 7692 13820 7744
rect 13872 7732 13878 7744
rect 13909 7735 13967 7741
rect 13909 7732 13921 7735
rect 13872 7704 13921 7732
rect 13872 7692 13878 7704
rect 13909 7701 13921 7704
rect 13955 7701 13967 7735
rect 13909 7695 13967 7701
rect 15010 7692 15016 7744
rect 15068 7732 15074 7744
rect 15105 7735 15163 7741
rect 15105 7732 15117 7735
rect 15068 7704 15117 7732
rect 15068 7692 15074 7704
rect 15105 7701 15117 7704
rect 15151 7701 15163 7735
rect 15672 7732 15700 7831
rect 15948 7812 15976 7842
rect 16132 7840 16555 7842
rect 16543 7837 16555 7840
rect 16589 7837 16601 7871
rect 16543 7831 16601 7837
rect 16666 7828 16672 7880
rect 16724 7868 16730 7880
rect 17681 7871 17739 7877
rect 17681 7868 17693 7871
rect 16724 7840 17693 7868
rect 16724 7828 16730 7840
rect 17681 7837 17693 7840
rect 17727 7837 17739 7871
rect 17681 7831 17739 7837
rect 17770 7828 17776 7880
rect 17828 7828 17834 7880
rect 18141 7871 18199 7877
rect 18141 7837 18153 7871
rect 18187 7837 18199 7871
rect 18141 7831 18199 7837
rect 15930 7760 15936 7812
rect 15988 7760 15994 7812
rect 16206 7760 16212 7812
rect 16264 7760 16270 7812
rect 16942 7760 16948 7812
rect 17000 7800 17006 7812
rect 17788 7800 17816 7828
rect 17000 7772 17816 7800
rect 17000 7760 17006 7772
rect 16022 7732 16028 7744
rect 15672 7704 16028 7732
rect 15105 7695 15163 7701
rect 16022 7692 16028 7704
rect 16080 7692 16086 7744
rect 17218 7692 17224 7744
rect 17276 7732 17282 7744
rect 17313 7735 17371 7741
rect 17313 7732 17325 7735
rect 17276 7704 17325 7732
rect 17276 7692 17282 7704
rect 17313 7701 17325 7704
rect 17359 7701 17371 7735
rect 17313 7695 17371 7701
rect 17494 7692 17500 7744
rect 17552 7732 17558 7744
rect 17773 7735 17831 7741
rect 17773 7732 17785 7735
rect 17552 7704 17785 7732
rect 17552 7692 17558 7704
rect 17773 7701 17785 7704
rect 17819 7701 17831 7735
rect 18156 7732 18184 7831
rect 18506 7828 18512 7880
rect 18564 7828 18570 7880
rect 18877 7871 18935 7877
rect 18877 7837 18889 7871
rect 18923 7868 18935 7871
rect 20714 7868 20720 7880
rect 18923 7840 20720 7868
rect 18923 7837 18935 7840
rect 18877 7831 18935 7837
rect 20714 7828 20720 7840
rect 20772 7828 20778 7880
rect 21085 7871 21143 7877
rect 21085 7868 21097 7871
rect 20824 7840 21097 7868
rect 19334 7760 19340 7812
rect 19392 7800 19398 7812
rect 19674 7803 19732 7809
rect 19674 7800 19686 7803
rect 19392 7772 19686 7800
rect 19392 7760 19398 7772
rect 19674 7769 19686 7772
rect 19720 7800 19732 7803
rect 20824 7800 20852 7840
rect 21085 7837 21097 7840
rect 21131 7837 21143 7871
rect 21085 7831 21143 7837
rect 21361 7871 21419 7877
rect 21361 7837 21373 7871
rect 21407 7837 21419 7871
rect 21361 7831 21419 7837
rect 21376 7800 21404 7831
rect 19720 7772 20852 7800
rect 20916 7772 21404 7800
rect 19720 7769 19732 7772
rect 19674 7763 19732 7769
rect 19978 7732 19984 7744
rect 18156 7704 19984 7732
rect 17773 7695 17831 7701
rect 19978 7692 19984 7704
rect 20036 7692 20042 7744
rect 20806 7692 20812 7744
rect 20864 7692 20870 7744
rect 20916 7741 20944 7772
rect 20901 7735 20959 7741
rect 20901 7701 20913 7735
rect 20947 7701 20959 7735
rect 20901 7695 20959 7701
rect 1104 7642 22056 7664
rect 1104 7590 6148 7642
rect 6200 7590 6212 7642
rect 6264 7590 6276 7642
rect 6328 7590 6340 7642
rect 6392 7590 6404 7642
rect 6456 7590 11346 7642
rect 11398 7590 11410 7642
rect 11462 7590 11474 7642
rect 11526 7590 11538 7642
rect 11590 7590 11602 7642
rect 11654 7590 16544 7642
rect 16596 7590 16608 7642
rect 16660 7590 16672 7642
rect 16724 7590 16736 7642
rect 16788 7590 16800 7642
rect 16852 7590 21742 7642
rect 21794 7590 21806 7642
rect 21858 7590 21870 7642
rect 21922 7590 21934 7642
rect 21986 7590 21998 7642
rect 22050 7590 22056 7642
rect 1104 7568 22056 7590
rect 1854 7488 1860 7540
rect 1912 7488 1918 7540
rect 3881 7531 3939 7537
rect 3881 7497 3893 7531
rect 3927 7528 3939 7531
rect 4062 7528 4068 7540
rect 3927 7500 4068 7528
rect 3927 7497 3939 7500
rect 3881 7491 3939 7497
rect 4062 7488 4068 7500
rect 4120 7488 4126 7540
rect 4154 7488 4160 7540
rect 4212 7488 4218 7540
rect 4430 7488 4436 7540
rect 4488 7488 4494 7540
rect 5534 7488 5540 7540
rect 5592 7488 5598 7540
rect 5813 7531 5871 7537
rect 5813 7497 5825 7531
rect 5859 7528 5871 7531
rect 7374 7528 7380 7540
rect 5859 7500 7380 7528
rect 5859 7497 5871 7500
rect 5813 7491 5871 7497
rect 7374 7488 7380 7500
rect 7432 7488 7438 7540
rect 8294 7488 8300 7540
rect 8352 7528 8358 7540
rect 9401 7531 9459 7537
rect 9401 7528 9413 7531
rect 8352 7500 9413 7528
rect 8352 7488 8358 7500
rect 9401 7497 9413 7500
rect 9447 7497 9459 7531
rect 10502 7528 10508 7540
rect 9401 7491 9459 7497
rect 9692 7500 10508 7528
rect 1302 7420 1308 7472
rect 1360 7460 1366 7472
rect 1581 7463 1639 7469
rect 1581 7460 1593 7463
rect 1360 7432 1593 7460
rect 1360 7420 1366 7432
rect 1581 7429 1593 7432
rect 1627 7429 1639 7463
rect 4172 7460 4200 7488
rect 1581 7423 1639 7429
rect 4080 7432 4200 7460
rect 1486 7352 1492 7404
rect 1544 7392 1550 7404
rect 2041 7395 2099 7401
rect 2041 7392 2053 7395
rect 1544 7364 2053 7392
rect 1544 7352 1550 7364
rect 2041 7361 2053 7364
rect 2087 7361 2099 7395
rect 2041 7355 2099 7361
rect 3234 7352 3240 7404
rect 3292 7352 3298 7404
rect 3970 7352 3976 7404
rect 4028 7392 4034 7404
rect 4080 7392 4108 7432
rect 5350 7420 5356 7472
rect 5408 7460 5414 7472
rect 5552 7460 5580 7488
rect 7009 7463 7067 7469
rect 7009 7460 7021 7463
rect 5408 7420 5442 7460
rect 5552 7432 7021 7460
rect 7009 7429 7021 7432
rect 7055 7429 7067 7463
rect 7009 7423 7067 7429
rect 4028 7364 4108 7392
rect 4028 7352 4034 7364
rect 1302 7148 1308 7200
rect 1360 7188 1366 7200
rect 1504 7188 1532 7352
rect 1578 7284 1584 7336
rect 1636 7324 1642 7336
rect 2222 7324 2228 7336
rect 1636 7296 2228 7324
rect 1636 7284 1642 7296
rect 2222 7284 2228 7296
rect 2280 7284 2286 7336
rect 2961 7327 3019 7333
rect 2961 7324 2973 7327
rect 2792 7296 2973 7324
rect 2590 7216 2596 7268
rect 2648 7256 2654 7268
rect 2685 7259 2743 7265
rect 2685 7256 2697 7259
rect 2648 7228 2697 7256
rect 2648 7216 2654 7228
rect 2685 7225 2697 7228
rect 2731 7225 2743 7259
rect 2685 7219 2743 7225
rect 1360 7160 1532 7188
rect 1360 7148 1366 7160
rect 2314 7148 2320 7200
rect 2372 7188 2378 7200
rect 2792 7188 2820 7296
rect 2961 7293 2973 7296
rect 3007 7293 3019 7327
rect 2961 7287 3019 7293
rect 3099 7327 3157 7333
rect 3099 7293 3111 7327
rect 3145 7324 3157 7327
rect 4080 7324 4108 7364
rect 4157 7395 4215 7401
rect 4157 7361 4169 7395
rect 4203 7361 4215 7395
rect 4157 7355 4215 7361
rect 4341 7395 4399 7401
rect 4341 7361 4353 7395
rect 4387 7392 4399 7395
rect 4706 7392 4712 7404
rect 4387 7364 4712 7392
rect 4387 7361 4399 7364
rect 4341 7355 4399 7361
rect 3145 7296 4108 7324
rect 3145 7293 3157 7296
rect 3099 7287 3157 7293
rect 3878 7216 3884 7268
rect 3936 7256 3942 7268
rect 3973 7259 4031 7265
rect 3973 7256 3985 7259
rect 3936 7228 3985 7256
rect 3936 7216 3942 7228
rect 3973 7225 3985 7228
rect 4019 7225 4031 7259
rect 4172 7256 4200 7355
rect 4706 7352 4712 7364
rect 4764 7352 4770 7404
rect 4982 7352 4988 7404
rect 5040 7392 5046 7404
rect 5075 7395 5133 7401
rect 5075 7392 5087 7395
rect 5040 7364 5087 7392
rect 5040 7352 5046 7364
rect 5075 7361 5087 7364
rect 5121 7361 5133 7395
rect 5075 7355 5133 7361
rect 4522 7284 4528 7336
rect 4580 7324 4586 7336
rect 4801 7327 4859 7333
rect 4801 7324 4813 7327
rect 4580 7296 4813 7324
rect 4580 7284 4586 7296
rect 4801 7293 4813 7296
rect 4847 7293 4859 7327
rect 5414 7324 5442 7420
rect 5534 7352 5540 7404
rect 5592 7392 5598 7404
rect 6457 7395 6515 7401
rect 6457 7392 6469 7395
rect 5592 7364 6469 7392
rect 5592 7352 5598 7364
rect 6457 7361 6469 7364
rect 6503 7361 6515 7395
rect 6457 7355 6515 7361
rect 8754 7352 8760 7404
rect 8812 7352 8818 7404
rect 9692 7392 9720 7500
rect 10502 7488 10508 7500
rect 10560 7488 10566 7540
rect 11698 7488 11704 7540
rect 11756 7528 11762 7540
rect 11756 7500 11928 7528
rect 11756 7488 11762 7500
rect 11238 7420 11244 7472
rect 11296 7460 11302 7472
rect 11900 7460 11928 7500
rect 12342 7488 12348 7540
rect 12400 7528 12406 7540
rect 12529 7531 12587 7537
rect 12529 7528 12541 7531
rect 12400 7500 12541 7528
rect 12400 7488 12406 7500
rect 12529 7497 12541 7500
rect 12575 7497 12587 7531
rect 12529 7491 12587 7497
rect 12894 7488 12900 7540
rect 12952 7528 12958 7540
rect 15746 7528 15752 7540
rect 12952 7500 15752 7528
rect 12952 7488 12958 7500
rect 15746 7488 15752 7500
rect 15804 7488 15810 7540
rect 16022 7488 16028 7540
rect 16080 7488 16086 7540
rect 16114 7488 16120 7540
rect 16172 7488 16178 7540
rect 17218 7488 17224 7540
rect 17276 7488 17282 7540
rect 17494 7488 17500 7540
rect 17552 7488 17558 7540
rect 17954 7488 17960 7540
rect 18012 7488 18018 7540
rect 18046 7488 18052 7540
rect 18104 7528 18110 7540
rect 18230 7528 18236 7540
rect 18104 7500 18236 7528
rect 18104 7488 18110 7500
rect 18230 7488 18236 7500
rect 18288 7488 18294 7540
rect 18598 7488 18604 7540
rect 18656 7488 18662 7540
rect 19518 7488 19524 7540
rect 19576 7528 19582 7540
rect 21450 7528 21456 7540
rect 19576 7500 21456 7528
rect 19576 7488 19582 7500
rect 21450 7488 21456 7500
rect 21508 7488 21514 7540
rect 14829 7463 14887 7469
rect 14829 7460 14841 7463
rect 11296 7432 11834 7460
rect 11900 7432 14841 7460
rect 11296 7420 11302 7432
rect 9416 7364 9720 7392
rect 7561 7327 7619 7333
rect 5414 7296 6592 7324
rect 4801 7287 4859 7293
rect 4172 7228 4936 7256
rect 3973 7219 4031 7225
rect 4706 7188 4712 7200
rect 2372 7160 4712 7188
rect 2372 7148 2378 7160
rect 4706 7148 4712 7160
rect 4764 7148 4770 7200
rect 4908 7188 4936 7228
rect 5994 7188 6000 7200
rect 4908 7160 6000 7188
rect 5994 7148 6000 7160
rect 6052 7148 6058 7200
rect 6564 7197 6592 7296
rect 7561 7293 7573 7327
rect 7607 7293 7619 7327
rect 7561 7287 7619 7293
rect 7576 7256 7604 7287
rect 7742 7284 7748 7336
rect 7800 7284 7806 7336
rect 8294 7284 8300 7336
rect 8352 7324 8358 7336
rect 8481 7327 8539 7333
rect 8481 7324 8493 7327
rect 8352 7296 8493 7324
rect 8352 7284 8358 7296
rect 8481 7293 8493 7296
rect 8527 7293 8539 7327
rect 8481 7287 8539 7293
rect 8619 7327 8677 7333
rect 8619 7293 8631 7327
rect 8665 7324 8677 7327
rect 9416 7324 9444 7364
rect 10410 7352 10416 7404
rect 10468 7352 10474 7404
rect 10502 7352 10508 7404
rect 10560 7401 10566 7404
rect 10560 7395 10588 7401
rect 10576 7361 10588 7395
rect 10560 7355 10588 7361
rect 11517 7395 11575 7401
rect 11517 7361 11529 7395
rect 11563 7392 11575 7395
rect 11698 7392 11704 7404
rect 11563 7364 11704 7392
rect 11563 7361 11575 7364
rect 11517 7355 11575 7361
rect 10560 7352 10566 7355
rect 11698 7352 11704 7364
rect 11756 7352 11762 7404
rect 11806 7401 11834 7432
rect 14829 7429 14841 7432
rect 14875 7429 14887 7463
rect 14829 7423 14887 7429
rect 14921 7463 14979 7469
rect 14921 7429 14933 7463
rect 14967 7460 14979 7463
rect 15105 7463 15163 7469
rect 15105 7460 15117 7463
rect 14967 7432 15117 7460
rect 14967 7429 14979 7432
rect 14921 7423 14979 7429
rect 15105 7429 15117 7432
rect 15151 7429 15163 7463
rect 15105 7423 15163 7429
rect 16038 7460 16066 7488
rect 17236 7460 17264 7488
rect 16038 7432 17264 7460
rect 11791 7395 11849 7401
rect 11791 7361 11803 7395
rect 11837 7392 11849 7395
rect 12434 7392 12440 7404
rect 11837 7364 12440 7392
rect 11837 7361 11849 7364
rect 11791 7355 11849 7361
rect 12434 7352 12440 7364
rect 12492 7352 12498 7404
rect 13262 7352 13268 7404
rect 13320 7352 13326 7404
rect 14550 7352 14556 7404
rect 14608 7352 14614 7404
rect 14737 7395 14795 7401
rect 14737 7361 14749 7395
rect 14783 7392 14795 7395
rect 15010 7392 15016 7404
rect 14783 7364 15016 7392
rect 14783 7361 14795 7364
rect 14737 7355 14795 7361
rect 15010 7352 15016 7364
rect 15068 7352 15074 7404
rect 16038 7401 16066 7432
rect 15197 7395 15255 7401
rect 15197 7361 15209 7395
rect 15243 7392 15255 7395
rect 16015 7395 16073 7401
rect 15243 7364 15976 7392
rect 15243 7361 15255 7364
rect 15197 7355 15255 7361
rect 8665 7296 9444 7324
rect 9493 7327 9551 7333
rect 8665 7293 8677 7296
rect 8619 7287 8677 7293
rect 9493 7293 9505 7327
rect 9539 7293 9551 7327
rect 9493 7287 9551 7293
rect 7926 7256 7932 7268
rect 7576 7228 7932 7256
rect 7926 7216 7932 7228
rect 7984 7216 7990 7268
rect 8202 7216 8208 7268
rect 8260 7216 8266 7268
rect 9306 7216 9312 7268
rect 9364 7256 9370 7268
rect 9508 7256 9536 7287
rect 9674 7284 9680 7336
rect 9732 7324 9738 7336
rect 10042 7324 10048 7336
rect 9732 7296 10048 7324
rect 9732 7284 9738 7296
rect 10042 7284 10048 7296
rect 10100 7284 10106 7336
rect 10686 7284 10692 7336
rect 10744 7284 10750 7336
rect 13280 7324 13308 7352
rect 15838 7324 15844 7336
rect 13280 7296 15844 7324
rect 15838 7284 15844 7296
rect 15896 7284 15902 7336
rect 9364 7228 9536 7256
rect 9364 7216 9370 7228
rect 10134 7216 10140 7268
rect 10192 7216 10198 7268
rect 11164 7228 11652 7256
rect 6549 7191 6607 7197
rect 6549 7157 6561 7191
rect 6595 7157 6607 7191
rect 6549 7151 6607 7157
rect 6822 7148 6828 7200
rect 6880 7188 6886 7200
rect 7101 7191 7159 7197
rect 7101 7188 7113 7191
rect 6880 7160 7113 7188
rect 6880 7148 6886 7160
rect 7101 7157 7113 7160
rect 7147 7157 7159 7191
rect 7101 7151 7159 7157
rect 7742 7148 7748 7200
rect 7800 7188 7806 7200
rect 11164 7188 11192 7228
rect 7800 7160 11192 7188
rect 7800 7148 7806 7160
rect 11238 7148 11244 7200
rect 11296 7188 11302 7200
rect 11333 7191 11391 7197
rect 11333 7188 11345 7191
rect 11296 7160 11345 7188
rect 11296 7148 11302 7160
rect 11333 7157 11345 7160
rect 11379 7157 11391 7191
rect 11624 7188 11652 7228
rect 12434 7216 12440 7268
rect 12492 7256 12498 7268
rect 13906 7256 13912 7268
rect 12492 7228 13912 7256
rect 12492 7216 12498 7228
rect 13906 7216 13912 7228
rect 13964 7216 13970 7268
rect 14274 7216 14280 7268
rect 14332 7256 14338 7268
rect 15562 7256 15568 7268
rect 14332 7228 15568 7256
rect 14332 7216 14338 7228
rect 15562 7216 15568 7228
rect 15620 7216 15626 7268
rect 15948 7256 15976 7364
rect 16015 7361 16027 7395
rect 16061 7361 16073 7395
rect 16015 7355 16073 7361
rect 16209 7395 16267 7401
rect 16209 7361 16221 7395
rect 16255 7361 16267 7395
rect 16209 7355 16267 7361
rect 16022 7256 16028 7268
rect 15948 7228 16028 7256
rect 16022 7216 16028 7228
rect 16080 7216 16086 7268
rect 11882 7188 11888 7200
rect 11624 7160 11888 7188
rect 11333 7151 11391 7157
rect 11882 7148 11888 7160
rect 11940 7188 11946 7200
rect 15838 7188 15844 7200
rect 11940 7160 15844 7188
rect 11940 7148 11946 7160
rect 15838 7148 15844 7160
rect 15896 7148 15902 7200
rect 16224 7188 16252 7355
rect 16298 7352 16304 7404
rect 16356 7392 16362 7404
rect 16485 7395 16543 7401
rect 16485 7392 16497 7395
rect 16356 7364 16497 7392
rect 16356 7352 16362 7364
rect 16485 7361 16497 7364
rect 16531 7361 16543 7395
rect 16485 7355 16543 7361
rect 16853 7395 16911 7401
rect 16853 7361 16865 7395
rect 16899 7392 16911 7395
rect 17126 7392 17132 7404
rect 16899 7364 17132 7392
rect 16899 7361 16911 7364
rect 16853 7355 16911 7361
rect 17126 7352 17132 7364
rect 17184 7352 17190 7404
rect 17221 7395 17279 7401
rect 17221 7361 17233 7395
rect 17267 7392 17279 7395
rect 17512 7392 17540 7488
rect 18616 7460 18644 7488
rect 17604 7432 18644 7460
rect 17604 7401 17632 7432
rect 17267 7364 17540 7392
rect 17589 7395 17647 7401
rect 17267 7361 17279 7364
rect 17221 7355 17279 7361
rect 17589 7361 17601 7395
rect 17635 7361 17647 7395
rect 17589 7355 17647 7361
rect 17865 7395 17923 7401
rect 17865 7361 17877 7395
rect 17911 7361 17923 7395
rect 18325 7395 18383 7401
rect 18325 7392 18337 7395
rect 17865 7355 17923 7361
rect 18064 7364 18337 7392
rect 17880 7324 17908 7355
rect 18064 7336 18092 7364
rect 18325 7361 18337 7364
rect 18371 7361 18383 7395
rect 18325 7355 18383 7361
rect 18874 7352 18880 7404
rect 18932 7352 18938 7404
rect 19426 7352 19432 7404
rect 19484 7392 19490 7404
rect 19886 7392 19892 7404
rect 19484 7364 19892 7392
rect 19484 7352 19490 7364
rect 19886 7352 19892 7364
rect 19944 7392 19950 7404
rect 19981 7395 20039 7401
rect 19981 7392 19993 7395
rect 19944 7364 19993 7392
rect 19944 7352 19950 7364
rect 19981 7361 19993 7364
rect 20027 7361 20039 7395
rect 19981 7355 20039 7361
rect 20070 7352 20076 7404
rect 20128 7392 20134 7404
rect 20237 7395 20295 7401
rect 20237 7392 20249 7395
rect 20128 7364 20249 7392
rect 20128 7352 20134 7364
rect 20237 7361 20249 7364
rect 20283 7361 20295 7395
rect 20237 7355 20295 7361
rect 16316 7296 17908 7324
rect 16316 7265 16344 7296
rect 18046 7284 18052 7336
rect 18104 7284 18110 7336
rect 18601 7327 18659 7333
rect 18601 7324 18613 7327
rect 18340 7296 18613 7324
rect 18340 7268 18368 7296
rect 18601 7293 18613 7296
rect 18647 7293 18659 7327
rect 18601 7287 18659 7293
rect 19794 7284 19800 7336
rect 19852 7284 19858 7336
rect 16301 7259 16359 7265
rect 16301 7225 16313 7259
rect 16347 7225 16359 7259
rect 16301 7219 16359 7225
rect 16390 7216 16396 7268
rect 16448 7256 16454 7268
rect 17497 7259 17555 7265
rect 17497 7256 17509 7259
rect 16448 7228 17509 7256
rect 16448 7216 16454 7228
rect 17497 7225 17509 7228
rect 17543 7225 17555 7259
rect 18141 7259 18199 7265
rect 18141 7256 18153 7259
rect 17497 7219 17555 7225
rect 17604 7228 18153 7256
rect 17604 7188 17632 7228
rect 18141 7225 18153 7228
rect 18187 7225 18199 7259
rect 18141 7219 18199 7225
rect 18322 7216 18328 7268
rect 18380 7216 18386 7268
rect 19812 7256 19840 7284
rect 19306 7228 19840 7256
rect 16224 7160 17632 7188
rect 17770 7148 17776 7200
rect 17828 7188 17834 7200
rect 19306 7188 19334 7228
rect 17828 7160 19334 7188
rect 19613 7191 19671 7197
rect 17828 7148 17834 7160
rect 19613 7157 19625 7191
rect 19659 7188 19671 7191
rect 19978 7188 19984 7200
rect 19659 7160 19984 7188
rect 19659 7157 19671 7160
rect 19613 7151 19671 7157
rect 19978 7148 19984 7160
rect 20036 7148 20042 7200
rect 21358 7148 21364 7200
rect 21416 7148 21422 7200
rect 1104 7098 21896 7120
rect 1104 7046 3549 7098
rect 3601 7046 3613 7098
rect 3665 7046 3677 7098
rect 3729 7046 3741 7098
rect 3793 7046 3805 7098
rect 3857 7046 8747 7098
rect 8799 7046 8811 7098
rect 8863 7046 8875 7098
rect 8927 7046 8939 7098
rect 8991 7046 9003 7098
rect 9055 7046 13945 7098
rect 13997 7046 14009 7098
rect 14061 7046 14073 7098
rect 14125 7046 14137 7098
rect 14189 7046 14201 7098
rect 14253 7046 19143 7098
rect 19195 7046 19207 7098
rect 19259 7046 19271 7098
rect 19323 7046 19335 7098
rect 19387 7046 19399 7098
rect 19451 7046 21896 7098
rect 1104 7024 21896 7046
rect 3326 6944 3332 6996
rect 3384 6984 3390 6996
rect 6822 6984 6828 6996
rect 3384 6956 6828 6984
rect 3384 6944 3390 6956
rect 6822 6944 6828 6956
rect 6880 6944 6886 6996
rect 6914 6944 6920 6996
rect 6972 6944 6978 6996
rect 7101 6987 7159 6993
rect 7101 6953 7113 6987
rect 7147 6984 7159 6987
rect 8202 6984 8208 6996
rect 7147 6956 8208 6984
rect 7147 6953 7159 6956
rect 7101 6947 7159 6953
rect 8202 6944 8208 6956
rect 8260 6944 8266 6996
rect 8481 6987 8539 6993
rect 8481 6953 8493 6987
rect 8527 6984 8539 6987
rect 8662 6984 8668 6996
rect 8527 6956 8668 6984
rect 8527 6953 8539 6956
rect 8481 6947 8539 6953
rect 8662 6944 8668 6956
rect 8720 6944 8726 6996
rect 10410 6984 10416 6996
rect 8772 6956 10416 6984
rect 4065 6919 4123 6925
rect 4065 6885 4077 6919
rect 4111 6916 4123 6919
rect 4246 6916 4252 6928
rect 4111 6888 4252 6916
rect 4111 6885 4123 6888
rect 4065 6879 4123 6885
rect 4246 6876 4252 6888
rect 4304 6876 4310 6928
rect 4724 6888 4936 6916
rect 4724 6860 4752 6888
rect 1486 6808 1492 6860
rect 1544 6848 1550 6860
rect 1544 6820 2360 6848
rect 1544 6808 1550 6820
rect 1946 6780 1952 6792
rect 1504 6752 1952 6780
rect 1504 6721 1532 6752
rect 1946 6740 1952 6752
rect 2004 6740 2010 6792
rect 2332 6789 2360 6820
rect 4706 6808 4712 6860
rect 4764 6808 4770 6860
rect 4798 6808 4804 6860
rect 4856 6808 4862 6860
rect 4908 6848 4936 6888
rect 5994 6876 6000 6928
rect 6052 6876 6058 6928
rect 5077 6851 5135 6857
rect 5077 6848 5089 6851
rect 4908 6820 5089 6848
rect 5077 6817 5089 6820
rect 5123 6817 5135 6851
rect 5077 6811 5135 6817
rect 5215 6851 5273 6857
rect 5215 6817 5227 6851
rect 5261 6848 5273 6851
rect 5902 6848 5908 6860
rect 5261 6820 5908 6848
rect 5261 6817 5273 6820
rect 5215 6811 5273 6817
rect 5902 6808 5908 6820
rect 5960 6808 5966 6860
rect 6932 6848 6960 6944
rect 8294 6876 8300 6928
rect 8352 6916 8358 6928
rect 8772 6916 8800 6956
rect 10410 6944 10416 6956
rect 10468 6944 10474 6996
rect 10597 6987 10655 6993
rect 10597 6953 10609 6987
rect 10643 6984 10655 6987
rect 10686 6984 10692 6996
rect 10643 6956 10692 6984
rect 10643 6953 10655 6956
rect 10597 6947 10655 6953
rect 10686 6944 10692 6956
rect 10744 6944 10750 6996
rect 10980 6956 11744 6984
rect 8352 6888 8800 6916
rect 8352 6876 8358 6888
rect 10980 6860 11008 6956
rect 11716 6928 11744 6956
rect 11790 6944 11796 6996
rect 11848 6984 11854 6996
rect 11977 6987 12035 6993
rect 11977 6984 11989 6987
rect 11848 6956 11989 6984
rect 11848 6944 11854 6956
rect 11977 6953 11989 6956
rect 12023 6953 12035 6987
rect 11977 6947 12035 6953
rect 12894 6944 12900 6996
rect 12952 6944 12958 6996
rect 13817 6987 13875 6993
rect 13817 6953 13829 6987
rect 13863 6984 13875 6987
rect 14550 6984 14556 6996
rect 13863 6956 14556 6984
rect 13863 6953 13875 6956
rect 13817 6947 13875 6953
rect 14550 6944 14556 6956
rect 14608 6944 14614 6996
rect 15473 6987 15531 6993
rect 15473 6953 15485 6987
rect 15519 6953 15531 6987
rect 15473 6947 15531 6953
rect 11698 6876 11704 6928
rect 11756 6916 11762 6928
rect 12912 6916 12940 6944
rect 11756 6888 12940 6916
rect 15488 6916 15516 6947
rect 15838 6944 15844 6996
rect 15896 6984 15902 6996
rect 17957 6987 18015 6993
rect 15896 6956 17540 6984
rect 15896 6944 15902 6956
rect 16022 6916 16028 6928
rect 15488 6888 16028 6916
rect 11756 6876 11762 6888
rect 16022 6876 16028 6888
rect 16080 6876 16086 6928
rect 17512 6916 17540 6956
rect 17957 6953 17969 6987
rect 18003 6984 18015 6987
rect 18046 6984 18052 6996
rect 18003 6956 18052 6984
rect 18003 6953 18015 6956
rect 17957 6947 18015 6953
rect 18046 6944 18052 6956
rect 18104 6944 18110 6996
rect 18506 6944 18512 6996
rect 18564 6984 18570 6996
rect 18693 6987 18751 6993
rect 18693 6984 18705 6987
rect 18564 6956 18705 6984
rect 18564 6944 18570 6956
rect 18693 6953 18705 6956
rect 18739 6953 18751 6987
rect 18693 6947 18751 6953
rect 18782 6956 20576 6984
rect 18782 6916 18810 6956
rect 17512 6888 18810 6916
rect 18877 6919 18935 6925
rect 18877 6885 18889 6919
rect 18923 6916 18935 6919
rect 19242 6916 19248 6928
rect 18923 6888 19248 6916
rect 18923 6885 18935 6888
rect 18877 6879 18935 6885
rect 19242 6876 19248 6888
rect 19300 6876 19306 6928
rect 20070 6916 20076 6928
rect 19352 6888 20076 6916
rect 7469 6851 7527 6857
rect 7469 6848 7481 6851
rect 6932 6820 7481 6848
rect 7469 6817 7481 6820
rect 7515 6817 7527 6851
rect 7469 6811 7527 6817
rect 2317 6783 2375 6789
rect 2317 6749 2329 6783
rect 2363 6749 2375 6783
rect 2317 6743 2375 6749
rect 2591 6783 2649 6789
rect 2591 6749 2603 6783
rect 2637 6780 2649 6783
rect 3326 6780 3332 6792
rect 2637 6752 3332 6780
rect 2637 6749 2649 6752
rect 2591 6743 2649 6749
rect 1489 6715 1547 6721
rect 1489 6681 1501 6715
rect 1535 6681 1547 6715
rect 2332 6712 2360 6743
rect 3326 6740 3332 6752
rect 3384 6740 3390 6792
rect 3694 6740 3700 6792
rect 3752 6740 3758 6792
rect 4157 6783 4215 6789
rect 4157 6749 4169 6783
rect 4203 6780 4215 6783
rect 4246 6780 4252 6792
rect 4203 6752 4252 6780
rect 4203 6749 4215 6752
rect 4157 6743 4215 6749
rect 4246 6740 4252 6752
rect 4304 6740 4310 6792
rect 4341 6783 4399 6789
rect 4341 6749 4353 6783
rect 4387 6780 4399 6783
rect 4522 6780 4528 6792
rect 4387 6752 4528 6780
rect 4387 6749 4399 6752
rect 4341 6743 4399 6749
rect 4522 6740 4528 6752
rect 4580 6740 4586 6792
rect 5350 6740 5356 6792
rect 5408 6740 5414 6792
rect 3712 6712 3740 6740
rect 2332 6684 3740 6712
rect 3881 6715 3939 6721
rect 1489 6675 1547 6681
rect 3881 6681 3893 6715
rect 3927 6681 3939 6715
rect 5920 6712 5948 6808
rect 6086 6740 6092 6792
rect 6144 6740 6150 6792
rect 6363 6783 6421 6789
rect 6363 6749 6375 6783
rect 6409 6780 6421 6783
rect 6730 6780 6736 6792
rect 6409 6752 6736 6780
rect 6409 6749 6421 6752
rect 6363 6743 6421 6749
rect 6730 6740 6736 6752
rect 6788 6740 6794 6792
rect 7374 6712 7380 6724
rect 5920 6684 7380 6712
rect 3881 6675 3939 6681
rect 1765 6647 1823 6653
rect 1765 6613 1777 6647
rect 1811 6644 1823 6647
rect 2498 6644 2504 6656
rect 1811 6616 2504 6644
rect 1811 6613 1823 6616
rect 1765 6607 1823 6613
rect 2498 6604 2504 6616
rect 2556 6604 2562 6656
rect 3329 6647 3387 6653
rect 3329 6613 3341 6647
rect 3375 6644 3387 6647
rect 3418 6644 3424 6656
rect 3375 6616 3424 6644
rect 3375 6613 3387 6616
rect 3329 6607 3387 6613
rect 3418 6604 3424 6616
rect 3476 6604 3482 6656
rect 3896 6644 3924 6675
rect 7374 6672 7380 6684
rect 7432 6672 7438 6724
rect 7484 6712 7512 6811
rect 8478 6808 8484 6860
rect 8536 6848 8542 6860
rect 9306 6848 9312 6860
rect 8536 6820 9312 6848
rect 8536 6808 8542 6820
rect 9306 6808 9312 6820
rect 9364 6848 9370 6860
rect 9585 6851 9643 6857
rect 9585 6848 9597 6851
rect 9364 6820 9597 6848
rect 9364 6808 9370 6820
rect 9585 6817 9597 6820
rect 9631 6817 9643 6851
rect 9585 6811 9643 6817
rect 10962 6808 10968 6860
rect 11020 6808 11026 6860
rect 18966 6848 18972 6860
rect 18340 6820 18972 6848
rect 7743 6783 7801 6789
rect 7743 6749 7755 6783
rect 7789 6780 7801 6783
rect 9859 6783 9917 6789
rect 7789 6752 9536 6780
rect 7789 6749 7801 6752
rect 7743 6743 7801 6749
rect 9508 6712 9536 6752
rect 9859 6749 9871 6783
rect 9905 6780 9917 6783
rect 9950 6780 9956 6792
rect 9905 6752 9956 6780
rect 9905 6749 9917 6752
rect 9859 6743 9917 6749
rect 9950 6740 9956 6752
rect 10008 6780 10014 6792
rect 10778 6780 10784 6792
rect 10008 6752 10784 6780
rect 10008 6740 10014 6752
rect 10778 6740 10784 6752
rect 10836 6740 10842 6792
rect 11239 6783 11297 6789
rect 11239 6749 11251 6783
rect 11285 6780 11297 6783
rect 12250 6780 12256 6792
rect 11285 6752 12256 6780
rect 11285 6749 11297 6752
rect 11239 6743 11297 6749
rect 12250 6740 12256 6752
rect 12308 6740 12314 6792
rect 13722 6740 13728 6792
rect 13780 6740 13786 6792
rect 14090 6740 14096 6792
rect 14148 6740 14154 6792
rect 14335 6783 14393 6789
rect 14335 6780 14347 6783
rect 14200 6752 14347 6780
rect 13262 6712 13268 6724
rect 7484 6684 7786 6712
rect 9508 6684 13268 6712
rect 4982 6644 4988 6656
rect 3896 6616 4988 6644
rect 4982 6604 4988 6616
rect 5040 6644 5046 6656
rect 7650 6644 7656 6656
rect 5040 6616 7656 6644
rect 5040 6604 5046 6616
rect 7650 6604 7656 6616
rect 7708 6604 7714 6656
rect 7758 6644 7786 6684
rect 13262 6672 13268 6684
rect 13320 6672 13326 6724
rect 10962 6644 10968 6656
rect 7758 6616 10968 6644
rect 10962 6604 10968 6616
rect 11020 6604 11026 6656
rect 11882 6604 11888 6656
rect 11940 6644 11946 6656
rect 14200 6644 14228 6752
rect 14335 6749 14347 6752
rect 14381 6780 14393 6783
rect 14458 6780 14464 6792
rect 14381 6752 14464 6780
rect 14381 6749 14393 6752
rect 14335 6743 14393 6749
rect 14458 6740 14464 6752
rect 14516 6740 14522 6792
rect 15654 6740 15660 6792
rect 15712 6740 15718 6792
rect 16577 6783 16635 6789
rect 16577 6749 16589 6783
rect 16623 6780 16635 6783
rect 16623 6752 16988 6780
rect 16623 6749 16635 6752
rect 16577 6743 16635 6749
rect 16298 6672 16304 6724
rect 16356 6712 16362 6724
rect 16822 6715 16880 6721
rect 16822 6712 16834 6715
rect 16356 6684 16834 6712
rect 16356 6672 16362 6684
rect 16822 6681 16834 6684
rect 16868 6681 16880 6715
rect 16822 6675 16880 6681
rect 16960 6656 16988 6752
rect 18230 6740 18236 6792
rect 18288 6740 18294 6792
rect 18340 6789 18368 6820
rect 18966 6808 18972 6820
rect 19024 6808 19030 6860
rect 19352 6792 19380 6888
rect 20070 6876 20076 6888
rect 20128 6876 20134 6928
rect 20548 6925 20576 6956
rect 20533 6919 20591 6925
rect 20533 6885 20545 6919
rect 20579 6885 20591 6919
rect 20533 6879 20591 6885
rect 19521 6851 19579 6857
rect 19521 6817 19533 6851
rect 19567 6848 19579 6851
rect 20993 6851 21051 6857
rect 20993 6848 21005 6851
rect 19567 6820 20116 6848
rect 19567 6817 19579 6820
rect 19521 6811 19579 6817
rect 18325 6783 18383 6789
rect 18325 6749 18337 6783
rect 18371 6749 18383 6783
rect 18325 6743 18383 6749
rect 18601 6783 18659 6789
rect 18601 6749 18613 6783
rect 18647 6749 18659 6783
rect 18601 6743 18659 6749
rect 19061 6783 19119 6789
rect 19061 6749 19073 6783
rect 19107 6780 19119 6783
rect 19334 6780 19340 6792
rect 19107 6752 19340 6780
rect 19107 6749 19119 6752
rect 19061 6743 19119 6749
rect 18616 6712 18644 6743
rect 19334 6740 19340 6752
rect 19392 6740 19398 6792
rect 19429 6783 19487 6789
rect 19429 6749 19441 6783
rect 19475 6749 19487 6783
rect 19429 6743 19487 6749
rect 18616 6684 19012 6712
rect 11940 6616 14228 6644
rect 11940 6604 11946 6616
rect 14642 6604 14648 6656
rect 14700 6644 14706 6656
rect 15105 6647 15163 6653
rect 15105 6644 15117 6647
rect 14700 6616 15117 6644
rect 14700 6604 14706 6616
rect 15105 6613 15117 6616
rect 15151 6613 15163 6647
rect 15105 6607 15163 6613
rect 16942 6604 16948 6656
rect 17000 6604 17006 6656
rect 18046 6604 18052 6656
rect 18104 6604 18110 6656
rect 18509 6647 18567 6653
rect 18509 6613 18521 6647
rect 18555 6644 18567 6647
rect 18690 6644 18696 6656
rect 18555 6616 18696 6644
rect 18555 6613 18567 6616
rect 18509 6607 18567 6613
rect 18690 6604 18696 6616
rect 18748 6604 18754 6656
rect 18984 6644 19012 6684
rect 19242 6672 19248 6724
rect 19300 6712 19306 6724
rect 19444 6712 19472 6743
rect 19610 6740 19616 6792
rect 19668 6780 19674 6792
rect 20088 6789 20116 6820
rect 20640 6820 21005 6848
rect 20640 6789 20668 6820
rect 20993 6817 21005 6820
rect 21039 6817 21051 6851
rect 20993 6811 21051 6817
rect 21174 6808 21180 6860
rect 21232 6848 21238 6860
rect 21232 6820 21404 6848
rect 21232 6808 21238 6820
rect 19705 6783 19763 6789
rect 19705 6780 19717 6783
rect 19668 6752 19717 6780
rect 19668 6740 19674 6752
rect 19705 6749 19717 6752
rect 19751 6749 19763 6783
rect 19705 6743 19763 6749
rect 20073 6783 20131 6789
rect 20073 6749 20085 6783
rect 20119 6749 20131 6783
rect 20073 6743 20131 6749
rect 20625 6783 20683 6789
rect 20625 6749 20637 6783
rect 20671 6749 20683 6783
rect 20901 6783 20959 6789
rect 20901 6780 20913 6783
rect 20625 6743 20683 6749
rect 20732 6752 20913 6780
rect 19300 6684 19472 6712
rect 19720 6712 19748 6743
rect 20732 6712 20760 6752
rect 20901 6749 20913 6752
rect 20947 6749 20959 6783
rect 20901 6743 20959 6749
rect 21082 6740 21088 6792
rect 21140 6740 21146 6792
rect 21376 6789 21404 6820
rect 21361 6783 21419 6789
rect 21361 6749 21373 6783
rect 21407 6749 21419 6783
rect 21361 6743 21419 6749
rect 19720 6684 20760 6712
rect 19300 6672 19306 6684
rect 19058 6644 19064 6656
rect 18984 6616 19064 6644
rect 19058 6604 19064 6616
rect 19116 6604 19122 6656
rect 19150 6604 19156 6656
rect 19208 6644 19214 6656
rect 20898 6644 20904 6656
rect 19208 6616 20904 6644
rect 19208 6604 19214 6616
rect 20898 6604 20904 6616
rect 20956 6604 20962 6656
rect 21177 6647 21235 6653
rect 21177 6613 21189 6647
rect 21223 6644 21235 6647
rect 21266 6644 21272 6656
rect 21223 6616 21272 6644
rect 21223 6613 21235 6616
rect 21177 6607 21235 6613
rect 21266 6604 21272 6616
rect 21324 6604 21330 6656
rect 1104 6554 22056 6576
rect 1104 6502 6148 6554
rect 6200 6502 6212 6554
rect 6264 6502 6276 6554
rect 6328 6502 6340 6554
rect 6392 6502 6404 6554
rect 6456 6502 11346 6554
rect 11398 6502 11410 6554
rect 11462 6502 11474 6554
rect 11526 6502 11538 6554
rect 11590 6502 11602 6554
rect 11654 6502 16544 6554
rect 16596 6502 16608 6554
rect 16660 6502 16672 6554
rect 16724 6502 16736 6554
rect 16788 6502 16800 6554
rect 16852 6502 21742 6554
rect 21794 6502 21806 6554
rect 21858 6502 21870 6554
rect 21922 6502 21934 6554
rect 21986 6502 21998 6554
rect 22050 6502 22056 6554
rect 1104 6480 22056 6502
rect 1210 6400 1216 6452
rect 1268 6440 1274 6452
rect 2501 6443 2559 6449
rect 1268 6412 1808 6440
rect 1268 6400 1274 6412
rect 1780 6343 1808 6412
rect 2501 6409 2513 6443
rect 2547 6440 2559 6443
rect 3142 6440 3148 6452
rect 2547 6412 3148 6440
rect 2547 6409 2559 6412
rect 2501 6403 2559 6409
rect 3142 6400 3148 6412
rect 3200 6400 3206 6452
rect 3421 6443 3479 6449
rect 3421 6409 3433 6443
rect 3467 6440 3479 6443
rect 3510 6440 3516 6452
rect 3467 6412 3516 6440
rect 3467 6409 3479 6412
rect 3421 6403 3479 6409
rect 3510 6400 3516 6412
rect 3568 6400 3574 6452
rect 3973 6443 4031 6449
rect 3973 6409 3985 6443
rect 4019 6440 4031 6443
rect 4154 6440 4160 6452
rect 4019 6412 4160 6440
rect 4019 6409 4031 6412
rect 3973 6403 4031 6409
rect 4154 6400 4160 6412
rect 4212 6400 4218 6452
rect 5074 6400 5080 6452
rect 5132 6440 5138 6452
rect 5353 6443 5411 6449
rect 5353 6440 5365 6443
rect 5132 6412 5365 6440
rect 5132 6400 5138 6412
rect 5353 6409 5365 6412
rect 5399 6409 5411 6443
rect 5353 6403 5411 6409
rect 5534 6400 5540 6452
rect 5592 6400 5598 6452
rect 5828 6412 8156 6440
rect 5552 6372 5580 6400
rect 5828 6381 5856 6412
rect 8128 6384 8156 6412
rect 10134 6400 10140 6452
rect 10192 6440 10198 6452
rect 10321 6443 10379 6449
rect 10321 6440 10333 6443
rect 10192 6412 10333 6440
rect 10192 6400 10198 6412
rect 10321 6409 10333 6412
rect 10367 6409 10379 6443
rect 10321 6403 10379 6409
rect 11054 6400 11060 6452
rect 11112 6400 11118 6452
rect 11238 6400 11244 6452
rect 11296 6400 11302 6452
rect 13262 6400 13268 6452
rect 13320 6440 13326 6452
rect 13538 6440 13544 6452
rect 13320 6412 13544 6440
rect 13320 6400 13326 6412
rect 13538 6400 13544 6412
rect 13596 6400 13602 6452
rect 13722 6400 13728 6452
rect 13780 6440 13786 6452
rect 14001 6443 14059 6449
rect 14001 6440 14013 6443
rect 13780 6412 14013 6440
rect 13780 6400 13786 6412
rect 14001 6409 14013 6412
rect 14047 6409 14059 6443
rect 14001 6403 14059 6409
rect 14182 6400 14188 6452
rect 14240 6440 14246 6452
rect 14240 6412 15516 6440
rect 14240 6400 14246 6412
rect 1747 6337 1808 6343
rect 1486 6264 1492 6316
rect 1544 6264 1550 6316
rect 1747 6303 1759 6337
rect 1793 6306 1808 6337
rect 2148 6344 5580 6372
rect 5813 6375 5871 6381
rect 1793 6303 1805 6306
rect 1747 6297 1805 6303
rect 1486 6060 1492 6112
rect 1544 6100 1550 6112
rect 2148 6100 2176 6344
rect 5813 6341 5825 6375
rect 5859 6341 5871 6375
rect 5813 6335 5871 6341
rect 6549 6375 6607 6381
rect 6549 6341 6561 6375
rect 6595 6372 6607 6375
rect 7558 6372 7564 6384
rect 6595 6344 7564 6372
rect 6595 6341 6607 6344
rect 6549 6335 6607 6341
rect 7558 6332 7564 6344
rect 7616 6332 7622 6384
rect 7650 6332 7656 6384
rect 7708 6332 7714 6384
rect 8110 6332 8116 6384
rect 8168 6332 8174 6384
rect 9766 6372 9772 6384
rect 9598 6344 9772 6372
rect 9598 6343 9626 6344
rect 9567 6337 9626 6343
rect 3145 6307 3203 6313
rect 3145 6273 3157 6307
rect 3191 6304 3203 6307
rect 3605 6307 3663 6313
rect 3605 6304 3617 6307
rect 3191 6276 3617 6304
rect 3191 6273 3203 6276
rect 3145 6267 3203 6273
rect 3605 6273 3617 6276
rect 3651 6304 3663 6307
rect 3786 6304 3792 6316
rect 3651 6276 3792 6304
rect 3651 6273 3663 6276
rect 3605 6267 3663 6273
rect 3786 6264 3792 6276
rect 3844 6264 3850 6316
rect 3881 6307 3939 6313
rect 3881 6273 3893 6307
rect 3927 6273 3939 6307
rect 3881 6267 3939 6273
rect 3418 6196 3424 6248
rect 3476 6236 3482 6248
rect 3896 6236 3924 6267
rect 4338 6264 4344 6316
rect 4396 6264 4402 6316
rect 4615 6307 4673 6313
rect 4615 6273 4627 6307
rect 4661 6304 4673 6307
rect 5074 6304 5080 6316
rect 4661 6276 5080 6304
rect 4661 6273 4673 6276
rect 4615 6267 4673 6273
rect 5074 6264 5080 6276
rect 5132 6264 5138 6316
rect 6822 6264 6828 6316
rect 6880 6264 6886 6316
rect 6914 6264 6920 6316
rect 6972 6264 6978 6316
rect 7282 6264 7288 6316
rect 7340 6264 7346 6316
rect 7374 6264 7380 6316
rect 7432 6304 7438 6316
rect 7432 6276 7694 6304
rect 7432 6264 7438 6276
rect 3476 6208 3924 6236
rect 6368 6248 6420 6254
rect 3476 6196 3482 6208
rect 6368 6190 6420 6196
rect 3694 6128 3700 6180
rect 3752 6168 3758 6180
rect 4338 6168 4344 6180
rect 3752 6140 4344 6168
rect 3752 6128 3758 6140
rect 4338 6128 4344 6140
rect 4396 6128 4402 6180
rect 7666 6168 7694 6276
rect 9306 6264 9312 6316
rect 9364 6264 9370 6316
rect 9567 6303 9579 6337
rect 9613 6306 9626 6337
rect 9766 6332 9772 6344
rect 9824 6332 9830 6384
rect 9613 6303 9625 6306
rect 9567 6297 9625 6303
rect 9784 6304 9812 6332
rect 10873 6307 10931 6313
rect 9784 6276 9996 6304
rect 7837 6171 7895 6177
rect 7837 6168 7849 6171
rect 7666 6140 7849 6168
rect 7837 6137 7849 6140
rect 7883 6137 7895 6171
rect 9968 6168 9996 6276
rect 10873 6273 10885 6307
rect 10919 6304 10931 6307
rect 11072 6304 11100 6400
rect 10919 6276 11100 6304
rect 11149 6307 11207 6313
rect 10919 6273 10931 6276
rect 10873 6267 10931 6273
rect 11149 6273 11161 6307
rect 11195 6304 11207 6307
rect 11256 6304 11284 6400
rect 12894 6332 12900 6384
rect 12952 6372 12958 6384
rect 14090 6372 14096 6384
rect 12952 6344 14096 6372
rect 12952 6332 12958 6344
rect 14090 6332 14096 6344
rect 14148 6372 14154 6384
rect 14366 6372 14372 6384
rect 14148 6344 14372 6372
rect 14148 6332 14154 6344
rect 14366 6332 14372 6344
rect 14424 6372 14430 6384
rect 15488 6372 15516 6412
rect 15654 6400 15660 6452
rect 15712 6400 15718 6452
rect 16022 6400 16028 6452
rect 16080 6440 16086 6452
rect 17494 6440 17500 6452
rect 16080 6412 17500 6440
rect 16080 6400 16086 6412
rect 17494 6400 17500 6412
rect 17552 6400 17558 6452
rect 18141 6443 18199 6449
rect 18141 6409 18153 6443
rect 18187 6440 18199 6443
rect 18690 6440 18696 6452
rect 18187 6412 18696 6440
rect 18187 6409 18199 6412
rect 18141 6403 18199 6409
rect 18690 6400 18696 6412
rect 18748 6400 18754 6452
rect 19242 6400 19248 6452
rect 19300 6440 19306 6452
rect 20714 6440 20720 6452
rect 19300 6412 20720 6440
rect 19300 6400 19306 6412
rect 20714 6400 20720 6412
rect 20772 6400 20778 6452
rect 20806 6400 20812 6452
rect 20864 6400 20870 6452
rect 20898 6400 20904 6452
rect 20956 6440 20962 6452
rect 21269 6443 21327 6449
rect 21269 6440 21281 6443
rect 20956 6412 21281 6440
rect 20956 6400 20962 6412
rect 21269 6409 21281 6412
rect 21315 6409 21327 6443
rect 21269 6403 21327 6409
rect 21361 6443 21419 6449
rect 21361 6409 21373 6443
rect 21407 6440 21419 6443
rect 21450 6440 21456 6452
rect 21407 6412 21456 6440
rect 21407 6409 21419 6412
rect 21361 6403 21419 6409
rect 21450 6400 21456 6412
rect 21508 6400 21514 6452
rect 20162 6381 20168 6384
rect 17773 6375 17831 6381
rect 17773 6372 17785 6375
rect 14424 6344 15424 6372
rect 15488 6344 17785 6372
rect 14424 6332 14430 6344
rect 11195 6276 11284 6304
rect 11609 6307 11667 6313
rect 11195 6273 11207 6276
rect 11149 6267 11207 6273
rect 11609 6273 11621 6307
rect 11655 6304 11667 6307
rect 12158 6304 12164 6316
rect 11655 6276 12164 6304
rect 11655 6273 11667 6276
rect 11609 6267 11667 6273
rect 12158 6264 12164 6276
rect 12216 6264 12222 6316
rect 14550 6313 14556 6316
rect 14185 6307 14243 6313
rect 14185 6273 14197 6307
rect 14231 6304 14243 6307
rect 14544 6304 14556 6313
rect 14231 6276 14556 6304
rect 14231 6273 14243 6276
rect 14185 6267 14243 6273
rect 14544 6267 14556 6276
rect 14550 6264 14556 6267
rect 14608 6264 14614 6316
rect 10042 6196 10048 6248
rect 10100 6236 10106 6248
rect 10100 6208 14228 6236
rect 10100 6196 10106 6208
rect 14200 6180 14228 6208
rect 14274 6196 14280 6248
rect 14332 6196 14338 6248
rect 15396 6236 15424 6344
rect 17773 6341 17785 6344
rect 17819 6341 17831 6375
rect 20156 6372 20168 6381
rect 17773 6335 17831 6341
rect 17972 6344 19334 6372
rect 20123 6344 20168 6372
rect 15654 6264 15660 6316
rect 15712 6304 15718 6316
rect 15749 6307 15807 6313
rect 15749 6304 15761 6307
rect 15712 6276 15761 6304
rect 15712 6264 15718 6276
rect 15749 6273 15761 6276
rect 15795 6273 15807 6307
rect 15749 6267 15807 6273
rect 15838 6264 15844 6316
rect 15896 6304 15902 6316
rect 15933 6307 15991 6313
rect 15933 6304 15945 6307
rect 15896 6276 15945 6304
rect 15896 6264 15902 6276
rect 15933 6273 15945 6276
rect 15979 6273 15991 6307
rect 15933 6267 15991 6273
rect 17034 6264 17040 6316
rect 17092 6264 17098 6316
rect 17494 6264 17500 6316
rect 17552 6264 17558 6316
rect 17972 6313 18000 6344
rect 17957 6307 18015 6313
rect 17957 6273 17969 6307
rect 18003 6273 18015 6307
rect 17957 6267 18015 6273
rect 18141 6307 18199 6313
rect 18141 6273 18153 6307
rect 18187 6304 18199 6307
rect 18230 6304 18236 6316
rect 18187 6276 18236 6304
rect 18187 6273 18199 6276
rect 18141 6267 18199 6273
rect 18230 6264 18236 6276
rect 18288 6264 18294 6316
rect 18414 6264 18420 6316
rect 18472 6264 18478 6316
rect 18782 6264 18788 6316
rect 18840 6264 18846 6316
rect 19306 6304 19334 6344
rect 20156 6335 20168 6344
rect 20162 6332 20168 6335
rect 20220 6332 20226 6384
rect 19306 6276 19564 6304
rect 16853 6239 16911 6245
rect 15396 6208 15774 6236
rect 11882 6168 11888 6180
rect 9968 6140 11888 6168
rect 7837 6131 7895 6137
rect 11882 6128 11888 6140
rect 11940 6128 11946 6180
rect 14182 6128 14188 6180
rect 14240 6128 14246 6180
rect 15654 6168 15660 6180
rect 15212 6140 15660 6168
rect 1544 6072 2176 6100
rect 1544 6060 1550 6072
rect 2866 6060 2872 6112
rect 2924 6100 2930 6112
rect 3142 6100 3148 6112
rect 2924 6072 3148 6100
rect 2924 6060 2930 6072
rect 3142 6060 3148 6072
rect 3200 6060 3206 6112
rect 4062 6060 4068 6112
rect 4120 6100 4126 6112
rect 5905 6103 5963 6109
rect 5905 6100 5917 6103
rect 4120 6072 5917 6100
rect 4120 6060 4126 6072
rect 5905 6069 5917 6072
rect 5951 6069 5963 6103
rect 5905 6063 5963 6069
rect 5994 6060 6000 6112
rect 6052 6100 6058 6112
rect 6546 6100 6552 6112
rect 6052 6072 6552 6100
rect 6052 6060 6058 6072
rect 6546 6060 6552 6072
rect 6604 6060 6610 6112
rect 9674 6060 9680 6112
rect 9732 6100 9738 6112
rect 10689 6103 10747 6109
rect 10689 6100 10701 6103
rect 9732 6072 10701 6100
rect 9732 6060 9738 6072
rect 10689 6069 10701 6072
rect 10735 6069 10747 6103
rect 10689 6063 10747 6069
rect 10962 6060 10968 6112
rect 11020 6060 11026 6112
rect 11790 6060 11796 6112
rect 11848 6060 11854 6112
rect 14642 6060 14648 6112
rect 14700 6100 14706 6112
rect 15212 6100 15240 6140
rect 15654 6128 15660 6140
rect 15712 6128 15718 6180
rect 15746 6168 15774 6208
rect 16853 6205 16865 6239
rect 16899 6236 16911 6239
rect 17126 6236 17132 6248
rect 16899 6208 17132 6236
rect 16899 6205 16911 6208
rect 16853 6199 16911 6205
rect 17126 6196 17132 6208
rect 17184 6196 17190 6248
rect 18506 6196 18512 6248
rect 18564 6196 18570 6248
rect 18524 6168 18552 6196
rect 15746 6140 18552 6168
rect 19334 6128 19340 6180
rect 19392 6128 19398 6180
rect 14700 6072 15240 6100
rect 14700 6060 14706 6072
rect 15286 6060 15292 6112
rect 15344 6100 15350 6112
rect 15841 6103 15899 6109
rect 15841 6100 15853 6103
rect 15344 6072 15853 6100
rect 15344 6060 15350 6072
rect 15841 6069 15853 6072
rect 15887 6069 15899 6103
rect 15841 6063 15899 6069
rect 18233 6103 18291 6109
rect 18233 6069 18245 6103
rect 18279 6100 18291 6103
rect 19352 6100 19380 6128
rect 19536 6109 19564 6276
rect 19886 6264 19892 6316
rect 19944 6264 19950 6316
rect 20824 6304 20852 6400
rect 21545 6307 21603 6313
rect 21545 6304 21557 6307
rect 20824 6276 21557 6304
rect 21545 6273 21557 6276
rect 21591 6273 21603 6307
rect 21545 6267 21603 6273
rect 18279 6072 19380 6100
rect 19521 6103 19579 6109
rect 18279 6069 18291 6072
rect 18233 6063 18291 6069
rect 19521 6069 19533 6103
rect 19567 6100 19579 6103
rect 20898 6100 20904 6112
rect 19567 6072 20904 6100
rect 19567 6069 19579 6072
rect 19521 6063 19579 6069
rect 20898 6060 20904 6072
rect 20956 6060 20962 6112
rect 1104 6010 21896 6032
rect 1104 5958 3549 6010
rect 3601 5958 3613 6010
rect 3665 5958 3677 6010
rect 3729 5958 3741 6010
rect 3793 5958 3805 6010
rect 3857 5958 8747 6010
rect 8799 5958 8811 6010
rect 8863 5958 8875 6010
rect 8927 5958 8939 6010
rect 8991 5958 9003 6010
rect 9055 5958 13945 6010
rect 13997 5958 14009 6010
rect 14061 5958 14073 6010
rect 14125 5958 14137 6010
rect 14189 5958 14201 6010
rect 14253 5958 19143 6010
rect 19195 5958 19207 6010
rect 19259 5958 19271 6010
rect 19323 5958 19335 6010
rect 19387 5958 19399 6010
rect 19451 5958 21896 6010
rect 1104 5936 21896 5958
rect 1486 5856 1492 5908
rect 1544 5856 1550 5908
rect 1872 5868 4016 5896
rect 1302 5720 1308 5772
rect 1360 5760 1366 5772
rect 1765 5763 1823 5769
rect 1765 5760 1777 5763
rect 1360 5732 1777 5760
rect 1360 5720 1366 5732
rect 1765 5729 1777 5732
rect 1811 5729 1823 5763
rect 1765 5723 1823 5729
rect 1578 5652 1584 5704
rect 1636 5652 1642 5704
rect 1673 5695 1731 5701
rect 1673 5661 1685 5695
rect 1719 5692 1731 5695
rect 1872 5692 1900 5868
rect 3988 5828 4016 5868
rect 4062 5856 4068 5908
rect 4120 5896 4126 5908
rect 5626 5896 5632 5908
rect 4120 5868 5632 5896
rect 4120 5856 4126 5868
rect 5626 5856 5632 5868
rect 5684 5856 5690 5908
rect 5902 5856 5908 5908
rect 5960 5856 5966 5908
rect 6178 5856 6184 5908
rect 6236 5856 6242 5908
rect 6638 5856 6644 5908
rect 6696 5856 6702 5908
rect 6914 5856 6920 5908
rect 6972 5896 6978 5908
rect 7561 5899 7619 5905
rect 7561 5896 7573 5899
rect 6972 5868 7573 5896
rect 6972 5856 6978 5868
rect 7561 5865 7573 5868
rect 7607 5865 7619 5899
rect 7561 5859 7619 5865
rect 9858 5856 9864 5908
rect 9916 5856 9922 5908
rect 11698 5856 11704 5908
rect 11756 5896 11762 5908
rect 15102 5896 15108 5908
rect 11756 5868 15108 5896
rect 11756 5856 11762 5868
rect 15102 5856 15108 5868
rect 15160 5856 15166 5908
rect 15286 5856 15292 5908
rect 15344 5856 15350 5908
rect 15381 5899 15439 5905
rect 15381 5865 15393 5899
rect 15427 5896 15439 5899
rect 15470 5896 15476 5908
rect 15427 5868 15476 5896
rect 15427 5865 15439 5868
rect 15381 5859 15439 5865
rect 15470 5856 15476 5868
rect 15528 5856 15534 5908
rect 15565 5899 15623 5905
rect 15565 5865 15577 5899
rect 15611 5896 15623 5899
rect 15838 5896 15844 5908
rect 15611 5868 15844 5896
rect 15611 5865 15623 5868
rect 15565 5859 15623 5865
rect 15838 5856 15844 5868
rect 15896 5856 15902 5908
rect 15933 5899 15991 5905
rect 15933 5865 15945 5899
rect 15979 5896 15991 5899
rect 17034 5896 17040 5908
rect 15979 5868 17040 5896
rect 15979 5865 15991 5868
rect 15933 5859 15991 5865
rect 17034 5856 17040 5868
rect 17092 5856 17098 5908
rect 17126 5856 17132 5908
rect 17184 5856 17190 5908
rect 18046 5856 18052 5908
rect 18104 5896 18110 5908
rect 18104 5868 20852 5896
rect 18104 5856 18110 5868
rect 4154 5828 4160 5840
rect 2332 5800 2544 5828
rect 3988 5800 4160 5828
rect 2332 5772 2360 5800
rect 2314 5720 2320 5772
rect 2372 5720 2378 5772
rect 2406 5720 2412 5772
rect 2464 5720 2470 5772
rect 2516 5760 2544 5800
rect 4154 5788 4160 5800
rect 4212 5788 4218 5840
rect 4246 5788 4252 5840
rect 4304 5788 4310 5840
rect 4430 5788 4436 5840
rect 4488 5828 4494 5840
rect 4709 5831 4767 5837
rect 4709 5828 4721 5831
rect 4488 5800 4721 5828
rect 4488 5788 4494 5800
rect 4709 5797 4721 5800
rect 4755 5797 4767 5831
rect 4709 5791 4767 5797
rect 2685 5763 2743 5769
rect 2685 5760 2697 5763
rect 2516 5732 2697 5760
rect 2685 5729 2697 5732
rect 2731 5729 2743 5763
rect 2685 5723 2743 5729
rect 2823 5763 2881 5769
rect 2823 5729 2835 5763
rect 2869 5760 2881 5763
rect 3878 5760 3884 5772
rect 2869 5732 3884 5760
rect 2869 5729 2881 5732
rect 2823 5723 2881 5729
rect 3878 5720 3884 5732
rect 3936 5720 3942 5772
rect 4065 5763 4123 5769
rect 4065 5729 4077 5763
rect 4111 5760 4123 5763
rect 4264 5760 4292 5788
rect 4111 5732 4292 5760
rect 4111 5729 4123 5732
rect 4065 5723 4123 5729
rect 4614 5720 4620 5772
rect 4672 5760 4678 5772
rect 5123 5763 5181 5769
rect 4672 5732 5028 5760
rect 4672 5720 4678 5732
rect 1719 5664 1900 5692
rect 1949 5695 2007 5701
rect 1719 5661 1731 5664
rect 1673 5655 1731 5661
rect 1949 5661 1961 5695
rect 1995 5661 2007 5695
rect 1949 5655 2007 5661
rect 1596 5624 1624 5652
rect 1964 5624 1992 5655
rect 2958 5652 2964 5704
rect 3016 5652 3022 5704
rect 3786 5652 3792 5704
rect 3844 5652 3850 5704
rect 3973 5695 4031 5701
rect 3973 5661 3985 5695
rect 4019 5692 4031 5695
rect 4154 5692 4160 5704
rect 4019 5664 4160 5692
rect 4019 5661 4031 5664
rect 3973 5655 4031 5661
rect 4154 5652 4160 5664
rect 4212 5652 4218 5704
rect 5000 5701 5028 5732
rect 5123 5729 5135 5763
rect 5169 5760 5181 5763
rect 5920 5760 5948 5856
rect 6656 5828 6684 5856
rect 6564 5800 6684 5828
rect 9876 5828 9904 5856
rect 14461 5831 14519 5837
rect 14461 5828 14473 5831
rect 9876 5800 14473 5828
rect 6564 5769 6592 5800
rect 14461 5797 14473 5800
rect 14507 5797 14519 5831
rect 14461 5791 14519 5797
rect 5169 5732 5948 5760
rect 6549 5763 6607 5769
rect 5169 5729 5181 5732
rect 5123 5723 5181 5729
rect 6549 5729 6561 5763
rect 6595 5729 6607 5763
rect 6549 5723 6607 5729
rect 7558 5720 7564 5772
rect 7616 5760 7622 5772
rect 12526 5760 12532 5772
rect 7616 5732 12532 5760
rect 7616 5720 7622 5732
rect 4249 5695 4307 5701
rect 4249 5661 4261 5695
rect 4295 5661 4307 5695
rect 4249 5655 4307 5661
rect 4985 5695 5043 5701
rect 4985 5661 4997 5695
rect 5031 5661 5043 5695
rect 4985 5655 5043 5661
rect 1596 5596 1992 5624
rect 3804 5624 3832 5652
rect 4264 5624 4292 5655
rect 5258 5652 5264 5704
rect 5316 5652 5322 5704
rect 5905 5695 5963 5701
rect 5905 5661 5917 5695
rect 5951 5692 5963 5695
rect 6454 5692 6460 5704
rect 5951 5664 6460 5692
rect 5951 5661 5963 5664
rect 5905 5655 5963 5661
rect 6454 5652 6460 5664
rect 6512 5652 6518 5704
rect 6791 5695 6849 5701
rect 6791 5692 6803 5695
rect 6564 5664 6803 5692
rect 3804 5596 4292 5624
rect 6089 5627 6147 5633
rect 6089 5593 6101 5627
rect 6135 5624 6147 5627
rect 6270 5624 6276 5636
rect 6135 5596 6276 5624
rect 6135 5593 6147 5596
rect 6089 5587 6147 5593
rect 6270 5584 6276 5596
rect 6328 5584 6334 5636
rect 1578 5516 1584 5568
rect 1636 5556 1642 5568
rect 3605 5559 3663 5565
rect 3605 5556 3617 5559
rect 1636 5528 3617 5556
rect 1636 5516 1642 5528
rect 3605 5525 3617 5528
rect 3651 5525 3663 5559
rect 3605 5519 3663 5525
rect 3789 5559 3847 5565
rect 3789 5525 3801 5559
rect 3835 5556 3847 5559
rect 3970 5556 3976 5568
rect 3835 5528 3976 5556
rect 3835 5525 3847 5528
rect 3789 5519 3847 5525
rect 3970 5516 3976 5528
rect 4028 5516 4034 5568
rect 4614 5516 4620 5568
rect 4672 5556 4678 5568
rect 4890 5556 4896 5568
rect 4672 5528 4896 5556
rect 4672 5516 4678 5528
rect 4890 5516 4896 5528
rect 4948 5556 4954 5568
rect 6564 5556 6592 5664
rect 6791 5661 6803 5664
rect 6837 5661 6849 5695
rect 6791 5655 6849 5661
rect 8018 5652 8024 5704
rect 8076 5692 8082 5704
rect 8113 5695 8171 5701
rect 8113 5692 8125 5695
rect 8076 5664 8125 5692
rect 8076 5652 8082 5664
rect 8113 5661 8125 5664
rect 8159 5661 8171 5695
rect 8113 5655 8171 5661
rect 8202 5652 8208 5704
rect 8260 5692 8266 5704
rect 9766 5692 9772 5704
rect 8260 5664 9772 5692
rect 8260 5652 8266 5664
rect 9766 5652 9772 5664
rect 9824 5652 9830 5704
rect 10612 5701 10640 5732
rect 12526 5720 12532 5732
rect 12584 5720 12590 5772
rect 13817 5763 13875 5769
rect 13817 5729 13829 5763
rect 13863 5760 13875 5763
rect 13863 5732 14504 5760
rect 13863 5729 13875 5732
rect 13817 5723 13875 5729
rect 14476 5701 14504 5732
rect 14642 5720 14648 5772
rect 14700 5720 14706 5772
rect 15304 5760 15332 5856
rect 18322 5788 18328 5840
rect 18380 5788 18386 5840
rect 19061 5831 19119 5837
rect 19061 5797 19073 5831
rect 19107 5828 19119 5831
rect 19150 5828 19156 5840
rect 19107 5800 19156 5828
rect 19107 5797 19119 5800
rect 19061 5791 19119 5797
rect 19150 5788 19156 5800
rect 19208 5788 19214 5840
rect 14844 5732 15332 5760
rect 15580 5732 16068 5760
rect 14844 5701 14872 5732
rect 15580 5704 15608 5732
rect 10597 5695 10655 5701
rect 10597 5661 10609 5695
rect 10643 5692 10655 5695
rect 13725 5695 13783 5701
rect 10643 5664 10677 5692
rect 10643 5661 10655 5664
rect 10597 5655 10655 5661
rect 13725 5661 13737 5695
rect 13771 5661 13783 5695
rect 13725 5655 13783 5661
rect 14461 5695 14519 5701
rect 14461 5661 14473 5695
rect 14507 5661 14519 5695
rect 14461 5655 14519 5661
rect 14829 5695 14887 5701
rect 14829 5661 14841 5695
rect 14875 5661 14887 5695
rect 14829 5655 14887 5661
rect 12158 5624 12164 5636
rect 7024 5596 12164 5624
rect 4948 5528 6592 5556
rect 4948 5516 4954 5528
rect 6822 5516 6828 5568
rect 6880 5556 6886 5568
rect 7024 5556 7052 5596
rect 12158 5584 12164 5596
rect 12216 5584 12222 5636
rect 13740 5624 13768 5655
rect 14918 5652 14924 5704
rect 14976 5652 14982 5704
rect 15105 5695 15163 5701
rect 15105 5661 15117 5695
rect 15151 5692 15163 5695
rect 15151 5664 15424 5692
rect 15151 5661 15163 5664
rect 15105 5655 15163 5661
rect 15286 5624 15292 5636
rect 13740 5596 15292 5624
rect 15286 5584 15292 5596
rect 15344 5584 15350 5636
rect 6880 5528 7052 5556
rect 6880 5516 6886 5528
rect 7098 5516 7104 5568
rect 7156 5556 7162 5568
rect 7929 5559 7987 5565
rect 7929 5556 7941 5559
rect 7156 5528 7941 5556
rect 7156 5516 7162 5528
rect 7929 5525 7941 5528
rect 7975 5525 7987 5559
rect 7929 5519 7987 5525
rect 10410 5516 10416 5568
rect 10468 5516 10474 5568
rect 10686 5516 10692 5568
rect 10744 5556 10750 5568
rect 12710 5556 12716 5568
rect 10744 5528 12716 5556
rect 10744 5516 10750 5528
rect 12710 5516 12716 5528
rect 12768 5516 12774 5568
rect 13538 5516 13544 5568
rect 13596 5556 13602 5568
rect 14734 5556 14740 5568
rect 13596 5528 14740 5556
rect 13596 5516 13602 5528
rect 14734 5516 14740 5528
rect 14792 5516 14798 5568
rect 15396 5556 15424 5664
rect 15562 5652 15568 5704
rect 15620 5652 15626 5704
rect 15746 5652 15752 5704
rect 15804 5652 15810 5704
rect 15841 5695 15899 5701
rect 15841 5661 15853 5695
rect 15887 5692 15899 5695
rect 16040 5692 16068 5732
rect 16114 5720 16120 5772
rect 16172 5720 16178 5772
rect 17586 5720 17592 5772
rect 17644 5760 17650 5772
rect 17644 5732 18442 5760
rect 17644 5720 17650 5732
rect 16359 5695 16417 5701
rect 16359 5692 16371 5695
rect 15887 5664 15976 5692
rect 16040 5664 16371 5692
rect 15887 5661 15899 5664
rect 15841 5655 15899 5661
rect 15473 5627 15531 5633
rect 15473 5593 15485 5627
rect 15519 5624 15531 5627
rect 15654 5624 15660 5636
rect 15519 5596 15660 5624
rect 15519 5593 15531 5596
rect 15473 5587 15531 5593
rect 15654 5584 15660 5596
rect 15712 5584 15718 5636
rect 15948 5624 15976 5664
rect 16359 5661 16371 5664
rect 16405 5661 16417 5695
rect 17865 5695 17923 5701
rect 17865 5692 17877 5695
rect 16359 5655 16417 5661
rect 17144 5664 17877 5692
rect 17034 5624 17040 5636
rect 15948 5596 17040 5624
rect 17034 5584 17040 5596
rect 17092 5584 17098 5636
rect 16114 5556 16120 5568
rect 15396 5528 16120 5556
rect 16114 5516 16120 5528
rect 16172 5516 16178 5568
rect 16206 5516 16212 5568
rect 16264 5556 16270 5568
rect 17144 5556 17172 5664
rect 17865 5661 17877 5664
rect 17911 5661 17923 5695
rect 17865 5655 17923 5661
rect 18325 5695 18383 5701
rect 18325 5661 18337 5695
rect 18371 5661 18383 5695
rect 18325 5655 18383 5661
rect 17218 5584 17224 5636
rect 17276 5624 17282 5636
rect 18340 5624 18368 5655
rect 17276 5596 18368 5624
rect 17276 5584 17282 5596
rect 16264 5528 17172 5556
rect 18414 5556 18442 5732
rect 18506 5720 18512 5772
rect 18564 5760 18570 5772
rect 19245 5763 19303 5769
rect 19245 5760 19257 5763
rect 18564 5732 19257 5760
rect 18564 5720 18570 5732
rect 18800 5704 18828 5732
rect 19245 5729 19257 5732
rect 19291 5729 19303 5763
rect 19245 5723 19303 5729
rect 18782 5652 18788 5704
rect 18840 5652 18846 5704
rect 18874 5652 18880 5704
rect 18932 5652 18938 5704
rect 19487 5695 19545 5701
rect 19168 5692 19288 5694
rect 19487 5692 19499 5695
rect 18984 5666 19499 5692
rect 18984 5664 19196 5666
rect 19260 5664 19499 5666
rect 18690 5584 18696 5636
rect 18748 5624 18754 5636
rect 18984 5624 19012 5664
rect 19487 5661 19499 5664
rect 19533 5661 19545 5695
rect 19487 5655 19545 5661
rect 19978 5652 19984 5704
rect 20036 5692 20042 5704
rect 20824 5701 20852 5868
rect 21082 5856 21088 5908
rect 21140 5896 21146 5908
rect 21361 5899 21419 5905
rect 21361 5896 21373 5899
rect 21140 5868 21373 5896
rect 21140 5856 21146 5868
rect 21361 5865 21373 5868
rect 21407 5865 21419 5899
rect 21361 5859 21419 5865
rect 20990 5720 20996 5772
rect 21048 5760 21054 5772
rect 21048 5732 21128 5760
rect 21048 5720 21054 5732
rect 21100 5701 21128 5732
rect 20625 5695 20683 5701
rect 20625 5692 20637 5695
rect 20036 5664 20637 5692
rect 20036 5652 20042 5664
rect 20625 5661 20637 5664
rect 20671 5661 20683 5695
rect 20625 5655 20683 5661
rect 20809 5695 20867 5701
rect 20809 5661 20821 5695
rect 20855 5661 20867 5695
rect 20809 5655 20867 5661
rect 21085 5695 21143 5701
rect 21085 5661 21097 5695
rect 21131 5661 21143 5695
rect 21085 5655 21143 5661
rect 21358 5652 21364 5704
rect 21416 5692 21422 5704
rect 21545 5695 21603 5701
rect 21545 5692 21557 5695
rect 21416 5664 21557 5692
rect 21416 5652 21422 5664
rect 21545 5661 21557 5664
rect 21591 5661 21603 5695
rect 21545 5655 21603 5661
rect 18748 5596 19012 5624
rect 18748 5584 18754 5596
rect 19058 5584 19064 5636
rect 19116 5624 19122 5636
rect 19116 5596 20944 5624
rect 19116 5584 19122 5596
rect 20257 5559 20315 5565
rect 20257 5556 20269 5559
rect 18414 5528 20269 5556
rect 16264 5516 16270 5528
rect 20257 5525 20269 5528
rect 20303 5525 20315 5559
rect 20257 5519 20315 5525
rect 20806 5516 20812 5568
rect 20864 5516 20870 5568
rect 20916 5565 20944 5596
rect 20901 5559 20959 5565
rect 20901 5525 20913 5559
rect 20947 5525 20959 5559
rect 20901 5519 20959 5525
rect 1104 5466 22056 5488
rect 1104 5414 6148 5466
rect 6200 5414 6212 5466
rect 6264 5414 6276 5466
rect 6328 5414 6340 5466
rect 6392 5414 6404 5466
rect 6456 5414 11346 5466
rect 11398 5414 11410 5466
rect 11462 5414 11474 5466
rect 11526 5414 11538 5466
rect 11590 5414 11602 5466
rect 11654 5414 16544 5466
rect 16596 5414 16608 5466
rect 16660 5414 16672 5466
rect 16724 5414 16736 5466
rect 16788 5414 16800 5466
rect 16852 5414 21742 5466
rect 21794 5414 21806 5466
rect 21858 5414 21870 5466
rect 21922 5414 21934 5466
rect 21986 5414 21998 5466
rect 22050 5414 22056 5466
rect 1104 5392 22056 5414
rect 1762 5312 1768 5364
rect 1820 5312 1826 5364
rect 2038 5312 2044 5364
rect 2096 5312 2102 5364
rect 2314 5312 2320 5364
rect 2372 5352 2378 5364
rect 2682 5352 2688 5364
rect 2372 5324 2688 5352
rect 2372 5312 2378 5324
rect 2682 5312 2688 5324
rect 2740 5312 2746 5364
rect 3050 5312 3056 5364
rect 3108 5352 3114 5364
rect 3145 5355 3203 5361
rect 3145 5352 3157 5355
rect 3108 5324 3157 5352
rect 3108 5312 3114 5324
rect 3145 5321 3157 5324
rect 3191 5321 3203 5355
rect 3145 5315 3203 5321
rect 4525 5355 4583 5361
rect 4525 5321 4537 5355
rect 4571 5352 4583 5355
rect 5350 5352 5356 5364
rect 4571 5324 5356 5352
rect 4571 5321 4583 5324
rect 4525 5315 4583 5321
rect 5350 5312 5356 5324
rect 5408 5312 5414 5364
rect 8478 5352 8484 5364
rect 5460 5324 8484 5352
rect 1486 5244 1492 5296
rect 1544 5244 1550 5296
rect 2056 5284 2084 5312
rect 3878 5284 3884 5296
rect 2056 5256 3464 5284
rect 2407 5219 2465 5225
rect 2407 5185 2419 5219
rect 2453 5216 2465 5219
rect 3050 5216 3056 5228
rect 2453 5188 3056 5216
rect 2453 5185 2465 5188
rect 2407 5179 2465 5185
rect 3050 5176 3056 5188
rect 3108 5176 3114 5228
rect 2130 5108 2136 5160
rect 2188 5108 2194 5160
rect 1946 4972 1952 5024
rect 2004 5012 2010 5024
rect 2498 5012 2504 5024
rect 2004 4984 2504 5012
rect 2004 4972 2010 4984
rect 2498 4972 2504 4984
rect 2556 4972 2562 5024
rect 3436 5012 3464 5256
rect 3528 5256 3884 5284
rect 3528 5225 3556 5256
rect 3878 5244 3884 5256
rect 3936 5284 3942 5296
rect 4338 5284 4344 5296
rect 3936 5256 4344 5284
rect 3936 5244 3942 5256
rect 4338 5244 4344 5256
rect 4396 5284 4402 5296
rect 5460 5284 5488 5324
rect 8478 5312 8484 5324
rect 8536 5312 8542 5364
rect 12986 5352 12992 5364
rect 9140 5324 12992 5352
rect 9140 5284 9168 5324
rect 12986 5312 12992 5324
rect 13044 5312 13050 5364
rect 13909 5355 13967 5361
rect 13909 5321 13921 5355
rect 13955 5352 13967 5355
rect 14918 5352 14924 5364
rect 13955 5324 14924 5352
rect 13955 5321 13967 5324
rect 13909 5315 13967 5321
rect 14918 5312 14924 5324
rect 14976 5352 14982 5364
rect 15562 5352 15568 5364
rect 14976 5324 15568 5352
rect 14976 5312 14982 5324
rect 15562 5312 15568 5324
rect 15620 5312 15626 5364
rect 15657 5355 15715 5361
rect 15657 5321 15669 5355
rect 15703 5352 15715 5355
rect 15746 5352 15752 5364
rect 15703 5324 15752 5352
rect 15703 5321 15715 5324
rect 15657 5315 15715 5321
rect 15746 5312 15752 5324
rect 15804 5312 15810 5364
rect 15838 5312 15844 5364
rect 15896 5352 15902 5364
rect 16393 5355 16451 5361
rect 16393 5352 16405 5355
rect 15896 5324 16405 5352
rect 15896 5312 15902 5324
rect 16393 5321 16405 5324
rect 16439 5321 16451 5355
rect 16393 5315 16451 5321
rect 16574 5312 16580 5364
rect 16632 5352 16638 5364
rect 17586 5352 17592 5364
rect 16632 5324 17592 5352
rect 16632 5312 16638 5324
rect 17586 5312 17592 5324
rect 17644 5312 17650 5364
rect 17678 5312 17684 5364
rect 17736 5352 17742 5364
rect 17862 5352 17868 5364
rect 17736 5324 17868 5352
rect 17736 5312 17742 5324
rect 17862 5312 17868 5324
rect 17920 5312 17926 5364
rect 18138 5312 18144 5364
rect 18196 5352 18202 5364
rect 18506 5352 18512 5364
rect 18196 5324 18512 5352
rect 18196 5312 18202 5324
rect 18506 5312 18512 5324
rect 18564 5312 18570 5364
rect 18690 5312 18696 5364
rect 18748 5352 18754 5364
rect 19153 5355 19211 5361
rect 19153 5352 19165 5355
rect 18748 5324 19165 5352
rect 18748 5312 18754 5324
rect 19153 5321 19165 5324
rect 19199 5321 19211 5355
rect 19153 5315 19211 5321
rect 4396 5256 5488 5284
rect 5920 5256 9168 5284
rect 4396 5244 4402 5256
rect 5920 5228 5948 5256
rect 10042 5244 10048 5296
rect 10100 5284 10106 5296
rect 12434 5284 12440 5296
rect 10100 5256 12440 5284
rect 10100 5244 10106 5256
rect 12434 5244 12440 5256
rect 12492 5244 12498 5296
rect 14476 5256 16712 5284
rect 3513 5219 3571 5225
rect 3513 5185 3525 5219
rect 3559 5185 3571 5219
rect 3513 5179 3571 5185
rect 3787 5219 3845 5225
rect 3787 5185 3799 5219
rect 3833 5216 3845 5219
rect 4614 5216 4620 5228
rect 3833 5188 4620 5216
rect 3833 5185 3845 5188
rect 3787 5179 3845 5185
rect 4614 5176 4620 5188
rect 4672 5176 4678 5228
rect 5074 5176 5080 5228
rect 5132 5216 5138 5228
rect 5167 5219 5225 5225
rect 5167 5216 5179 5219
rect 5132 5188 5179 5216
rect 5132 5176 5138 5188
rect 5167 5185 5179 5188
rect 5213 5216 5225 5219
rect 5213 5188 5856 5216
rect 5213 5185 5225 5188
rect 5167 5179 5225 5185
rect 4890 5108 4896 5160
rect 4948 5108 4954 5160
rect 5828 5148 5856 5188
rect 5902 5176 5908 5228
rect 5960 5176 5966 5228
rect 5994 5176 6000 5228
rect 6052 5176 6058 5228
rect 6546 5176 6552 5228
rect 6604 5176 6610 5228
rect 6638 5176 6644 5228
rect 6696 5216 6702 5228
rect 12728 5216 12940 5220
rect 13171 5219 13229 5225
rect 13171 5216 13183 5219
rect 6696 5192 13183 5216
rect 6696 5188 12756 5192
rect 12912 5188 13183 5192
rect 6696 5176 6702 5188
rect 13171 5185 13183 5188
rect 13217 5216 13229 5219
rect 13217 5188 13584 5216
rect 13217 5185 13229 5188
rect 13171 5179 13229 5185
rect 6012 5148 6040 5176
rect 5828 5120 6040 5148
rect 5905 5083 5963 5089
rect 5905 5049 5917 5083
rect 5951 5080 5963 5083
rect 6564 5080 6592 5176
rect 6914 5108 6920 5160
rect 6972 5148 6978 5160
rect 11146 5148 11152 5160
rect 6972 5120 11152 5148
rect 6972 5108 6978 5120
rect 11146 5108 11152 5120
rect 11204 5108 11210 5160
rect 12894 5108 12900 5160
rect 12952 5108 12958 5160
rect 5951 5052 6592 5080
rect 5951 5049 5963 5052
rect 5905 5043 5963 5049
rect 10318 5012 10324 5024
rect 3436 4984 10324 5012
rect 10318 4972 10324 4984
rect 10376 4972 10382 5024
rect 13556 5012 13584 5188
rect 14274 5176 14280 5228
rect 14332 5216 14338 5228
rect 14476 5216 14504 5256
rect 14332 5188 14504 5216
rect 14544 5219 14602 5225
rect 14332 5176 14338 5188
rect 14544 5185 14556 5219
rect 14590 5216 14602 5219
rect 15930 5216 15936 5228
rect 14590 5188 15936 5216
rect 14590 5185 14602 5188
rect 14544 5179 14602 5185
rect 15930 5176 15936 5188
rect 15988 5176 15994 5228
rect 16025 5219 16083 5225
rect 16025 5185 16037 5219
rect 16071 5216 16083 5219
rect 16301 5219 16359 5225
rect 16071 5188 16252 5216
rect 16071 5185 16083 5188
rect 16025 5179 16083 5185
rect 16114 5108 16120 5160
rect 16172 5108 16178 5160
rect 16224 5080 16252 5188
rect 16301 5185 16313 5219
rect 16347 5185 16359 5219
rect 16301 5179 16359 5185
rect 16485 5219 16543 5225
rect 16485 5185 16497 5219
rect 16531 5185 16543 5219
rect 16485 5179 16543 5185
rect 15212 5052 16252 5080
rect 14458 5012 14464 5024
rect 13556 4984 14464 5012
rect 14458 4972 14464 4984
rect 14516 4972 14522 5024
rect 14642 4972 14648 5024
rect 14700 5012 14706 5024
rect 15212 5012 15240 5052
rect 14700 4984 15240 5012
rect 14700 4972 14706 4984
rect 15286 4972 15292 5024
rect 15344 5012 15350 5024
rect 15749 5015 15807 5021
rect 15749 5012 15761 5015
rect 15344 4984 15761 5012
rect 15344 4972 15350 4984
rect 15749 4981 15761 4984
rect 15795 4981 15807 5015
rect 15749 4975 15807 4981
rect 15838 4972 15844 5024
rect 15896 5012 15902 5024
rect 16316 5012 16344 5179
rect 16390 5108 16396 5160
rect 16448 5148 16454 5160
rect 16500 5148 16528 5179
rect 16684 5160 16712 5256
rect 18414 5255 18420 5296
rect 18399 5249 18420 5255
rect 16758 5176 16764 5228
rect 16816 5216 16822 5228
rect 16925 5219 16983 5225
rect 16925 5216 16937 5219
rect 16816 5188 16937 5216
rect 16816 5176 16822 5188
rect 16925 5185 16937 5188
rect 16971 5185 16983 5219
rect 18399 5215 18411 5249
rect 18472 5244 18478 5296
rect 20714 5244 20720 5296
rect 20772 5284 20778 5296
rect 21453 5287 21511 5293
rect 21453 5284 21465 5287
rect 20772 5256 21465 5284
rect 20772 5244 20778 5256
rect 21453 5253 21465 5256
rect 21499 5253 21511 5287
rect 21453 5247 21511 5253
rect 18445 5218 18460 5244
rect 19795 5219 19853 5225
rect 18445 5215 18457 5218
rect 18399 5209 18457 5215
rect 16925 5179 16983 5185
rect 19795 5185 19807 5219
rect 19841 5216 19853 5219
rect 20254 5216 20260 5228
rect 19841 5188 20260 5216
rect 19841 5185 19853 5188
rect 19795 5179 19853 5185
rect 20254 5176 20260 5188
rect 20312 5176 20318 5228
rect 20898 5176 20904 5228
rect 20956 5176 20962 5228
rect 21082 5176 21088 5228
rect 21140 5176 21146 5228
rect 21174 5176 21180 5228
rect 21232 5216 21238 5228
rect 21361 5219 21419 5225
rect 21361 5216 21373 5219
rect 21232 5188 21373 5216
rect 21232 5176 21238 5188
rect 21361 5185 21373 5188
rect 21407 5185 21419 5219
rect 21361 5179 21419 5185
rect 16448 5120 16528 5148
rect 16448 5108 16454 5120
rect 16666 5108 16672 5160
rect 16724 5108 16730 5160
rect 18141 5151 18199 5157
rect 18141 5117 18153 5151
rect 18187 5117 18199 5151
rect 18141 5111 18199 5117
rect 18156 5080 18184 5111
rect 19518 5108 19524 5160
rect 19576 5108 19582 5160
rect 18156 5052 18276 5080
rect 18248 5024 18276 5052
rect 15896 4984 16344 5012
rect 15896 4972 15902 4984
rect 17678 4972 17684 5024
rect 17736 5012 17742 5024
rect 18049 5015 18107 5021
rect 18049 5012 18061 5015
rect 17736 4984 18061 5012
rect 17736 4972 17742 4984
rect 18049 4981 18061 4984
rect 18095 4981 18107 5015
rect 18049 4975 18107 4981
rect 18230 4972 18236 5024
rect 18288 4972 18294 5024
rect 19058 4972 19064 5024
rect 19116 5012 19122 5024
rect 20533 5015 20591 5021
rect 20533 5012 20545 5015
rect 19116 4984 20545 5012
rect 19116 4972 19122 4984
rect 20533 4981 20545 4984
rect 20579 4981 20591 5015
rect 20533 4975 20591 4981
rect 1104 4922 21896 4944
rect 1104 4870 3549 4922
rect 3601 4870 3613 4922
rect 3665 4870 3677 4922
rect 3729 4870 3741 4922
rect 3793 4870 3805 4922
rect 3857 4870 8747 4922
rect 8799 4870 8811 4922
rect 8863 4870 8875 4922
rect 8927 4870 8939 4922
rect 8991 4870 9003 4922
rect 9055 4870 13945 4922
rect 13997 4870 14009 4922
rect 14061 4870 14073 4922
rect 14125 4870 14137 4922
rect 14189 4870 14201 4922
rect 14253 4870 19143 4922
rect 19195 4870 19207 4922
rect 19259 4870 19271 4922
rect 19323 4870 19335 4922
rect 19387 4870 19399 4922
rect 19451 4870 21896 4922
rect 1104 4848 21896 4870
rect 2133 4811 2191 4817
rect 2133 4777 2145 4811
rect 2179 4808 2191 4811
rect 3142 4808 3148 4820
rect 2179 4780 3148 4808
rect 2179 4777 2191 4780
rect 2133 4771 2191 4777
rect 3142 4768 3148 4780
rect 3200 4768 3206 4820
rect 3329 4811 3387 4817
rect 3329 4777 3341 4811
rect 3375 4808 3387 4811
rect 3375 4780 3648 4808
rect 3375 4777 3387 4780
rect 3329 4771 3387 4777
rect 3620 4752 3648 4780
rect 4706 4768 4712 4820
rect 4764 4768 4770 4820
rect 4798 4768 4804 4820
rect 4856 4808 4862 4820
rect 4893 4811 4951 4817
rect 4893 4808 4905 4811
rect 4856 4780 4905 4808
rect 4856 4768 4862 4780
rect 4893 4777 4905 4780
rect 4939 4777 4951 4811
rect 6273 4811 6331 4817
rect 6273 4808 6285 4811
rect 4893 4771 4951 4777
rect 5368 4780 6285 4808
rect 3602 4700 3608 4752
rect 3660 4700 3666 4752
rect 4724 4740 4752 4768
rect 5368 4740 5396 4780
rect 6273 4777 6285 4780
rect 6319 4777 6331 4811
rect 6273 4771 6331 4777
rect 12802 4768 12808 4820
rect 12860 4808 12866 4820
rect 15194 4808 15200 4820
rect 12860 4780 15200 4808
rect 12860 4768 12866 4780
rect 15194 4768 15200 4780
rect 15252 4768 15258 4820
rect 15657 4811 15715 4817
rect 15657 4777 15669 4811
rect 15703 4808 15715 4811
rect 16298 4808 16304 4820
rect 15703 4780 16304 4808
rect 15703 4777 15715 4780
rect 15657 4771 15715 4777
rect 16298 4768 16304 4780
rect 16356 4768 16362 4820
rect 16393 4811 16451 4817
rect 16393 4777 16405 4811
rect 16439 4808 16451 4811
rect 16850 4808 16856 4820
rect 16439 4780 16856 4808
rect 16439 4777 16451 4780
rect 16393 4771 16451 4777
rect 16850 4768 16856 4780
rect 16908 4768 16914 4820
rect 16945 4811 17003 4817
rect 16945 4777 16957 4811
rect 16991 4808 17003 4811
rect 17494 4808 17500 4820
rect 16991 4780 17500 4808
rect 16991 4777 17003 4780
rect 16945 4771 17003 4777
rect 17494 4768 17500 4780
rect 17552 4768 17558 4820
rect 18248 4780 19288 4808
rect 18248 4752 18276 4780
rect 4724 4712 5396 4740
rect 15565 4743 15623 4749
rect 15565 4709 15577 4743
rect 15611 4709 15623 4743
rect 15565 4703 15623 4709
rect 16209 4743 16267 4749
rect 16209 4709 16221 4743
rect 16255 4740 16267 4743
rect 16482 4740 16488 4752
rect 16255 4712 16488 4740
rect 16255 4709 16267 4712
rect 16209 4703 16267 4709
rect 2130 4632 2136 4684
rect 2188 4672 2194 4684
rect 2317 4675 2375 4681
rect 2317 4672 2329 4675
rect 2188 4644 2329 4672
rect 2188 4632 2194 4644
rect 2317 4641 2329 4644
rect 2363 4641 2375 4675
rect 2317 4635 2375 4641
rect 1578 4564 1584 4616
rect 1636 4564 1642 4616
rect 1854 4564 1860 4616
rect 1912 4564 1918 4616
rect 2332 4536 2360 4635
rect 3878 4632 3884 4684
rect 3936 4632 3942 4684
rect 2498 4564 2504 4616
rect 2556 4604 2562 4616
rect 2591 4607 2649 4613
rect 2591 4604 2603 4607
rect 2556 4576 2603 4604
rect 2556 4564 2562 4576
rect 2591 4573 2603 4576
rect 2637 4573 2649 4607
rect 2591 4567 2649 4573
rect 4155 4607 4213 4613
rect 4155 4573 4167 4607
rect 4201 4604 4213 4607
rect 5074 4604 5080 4616
rect 4201 4576 5080 4604
rect 4201 4573 4213 4576
rect 4155 4567 4213 4573
rect 5074 4564 5080 4576
rect 5132 4564 5138 4616
rect 5261 4607 5319 4613
rect 5261 4573 5273 4607
rect 5307 4573 5319 4607
rect 5261 4567 5319 4573
rect 5535 4607 5593 4613
rect 5535 4573 5547 4607
rect 5581 4604 5593 4607
rect 6822 4604 6828 4616
rect 5581 4576 6828 4604
rect 5581 4573 5593 4576
rect 5535 4567 5593 4573
rect 3786 4536 3792 4548
rect 2332 4508 3792 4536
rect 3786 4496 3792 4508
rect 3844 4536 3850 4548
rect 4338 4536 4344 4548
rect 3844 4508 4344 4536
rect 3844 4496 3850 4508
rect 4338 4496 4344 4508
rect 4396 4536 4402 4548
rect 5276 4536 5304 4567
rect 6822 4564 6828 4576
rect 6880 4564 6886 4616
rect 14185 4607 14243 4613
rect 14185 4573 14197 4607
rect 14231 4604 14243 4607
rect 14274 4604 14280 4616
rect 14231 4576 14280 4604
rect 14231 4573 14243 4576
rect 14185 4567 14243 4573
rect 14274 4564 14280 4576
rect 14332 4564 14338 4616
rect 14458 4613 14464 4616
rect 14441 4607 14464 4613
rect 14441 4573 14453 4607
rect 14441 4567 14464 4573
rect 14458 4564 14464 4567
rect 14516 4564 14522 4616
rect 15580 4604 15608 4703
rect 16482 4700 16488 4712
rect 16540 4700 16546 4752
rect 16577 4743 16635 4749
rect 16577 4709 16589 4743
rect 16623 4740 16635 4743
rect 17034 4740 17040 4752
rect 16623 4712 17040 4740
rect 16623 4709 16635 4712
rect 16577 4703 16635 4709
rect 17034 4700 17040 4712
rect 17092 4700 17098 4752
rect 18230 4700 18236 4752
rect 18288 4700 18294 4752
rect 19058 4740 19064 4752
rect 18892 4712 19064 4740
rect 16666 4672 16672 4684
rect 16224 4644 16672 4672
rect 16224 4616 16252 4644
rect 16666 4632 16672 4644
rect 16724 4672 16730 4684
rect 17129 4675 17187 4681
rect 17129 4672 17141 4675
rect 16724 4644 17141 4672
rect 16724 4632 16730 4644
rect 17129 4641 17141 4644
rect 17175 4641 17187 4675
rect 17129 4635 17187 4641
rect 15841 4607 15899 4613
rect 15841 4604 15853 4607
rect 15580 4576 15853 4604
rect 15841 4573 15853 4576
rect 15887 4573 15899 4607
rect 15841 4567 15899 4573
rect 15930 4564 15936 4616
rect 15988 4604 15994 4616
rect 16025 4607 16083 4613
rect 16025 4604 16037 4607
rect 15988 4576 16037 4604
rect 15988 4564 15994 4576
rect 16025 4573 16037 4576
rect 16071 4573 16083 4607
rect 16025 4567 16083 4573
rect 16206 4564 16212 4616
rect 16264 4564 16270 4616
rect 16301 4607 16359 4613
rect 16301 4573 16313 4607
rect 16347 4604 16359 4607
rect 16390 4604 16396 4616
rect 16347 4576 16396 4604
rect 16347 4573 16359 4576
rect 16301 4567 16359 4573
rect 16390 4564 16396 4576
rect 16448 4564 16454 4616
rect 16485 4607 16543 4613
rect 16485 4573 16497 4607
rect 16531 4573 16543 4607
rect 16485 4567 16543 4573
rect 4396 4508 5304 4536
rect 4396 4496 4402 4508
rect 5350 4496 5356 4548
rect 5408 4536 5414 4548
rect 7282 4536 7288 4548
rect 5408 4508 7288 4536
rect 5408 4496 5414 4508
rect 7282 4496 7288 4508
rect 7340 4496 7346 4548
rect 16500 4536 16528 4567
rect 16758 4564 16764 4616
rect 16816 4564 16822 4616
rect 16853 4607 16911 4613
rect 16853 4573 16865 4607
rect 16899 4573 16911 4607
rect 16853 4567 16911 4573
rect 16666 4536 16672 4548
rect 16500 4508 16672 4536
rect 16666 4496 16672 4508
rect 16724 4496 16730 4548
rect 1397 4471 1455 4477
rect 1397 4437 1409 4471
rect 1443 4468 1455 4471
rect 3418 4468 3424 4480
rect 1443 4440 3424 4468
rect 1443 4437 1455 4440
rect 1397 4431 1455 4437
rect 3418 4428 3424 4440
rect 3476 4428 3482 4480
rect 5166 4428 5172 4480
rect 5224 4468 5230 4480
rect 5534 4468 5540 4480
rect 5224 4440 5540 4468
rect 5224 4428 5230 4440
rect 5534 4428 5540 4440
rect 5592 4428 5598 4480
rect 10594 4428 10600 4480
rect 10652 4468 10658 4480
rect 14734 4468 14740 4480
rect 10652 4440 14740 4468
rect 10652 4428 10658 4440
rect 14734 4428 14740 4440
rect 14792 4428 14798 4480
rect 16298 4428 16304 4480
rect 16356 4468 16362 4480
rect 16776 4468 16804 4564
rect 16868 4536 16896 4567
rect 17034 4564 17040 4616
rect 17092 4564 17098 4616
rect 17218 4564 17224 4616
rect 17276 4564 17282 4616
rect 18892 4613 18920 4712
rect 19058 4700 19064 4712
rect 19116 4700 19122 4752
rect 19260 4749 19288 4780
rect 19518 4768 19524 4820
rect 19576 4808 19582 4820
rect 21174 4808 21180 4820
rect 19576 4780 21180 4808
rect 19576 4768 19582 4780
rect 21174 4768 21180 4780
rect 21232 4768 21238 4820
rect 19245 4743 19303 4749
rect 19245 4709 19257 4743
rect 19291 4740 19303 4743
rect 19291 4712 19656 4740
rect 19291 4709 19303 4712
rect 19245 4703 19303 4709
rect 19334 4672 19340 4684
rect 19076 4644 19340 4672
rect 19076 4613 19104 4644
rect 19334 4632 19340 4644
rect 19392 4632 19398 4684
rect 18785 4607 18843 4613
rect 18785 4604 18797 4607
rect 18524 4576 18797 4604
rect 17126 4536 17132 4548
rect 16868 4508 17132 4536
rect 17126 4496 17132 4508
rect 17184 4496 17190 4548
rect 16356 4440 16804 4468
rect 16356 4428 16362 4440
rect 16850 4428 16856 4480
rect 16908 4468 16914 4480
rect 17236 4468 17264 4564
rect 17396 4539 17454 4545
rect 17396 4505 17408 4539
rect 17442 4505 17454 4539
rect 17396 4499 17454 4505
rect 16908 4440 17264 4468
rect 17420 4468 17448 4499
rect 17494 4496 17500 4548
rect 17552 4536 17558 4548
rect 17862 4536 17868 4548
rect 17552 4508 17868 4536
rect 17552 4496 17558 4508
rect 17862 4496 17868 4508
rect 17920 4496 17926 4548
rect 17586 4468 17592 4480
rect 17420 4440 17592 4468
rect 16908 4428 16914 4440
rect 17586 4428 17592 4440
rect 17644 4428 17650 4480
rect 18524 4477 18552 4576
rect 18785 4573 18797 4576
rect 18831 4573 18843 4607
rect 18785 4567 18843 4573
rect 18877 4607 18935 4613
rect 18877 4573 18889 4607
rect 18923 4573 18935 4607
rect 18877 4567 18935 4573
rect 19061 4607 19119 4613
rect 19061 4573 19073 4607
rect 19107 4573 19119 4607
rect 19061 4567 19119 4573
rect 18509 4471 18567 4477
rect 18509 4437 18521 4471
rect 18555 4437 18567 4471
rect 18509 4431 18567 4437
rect 18598 4428 18604 4480
rect 18656 4428 18662 4480
rect 18892 4468 18920 4567
rect 19242 4564 19248 4616
rect 19300 4604 19306 4616
rect 19429 4607 19487 4613
rect 19429 4604 19441 4607
rect 19300 4576 19441 4604
rect 19300 4564 19306 4576
rect 19429 4573 19441 4576
rect 19475 4573 19487 4607
rect 19429 4567 19487 4573
rect 19518 4564 19524 4616
rect 19576 4564 19582 4616
rect 19628 4604 19656 4712
rect 19886 4632 19892 4684
rect 19944 4672 19950 4684
rect 19981 4675 20039 4681
rect 19981 4672 19993 4675
rect 19944 4644 19993 4672
rect 19944 4632 19950 4644
rect 19981 4641 19993 4644
rect 20027 4641 20039 4675
rect 19981 4635 20039 4641
rect 20237 4607 20295 4613
rect 20237 4604 20249 4607
rect 19628 4576 20249 4604
rect 20237 4573 20249 4576
rect 20283 4573 20295 4607
rect 20237 4567 20295 4573
rect 18969 4539 19027 4545
rect 18969 4505 18981 4539
rect 19015 4536 19027 4539
rect 19015 4508 19564 4536
rect 19015 4505 19027 4508
rect 18969 4499 19027 4505
rect 19536 4480 19564 4508
rect 19058 4468 19064 4480
rect 18892 4440 19064 4468
rect 19058 4428 19064 4440
rect 19116 4428 19122 4480
rect 19518 4428 19524 4480
rect 19576 4428 19582 4480
rect 19610 4428 19616 4480
rect 19668 4428 19674 4480
rect 21358 4428 21364 4480
rect 21416 4428 21422 4480
rect 1104 4378 22056 4400
rect 1104 4326 6148 4378
rect 6200 4326 6212 4378
rect 6264 4326 6276 4378
rect 6328 4326 6340 4378
rect 6392 4326 6404 4378
rect 6456 4326 11346 4378
rect 11398 4326 11410 4378
rect 11462 4326 11474 4378
rect 11526 4326 11538 4378
rect 11590 4326 11602 4378
rect 11654 4326 16544 4378
rect 16596 4326 16608 4378
rect 16660 4326 16672 4378
rect 16724 4326 16736 4378
rect 16788 4326 16800 4378
rect 16852 4326 21742 4378
rect 21794 4326 21806 4378
rect 21858 4326 21870 4378
rect 21922 4326 21934 4378
rect 21986 4326 21998 4378
rect 22050 4326 22056 4378
rect 1104 4304 22056 4326
rect 2593 4267 2651 4273
rect 2593 4233 2605 4267
rect 2639 4264 2651 4267
rect 2682 4264 2688 4276
rect 2639 4236 2688 4264
rect 2639 4233 2651 4236
rect 2593 4227 2651 4233
rect 2682 4224 2688 4236
rect 2740 4224 2746 4276
rect 3970 4264 3976 4276
rect 2792 4236 3976 4264
rect 1946 4156 1952 4208
rect 2004 4196 2010 4208
rect 2792 4196 2820 4236
rect 3970 4224 3976 4236
rect 4028 4224 4034 4276
rect 4798 4224 4804 4276
rect 4856 4264 4862 4276
rect 11974 4264 11980 4276
rect 4856 4236 11980 4264
rect 4856 4224 4862 4236
rect 11974 4224 11980 4236
rect 12032 4224 12038 4276
rect 14461 4267 14519 4273
rect 14461 4233 14473 4267
rect 14507 4264 14519 4267
rect 14642 4264 14648 4276
rect 14507 4236 14648 4264
rect 14507 4233 14519 4236
rect 14461 4227 14519 4233
rect 14642 4224 14648 4236
rect 14700 4224 14706 4276
rect 14826 4224 14832 4276
rect 14884 4224 14890 4276
rect 14921 4267 14979 4273
rect 14921 4233 14933 4267
rect 14967 4264 14979 4267
rect 15102 4264 15108 4276
rect 14967 4236 15108 4264
rect 14967 4233 14979 4236
rect 14921 4227 14979 4233
rect 15102 4224 15108 4236
rect 15160 4224 15166 4276
rect 15289 4267 15347 4273
rect 15289 4233 15301 4267
rect 15335 4264 15347 4267
rect 16022 4264 16028 4276
rect 15335 4236 16028 4264
rect 15335 4233 15347 4236
rect 15289 4227 15347 4233
rect 16022 4224 16028 4236
rect 16080 4224 16086 4276
rect 17218 4264 17224 4276
rect 16500 4236 17224 4264
rect 3050 4196 3056 4208
rect 2004 4168 2820 4196
rect 2976 4168 3056 4196
rect 2004 4156 2010 4168
rect 1855 4131 1913 4137
rect 1855 4097 1867 4131
rect 1901 4128 1913 4131
rect 2222 4128 2228 4140
rect 1901 4100 2228 4128
rect 1901 4097 1913 4100
rect 1855 4091 1913 4097
rect 2222 4088 2228 4100
rect 2280 4088 2286 4140
rect 2976 4137 3004 4168
rect 3050 4156 3056 4168
rect 3108 4196 3114 4208
rect 3108 4168 3924 4196
rect 3108 4156 3114 4168
rect 3896 4140 3924 4168
rect 4338 4156 4344 4208
rect 4396 4196 4402 4208
rect 5810 4196 5816 4208
rect 4396 4168 5816 4196
rect 4396 4156 4402 4168
rect 5810 4156 5816 4168
rect 5868 4156 5874 4208
rect 6086 4156 6092 4208
rect 6144 4196 6150 4208
rect 6730 4196 6736 4208
rect 6144 4168 6736 4196
rect 6144 4156 6150 4168
rect 6730 4156 6736 4168
rect 6788 4156 6794 4208
rect 13078 4196 13084 4208
rect 12820 4168 13084 4196
rect 2961 4131 3019 4137
rect 2961 4097 2973 4131
rect 3007 4097 3019 4131
rect 2961 4091 3019 4097
rect 3235 4131 3293 4137
rect 3235 4097 3247 4131
rect 3281 4128 3293 4131
rect 3694 4128 3700 4140
rect 3281 4100 3700 4128
rect 3281 4097 3293 4100
rect 3235 4091 3293 4097
rect 3694 4088 3700 4100
rect 3752 4088 3758 4140
rect 3878 4088 3884 4140
rect 3936 4088 3942 4140
rect 4154 4088 4160 4140
rect 4212 4128 4218 4140
rect 4583 4131 4641 4137
rect 4583 4128 4595 4131
rect 4212 4100 4595 4128
rect 4212 4088 4218 4100
rect 4583 4097 4595 4100
rect 4629 4097 4641 4131
rect 5442 4128 5448 4140
rect 4583 4091 4641 4097
rect 5184 4100 5448 4128
rect 1578 4020 1584 4072
rect 1636 4020 1642 4072
rect 3786 4020 3792 4072
rect 3844 4060 3850 4072
rect 4341 4063 4399 4069
rect 4341 4060 4353 4063
rect 3844 4032 4353 4060
rect 3844 4020 3850 4032
rect 4341 4029 4353 4032
rect 4387 4029 4399 4063
rect 4341 4023 4399 4029
rect 3234 3884 3240 3936
rect 3292 3924 3298 3936
rect 3973 3927 4031 3933
rect 3973 3924 3985 3927
rect 3292 3896 3985 3924
rect 3292 3884 3298 3896
rect 3973 3893 3985 3896
rect 4019 3893 4031 3927
rect 3973 3887 4031 3893
rect 4614 3884 4620 3936
rect 4672 3924 4678 3936
rect 5184 3924 5212 4100
rect 5442 4088 5448 4100
rect 5500 4088 5506 4140
rect 5718 4088 5724 4140
rect 5776 4128 5782 4140
rect 5905 4131 5963 4137
rect 5905 4128 5917 4131
rect 5776 4100 5917 4128
rect 5776 4088 5782 4100
rect 5905 4097 5917 4100
rect 5951 4097 5963 4131
rect 5905 4091 5963 4097
rect 6546 4088 6552 4140
rect 6604 4128 6610 4140
rect 12820 4128 12848 4168
rect 13078 4156 13084 4168
rect 13136 4156 13142 4208
rect 14844 4196 14872 4224
rect 16500 4196 16528 4236
rect 17218 4224 17224 4236
rect 17276 4224 17282 4276
rect 17678 4224 17684 4276
rect 17736 4224 17742 4276
rect 18046 4224 18052 4276
rect 18104 4264 18110 4276
rect 18104 4236 19104 4264
rect 18104 4224 18110 4236
rect 17586 4196 17592 4208
rect 14844 4168 16528 4196
rect 16592 4168 17592 4196
rect 16592 4140 16620 4168
rect 17586 4156 17592 4168
rect 17644 4156 17650 4208
rect 13814 4128 13820 4140
rect 6604 4100 12848 4128
rect 12912 4100 13820 4128
rect 6604 4088 6610 4100
rect 5258 4020 5264 4072
rect 5316 4020 5322 4072
rect 5810 4020 5816 4072
rect 5868 4060 5874 4072
rect 7834 4060 7840 4072
rect 5868 4032 7840 4060
rect 5868 4020 5874 4032
rect 7834 4020 7840 4032
rect 7892 4020 7898 4072
rect 4672 3896 5212 3924
rect 5276 3924 5304 4020
rect 5442 3952 5448 4004
rect 5500 3992 5506 4004
rect 12912 3992 12940 4100
rect 13814 4088 13820 4100
rect 13872 4088 13878 4140
rect 14366 4088 14372 4140
rect 14424 4088 14430 4140
rect 14645 4131 14703 4137
rect 14645 4097 14657 4131
rect 14691 4097 14703 4131
rect 14645 4091 14703 4097
rect 14458 4060 14464 4072
rect 5500 3964 12940 3992
rect 13004 4032 14464 4060
rect 5500 3952 5506 3964
rect 13004 3936 13032 4032
rect 14458 4020 14464 4032
rect 14516 4060 14522 4072
rect 14660 4060 14688 4091
rect 14918 4088 14924 4140
rect 14976 4128 14982 4140
rect 15105 4131 15163 4137
rect 15105 4128 15117 4131
rect 14976 4100 15117 4128
rect 14976 4088 14982 4100
rect 15105 4097 15117 4100
rect 15151 4097 15163 4131
rect 15105 4091 15163 4097
rect 15194 4088 15200 4140
rect 15252 4088 15258 4140
rect 15473 4131 15531 4137
rect 15473 4097 15485 4131
rect 15519 4097 15531 4131
rect 15473 4091 15531 4097
rect 14516 4032 14688 4060
rect 14516 4020 14522 4032
rect 15010 4020 15016 4072
rect 15068 4060 15074 4072
rect 15488 4060 15516 4091
rect 15562 4088 15568 4140
rect 15620 4088 15626 4140
rect 15933 4131 15991 4137
rect 15933 4097 15945 4131
rect 15979 4128 15991 4131
rect 16022 4128 16028 4140
rect 15979 4100 16028 4128
rect 15979 4097 15991 4100
rect 15933 4091 15991 4097
rect 16022 4088 16028 4100
rect 16080 4088 16086 4140
rect 16114 4088 16120 4140
rect 16172 4088 16178 4140
rect 16209 4131 16267 4137
rect 16209 4097 16221 4131
rect 16255 4097 16267 4131
rect 16209 4091 16267 4097
rect 16132 4060 16160 4088
rect 15068 4032 15516 4060
rect 15948 4032 16160 4060
rect 16224 4060 16252 4091
rect 16482 4088 16488 4140
rect 16540 4088 16546 4140
rect 16574 4088 16580 4140
rect 16632 4088 16638 4140
rect 17037 4131 17095 4137
rect 17037 4097 17049 4131
rect 17083 4128 17095 4131
rect 17218 4128 17224 4140
rect 17083 4100 17224 4128
rect 17083 4097 17095 4100
rect 17037 4091 17095 4097
rect 17218 4088 17224 4100
rect 17276 4088 17282 4140
rect 17313 4131 17371 4137
rect 17313 4097 17325 4131
rect 17359 4128 17371 4131
rect 17696 4128 17724 4224
rect 18156 4168 18552 4196
rect 17359 4100 17724 4128
rect 17359 4097 17371 4100
rect 17313 4091 17371 4097
rect 17862 4088 17868 4140
rect 17920 4088 17926 4140
rect 16758 4060 16764 4072
rect 16224 4032 16764 4060
rect 15068 4020 15074 4032
rect 14185 3995 14243 4001
rect 14185 3961 14197 3995
rect 14231 3992 14243 3995
rect 15948 3992 15976 4032
rect 16758 4020 16764 4032
rect 16816 4020 16822 4072
rect 17681 4063 17739 4069
rect 16868 4032 17632 4060
rect 14231 3964 15976 3992
rect 16025 3995 16083 4001
rect 14231 3961 14243 3964
rect 14185 3955 14243 3961
rect 16025 3961 16037 3995
rect 16071 3992 16083 3995
rect 16868 3992 16896 4032
rect 16071 3964 16896 3992
rect 16071 3961 16083 3964
rect 16025 3955 16083 3961
rect 16942 3952 16948 4004
rect 17000 3992 17006 4004
rect 17129 3995 17187 4001
rect 17129 3992 17141 3995
rect 17000 3964 17141 3992
rect 17000 3952 17006 3964
rect 17129 3961 17141 3964
rect 17175 3961 17187 3995
rect 17604 3992 17632 4032
rect 17681 4029 17693 4063
rect 17727 4060 17739 4063
rect 18156 4060 18184 4168
rect 18230 4088 18236 4140
rect 18288 4088 18294 4140
rect 18417 4131 18475 4137
rect 18417 4097 18429 4131
rect 18463 4097 18475 4131
rect 18524 4128 18552 4168
rect 18598 4156 18604 4208
rect 18656 4196 18662 4208
rect 19076 4196 19104 4236
rect 19150 4224 19156 4276
rect 19208 4224 19214 4276
rect 19334 4224 19340 4276
rect 19392 4264 19398 4276
rect 21085 4267 21143 4273
rect 21085 4264 21097 4267
rect 19392 4236 21097 4264
rect 19392 4224 19398 4236
rect 21085 4233 21097 4236
rect 21131 4233 21143 4267
rect 21085 4227 21143 4233
rect 19702 4196 19708 4208
rect 18656 4168 18920 4196
rect 19076 4168 19708 4196
rect 18656 4156 18662 4168
rect 18690 4128 18696 4140
rect 18524 4100 18696 4128
rect 18417 4091 18475 4097
rect 17727 4032 18184 4060
rect 17727 4029 17739 4032
rect 17681 4023 17739 4029
rect 18138 3992 18144 4004
rect 17604 3964 18144 3992
rect 17129 3955 17187 3961
rect 18138 3952 18144 3964
rect 18196 3952 18202 4004
rect 18248 3992 18276 4088
rect 18432 4060 18460 4091
rect 18690 4088 18696 4100
rect 18748 4088 18754 4140
rect 18892 4137 18920 4168
rect 19702 4156 19708 4168
rect 19760 4156 19766 4208
rect 19880 4199 19938 4205
rect 19880 4165 19892 4199
rect 19926 4196 19938 4199
rect 19978 4196 19984 4208
rect 19926 4168 19984 4196
rect 19926 4165 19938 4168
rect 19880 4159 19938 4165
rect 19978 4156 19984 4168
rect 20036 4156 20042 4208
rect 18877 4131 18935 4137
rect 18877 4097 18889 4131
rect 18923 4097 18935 4131
rect 18877 4091 18935 4097
rect 18966 4088 18972 4140
rect 19024 4088 19030 4140
rect 19429 4131 19487 4137
rect 19429 4097 19441 4131
rect 19475 4128 19487 4131
rect 21082 4128 21088 4140
rect 19475 4100 21088 4128
rect 19475 4097 19487 4100
rect 19429 4091 19487 4097
rect 21082 4088 21088 4100
rect 21140 4088 21146 4140
rect 21266 4088 21272 4140
rect 21324 4088 21330 4140
rect 21545 4131 21603 4137
rect 21545 4097 21557 4131
rect 21591 4097 21603 4131
rect 21545 4091 21603 4097
rect 18785 4063 18843 4069
rect 18785 4060 18797 4063
rect 18432 4032 18797 4060
rect 18785 4029 18797 4032
rect 18831 4029 18843 4063
rect 18785 4023 18843 4029
rect 19613 4063 19671 4069
rect 19613 4029 19625 4063
rect 19659 4029 19671 4063
rect 19613 4023 19671 4029
rect 18325 3995 18383 4001
rect 18325 3992 18337 3995
rect 18248 3964 18337 3992
rect 18325 3961 18337 3964
rect 18371 3961 18383 3995
rect 18325 3955 18383 3961
rect 18414 3952 18420 4004
rect 18472 3992 18478 4004
rect 19245 3995 19303 4001
rect 19245 3992 19257 3995
rect 18472 3964 19257 3992
rect 18472 3952 18478 3964
rect 19245 3961 19257 3964
rect 19291 3961 19303 3995
rect 19245 3955 19303 3961
rect 5353 3927 5411 3933
rect 5353 3924 5365 3927
rect 5276 3896 5365 3924
rect 4672 3884 4678 3896
rect 5353 3893 5365 3896
rect 5399 3893 5411 3927
rect 5353 3887 5411 3893
rect 5718 3884 5724 3936
rect 5776 3884 5782 3936
rect 6730 3884 6736 3936
rect 6788 3924 6794 3936
rect 9674 3924 9680 3936
rect 6788 3896 9680 3924
rect 6788 3884 6794 3896
rect 9674 3884 9680 3896
rect 9732 3884 9738 3936
rect 12986 3884 12992 3936
rect 13044 3884 13050 3936
rect 15746 3884 15752 3936
rect 15804 3884 15810 3936
rect 16298 3884 16304 3936
rect 16356 3884 16362 3936
rect 16853 3927 16911 3933
rect 16853 3893 16865 3927
rect 16899 3924 16911 3927
rect 18782 3924 18788 3936
rect 16899 3896 18788 3924
rect 16899 3893 16911 3896
rect 16853 3887 16911 3893
rect 18782 3884 18788 3896
rect 18840 3884 18846 3936
rect 19628 3924 19656 4023
rect 21560 3992 21588 4091
rect 20548 3964 21588 3992
rect 19886 3924 19892 3936
rect 19628 3896 19892 3924
rect 19886 3884 19892 3896
rect 19944 3884 19950 3936
rect 20254 3884 20260 3936
rect 20312 3924 20318 3936
rect 20548 3924 20576 3964
rect 20312 3896 20576 3924
rect 20312 3884 20318 3896
rect 20990 3884 20996 3936
rect 21048 3884 21054 3936
rect 21358 3884 21364 3936
rect 21416 3884 21422 3936
rect 1104 3834 21896 3856
rect 1104 3782 3549 3834
rect 3601 3782 3613 3834
rect 3665 3782 3677 3834
rect 3729 3782 3741 3834
rect 3793 3782 3805 3834
rect 3857 3782 8747 3834
rect 8799 3782 8811 3834
rect 8863 3782 8875 3834
rect 8927 3782 8939 3834
rect 8991 3782 9003 3834
rect 9055 3782 13945 3834
rect 13997 3782 14009 3834
rect 14061 3782 14073 3834
rect 14125 3782 14137 3834
rect 14189 3782 14201 3834
rect 14253 3782 19143 3834
rect 19195 3782 19207 3834
rect 19259 3782 19271 3834
rect 19323 3782 19335 3834
rect 19387 3782 19399 3834
rect 19451 3782 21896 3834
rect 1104 3760 21896 3782
rect 2593 3723 2651 3729
rect 2593 3689 2605 3723
rect 2639 3720 2651 3723
rect 2866 3720 2872 3732
rect 2639 3692 2872 3720
rect 2639 3689 2651 3692
rect 2593 3683 2651 3689
rect 2866 3680 2872 3692
rect 2924 3680 2930 3732
rect 3326 3680 3332 3732
rect 3384 3680 3390 3732
rect 5537 3723 5595 3729
rect 3804 3692 4844 3720
rect 2406 3612 2412 3664
rect 2464 3652 2470 3664
rect 3804 3652 3832 3692
rect 4816 3661 4844 3692
rect 5537 3689 5549 3723
rect 5583 3720 5595 3723
rect 5626 3720 5632 3732
rect 5583 3692 5632 3720
rect 5583 3689 5595 3692
rect 5537 3683 5595 3689
rect 5626 3680 5632 3692
rect 5684 3680 5690 3732
rect 5721 3723 5779 3729
rect 5721 3689 5733 3723
rect 5767 3689 5779 3723
rect 5721 3683 5779 3689
rect 8941 3723 8999 3729
rect 8941 3689 8953 3723
rect 8987 3720 8999 3723
rect 11606 3720 11612 3732
rect 8987 3692 11612 3720
rect 8987 3689 8999 3692
rect 8941 3683 8999 3689
rect 2464 3624 3832 3652
rect 4801 3655 4859 3661
rect 2464 3612 2470 3624
rect 4801 3621 4813 3655
rect 4847 3621 4859 3655
rect 4801 3615 4859 3621
rect 1578 3544 1584 3596
rect 1636 3544 1642 3596
rect 3786 3544 3792 3596
rect 3844 3544 3850 3596
rect 5626 3544 5632 3596
rect 5684 3584 5690 3596
rect 5736 3584 5764 3683
rect 11606 3680 11612 3692
rect 11664 3680 11670 3732
rect 11790 3680 11796 3732
rect 11848 3680 11854 3732
rect 14645 3723 14703 3729
rect 14645 3689 14657 3723
rect 14691 3720 14703 3723
rect 15194 3720 15200 3732
rect 14691 3692 15200 3720
rect 14691 3689 14703 3692
rect 14645 3683 14703 3689
rect 15194 3680 15200 3692
rect 15252 3680 15258 3732
rect 16390 3720 16396 3732
rect 15396 3692 16396 3720
rect 11808 3652 11836 3680
rect 13170 3652 13176 3664
rect 5684 3556 5764 3584
rect 5828 3624 11836 3652
rect 11900 3624 13176 3652
rect 5684 3544 5690 3556
rect 474 3476 480 3528
rect 532 3516 538 3528
rect 1823 3519 1881 3525
rect 1823 3516 1835 3519
rect 532 3488 1835 3516
rect 532 3476 538 3488
rect 1823 3485 1835 3488
rect 1869 3485 1881 3519
rect 5261 3519 5319 3525
rect 1823 3479 1881 3485
rect 2746 3489 4108 3516
rect 2746 3488 4059 3489
rect 1026 3408 1032 3460
rect 1084 3448 1090 3460
rect 2746 3448 2774 3488
rect 1084 3420 2774 3448
rect 1084 3408 1090 3420
rect 3234 3408 3240 3460
rect 3292 3408 3298 3460
rect 4047 3455 4059 3488
rect 4093 3458 4108 3489
rect 5261 3485 5273 3519
rect 5307 3516 5319 3519
rect 5828 3516 5856 3624
rect 6730 3544 6736 3596
rect 6788 3544 6794 3596
rect 6914 3544 6920 3596
rect 6972 3584 6978 3596
rect 7190 3584 7196 3596
rect 6972 3556 7196 3584
rect 6972 3544 6978 3556
rect 7190 3544 7196 3556
rect 7248 3544 7254 3596
rect 8662 3544 8668 3596
rect 8720 3584 8726 3596
rect 8720 3556 9168 3584
rect 8720 3544 8726 3556
rect 5307 3488 5856 3516
rect 5307 3485 5319 3488
rect 5261 3479 5319 3485
rect 5902 3476 5908 3528
rect 5960 3476 5966 3528
rect 4093 3455 4105 3458
rect 4047 3449 4105 3455
rect 6748 3448 6776 3544
rect 7650 3476 7656 3528
rect 7708 3476 7714 3528
rect 7742 3476 7748 3528
rect 7800 3516 7806 3528
rect 8021 3519 8079 3525
rect 8021 3516 8033 3519
rect 7800 3488 8033 3516
rect 7800 3476 7806 3488
rect 8021 3485 8033 3488
rect 8067 3485 8079 3519
rect 8021 3479 8079 3485
rect 8481 3519 8539 3525
rect 8481 3485 8493 3519
rect 8527 3485 8539 3519
rect 8481 3479 8539 3485
rect 7006 3448 7012 3460
rect 4172 3420 6776 3448
rect 6840 3420 7012 3448
rect 3142 3340 3148 3392
rect 3200 3380 3206 3392
rect 4172 3380 4200 3420
rect 3200 3352 4200 3380
rect 3200 3340 3206 3352
rect 4430 3340 4436 3392
rect 4488 3380 4494 3392
rect 6840 3380 6868 3420
rect 7006 3408 7012 3420
rect 7064 3408 7070 3460
rect 8496 3448 8524 3479
rect 8754 3476 8760 3528
rect 8812 3476 8818 3528
rect 9140 3525 9168 3556
rect 9766 3544 9772 3596
rect 9824 3584 9830 3596
rect 11900 3584 11928 3624
rect 13170 3612 13176 3624
rect 13228 3612 13234 3664
rect 13357 3655 13415 3661
rect 13357 3621 13369 3655
rect 13403 3652 13415 3655
rect 13722 3652 13728 3664
rect 13403 3624 13728 3652
rect 13403 3621 13415 3624
rect 13357 3615 13415 3621
rect 13722 3612 13728 3624
rect 13780 3612 13786 3664
rect 14277 3655 14335 3661
rect 14277 3621 14289 3655
rect 14323 3621 14335 3655
rect 14277 3615 14335 3621
rect 14369 3655 14427 3661
rect 14369 3621 14381 3655
rect 14415 3652 14427 3655
rect 15396 3652 15424 3692
rect 16390 3680 16396 3692
rect 16448 3680 16454 3732
rect 17681 3723 17739 3729
rect 17681 3689 17693 3723
rect 17727 3720 17739 3723
rect 17862 3720 17868 3732
rect 17727 3692 17868 3720
rect 17727 3689 17739 3692
rect 17681 3683 17739 3689
rect 17862 3680 17868 3692
rect 17920 3680 17926 3732
rect 18414 3680 18420 3732
rect 18472 3680 18478 3732
rect 18506 3680 18512 3732
rect 18564 3680 18570 3732
rect 18782 3680 18788 3732
rect 18840 3720 18846 3732
rect 20438 3720 20444 3732
rect 18840 3692 20444 3720
rect 18840 3680 18846 3692
rect 20438 3680 20444 3692
rect 20496 3680 20502 3732
rect 20625 3723 20683 3729
rect 20625 3689 20637 3723
rect 20671 3720 20683 3723
rect 21266 3720 21272 3732
rect 20671 3692 21272 3720
rect 20671 3689 20683 3692
rect 20625 3683 20683 3689
rect 21266 3680 21272 3692
rect 21324 3680 21330 3732
rect 22646 3680 22652 3732
rect 22704 3680 22710 3732
rect 14415 3624 15424 3652
rect 14415 3621 14427 3624
rect 14369 3615 14427 3621
rect 12618 3584 12624 3596
rect 9824 3556 11928 3584
rect 12406 3556 12624 3584
rect 9824 3544 9830 3556
rect 9125 3519 9183 3525
rect 9125 3485 9137 3519
rect 9171 3485 9183 3519
rect 9125 3479 9183 3485
rect 9398 3476 9404 3528
rect 9456 3516 9462 3528
rect 9677 3519 9735 3525
rect 9677 3516 9689 3519
rect 9456 3488 9689 3516
rect 9456 3476 9462 3488
rect 9677 3485 9689 3488
rect 9723 3485 9735 3519
rect 9677 3479 9735 3485
rect 10045 3519 10103 3525
rect 10045 3485 10057 3519
rect 10091 3516 10103 3519
rect 12406 3516 12434 3556
rect 12618 3544 12624 3556
rect 12676 3544 12682 3596
rect 14292 3584 14320 3615
rect 15838 3612 15844 3664
rect 15896 3652 15902 3664
rect 16761 3655 16819 3661
rect 16761 3652 16773 3655
rect 15896 3624 16773 3652
rect 15896 3612 15902 3624
rect 16761 3621 16773 3624
rect 16807 3621 16819 3655
rect 17402 3652 17408 3664
rect 16761 3615 16819 3621
rect 16868 3624 17408 3652
rect 16574 3584 16580 3596
rect 14292 3556 16580 3584
rect 16574 3544 16580 3556
rect 16632 3544 16638 3596
rect 16868 3584 16896 3624
rect 17402 3612 17408 3624
rect 17460 3612 17466 3664
rect 17310 3584 17316 3596
rect 16684 3556 16896 3584
rect 16960 3556 17316 3584
rect 10091 3488 12434 3516
rect 13081 3519 13139 3525
rect 10091 3485 10103 3488
rect 10045 3479 10103 3485
rect 13081 3485 13093 3519
rect 13127 3516 13139 3519
rect 13446 3516 13452 3528
rect 13127 3488 13452 3516
rect 13127 3485 13139 3488
rect 13081 3479 13139 3485
rect 13446 3476 13452 3488
rect 13504 3476 13510 3528
rect 13541 3519 13599 3525
rect 13541 3485 13553 3519
rect 13587 3516 13599 3519
rect 13814 3516 13820 3528
rect 13587 3488 13820 3516
rect 13587 3485 13599 3488
rect 13541 3479 13599 3485
rect 13814 3476 13820 3488
rect 13872 3476 13878 3528
rect 13909 3519 13967 3525
rect 13909 3485 13921 3519
rect 13955 3485 13967 3519
rect 13909 3479 13967 3485
rect 14093 3519 14151 3525
rect 14093 3485 14105 3519
rect 14139 3516 14151 3519
rect 14458 3516 14464 3528
rect 14139 3488 14464 3516
rect 14139 3485 14151 3488
rect 14093 3479 14151 3485
rect 9306 3448 9312 3460
rect 8496 3420 9312 3448
rect 9306 3408 9312 3420
rect 9364 3408 9370 3460
rect 13924 3448 13952 3479
rect 14458 3476 14464 3488
rect 14516 3476 14522 3528
rect 14553 3519 14611 3525
rect 14553 3485 14565 3519
rect 14599 3516 14611 3519
rect 14734 3516 14740 3528
rect 14599 3488 14740 3516
rect 14599 3485 14611 3488
rect 14553 3479 14611 3485
rect 14734 3476 14740 3488
rect 14792 3476 14798 3528
rect 14826 3476 14832 3528
rect 14884 3476 14890 3528
rect 15102 3476 15108 3528
rect 15160 3476 15166 3528
rect 15194 3476 15200 3528
rect 15252 3476 15258 3528
rect 15381 3519 15439 3525
rect 15381 3485 15393 3519
rect 15427 3516 15439 3519
rect 15562 3516 15568 3528
rect 15427 3488 15568 3516
rect 15427 3485 15439 3488
rect 15381 3479 15439 3485
rect 15562 3476 15568 3488
rect 15620 3476 15626 3528
rect 15654 3476 15660 3528
rect 15712 3476 15718 3528
rect 15930 3476 15936 3528
rect 15988 3516 15994 3528
rect 16482 3516 16488 3528
rect 15988 3488 16488 3516
rect 15988 3476 15994 3488
rect 16482 3476 16488 3488
rect 16540 3476 16546 3528
rect 16684 3525 16712 3556
rect 16960 3525 16988 3556
rect 17310 3544 17316 3556
rect 17368 3544 17374 3596
rect 17770 3584 17776 3596
rect 17512 3556 17776 3584
rect 16669 3519 16727 3525
rect 16669 3485 16681 3519
rect 16715 3485 16727 3519
rect 16669 3479 16727 3485
rect 16945 3519 17003 3525
rect 16945 3485 16957 3519
rect 16991 3485 17003 3519
rect 16945 3479 17003 3485
rect 17221 3519 17279 3525
rect 17221 3485 17233 3519
rect 17267 3516 17279 3519
rect 17402 3516 17408 3528
rect 17267 3488 17408 3516
rect 17267 3485 17279 3488
rect 17221 3479 17279 3485
rect 17402 3476 17408 3488
rect 17460 3476 17466 3528
rect 17512 3525 17540 3556
rect 17770 3544 17776 3556
rect 17828 3544 17834 3596
rect 17862 3544 17868 3596
rect 17920 3584 17926 3596
rect 17920 3556 18092 3584
rect 17920 3544 17926 3556
rect 18064 3525 18092 3556
rect 17497 3519 17555 3525
rect 17497 3485 17509 3519
rect 17543 3485 17555 3519
rect 17497 3479 17555 3485
rect 17589 3519 17647 3525
rect 17589 3485 17601 3519
rect 17635 3516 17647 3519
rect 18049 3519 18107 3525
rect 17635 3488 17908 3516
rect 17635 3485 17647 3488
rect 17589 3479 17647 3485
rect 14642 3448 14648 3460
rect 11624 3420 13860 3448
rect 13924 3420 14648 3448
rect 11624 3392 11652 3420
rect 4488 3352 6868 3380
rect 4488 3340 4494 3352
rect 6914 3340 6920 3392
rect 6972 3380 6978 3392
rect 7469 3383 7527 3389
rect 7469 3380 7481 3383
rect 6972 3352 7481 3380
rect 6972 3340 6978 3352
rect 7469 3349 7481 3352
rect 7515 3349 7527 3383
rect 7469 3343 7527 3349
rect 7558 3340 7564 3392
rect 7616 3380 7622 3392
rect 7837 3383 7895 3389
rect 7837 3380 7849 3383
rect 7616 3352 7849 3380
rect 7616 3340 7622 3352
rect 7837 3349 7849 3352
rect 7883 3349 7895 3383
rect 7837 3343 7895 3349
rect 8294 3340 8300 3392
rect 8352 3340 8358 3392
rect 8570 3340 8576 3392
rect 8628 3340 8634 3392
rect 9214 3340 9220 3392
rect 9272 3340 9278 3392
rect 9858 3340 9864 3392
rect 9916 3340 9922 3392
rect 11606 3340 11612 3392
rect 11664 3340 11670 3392
rect 12894 3340 12900 3392
rect 12952 3340 12958 3392
rect 13446 3340 13452 3392
rect 13504 3380 13510 3392
rect 13725 3383 13783 3389
rect 13725 3380 13737 3383
rect 13504 3352 13737 3380
rect 13504 3340 13510 3352
rect 13725 3349 13737 3352
rect 13771 3349 13783 3383
rect 13832 3380 13860 3420
rect 14642 3408 14648 3420
rect 14700 3408 14706 3460
rect 15212 3448 15240 3476
rect 14752 3420 15240 3448
rect 14458 3380 14464 3392
rect 13832 3352 14464 3380
rect 13725 3343 13783 3349
rect 14458 3340 14464 3352
rect 14516 3340 14522 3392
rect 14550 3340 14556 3392
rect 14608 3380 14614 3392
rect 14752 3380 14780 3420
rect 15286 3408 15292 3460
rect 15344 3448 15350 3460
rect 16025 3451 16083 3457
rect 15344 3420 15884 3448
rect 15344 3408 15350 3420
rect 14608 3352 14780 3380
rect 14608 3340 14614 3352
rect 14918 3340 14924 3392
rect 14976 3340 14982 3392
rect 15194 3340 15200 3392
rect 15252 3340 15258 3392
rect 15473 3383 15531 3389
rect 15473 3349 15485 3383
rect 15519 3380 15531 3383
rect 15746 3380 15752 3392
rect 15519 3352 15752 3380
rect 15519 3349 15531 3352
rect 15473 3343 15531 3349
rect 15746 3340 15752 3352
rect 15804 3340 15810 3392
rect 15856 3380 15884 3420
rect 16025 3417 16037 3451
rect 16071 3448 16083 3451
rect 16071 3420 17356 3448
rect 16071 3417 16083 3420
rect 16025 3411 16083 3417
rect 16117 3383 16175 3389
rect 16117 3380 16129 3383
rect 15856 3352 16129 3380
rect 16117 3349 16129 3352
rect 16163 3349 16175 3383
rect 16117 3343 16175 3349
rect 16390 3340 16396 3392
rect 16448 3380 16454 3392
rect 16485 3383 16543 3389
rect 16485 3380 16497 3383
rect 16448 3352 16497 3380
rect 16448 3340 16454 3352
rect 16485 3349 16497 3352
rect 16531 3349 16543 3383
rect 16485 3343 16543 3349
rect 16758 3340 16764 3392
rect 16816 3380 16822 3392
rect 17328 3389 17356 3420
rect 17880 3389 17908 3488
rect 18049 3485 18061 3519
rect 18095 3485 18107 3519
rect 18049 3479 18107 3485
rect 18322 3476 18328 3528
rect 18380 3476 18386 3528
rect 18432 3448 18460 3680
rect 18524 3652 18552 3680
rect 18877 3655 18935 3661
rect 18877 3652 18889 3655
rect 18524 3624 18889 3652
rect 18877 3621 18889 3624
rect 18923 3621 18935 3655
rect 18877 3615 18935 3621
rect 21361 3655 21419 3661
rect 21361 3621 21373 3655
rect 21407 3652 21419 3655
rect 22664 3652 22692 3680
rect 21407 3624 22692 3652
rect 21407 3621 21419 3624
rect 21361 3615 21419 3621
rect 20993 3587 21051 3593
rect 20993 3553 21005 3587
rect 21039 3584 21051 3587
rect 22462 3584 22468 3596
rect 21039 3556 22468 3584
rect 21039 3553 21051 3556
rect 20993 3547 21051 3553
rect 22462 3544 22468 3556
rect 22520 3544 22526 3596
rect 18598 3476 18604 3528
rect 18656 3476 18662 3528
rect 18690 3476 18696 3528
rect 18748 3476 18754 3528
rect 19245 3519 19303 3525
rect 19245 3485 19257 3519
rect 19291 3516 19303 3519
rect 19886 3516 19892 3528
rect 19291 3488 19892 3516
rect 19291 3485 19303 3488
rect 19245 3479 19303 3485
rect 19886 3476 19892 3488
rect 19944 3476 19950 3528
rect 20714 3476 20720 3528
rect 20772 3516 20778 3528
rect 20809 3519 20867 3525
rect 20809 3516 20821 3519
rect 20772 3488 20821 3516
rect 20772 3476 20778 3488
rect 20809 3485 20821 3488
rect 20855 3485 20867 3519
rect 20809 3479 20867 3485
rect 19490 3451 19548 3457
rect 19490 3448 19502 3451
rect 18432 3420 19502 3448
rect 19490 3417 19502 3420
rect 19536 3417 19548 3451
rect 19490 3411 19548 3417
rect 21177 3451 21235 3457
rect 21177 3417 21189 3451
rect 21223 3448 21235 3451
rect 21542 3448 21548 3460
rect 21223 3420 21548 3448
rect 21223 3417 21235 3420
rect 21177 3411 21235 3417
rect 21542 3408 21548 3420
rect 21600 3408 21606 3460
rect 17037 3383 17095 3389
rect 17037 3380 17049 3383
rect 16816 3352 17049 3380
rect 16816 3340 16822 3352
rect 17037 3349 17049 3352
rect 17083 3349 17095 3383
rect 17037 3343 17095 3349
rect 17313 3383 17371 3389
rect 17313 3349 17325 3383
rect 17359 3349 17371 3383
rect 17313 3343 17371 3349
rect 17865 3383 17923 3389
rect 17865 3349 17877 3383
rect 17911 3349 17923 3383
rect 17865 3343 17923 3349
rect 18046 3340 18052 3392
rect 18104 3380 18110 3392
rect 18141 3383 18199 3389
rect 18141 3380 18153 3383
rect 18104 3352 18153 3380
rect 18104 3340 18110 3352
rect 18141 3349 18153 3352
rect 18187 3349 18199 3383
rect 18141 3343 18199 3349
rect 18414 3340 18420 3392
rect 18472 3380 18478 3392
rect 19978 3380 19984 3392
rect 18472 3352 19984 3380
rect 18472 3340 18478 3352
rect 19978 3340 19984 3352
rect 20036 3340 20042 3392
rect 20898 3340 20904 3392
rect 20956 3380 20962 3392
rect 22554 3380 22560 3392
rect 20956 3352 22560 3380
rect 20956 3340 20962 3352
rect 22554 3340 22560 3352
rect 22612 3340 22618 3392
rect 1104 3290 22056 3312
rect 1104 3238 6148 3290
rect 6200 3238 6212 3290
rect 6264 3238 6276 3290
rect 6328 3238 6340 3290
rect 6392 3238 6404 3290
rect 6456 3238 11346 3290
rect 11398 3238 11410 3290
rect 11462 3238 11474 3290
rect 11526 3238 11538 3290
rect 11590 3238 11602 3290
rect 11654 3238 16544 3290
rect 16596 3238 16608 3290
rect 16660 3238 16672 3290
rect 16724 3238 16736 3290
rect 16788 3238 16800 3290
rect 16852 3238 21742 3290
rect 21794 3238 21806 3290
rect 21858 3238 21870 3290
rect 21922 3238 21934 3290
rect 21986 3238 21998 3290
rect 22050 3238 22056 3290
rect 1104 3216 22056 3238
rect 1578 3136 1584 3188
rect 1636 3176 1642 3188
rect 1636 3148 2452 3176
rect 1636 3136 1642 3148
rect 1688 3049 1716 3148
rect 1931 3073 1989 3079
rect 1673 3043 1731 3049
rect 1673 3009 1685 3043
rect 1719 3009 1731 3043
rect 1931 3039 1943 3073
rect 1977 3070 1989 3073
rect 1977 3040 1992 3070
rect 2314 3040 2320 3052
rect 1977 3039 2320 3040
rect 1931 3033 2320 3039
rect 1964 3012 2320 3033
rect 1673 3003 1731 3009
rect 2314 3000 2320 3012
rect 2372 3000 2378 3052
rect 2424 3040 2452 3148
rect 2590 3136 2596 3188
rect 2648 3176 2654 3188
rect 2685 3179 2743 3185
rect 2685 3176 2697 3179
rect 2648 3148 2697 3176
rect 2648 3136 2654 3148
rect 2685 3145 2697 3148
rect 2731 3145 2743 3179
rect 2685 3139 2743 3145
rect 3142 3136 3148 3188
rect 3200 3136 3206 3188
rect 3234 3136 3240 3188
rect 3292 3176 3298 3188
rect 4985 3179 5043 3185
rect 4985 3176 4997 3179
rect 3292 3148 4997 3176
rect 3292 3136 3298 3148
rect 4985 3145 4997 3148
rect 5031 3145 5043 3179
rect 4985 3139 5043 3145
rect 5261 3179 5319 3185
rect 5261 3145 5273 3179
rect 5307 3145 5319 3179
rect 5261 3139 5319 3145
rect 2498 3068 2504 3120
rect 2556 3108 2562 3120
rect 3160 3108 3188 3136
rect 2556 3080 3188 3108
rect 2556 3068 2562 3080
rect 3311 3073 3369 3079
rect 3050 3040 3056 3052
rect 2424 3012 3056 3040
rect 3050 3000 3056 3012
rect 3108 3000 3114 3052
rect 3311 3039 3323 3073
rect 3357 3070 3369 3073
rect 3357 3040 3372 3070
rect 3418 3068 3424 3120
rect 3476 3108 3482 3120
rect 4430 3108 4436 3120
rect 3476 3080 4436 3108
rect 3476 3068 3482 3080
rect 4430 3068 4436 3080
rect 4488 3068 4494 3120
rect 4525 3111 4583 3117
rect 4525 3077 4537 3111
rect 4571 3108 4583 3111
rect 5276 3108 5304 3139
rect 5994 3136 6000 3188
rect 6052 3136 6058 3188
rect 6549 3179 6607 3185
rect 6549 3145 6561 3179
rect 6595 3176 6607 3179
rect 6822 3176 6828 3188
rect 6595 3148 6828 3176
rect 6595 3145 6607 3148
rect 6549 3139 6607 3145
rect 6822 3136 6828 3148
rect 6880 3136 6886 3188
rect 7101 3179 7159 3185
rect 7101 3145 7113 3179
rect 7147 3176 7159 3179
rect 9766 3176 9772 3188
rect 7147 3148 9772 3176
rect 7147 3145 7159 3148
rect 7101 3139 7159 3145
rect 9766 3136 9772 3148
rect 9824 3136 9830 3188
rect 10410 3136 10416 3188
rect 10468 3136 10474 3188
rect 11517 3179 11575 3185
rect 11517 3145 11529 3179
rect 11563 3145 11575 3179
rect 11517 3139 11575 3145
rect 13265 3179 13323 3185
rect 13265 3145 13277 3179
rect 13311 3176 13323 3179
rect 13311 3148 13584 3176
rect 13311 3145 13323 3148
rect 13265 3139 13323 3145
rect 6012 3108 6040 3136
rect 10428 3108 10456 3136
rect 4571 3080 5304 3108
rect 5368 3080 6040 3108
rect 8680 3080 10456 3108
rect 4571 3077 4583 3080
rect 4525 3071 4583 3077
rect 5169 3043 5227 3049
rect 3357 3039 5120 3040
rect 3311 3033 5120 3039
rect 3344 3012 5120 3033
rect 2590 2932 2596 2984
rect 2648 2972 2654 2984
rect 2866 2972 2872 2984
rect 2648 2944 2872 2972
rect 2648 2932 2654 2944
rect 2866 2932 2872 2944
rect 2924 2932 2930 2984
rect 2958 2932 2964 2984
rect 3016 2932 3022 2984
rect 5092 2972 5120 3012
rect 5169 3009 5181 3043
rect 5215 3040 5227 3043
rect 5368 3040 5396 3080
rect 5215 3012 5396 3040
rect 5215 3009 5227 3012
rect 5169 3003 5227 3009
rect 5442 3000 5448 3052
rect 5500 3000 5506 3052
rect 6730 3000 6736 3052
rect 6788 3000 6794 3052
rect 7006 3000 7012 3052
rect 7064 3000 7070 3052
rect 7190 3000 7196 3052
rect 7248 3040 7254 3052
rect 7285 3043 7343 3049
rect 7285 3040 7297 3043
rect 7248 3012 7297 3040
rect 7248 3000 7254 3012
rect 7285 3009 7297 3012
rect 7331 3009 7343 3043
rect 7285 3003 7343 3009
rect 7374 3000 7380 3052
rect 7432 3040 7438 3052
rect 7561 3043 7619 3049
rect 7561 3040 7573 3043
rect 7432 3012 7573 3040
rect 7432 3000 7438 3012
rect 7561 3009 7573 3012
rect 7607 3009 7619 3043
rect 7561 3003 7619 3009
rect 7834 3000 7840 3052
rect 7892 3000 7898 3052
rect 8113 3043 8171 3049
rect 8113 3009 8125 3043
rect 8159 3040 8171 3043
rect 8294 3040 8300 3052
rect 8159 3012 8300 3040
rect 8159 3009 8171 3012
rect 8113 3003 8171 3009
rect 8294 3000 8300 3012
rect 8352 3000 8358 3052
rect 8386 3000 8392 3052
rect 8444 3000 8450 3052
rect 8680 3049 8708 3080
rect 8665 3043 8723 3049
rect 8665 3009 8677 3043
rect 8711 3009 8723 3043
rect 8665 3003 8723 3009
rect 8938 3000 8944 3052
rect 8996 3000 9002 3052
rect 9214 3000 9220 3052
rect 9272 3000 9278 3052
rect 9490 3000 9496 3052
rect 9548 3000 9554 3052
rect 9585 3043 9643 3049
rect 9585 3009 9597 3043
rect 9631 3009 9643 3043
rect 9585 3003 9643 3009
rect 6638 2972 6644 2984
rect 5092 2944 6644 2972
rect 6638 2932 6644 2944
rect 6696 2932 6702 2984
rect 8478 2932 8484 2984
rect 8536 2932 8542 2984
rect 9600 2972 9628 3003
rect 10226 3000 10232 3052
rect 10284 3000 10290 3052
rect 10689 3043 10747 3049
rect 10689 3009 10701 3043
rect 10735 3040 10747 3043
rect 10778 3040 10784 3052
rect 10735 3012 10784 3040
rect 10735 3009 10747 3012
rect 10689 3003 10747 3009
rect 10778 3000 10784 3012
rect 10836 3000 10842 3052
rect 11054 3000 11060 3052
rect 11112 3000 11118 3052
rect 11532 2972 11560 3139
rect 13354 3108 13360 3120
rect 12544 3080 13360 3108
rect 11701 3043 11759 3049
rect 11701 3009 11713 3043
rect 11747 3040 11759 3043
rect 12066 3040 12072 3052
rect 11747 3012 12072 3040
rect 11747 3009 11759 3012
rect 11701 3003 11759 3009
rect 12066 3000 12072 3012
rect 12124 3000 12130 3052
rect 12544 3049 12572 3080
rect 13354 3068 13360 3080
rect 13412 3068 13418 3120
rect 13556 3108 13584 3148
rect 13630 3136 13636 3188
rect 13688 3176 13694 3188
rect 13725 3179 13783 3185
rect 13725 3176 13737 3179
rect 13688 3148 13737 3176
rect 13688 3136 13694 3148
rect 13725 3145 13737 3148
rect 13771 3145 13783 3179
rect 13725 3139 13783 3145
rect 14090 3136 14096 3188
rect 14148 3136 14154 3188
rect 14550 3136 14556 3188
rect 14608 3136 14614 3188
rect 14645 3179 14703 3185
rect 14645 3145 14657 3179
rect 14691 3176 14703 3179
rect 15010 3176 15016 3188
rect 14691 3148 15016 3176
rect 14691 3145 14703 3148
rect 14645 3139 14703 3145
rect 15010 3136 15016 3148
rect 15068 3136 15074 3188
rect 15378 3136 15384 3188
rect 15436 3176 15442 3188
rect 16117 3179 16175 3185
rect 16117 3176 16129 3179
rect 15436 3148 16129 3176
rect 15436 3136 15442 3148
rect 16117 3145 16129 3148
rect 16163 3145 16175 3179
rect 16117 3139 16175 3145
rect 18049 3179 18107 3185
rect 18049 3145 18061 3179
rect 18095 3145 18107 3179
rect 18049 3139 18107 3145
rect 14568 3108 14596 3136
rect 15657 3111 15715 3117
rect 13556 3080 14596 3108
rect 14844 3080 15608 3108
rect 12529 3043 12587 3049
rect 12529 3009 12541 3043
rect 12575 3009 12587 3043
rect 12529 3003 12587 3009
rect 12802 3000 12808 3052
rect 12860 3000 12866 3052
rect 13556 3049 13584 3080
rect 14844 3052 14872 3080
rect 13541 3043 13599 3049
rect 13541 3009 13553 3043
rect 13587 3009 13599 3043
rect 13541 3003 13599 3009
rect 14001 3043 14059 3049
rect 14001 3009 14013 3043
rect 14047 3009 14059 3043
rect 14001 3003 14059 3009
rect 14277 3043 14335 3049
rect 14277 3009 14289 3043
rect 14323 3040 14335 3043
rect 14366 3040 14372 3052
rect 14323 3012 14372 3040
rect 14323 3009 14335 3012
rect 14277 3003 14335 3009
rect 9324 2944 9628 2972
rect 9692 2944 11560 2972
rect 14016 2972 14044 3003
rect 14366 3000 14372 3012
rect 14424 3000 14430 3052
rect 14553 3043 14611 3049
rect 14553 3009 14565 3043
rect 14599 3040 14611 3043
rect 14734 3040 14740 3052
rect 14599 3012 14740 3040
rect 14599 3009 14611 3012
rect 14553 3003 14611 3009
rect 14734 3000 14740 3012
rect 14792 3000 14798 3052
rect 14826 3000 14832 3052
rect 14884 3000 14890 3052
rect 15105 3043 15163 3049
rect 15105 3009 15117 3043
rect 15151 3009 15163 3043
rect 15105 3003 15163 3009
rect 14458 2972 14464 2984
rect 14016 2944 14464 2972
rect 2976 2836 3004 2932
rect 3970 2864 3976 2916
rect 4028 2904 4034 2916
rect 7098 2904 7104 2916
rect 4028 2876 7104 2904
rect 4028 2864 4034 2876
rect 7098 2864 7104 2876
rect 7156 2864 7162 2916
rect 8496 2904 8524 2932
rect 9324 2913 9352 2944
rect 7760 2876 8524 2904
rect 9309 2907 9367 2913
rect 7760 2848 7788 2876
rect 9309 2873 9321 2907
rect 9355 2873 9367 2907
rect 9309 2867 9367 2873
rect 9490 2864 9496 2916
rect 9548 2904 9554 2916
rect 9692 2904 9720 2944
rect 14458 2932 14464 2944
rect 14516 2932 14522 2984
rect 15120 2972 15148 3003
rect 15194 3000 15200 3052
rect 15252 3000 15258 3052
rect 15381 3043 15439 3049
rect 15381 3009 15393 3043
rect 15427 3040 15439 3043
rect 15470 3040 15476 3052
rect 15427 3012 15476 3040
rect 15427 3009 15439 3012
rect 15381 3003 15439 3009
rect 15470 3000 15476 3012
rect 15528 3000 15534 3052
rect 15580 3040 15608 3080
rect 15657 3077 15669 3111
rect 15703 3108 15715 3111
rect 15930 3108 15936 3120
rect 15703 3080 15936 3108
rect 15703 3077 15715 3080
rect 15657 3071 15715 3077
rect 15930 3068 15936 3080
rect 15988 3068 15994 3120
rect 17313 3111 17371 3117
rect 16224 3080 16896 3108
rect 16224 3040 16252 3080
rect 15580 3012 16252 3040
rect 16298 3000 16304 3052
rect 16356 3000 16362 3052
rect 16761 3043 16819 3049
rect 16761 3009 16773 3043
rect 16807 3009 16819 3043
rect 16761 3003 16819 3009
rect 14936 2944 15148 2972
rect 15212 2972 15240 3000
rect 16776 2972 16804 3003
rect 15212 2944 16804 2972
rect 16868 2972 16896 3080
rect 17313 3077 17325 3111
rect 17359 3108 17371 3111
rect 18064 3108 18092 3139
rect 18138 3136 18144 3188
rect 18196 3136 18202 3188
rect 18506 3136 18512 3188
rect 18564 3136 18570 3188
rect 19610 3176 19616 3188
rect 19168 3148 19616 3176
rect 17359 3080 18092 3108
rect 17359 3077 17371 3080
rect 17313 3071 17371 3077
rect 17954 3000 17960 3052
rect 18012 3000 18018 3052
rect 18046 2972 18052 2984
rect 16868 2944 18052 2972
rect 9548 2876 9720 2904
rect 9769 2907 9827 2913
rect 9548 2864 9554 2876
rect 9769 2873 9781 2907
rect 9815 2904 9827 2907
rect 10318 2904 10324 2916
rect 9815 2876 10324 2904
rect 9815 2873 9827 2876
rect 9769 2867 9827 2873
rect 10318 2864 10324 2876
rect 10376 2864 10382 2916
rect 11882 2904 11888 2916
rect 11256 2876 11888 2904
rect 4065 2839 4123 2845
rect 4065 2836 4077 2839
rect 2976 2808 4077 2836
rect 4065 2805 4077 2808
rect 4111 2805 4123 2839
rect 4065 2799 4123 2805
rect 4246 2796 4252 2848
rect 4304 2836 4310 2848
rect 4617 2839 4675 2845
rect 4617 2836 4629 2839
rect 4304 2808 4629 2836
rect 4304 2796 4310 2808
rect 4617 2805 4629 2808
rect 4663 2805 4675 2839
rect 4617 2799 4675 2805
rect 6822 2796 6828 2848
rect 6880 2796 6886 2848
rect 7374 2796 7380 2848
rect 7432 2796 7438 2848
rect 7650 2796 7656 2848
rect 7708 2796 7714 2848
rect 7742 2796 7748 2848
rect 7800 2796 7806 2848
rect 7926 2796 7932 2848
rect 7984 2796 7990 2848
rect 8202 2796 8208 2848
rect 8260 2796 8266 2848
rect 8478 2796 8484 2848
rect 8536 2796 8542 2848
rect 8570 2796 8576 2848
rect 8628 2836 8634 2848
rect 8757 2839 8815 2845
rect 8757 2836 8769 2839
rect 8628 2808 8769 2836
rect 8628 2796 8634 2808
rect 8757 2805 8769 2808
rect 8803 2805 8815 2839
rect 8757 2799 8815 2805
rect 9033 2839 9091 2845
rect 9033 2805 9045 2839
rect 9079 2836 9091 2839
rect 9122 2836 9128 2848
rect 9079 2808 9128 2836
rect 9079 2805 9091 2808
rect 9033 2799 9091 2805
rect 9122 2796 9128 2808
rect 9180 2796 9186 2848
rect 9674 2796 9680 2848
rect 9732 2836 9738 2848
rect 10045 2839 10103 2845
rect 10045 2836 10057 2839
rect 9732 2808 10057 2836
rect 9732 2796 9738 2808
rect 10045 2805 10057 2808
rect 10091 2805 10103 2839
rect 10045 2799 10103 2805
rect 10502 2796 10508 2848
rect 10560 2796 10566 2848
rect 11256 2845 11284 2876
rect 11882 2864 11888 2876
rect 11940 2864 11946 2916
rect 13630 2864 13636 2916
rect 13688 2904 13694 2916
rect 14936 2904 14964 2944
rect 18046 2932 18052 2944
rect 18104 2932 18110 2984
rect 18156 2972 18184 3136
rect 18230 3000 18236 3052
rect 18288 3000 18294 3052
rect 18414 3000 18420 3052
rect 18472 3000 18478 3052
rect 18877 3043 18935 3049
rect 18877 3009 18889 3043
rect 18923 3040 18935 3043
rect 19058 3040 19064 3052
rect 18923 3012 19064 3040
rect 18923 3009 18935 3012
rect 18877 3003 18935 3009
rect 19058 3000 19064 3012
rect 19116 3000 19122 3052
rect 19168 3049 19196 3148
rect 19610 3136 19616 3148
rect 19668 3136 19674 3188
rect 20070 3136 20076 3188
rect 20128 3136 20134 3188
rect 20441 3179 20499 3185
rect 20441 3145 20453 3179
rect 20487 3176 20499 3179
rect 20622 3176 20628 3188
rect 20487 3148 20628 3176
rect 20487 3145 20499 3148
rect 20441 3139 20499 3145
rect 20622 3136 20628 3148
rect 20680 3136 20686 3188
rect 20809 3179 20867 3185
rect 20809 3145 20821 3179
rect 20855 3176 20867 3179
rect 20898 3176 20904 3188
rect 20855 3148 20904 3176
rect 20855 3145 20867 3148
rect 20809 3139 20867 3145
rect 20898 3136 20904 3148
rect 20956 3136 20962 3188
rect 21358 3136 21364 3188
rect 21416 3136 21422 3188
rect 19981 3111 20039 3117
rect 19981 3077 19993 3111
rect 20027 3108 20039 3111
rect 21376 3108 21404 3136
rect 20027 3080 21404 3108
rect 20027 3077 20039 3080
rect 19981 3071 20039 3077
rect 19153 3043 19211 3049
rect 19153 3009 19165 3043
rect 19199 3009 19211 3043
rect 19153 3003 19211 3009
rect 19518 3000 19524 3052
rect 19576 3000 19582 3052
rect 20349 3043 20407 3049
rect 20349 3040 20361 3043
rect 19628 3012 20361 3040
rect 19628 2972 19656 3012
rect 20349 3009 20361 3012
rect 20395 3009 20407 3043
rect 20349 3003 20407 3009
rect 20438 3000 20444 3052
rect 20496 3040 20502 3052
rect 20717 3043 20775 3049
rect 20717 3040 20729 3043
rect 20496 3012 20729 3040
rect 20496 3000 20502 3012
rect 20717 3009 20729 3012
rect 20763 3009 20775 3043
rect 20717 3003 20775 3009
rect 20806 3000 20812 3052
rect 20864 3040 20870 3052
rect 21085 3043 21143 3049
rect 21085 3040 21097 3043
rect 20864 3012 21097 3040
rect 20864 3000 20870 3012
rect 21085 3009 21097 3012
rect 21131 3009 21143 3043
rect 21085 3003 21143 3009
rect 21545 3043 21603 3049
rect 21545 3009 21557 3043
rect 21591 3009 21603 3043
rect 21545 3003 21603 3009
rect 18156 2944 19656 2972
rect 19794 2932 19800 2984
rect 19852 2972 19858 2984
rect 21560 2972 21588 3003
rect 19852 2944 21588 2972
rect 19852 2932 19858 2944
rect 22186 2932 22192 2984
rect 22244 2932 22250 2984
rect 13688 2876 14964 2904
rect 13688 2864 13694 2876
rect 15010 2864 15016 2916
rect 15068 2904 15074 2916
rect 15068 2876 15792 2904
rect 15068 2864 15074 2876
rect 11241 2839 11299 2845
rect 11241 2805 11253 2839
rect 11287 2805 11299 2839
rect 11241 2799 11299 2805
rect 12066 2796 12072 2848
rect 12124 2836 12130 2848
rect 12345 2839 12403 2845
rect 12345 2836 12357 2839
rect 12124 2808 12357 2836
rect 12124 2796 12130 2808
rect 12345 2805 12357 2808
rect 12391 2805 12403 2839
rect 12345 2799 12403 2805
rect 12618 2796 12624 2848
rect 12676 2796 12682 2848
rect 13814 2796 13820 2848
rect 13872 2796 13878 2848
rect 14366 2796 14372 2848
rect 14424 2796 14430 2848
rect 14734 2796 14740 2848
rect 14792 2836 14798 2848
rect 14921 2839 14979 2845
rect 14921 2836 14933 2839
rect 14792 2808 14933 2836
rect 14792 2796 14798 2808
rect 14921 2805 14933 2808
rect 14967 2805 14979 2839
rect 14921 2799 14979 2805
rect 15197 2839 15255 2845
rect 15197 2805 15209 2839
rect 15243 2836 15255 2839
rect 15470 2836 15476 2848
rect 15243 2808 15476 2836
rect 15243 2805 15255 2808
rect 15197 2799 15255 2805
rect 15470 2796 15476 2808
rect 15528 2796 15534 2848
rect 15764 2845 15792 2876
rect 15838 2864 15844 2916
rect 15896 2904 15902 2916
rect 16945 2907 17003 2913
rect 16945 2904 16957 2907
rect 15896 2876 16957 2904
rect 15896 2864 15902 2876
rect 16945 2873 16957 2876
rect 16991 2873 17003 2907
rect 16945 2867 17003 2873
rect 17218 2864 17224 2916
rect 17276 2904 17282 2916
rect 19334 2904 19340 2916
rect 17276 2876 19340 2904
rect 17276 2864 17282 2876
rect 19334 2864 19340 2876
rect 19392 2864 19398 2916
rect 19521 2907 19579 2913
rect 19521 2873 19533 2907
rect 19567 2904 19579 2907
rect 20530 2904 20536 2916
rect 19567 2876 20536 2904
rect 19567 2873 19579 2876
rect 19521 2867 19579 2873
rect 20530 2864 20536 2876
rect 20588 2864 20594 2916
rect 21269 2907 21327 2913
rect 21269 2873 21281 2907
rect 21315 2904 21327 2907
rect 22204 2904 22232 2932
rect 21315 2876 22232 2904
rect 21315 2873 21327 2876
rect 21269 2867 21327 2873
rect 15749 2839 15807 2845
rect 15749 2805 15761 2839
rect 15795 2805 15807 2839
rect 15749 2799 15807 2805
rect 16022 2796 16028 2848
rect 16080 2836 16086 2848
rect 17405 2839 17463 2845
rect 17405 2836 17417 2839
rect 16080 2808 17417 2836
rect 16080 2796 16086 2808
rect 17405 2805 17417 2808
rect 17451 2805 17463 2839
rect 17405 2799 17463 2805
rect 17770 2796 17776 2848
rect 17828 2796 17834 2848
rect 18874 2796 18880 2848
rect 18932 2836 18938 2848
rect 19058 2836 19064 2848
rect 18932 2808 19064 2836
rect 18932 2796 18938 2808
rect 19058 2796 19064 2808
rect 19116 2796 19122 2848
rect 21358 2796 21364 2848
rect 21416 2796 21422 2848
rect 1104 2746 21896 2768
rect 1104 2694 3549 2746
rect 3601 2694 3613 2746
rect 3665 2694 3677 2746
rect 3729 2694 3741 2746
rect 3793 2694 3805 2746
rect 3857 2694 8747 2746
rect 8799 2694 8811 2746
rect 8863 2694 8875 2746
rect 8927 2694 8939 2746
rect 8991 2694 9003 2746
rect 9055 2694 13945 2746
rect 13997 2694 14009 2746
rect 14061 2694 14073 2746
rect 14125 2694 14137 2746
rect 14189 2694 14201 2746
rect 14253 2694 19143 2746
rect 19195 2694 19207 2746
rect 19259 2694 19271 2746
rect 19323 2694 19335 2746
rect 19387 2694 19399 2746
rect 19451 2694 21896 2746
rect 1104 2672 21896 2694
rect 2314 2592 2320 2644
rect 2372 2592 2378 2644
rect 3329 2635 3387 2641
rect 3329 2632 3341 2635
rect 2746 2604 3341 2632
rect 1302 2524 1308 2576
rect 1360 2564 1366 2576
rect 2746 2564 2774 2604
rect 3329 2601 3341 2604
rect 3375 2601 3387 2635
rect 3329 2595 3387 2601
rect 4154 2592 4160 2644
rect 4212 2592 4218 2644
rect 4522 2592 4528 2644
rect 4580 2592 4586 2644
rect 5166 2592 5172 2644
rect 5224 2592 5230 2644
rect 5350 2592 5356 2644
rect 5408 2632 5414 2644
rect 5445 2635 5503 2641
rect 5445 2632 5457 2635
rect 5408 2604 5457 2632
rect 5408 2592 5414 2604
rect 5445 2601 5457 2604
rect 5491 2601 5503 2635
rect 5445 2595 5503 2601
rect 7190 2592 7196 2644
rect 7248 2632 7254 2644
rect 7561 2635 7619 2641
rect 7561 2632 7573 2635
rect 7248 2604 7573 2632
rect 7248 2592 7254 2604
rect 7561 2601 7573 2604
rect 7607 2601 7619 2635
rect 7561 2595 7619 2601
rect 7926 2592 7932 2644
rect 7984 2592 7990 2644
rect 8665 2635 8723 2641
rect 8665 2601 8677 2635
rect 8711 2632 8723 2635
rect 10686 2632 10692 2644
rect 8711 2604 10692 2632
rect 8711 2601 8723 2604
rect 8665 2595 8723 2601
rect 10686 2592 10692 2604
rect 10744 2592 10750 2644
rect 10781 2635 10839 2641
rect 10781 2601 10793 2635
rect 10827 2632 10839 2635
rect 10962 2632 10968 2644
rect 10827 2604 10968 2632
rect 10827 2601 10839 2604
rect 10781 2595 10839 2601
rect 10962 2592 10968 2604
rect 11020 2592 11026 2644
rect 12529 2635 12587 2641
rect 12529 2632 12541 2635
rect 11900 2604 12541 2632
rect 1360 2536 2774 2564
rect 9309 2567 9367 2573
rect 1360 2524 1366 2536
rect 9309 2533 9321 2567
rect 9355 2564 9367 2567
rect 10870 2564 10876 2576
rect 9355 2536 10876 2564
rect 9355 2533 9367 2536
rect 9309 2527 9367 2533
rect 10870 2524 10876 2536
rect 10928 2524 10934 2576
rect 11054 2524 11060 2576
rect 11112 2564 11118 2576
rect 11900 2564 11928 2604
rect 12529 2601 12541 2604
rect 12575 2632 12587 2635
rect 12897 2635 12955 2641
rect 12897 2632 12909 2635
rect 12575 2604 12909 2632
rect 12575 2601 12587 2604
rect 12529 2595 12587 2601
rect 12897 2601 12909 2604
rect 12943 2601 12955 2635
rect 12897 2595 12955 2601
rect 14461 2635 14519 2641
rect 14461 2601 14473 2635
rect 14507 2632 14519 2635
rect 14826 2632 14832 2644
rect 14507 2604 14832 2632
rect 14507 2601 14519 2604
rect 14461 2595 14519 2601
rect 14826 2592 14832 2604
rect 14884 2592 14890 2644
rect 15562 2592 15568 2644
rect 15620 2592 15626 2644
rect 15654 2592 15660 2644
rect 15712 2632 15718 2644
rect 16669 2635 16727 2641
rect 16669 2632 16681 2635
rect 15712 2604 16681 2632
rect 15712 2592 15718 2604
rect 16669 2601 16681 2604
rect 16715 2601 16727 2635
rect 16669 2595 16727 2601
rect 18969 2635 19027 2641
rect 18969 2601 18981 2635
rect 19015 2632 19027 2635
rect 21634 2632 21640 2644
rect 19015 2604 21640 2632
rect 19015 2601 19027 2604
rect 18969 2595 19027 2601
rect 21634 2592 21640 2604
rect 21692 2592 21698 2644
rect 16574 2564 16580 2576
rect 11112 2536 11928 2564
rect 11112 2524 11118 2536
rect 1210 2456 1216 2508
rect 1268 2496 1274 2508
rect 2869 2499 2927 2505
rect 2869 2496 2881 2499
rect 1268 2468 2881 2496
rect 1268 2456 1274 2468
rect 2869 2465 2881 2468
rect 2915 2465 2927 2499
rect 8389 2499 8447 2505
rect 2869 2459 2927 2465
rect 3804 2468 4936 2496
rect 1673 2431 1731 2437
rect 1673 2397 1685 2431
rect 1719 2428 1731 2431
rect 2038 2428 2044 2440
rect 1719 2400 2044 2428
rect 1719 2397 1731 2400
rect 1673 2391 1731 2397
rect 2038 2388 2044 2400
rect 2096 2388 2102 2440
rect 2590 2388 2596 2440
rect 2648 2388 2654 2440
rect 3804 2428 3832 2468
rect 2700 2400 3832 2428
rect 658 2320 664 2372
rect 716 2360 722 2372
rect 2700 2360 2728 2400
rect 3878 2388 3884 2440
rect 3936 2388 3942 2440
rect 4154 2388 4160 2440
rect 4212 2388 4218 2440
rect 4341 2431 4399 2437
rect 4341 2397 4353 2431
rect 4387 2397 4399 2431
rect 4341 2391 4399 2397
rect 716 2332 2728 2360
rect 3237 2363 3295 2369
rect 716 2320 722 2332
rect 3237 2329 3249 2363
rect 3283 2360 3295 2363
rect 4172 2360 4200 2388
rect 3283 2332 4200 2360
rect 3283 2329 3295 2332
rect 3237 2323 3295 2329
rect 934 2252 940 2304
rect 992 2292 998 2304
rect 3694 2292 3700 2304
rect 992 2264 3700 2292
rect 992 2252 998 2264
rect 3694 2252 3700 2264
rect 3752 2252 3758 2304
rect 4154 2252 4160 2304
rect 4212 2292 4218 2304
rect 4356 2292 4384 2391
rect 4430 2388 4436 2440
rect 4488 2428 4494 2440
rect 4798 2428 4804 2440
rect 4488 2400 4804 2428
rect 4488 2388 4494 2400
rect 4798 2388 4804 2400
rect 4856 2388 4862 2440
rect 4908 2437 4936 2468
rect 8389 2465 8401 2499
rect 8435 2496 8447 2499
rect 10778 2496 10784 2508
rect 8435 2468 10784 2496
rect 8435 2465 8447 2468
rect 8389 2459 8447 2465
rect 10778 2456 10784 2468
rect 10836 2456 10842 2508
rect 11241 2499 11299 2505
rect 11241 2496 11253 2499
rect 10870 2468 11253 2496
rect 4893 2431 4951 2437
rect 4893 2397 4905 2431
rect 4939 2397 4951 2431
rect 4893 2391 4951 2397
rect 4985 2431 5043 2437
rect 4985 2397 4997 2431
rect 5031 2397 5043 2431
rect 4985 2391 5043 2397
rect 4614 2320 4620 2372
rect 4672 2360 4678 2372
rect 5000 2360 5028 2391
rect 5626 2388 5632 2440
rect 5684 2388 5690 2440
rect 5828 2400 6592 2428
rect 4672 2332 5028 2360
rect 4672 2320 4678 2332
rect 4212 2264 4384 2292
rect 4709 2295 4767 2301
rect 4212 2252 4218 2264
rect 4709 2261 4721 2295
rect 4755 2292 4767 2295
rect 5828 2292 5856 2400
rect 5902 2320 5908 2372
rect 5960 2360 5966 2372
rect 6089 2363 6147 2369
rect 6089 2360 6101 2363
rect 5960 2332 6101 2360
rect 5960 2320 5966 2332
rect 6089 2329 6101 2332
rect 6135 2329 6147 2363
rect 6089 2323 6147 2329
rect 6270 2320 6276 2372
rect 6328 2320 6334 2372
rect 6457 2363 6515 2369
rect 6457 2329 6469 2363
rect 6503 2329 6515 2363
rect 6457 2323 6515 2329
rect 4755 2264 5856 2292
rect 4755 2261 4767 2264
rect 4709 2255 4767 2261
rect 5994 2252 6000 2304
rect 6052 2292 6058 2304
rect 6472 2292 6500 2323
rect 6052 2264 6500 2292
rect 6564 2292 6592 2400
rect 6914 2388 6920 2440
rect 6972 2388 6978 2440
rect 7469 2431 7527 2437
rect 7469 2397 7481 2431
rect 7515 2428 7527 2431
rect 7558 2428 7564 2440
rect 7515 2400 7564 2428
rect 7515 2397 7527 2400
rect 7469 2391 7527 2397
rect 7558 2388 7564 2400
rect 7616 2388 7622 2440
rect 7650 2388 7656 2440
rect 7708 2428 7714 2440
rect 7745 2431 7803 2437
rect 7745 2428 7757 2431
rect 7708 2400 7757 2428
rect 7708 2388 7714 2400
rect 7745 2397 7757 2400
rect 7791 2397 7803 2431
rect 7745 2391 7803 2397
rect 8202 2388 8208 2440
rect 8260 2388 8266 2440
rect 8481 2431 8539 2437
rect 8481 2397 8493 2431
rect 8527 2428 8539 2431
rect 8570 2428 8576 2440
rect 8527 2400 8576 2428
rect 8527 2397 8539 2400
rect 8481 2391 8539 2397
rect 8570 2388 8576 2400
rect 8628 2388 8634 2440
rect 9582 2388 9588 2440
rect 9640 2388 9646 2440
rect 9677 2431 9735 2437
rect 9677 2397 9689 2431
rect 9723 2428 9735 2431
rect 10137 2431 10195 2437
rect 10137 2428 10149 2431
rect 9723 2400 10149 2428
rect 9723 2397 9735 2400
rect 9677 2391 9735 2397
rect 6641 2363 6699 2369
rect 6641 2329 6653 2363
rect 6687 2360 6699 2363
rect 9600 2360 9628 2388
rect 9784 2372 9812 2400
rect 10137 2397 10149 2400
rect 10183 2397 10195 2431
rect 10137 2391 10195 2397
rect 10413 2431 10471 2437
rect 10413 2397 10425 2431
rect 10459 2428 10471 2431
rect 10594 2428 10600 2440
rect 10459 2400 10600 2428
rect 10459 2397 10471 2400
rect 10413 2391 10471 2397
rect 10594 2388 10600 2400
rect 10652 2388 10658 2440
rect 10689 2431 10747 2437
rect 10689 2397 10701 2431
rect 10735 2428 10747 2431
rect 10870 2428 10898 2468
rect 11241 2465 11253 2468
rect 11287 2465 11299 2499
rect 11241 2459 11299 2465
rect 10735 2400 10898 2428
rect 10965 2431 11023 2437
rect 10735 2397 10747 2400
rect 10689 2391 10747 2397
rect 10965 2397 10977 2431
rect 11011 2397 11023 2431
rect 10965 2391 11023 2397
rect 6687 2332 9628 2360
rect 6687 2329 6699 2332
rect 6641 2323 6699 2329
rect 9766 2320 9772 2372
rect 9824 2320 9830 2372
rect 10704 2360 10732 2391
rect 9876 2332 10732 2360
rect 6914 2292 6920 2304
rect 6564 2264 6920 2292
rect 6052 2252 6058 2264
rect 6914 2252 6920 2264
rect 6972 2252 6978 2304
rect 7006 2252 7012 2304
rect 7064 2252 7070 2304
rect 7190 2252 7196 2304
rect 7248 2292 7254 2304
rect 9876 2292 9904 2332
rect 10870 2320 10876 2372
rect 10928 2360 10934 2372
rect 10980 2360 11008 2391
rect 11606 2388 11612 2440
rect 11664 2388 11670 2440
rect 11900 2437 11928 2536
rect 14568 2536 16580 2564
rect 11885 2431 11943 2437
rect 11885 2397 11897 2431
rect 11931 2397 11943 2431
rect 12253 2431 12311 2437
rect 12253 2428 12265 2431
rect 11885 2391 11943 2397
rect 11992 2400 12265 2428
rect 10928 2332 11836 2360
rect 10928 2320 10934 2332
rect 11808 2304 11836 2332
rect 11992 2304 12020 2400
rect 12253 2397 12265 2400
rect 12299 2397 12311 2431
rect 12253 2391 12311 2397
rect 13357 2431 13415 2437
rect 13357 2397 13369 2431
rect 13403 2428 13415 2431
rect 13817 2431 13875 2437
rect 13817 2428 13829 2431
rect 13403 2400 13829 2428
rect 13403 2397 13415 2400
rect 13357 2391 13415 2397
rect 13817 2397 13829 2400
rect 13863 2428 13875 2431
rect 14568 2428 14596 2536
rect 16574 2524 16580 2536
rect 16632 2524 16638 2576
rect 18046 2524 18052 2576
rect 18104 2564 18110 2576
rect 18104 2536 20392 2564
rect 18104 2524 18110 2536
rect 15102 2456 15108 2508
rect 15160 2496 15166 2508
rect 15160 2468 15516 2496
rect 15160 2456 15166 2468
rect 13863 2400 14596 2428
rect 14645 2431 14703 2437
rect 13863 2397 13875 2400
rect 13817 2391 13875 2397
rect 14645 2397 14657 2431
rect 14691 2397 14703 2431
rect 14645 2391 14703 2397
rect 14829 2431 14887 2437
rect 14829 2397 14841 2431
rect 14875 2428 14887 2431
rect 15378 2428 15384 2440
rect 14875 2400 15384 2428
rect 14875 2397 14887 2400
rect 14829 2391 14887 2397
rect 12268 2360 12296 2391
rect 14277 2363 14335 2369
rect 14277 2360 14289 2363
rect 12268 2332 14289 2360
rect 14277 2329 14289 2332
rect 14323 2329 14335 2363
rect 14660 2360 14688 2391
rect 15378 2388 15384 2400
rect 15436 2388 15442 2440
rect 15488 2369 15516 2468
rect 16114 2456 16120 2508
rect 16172 2496 16178 2508
rect 16172 2468 16620 2496
rect 16172 2456 16178 2468
rect 16592 2437 16620 2468
rect 17586 2456 17592 2508
rect 17644 2456 17650 2508
rect 17678 2456 17684 2508
rect 17736 2496 17742 2508
rect 17736 2468 19288 2496
rect 17736 2456 17742 2468
rect 16007 2431 16065 2437
rect 16007 2397 16019 2431
rect 16053 2428 16065 2431
rect 16577 2431 16635 2437
rect 16053 2424 16068 2428
rect 16053 2397 16342 2424
rect 16007 2396 16342 2397
rect 16007 2391 16065 2396
rect 15473 2363 15531 2369
rect 14660 2332 15424 2360
rect 14277 2323 14335 2329
rect 7248 2264 9904 2292
rect 7248 2252 7254 2264
rect 9950 2252 9956 2304
rect 10008 2252 10014 2304
rect 10226 2252 10232 2304
rect 10284 2252 10290 2304
rect 10502 2252 10508 2304
rect 10560 2252 10566 2304
rect 11238 2252 11244 2304
rect 11296 2292 11302 2304
rect 11425 2295 11483 2301
rect 11425 2292 11437 2295
rect 11296 2264 11437 2292
rect 11296 2252 11302 2264
rect 11425 2261 11437 2264
rect 11471 2261 11483 2295
rect 11425 2255 11483 2261
rect 11698 2252 11704 2304
rect 11756 2252 11762 2304
rect 11790 2252 11796 2304
rect 11848 2252 11854 2304
rect 11974 2252 11980 2304
rect 12032 2252 12038 2304
rect 12069 2295 12127 2301
rect 12069 2261 12081 2295
rect 12115 2292 12127 2295
rect 12434 2292 12440 2304
rect 12115 2264 12440 2292
rect 12115 2261 12127 2264
rect 12069 2255 12127 2261
rect 12434 2252 12440 2264
rect 12492 2252 12498 2304
rect 13630 2252 13636 2304
rect 13688 2252 13694 2304
rect 15013 2295 15071 2301
rect 15013 2261 15025 2295
rect 15059 2292 15071 2295
rect 15102 2292 15108 2304
rect 15059 2264 15108 2292
rect 15059 2261 15071 2264
rect 15013 2255 15071 2261
rect 15102 2252 15108 2264
rect 15160 2252 15166 2304
rect 15396 2292 15424 2332
rect 15473 2329 15485 2363
rect 15519 2329 15531 2363
rect 16314 2360 16342 2396
rect 16577 2397 16589 2431
rect 16623 2397 16635 2431
rect 16577 2391 16635 2397
rect 17218 2388 17224 2440
rect 17276 2388 17282 2440
rect 17770 2388 17776 2440
rect 17828 2388 17834 2440
rect 18506 2388 18512 2440
rect 18564 2388 18570 2440
rect 18690 2388 18696 2440
rect 18748 2428 18754 2440
rect 19260 2437 19288 2468
rect 20070 2456 20076 2508
rect 20128 2456 20134 2508
rect 20364 2437 20392 2536
rect 21174 2456 21180 2508
rect 21232 2456 21238 2508
rect 18877 2431 18935 2437
rect 18877 2428 18889 2431
rect 18748 2400 18889 2428
rect 18748 2388 18754 2400
rect 18877 2397 18889 2400
rect 18923 2397 18935 2431
rect 18877 2391 18935 2397
rect 19245 2431 19303 2437
rect 19245 2397 19257 2431
rect 19291 2397 19303 2431
rect 19245 2391 19303 2397
rect 20349 2431 20407 2437
rect 20349 2397 20361 2431
rect 20395 2397 20407 2431
rect 20349 2391 20407 2397
rect 17788 2360 17816 2388
rect 20162 2360 20168 2372
rect 15473 2323 15531 2329
rect 16040 2332 16252 2360
rect 16314 2332 17816 2360
rect 17880 2332 20168 2360
rect 16040 2292 16068 2332
rect 15396 2264 16068 2292
rect 16114 2252 16120 2304
rect 16172 2252 16178 2304
rect 16224 2292 16252 2332
rect 17880 2292 17908 2332
rect 20162 2320 20168 2332
rect 20220 2320 20226 2372
rect 16224 2264 17908 2292
rect 18322 2252 18328 2304
rect 18380 2252 18386 2304
rect 1104 2202 22056 2224
rect 1104 2150 6148 2202
rect 6200 2150 6212 2202
rect 6264 2150 6276 2202
rect 6328 2150 6340 2202
rect 6392 2150 6404 2202
rect 6456 2150 11346 2202
rect 11398 2150 11410 2202
rect 11462 2150 11474 2202
rect 11526 2150 11538 2202
rect 11590 2150 11602 2202
rect 11654 2150 16544 2202
rect 16596 2150 16608 2202
rect 16660 2150 16672 2202
rect 16724 2150 16736 2202
rect 16788 2150 16800 2202
rect 16852 2150 21742 2202
rect 21794 2150 21806 2202
rect 21858 2150 21870 2202
rect 21922 2150 21934 2202
rect 21986 2150 21998 2202
rect 22050 2150 22056 2202
rect 1104 2128 22056 2150
rect 1394 2048 1400 2100
rect 1452 2088 1458 2100
rect 1581 2091 1639 2097
rect 1581 2088 1593 2091
rect 1452 2060 1593 2088
rect 1452 2048 1458 2060
rect 1581 2057 1593 2060
rect 1627 2057 1639 2091
rect 1581 2051 1639 2057
rect 2590 2048 2596 2100
rect 2648 2048 2654 2100
rect 2866 2048 2872 2100
rect 2924 2048 2930 2100
rect 3421 2091 3479 2097
rect 3421 2057 3433 2091
rect 3467 2057 3479 2091
rect 3421 2051 3479 2057
rect 1486 1980 1492 2032
rect 1544 1980 1550 2032
rect 1946 1980 1952 2032
rect 2004 2020 2010 2032
rect 2041 2023 2099 2029
rect 2041 2020 2053 2023
rect 2004 1992 2053 2020
rect 2004 1980 2010 1992
rect 2041 1989 2053 1992
rect 2087 1989 2099 2023
rect 2041 1983 2099 1989
rect 2409 2023 2467 2029
rect 2409 1989 2421 2023
rect 2455 2020 2467 2023
rect 2608 2020 2636 2048
rect 2455 1992 2636 2020
rect 3436 2020 3464 2051
rect 3970 2048 3976 2100
rect 4028 2088 4034 2100
rect 4341 2091 4399 2097
rect 4341 2088 4353 2091
rect 4028 2060 4353 2088
rect 4028 2048 4034 2060
rect 4341 2057 4353 2060
rect 4387 2057 4399 2091
rect 4341 2051 4399 2057
rect 4522 2048 4528 2100
rect 4580 2048 4586 2100
rect 4709 2091 4767 2097
rect 4709 2057 4721 2091
rect 4755 2088 4767 2091
rect 4798 2088 4804 2100
rect 4755 2060 4804 2088
rect 4755 2057 4767 2060
rect 4709 2051 4767 2057
rect 4798 2048 4804 2060
rect 4856 2048 4862 2100
rect 5718 2048 5724 2100
rect 5776 2088 5782 2100
rect 6825 2091 6883 2097
rect 6825 2088 6837 2091
rect 5776 2060 6837 2088
rect 5776 2048 5782 2060
rect 6825 2057 6837 2060
rect 6871 2057 6883 2091
rect 7190 2088 7196 2100
rect 6825 2051 6883 2057
rect 7024 2060 7196 2088
rect 4540 2020 4568 2048
rect 7024 2020 7052 2060
rect 7190 2048 7196 2060
rect 7248 2048 7254 2100
rect 8018 2088 8024 2100
rect 7484 2060 8024 2088
rect 3436 1992 4568 2020
rect 4816 1992 7052 2020
rect 7101 2023 7159 2029
rect 2455 1989 2467 1992
rect 2409 1983 2467 1989
rect 4816 1964 4844 1992
rect 7101 1989 7113 2023
rect 7147 2020 7159 2023
rect 7374 2020 7380 2032
rect 7147 1992 7380 2020
rect 7147 1989 7159 1992
rect 7101 1983 7159 1989
rect 7374 1980 7380 1992
rect 7432 1980 7438 2032
rect 7484 2029 7512 2060
rect 8018 2048 8024 2060
rect 8076 2048 8082 2100
rect 8665 2091 8723 2097
rect 8665 2057 8677 2091
rect 8711 2088 8723 2091
rect 9398 2088 9404 2100
rect 8711 2060 9404 2088
rect 8711 2057 8723 2060
rect 8665 2051 8723 2057
rect 9398 2048 9404 2060
rect 9456 2048 9462 2100
rect 9950 2048 9956 2100
rect 10008 2088 10014 2100
rect 10008 2060 11008 2088
rect 10008 2048 10014 2060
rect 7469 2023 7527 2029
rect 7469 1989 7481 2023
rect 7515 1989 7527 2023
rect 7469 1983 7527 1989
rect 7834 1980 7840 2032
rect 7892 1980 7898 2032
rect 8202 1980 8208 2032
rect 8260 1980 8266 2032
rect 9122 2020 9128 2032
rect 8496 1992 9128 2020
rect 2498 1912 2504 1964
rect 2556 1952 2562 1964
rect 2593 1955 2651 1961
rect 2593 1952 2605 1955
rect 2556 1924 2605 1952
rect 2556 1912 2562 1924
rect 2593 1921 2605 1924
rect 2639 1921 2651 1955
rect 2593 1915 2651 1921
rect 3234 1912 3240 1964
rect 3292 1912 3298 1964
rect 3418 1912 3424 1964
rect 3476 1952 3482 1964
rect 3697 1955 3755 1961
rect 3697 1952 3709 1955
rect 3476 1924 3709 1952
rect 3476 1912 3482 1924
rect 3697 1921 3709 1924
rect 3743 1921 3755 1955
rect 3697 1915 3755 1921
rect 3878 1912 3884 1964
rect 3936 1952 3942 1964
rect 4157 1955 4215 1961
rect 4157 1952 4169 1955
rect 3936 1924 4169 1952
rect 3936 1912 3942 1924
rect 4157 1921 4169 1924
rect 4203 1921 4215 1955
rect 4157 1915 4215 1921
rect 4614 1912 4620 1964
rect 4672 1912 4678 1964
rect 4798 1912 4804 1964
rect 4856 1912 4862 1964
rect 4890 1912 4896 1964
rect 4948 1912 4954 1964
rect 5537 1955 5595 1961
rect 5537 1921 5549 1955
rect 5583 1952 5595 1955
rect 6546 1952 6552 1964
rect 5583 1924 6552 1952
rect 5583 1921 5595 1924
rect 5537 1915 5595 1921
rect 6546 1912 6552 1924
rect 6604 1912 6610 1964
rect 6641 1955 6699 1961
rect 6641 1921 6653 1955
rect 6687 1952 6699 1955
rect 6822 1952 6828 1964
rect 6687 1924 6828 1952
rect 6687 1921 6699 1924
rect 6641 1915 6699 1921
rect 6822 1912 6828 1924
rect 6880 1912 6886 1964
rect 8496 1961 8524 1992
rect 9122 1980 9128 1992
rect 9180 1980 9186 2032
rect 9309 2023 9367 2029
rect 9309 1989 9321 2023
rect 9355 2020 9367 2023
rect 9674 2020 9680 2032
rect 9355 1992 9680 2020
rect 9355 1989 9367 1992
rect 9309 1983 9367 1989
rect 9674 1980 9680 1992
rect 9732 1980 9738 2032
rect 10410 1980 10416 2032
rect 10468 1980 10474 2032
rect 10980 2029 11008 2060
rect 12986 2048 12992 2100
rect 13044 2048 13050 2100
rect 13832 2060 15332 2088
rect 10965 2023 11023 2029
rect 10965 1989 10977 2023
rect 11011 1989 11023 2023
rect 10965 1983 11023 1989
rect 11238 1980 11244 2032
rect 11296 2020 11302 2032
rect 11609 2023 11667 2029
rect 11609 2020 11621 2023
rect 11296 1992 11621 2020
rect 11296 1980 11302 1992
rect 11609 1989 11621 1992
rect 11655 1989 11667 2023
rect 13630 2020 13636 2032
rect 11609 1983 11667 1989
rect 11716 1992 13636 2020
rect 8481 1955 8539 1961
rect 8481 1921 8493 1955
rect 8527 1921 8539 1955
rect 8481 1915 8539 1921
rect 8849 1955 8907 1961
rect 8849 1921 8861 1955
rect 8895 1921 8907 1955
rect 8849 1915 8907 1921
rect 9861 1955 9919 1961
rect 9861 1921 9873 1955
rect 9907 1952 9919 1955
rect 11716 1952 11744 1992
rect 13630 1980 13636 1992
rect 13688 1980 13694 2032
rect 13832 2029 13860 2060
rect 13817 2023 13875 2029
rect 13817 1989 13829 2023
rect 13863 1989 13875 2023
rect 13817 1983 13875 1989
rect 14369 2023 14427 2029
rect 14369 1989 14381 2023
rect 14415 2020 14427 2023
rect 15194 2020 15200 2032
rect 14415 1992 15200 2020
rect 14415 1989 14427 1992
rect 14369 1983 14427 1989
rect 15194 1980 15200 1992
rect 15252 1980 15258 2032
rect 9907 1924 11744 1952
rect 12161 1955 12219 1961
rect 9907 1921 9919 1924
rect 9861 1915 9919 1921
rect 12161 1921 12173 1955
rect 12207 1921 12219 1955
rect 12161 1915 12219 1921
rect 566 1844 572 1896
rect 624 1884 630 1896
rect 624 1856 5120 1884
rect 624 1844 630 1856
rect 290 1776 296 1828
rect 348 1816 354 1828
rect 3142 1816 3148 1828
rect 348 1788 3148 1816
rect 348 1776 354 1788
rect 3142 1776 3148 1788
rect 3200 1776 3206 1828
rect 3694 1776 3700 1828
rect 3752 1776 3758 1828
rect 3973 1819 4031 1825
rect 3973 1785 3985 1819
rect 4019 1816 4031 1819
rect 4982 1816 4988 1828
rect 4019 1788 4988 1816
rect 4019 1785 4031 1788
rect 3973 1779 4031 1785
rect 4982 1776 4988 1788
rect 5040 1776 5046 1828
rect 5092 1825 5120 1856
rect 5258 1844 5264 1896
rect 5316 1844 5322 1896
rect 5442 1844 5448 1896
rect 5500 1884 5506 1896
rect 7653 1887 7711 1893
rect 7653 1884 7665 1887
rect 5500 1856 7665 1884
rect 5500 1844 5506 1856
rect 7653 1853 7665 1856
rect 7699 1853 7711 1887
rect 7653 1847 7711 1853
rect 8018 1844 8024 1896
rect 8076 1884 8082 1896
rect 8864 1884 8892 1915
rect 10134 1884 10140 1896
rect 8076 1856 8892 1884
rect 8956 1856 10140 1884
rect 8076 1844 8082 1856
rect 5077 1819 5135 1825
rect 5077 1785 5089 1819
rect 5123 1785 5135 1819
rect 8956 1816 8984 1856
rect 10134 1844 10140 1856
rect 10192 1844 10198 1896
rect 10502 1844 10508 1896
rect 10560 1884 10566 1896
rect 12176 1884 12204 1915
rect 12710 1912 12716 1964
rect 12768 1952 12774 1964
rect 12805 1955 12863 1961
rect 12805 1952 12817 1955
rect 12768 1924 12817 1952
rect 12768 1912 12774 1924
rect 12805 1921 12817 1924
rect 12851 1921 12863 1955
rect 12805 1915 12863 1921
rect 12894 1912 12900 1964
rect 12952 1952 12958 1964
rect 13265 1955 13323 1961
rect 13265 1952 13277 1955
rect 12952 1924 13277 1952
rect 12952 1912 12958 1924
rect 13265 1921 13277 1924
rect 13311 1921 13323 1955
rect 13265 1915 13323 1921
rect 14918 1912 14924 1964
rect 14976 1912 14982 1964
rect 14458 1884 14464 1896
rect 10560 1856 12204 1884
rect 12406 1856 14464 1884
rect 10560 1844 10566 1856
rect 5077 1779 5135 1785
rect 7116 1788 8984 1816
rect 9033 1819 9091 1825
rect 3712 1748 3740 1776
rect 7116 1748 7144 1788
rect 9033 1785 9045 1819
rect 9079 1816 9091 1819
rect 10042 1816 10048 1828
rect 9079 1788 10048 1816
rect 9079 1785 9091 1788
rect 9033 1779 9091 1785
rect 10042 1776 10048 1788
rect 10100 1776 10106 1828
rect 10594 1816 10600 1828
rect 10244 1788 10600 1816
rect 10244 1760 10272 1788
rect 10594 1776 10600 1788
rect 10652 1776 10658 1828
rect 10778 1776 10784 1828
rect 10836 1816 10842 1828
rect 12406 1816 12434 1856
rect 14458 1844 14464 1856
rect 14516 1844 14522 1896
rect 15304 1884 15332 2060
rect 17126 2048 17132 2100
rect 17184 2088 17190 2100
rect 18874 2088 18880 2100
rect 17184 2060 18880 2088
rect 17184 2048 17190 2060
rect 18874 2048 18880 2060
rect 18932 2048 18938 2100
rect 20901 2091 20959 2097
rect 20901 2057 20913 2091
rect 20947 2088 20959 2091
rect 20990 2088 20996 2100
rect 20947 2060 20996 2088
rect 20947 2057 20959 2060
rect 20901 2051 20959 2057
rect 20990 2048 20996 2060
rect 21048 2048 21054 2100
rect 21269 2091 21327 2097
rect 21269 2057 21281 2091
rect 21315 2088 21327 2091
rect 21358 2088 21364 2100
rect 21315 2060 21364 2088
rect 21315 2057 21327 2060
rect 21269 2051 21327 2057
rect 21358 2048 21364 2060
rect 21416 2048 21422 2100
rect 15470 1980 15476 2032
rect 15528 1980 15534 2032
rect 15746 1980 15752 2032
rect 15804 2020 15810 2032
rect 16025 2023 16083 2029
rect 16025 2020 16037 2023
rect 15804 1992 16037 2020
rect 15804 1980 15810 1992
rect 16025 1989 16037 1992
rect 16071 1989 16083 2023
rect 16025 1983 16083 1989
rect 17034 1980 17040 2032
rect 17092 2020 17098 2032
rect 18782 2020 18788 2032
rect 17092 1992 18788 2020
rect 17092 1980 17098 1992
rect 18782 1980 18788 1992
rect 18840 1980 18846 2032
rect 20346 1980 20352 2032
rect 20404 2020 20410 2032
rect 20441 2023 20499 2029
rect 20441 2020 20453 2023
rect 20404 1992 20453 2020
rect 20404 1980 20410 1992
rect 20441 1989 20453 1992
rect 20487 1989 20499 2023
rect 20441 1983 20499 1989
rect 20809 2023 20867 2029
rect 20809 1989 20821 2023
rect 20855 2020 20867 2023
rect 21450 2020 21456 2032
rect 20855 1992 21456 2020
rect 20855 1989 20867 1992
rect 20809 1983 20867 1989
rect 21450 1980 21456 1992
rect 21508 1980 21514 2032
rect 16669 1955 16727 1961
rect 16669 1921 16681 1955
rect 16715 1952 16727 1955
rect 16850 1952 16856 1964
rect 16715 1924 16856 1952
rect 16715 1921 16727 1924
rect 16669 1915 16727 1921
rect 16850 1912 16856 1924
rect 16908 1912 16914 1964
rect 17126 1912 17132 1964
rect 17184 1952 17190 1964
rect 17773 1955 17831 1961
rect 17773 1952 17785 1955
rect 17184 1924 17785 1952
rect 17184 1912 17190 1924
rect 17773 1921 17785 1924
rect 17819 1921 17831 1955
rect 17773 1915 17831 1921
rect 17862 1912 17868 1964
rect 17920 1952 17926 1964
rect 19613 1955 19671 1961
rect 19613 1952 19625 1955
rect 17920 1924 19625 1952
rect 17920 1912 17926 1924
rect 19613 1921 19625 1924
rect 19659 1921 19671 1955
rect 19613 1915 19671 1921
rect 20714 1912 20720 1964
rect 20772 1952 20778 1964
rect 21177 1955 21235 1961
rect 21177 1952 21189 1955
rect 20772 1924 21189 1952
rect 20772 1912 20778 1924
rect 21177 1921 21189 1924
rect 21223 1921 21235 1955
rect 21177 1915 21235 1921
rect 15304 1856 16252 1884
rect 10836 1788 12434 1816
rect 10836 1776 10842 1788
rect 14366 1776 14372 1828
rect 14424 1816 14430 1828
rect 14424 1788 14596 1816
rect 14424 1776 14430 1788
rect 3712 1720 7144 1748
rect 7190 1708 7196 1760
rect 7248 1708 7254 1760
rect 7650 1708 7656 1760
rect 7708 1748 7714 1760
rect 7929 1751 7987 1757
rect 7929 1748 7941 1751
rect 7708 1720 7941 1748
rect 7708 1708 7714 1720
rect 7929 1717 7941 1720
rect 7975 1717 7987 1751
rect 7929 1711 7987 1717
rect 8297 1751 8355 1757
rect 8297 1717 8309 1751
rect 8343 1748 8355 1751
rect 8754 1748 8760 1760
rect 8343 1720 8760 1748
rect 8343 1717 8355 1720
rect 8297 1711 8355 1717
rect 8754 1708 8760 1720
rect 8812 1708 8818 1760
rect 9582 1708 9588 1760
rect 9640 1708 9646 1760
rect 10134 1708 10140 1760
rect 10192 1708 10198 1760
rect 10226 1708 10232 1760
rect 10284 1708 10290 1760
rect 10502 1708 10508 1760
rect 10560 1708 10566 1760
rect 11054 1708 11060 1760
rect 11112 1708 11118 1760
rect 11238 1708 11244 1760
rect 11296 1748 11302 1760
rect 11701 1751 11759 1757
rect 11701 1748 11713 1751
rect 11296 1720 11713 1748
rect 11296 1708 11302 1720
rect 11701 1717 11713 1720
rect 11747 1717 11759 1751
rect 11701 1711 11759 1717
rect 11974 1708 11980 1760
rect 12032 1748 12038 1760
rect 12253 1751 12311 1757
rect 12253 1748 12265 1751
rect 12032 1720 12265 1748
rect 12032 1708 12038 1720
rect 12253 1717 12265 1720
rect 12299 1717 12311 1751
rect 12253 1711 12311 1717
rect 13078 1708 13084 1760
rect 13136 1748 13142 1760
rect 13357 1751 13415 1757
rect 13357 1748 13369 1751
rect 13136 1720 13369 1748
rect 13136 1708 13142 1720
rect 13357 1717 13369 1720
rect 13403 1717 13415 1751
rect 13357 1711 13415 1717
rect 13446 1708 13452 1760
rect 13504 1748 13510 1760
rect 13909 1751 13967 1757
rect 13909 1748 13921 1751
rect 13504 1720 13921 1748
rect 13504 1708 13510 1720
rect 13909 1717 13921 1720
rect 13955 1717 13967 1751
rect 13909 1711 13967 1717
rect 14090 1708 14096 1760
rect 14148 1748 14154 1760
rect 14461 1751 14519 1757
rect 14461 1748 14473 1751
rect 14148 1720 14473 1748
rect 14148 1708 14154 1720
rect 14461 1717 14473 1720
rect 14507 1717 14519 1751
rect 14568 1748 14596 1788
rect 14642 1776 14648 1828
rect 14700 1816 14706 1828
rect 14700 1788 15608 1816
rect 14700 1776 14706 1788
rect 15580 1757 15608 1788
rect 15013 1751 15071 1757
rect 15013 1748 15025 1751
rect 14568 1720 15025 1748
rect 14461 1711 14519 1717
rect 15013 1717 15025 1720
rect 15059 1717 15071 1751
rect 15013 1711 15071 1717
rect 15565 1751 15623 1757
rect 15565 1717 15577 1751
rect 15611 1717 15623 1751
rect 15565 1711 15623 1717
rect 15746 1708 15752 1760
rect 15804 1748 15810 1760
rect 16117 1751 16175 1757
rect 16117 1748 16129 1751
rect 15804 1720 16129 1748
rect 15804 1708 15810 1720
rect 16117 1717 16129 1720
rect 16163 1717 16175 1751
rect 16224 1748 16252 1856
rect 17034 1844 17040 1896
rect 17092 1844 17098 1896
rect 18322 1844 18328 1896
rect 18380 1844 18386 1896
rect 19521 1887 19579 1893
rect 19521 1853 19533 1887
rect 19567 1884 19579 1887
rect 22830 1884 22836 1896
rect 19567 1856 22836 1884
rect 19567 1853 19579 1856
rect 19521 1847 19579 1853
rect 22830 1844 22836 1856
rect 22888 1844 22894 1896
rect 18340 1748 18368 1844
rect 16224 1720 18368 1748
rect 16117 1711 16175 1717
rect 1104 1658 21896 1680
rect 1104 1606 3549 1658
rect 3601 1606 3613 1658
rect 3665 1606 3677 1658
rect 3729 1606 3741 1658
rect 3793 1606 3805 1658
rect 3857 1606 8747 1658
rect 8799 1606 8811 1658
rect 8863 1606 8875 1658
rect 8927 1606 8939 1658
rect 8991 1606 9003 1658
rect 9055 1606 13945 1658
rect 13997 1606 14009 1658
rect 14061 1606 14073 1658
rect 14125 1606 14137 1658
rect 14189 1606 14201 1658
rect 14253 1606 19143 1658
rect 19195 1606 19207 1658
rect 19259 1606 19271 1658
rect 19323 1606 19335 1658
rect 19387 1606 19399 1658
rect 19451 1606 21896 1658
rect 1104 1584 21896 1606
rect 1578 1504 1584 1556
rect 1636 1504 1642 1556
rect 5353 1547 5411 1553
rect 5353 1544 5365 1547
rect 2608 1516 5365 1544
rect 382 1300 388 1352
rect 440 1340 446 1352
rect 2608 1340 2636 1516
rect 5353 1513 5365 1516
rect 5399 1513 5411 1547
rect 5353 1507 5411 1513
rect 5810 1504 5816 1556
rect 5868 1544 5874 1556
rect 6089 1547 6147 1553
rect 6089 1544 6101 1547
rect 5868 1516 6101 1544
rect 5868 1504 5874 1516
rect 6089 1513 6101 1516
rect 6135 1513 6147 1547
rect 6089 1507 6147 1513
rect 6638 1504 6644 1556
rect 6696 1504 6702 1556
rect 7098 1504 7104 1556
rect 7156 1544 7162 1556
rect 7558 1544 7564 1556
rect 7156 1516 7564 1544
rect 7156 1504 7162 1516
rect 7558 1504 7564 1516
rect 7616 1504 7622 1556
rect 8018 1504 8024 1556
rect 8076 1504 8082 1556
rect 9030 1504 9036 1556
rect 9088 1544 9094 1556
rect 9306 1544 9312 1556
rect 9088 1516 9312 1544
rect 9088 1504 9094 1516
rect 9306 1504 9312 1516
rect 9364 1504 9370 1556
rect 10962 1544 10968 1556
rect 9600 1516 10968 1544
rect 3142 1436 3148 1488
rect 3200 1476 3206 1488
rect 9600 1476 9628 1516
rect 10962 1504 10968 1516
rect 11020 1504 11026 1556
rect 12342 1504 12348 1556
rect 12400 1544 12406 1556
rect 12437 1547 12495 1553
rect 12437 1544 12449 1547
rect 12400 1516 12449 1544
rect 12400 1504 12406 1516
rect 12437 1513 12449 1516
rect 12483 1513 12495 1547
rect 12437 1507 12495 1513
rect 13262 1504 13268 1556
rect 13320 1544 13326 1556
rect 14277 1547 14335 1553
rect 14277 1544 14289 1547
rect 13320 1516 14289 1544
rect 13320 1504 13326 1516
rect 14277 1513 14289 1516
rect 14323 1513 14335 1547
rect 14277 1507 14335 1513
rect 14829 1547 14887 1553
rect 14829 1513 14841 1547
rect 14875 1513 14887 1547
rect 14829 1507 14887 1513
rect 3200 1448 9628 1476
rect 9677 1479 9735 1485
rect 3200 1436 3206 1448
rect 9677 1445 9689 1479
rect 9723 1476 9735 1479
rect 9723 1448 11008 1476
rect 9723 1445 9735 1448
rect 9677 1439 9735 1445
rect 3326 1408 3332 1420
rect 2976 1380 3332 1408
rect 2774 1340 2780 1352
rect 440 1312 2636 1340
rect 2700 1312 2780 1340
rect 440 1300 446 1312
rect 1486 1232 1492 1284
rect 1544 1232 1550 1284
rect 2317 1275 2375 1281
rect 2317 1241 2329 1275
rect 2363 1272 2375 1275
rect 2590 1272 2596 1284
rect 2363 1244 2596 1272
rect 2363 1241 2375 1244
rect 2317 1235 2375 1241
rect 2590 1232 2596 1244
rect 2648 1232 2654 1284
rect 2700 1281 2728 1312
rect 2774 1300 2780 1312
rect 2832 1300 2838 1352
rect 2869 1343 2927 1349
rect 2869 1309 2881 1343
rect 2915 1340 2927 1343
rect 2976 1340 3004 1380
rect 3326 1368 3332 1380
rect 3384 1368 3390 1420
rect 4246 1368 4252 1420
rect 4304 1408 4310 1420
rect 4341 1411 4399 1417
rect 4341 1408 4353 1411
rect 4304 1380 4353 1408
rect 4304 1368 4310 1380
rect 4341 1377 4353 1380
rect 4387 1377 4399 1411
rect 4341 1371 4399 1377
rect 8665 1411 8723 1417
rect 8665 1377 8677 1411
rect 8711 1408 8723 1411
rect 10042 1408 10048 1420
rect 8711 1380 10048 1408
rect 8711 1377 8723 1380
rect 8665 1371 8723 1377
rect 10042 1368 10048 1380
rect 10100 1368 10106 1420
rect 10229 1411 10287 1417
rect 10229 1377 10241 1411
rect 10275 1408 10287 1411
rect 10410 1408 10416 1420
rect 10275 1380 10416 1408
rect 10275 1377 10287 1380
rect 10229 1371 10287 1377
rect 10410 1368 10416 1380
rect 10468 1368 10474 1420
rect 3694 1340 3700 1352
rect 2915 1312 3004 1340
rect 3068 1312 3700 1340
rect 2915 1309 2927 1312
rect 2869 1303 2927 1309
rect 3068 1281 3096 1312
rect 3694 1300 3700 1312
rect 3752 1300 3758 1352
rect 4433 1343 4491 1349
rect 4433 1309 4445 1343
rect 4479 1340 4491 1343
rect 4522 1340 4528 1352
rect 4479 1312 4528 1340
rect 4479 1309 4491 1312
rect 4433 1303 4491 1309
rect 4522 1300 4528 1312
rect 4580 1300 4586 1352
rect 4982 1340 4988 1352
rect 4816 1312 4988 1340
rect 2685 1275 2743 1281
rect 2685 1241 2697 1275
rect 2731 1241 2743 1275
rect 2685 1235 2743 1241
rect 3053 1275 3111 1281
rect 3053 1241 3065 1275
rect 3099 1241 3111 1275
rect 3053 1235 3111 1241
rect 3237 1275 3295 1281
rect 3237 1241 3249 1275
rect 3283 1272 3295 1275
rect 3326 1272 3332 1284
rect 3283 1244 3332 1272
rect 3283 1241 3295 1244
rect 3237 1235 3295 1241
rect 3326 1232 3332 1244
rect 3384 1232 3390 1284
rect 3421 1275 3479 1281
rect 3421 1241 3433 1275
rect 3467 1272 3479 1275
rect 4157 1275 4215 1281
rect 3467 1244 4108 1272
rect 3467 1241 3479 1244
rect 3421 1235 3479 1241
rect 2409 1207 2467 1213
rect 2409 1173 2421 1207
rect 2455 1204 2467 1207
rect 2498 1204 2504 1216
rect 2455 1176 2504 1204
rect 2455 1173 2467 1176
rect 2409 1167 2467 1173
rect 2498 1164 2504 1176
rect 2556 1164 2562 1216
rect 3510 1164 3516 1216
rect 3568 1164 3574 1216
rect 4080 1204 4108 1244
rect 4157 1241 4169 1275
rect 4203 1272 4215 1275
rect 4816 1272 4844 1312
rect 4982 1300 4988 1312
rect 5040 1300 5046 1352
rect 5074 1300 5080 1352
rect 5132 1300 5138 1352
rect 5184 1349 5304 1356
rect 5169 1343 5304 1349
rect 5169 1309 5181 1343
rect 5215 1340 5304 1343
rect 5350 1340 5356 1352
rect 5215 1328 5356 1340
rect 5215 1309 5227 1328
rect 5276 1312 5356 1328
rect 5169 1303 5227 1309
rect 5350 1300 5356 1312
rect 5408 1300 5414 1352
rect 5534 1300 5540 1352
rect 5592 1340 5598 1352
rect 5813 1343 5871 1349
rect 5813 1340 5825 1343
rect 5592 1312 5825 1340
rect 5592 1300 5598 1312
rect 5813 1309 5825 1312
rect 5859 1309 5871 1343
rect 6822 1340 6828 1352
rect 5813 1303 5871 1309
rect 5920 1312 6828 1340
rect 4203 1244 4844 1272
rect 4893 1275 4951 1281
rect 4203 1241 4215 1244
rect 4157 1235 4215 1241
rect 4893 1241 4905 1275
rect 4939 1272 4951 1275
rect 5442 1272 5448 1284
rect 4939 1244 5448 1272
rect 4939 1241 4951 1244
rect 4893 1235 4951 1241
rect 5442 1232 5448 1244
rect 5500 1232 5506 1284
rect 5629 1275 5687 1281
rect 5629 1241 5641 1275
rect 5675 1272 5687 1275
rect 5920 1272 5948 1312
rect 6822 1300 6828 1312
rect 6880 1300 6886 1352
rect 7098 1300 7104 1352
rect 7156 1300 7162 1352
rect 7374 1300 7380 1352
rect 7432 1300 7438 1352
rect 8202 1300 8208 1352
rect 8260 1300 8266 1352
rect 8570 1300 8576 1352
rect 8628 1340 8634 1352
rect 8941 1343 8999 1349
rect 8941 1340 8953 1343
rect 8628 1312 8953 1340
rect 8628 1300 8634 1312
rect 8941 1309 8953 1312
rect 8987 1309 8999 1343
rect 8941 1303 8999 1309
rect 9398 1300 9404 1352
rect 9456 1300 9462 1352
rect 9858 1300 9864 1352
rect 9916 1340 9922 1352
rect 9953 1343 10011 1349
rect 9953 1340 9965 1343
rect 9916 1312 9965 1340
rect 9916 1300 9922 1312
rect 9953 1309 9965 1312
rect 9999 1309 10011 1343
rect 9953 1303 10011 1309
rect 10594 1300 10600 1352
rect 10652 1340 10658 1352
rect 10781 1343 10839 1349
rect 10781 1340 10793 1343
rect 10652 1312 10793 1340
rect 10652 1300 10658 1312
rect 10781 1309 10793 1312
rect 10827 1309 10839 1343
rect 10781 1303 10839 1309
rect 5675 1244 5948 1272
rect 5997 1275 6055 1281
rect 5675 1241 5687 1244
rect 5629 1235 5687 1241
rect 5997 1241 6009 1275
rect 6043 1272 6055 1275
rect 6043 1244 6500 1272
rect 6043 1241 6055 1244
rect 5997 1235 6055 1241
rect 4246 1204 4252 1216
rect 4080 1176 4252 1204
rect 4246 1164 4252 1176
rect 4304 1164 4310 1216
rect 4617 1207 4675 1213
rect 4617 1173 4629 1207
rect 4663 1204 4675 1207
rect 4798 1204 4804 1216
rect 4663 1176 4804 1204
rect 4663 1173 4675 1176
rect 4617 1167 4675 1173
rect 4798 1164 4804 1176
rect 4856 1164 4862 1216
rect 6472 1204 6500 1244
rect 6546 1232 6552 1284
rect 6604 1232 6610 1284
rect 7282 1232 7288 1284
rect 7340 1272 7346 1284
rect 7834 1272 7840 1284
rect 7340 1244 7840 1272
rect 7340 1232 7346 1244
rect 7834 1232 7840 1244
rect 7892 1232 7898 1284
rect 8386 1232 8392 1284
rect 8444 1232 8450 1284
rect 8662 1232 8668 1284
rect 8720 1272 8726 1284
rect 9030 1272 9036 1284
rect 8720 1244 9036 1272
rect 8720 1232 8726 1244
rect 9030 1232 9036 1244
rect 9088 1232 9094 1284
rect 10686 1272 10692 1284
rect 9140 1244 10692 1272
rect 7190 1204 7196 1216
rect 6472 1176 7196 1204
rect 7190 1164 7196 1176
rect 7248 1164 7254 1216
rect 9140 1213 9168 1244
rect 10686 1232 10692 1244
rect 10744 1232 10750 1284
rect 10980 1272 11008 1448
rect 11698 1436 11704 1488
rect 11756 1476 11762 1488
rect 11756 1448 12388 1476
rect 11756 1436 11762 1448
rect 11057 1411 11115 1417
rect 11057 1377 11069 1411
rect 11103 1408 11115 1411
rect 11146 1408 11152 1420
rect 11103 1380 11152 1408
rect 11103 1377 11115 1380
rect 11057 1371 11115 1377
rect 11146 1368 11152 1380
rect 11204 1368 11210 1420
rect 11624 1380 12020 1408
rect 11517 1343 11575 1349
rect 11517 1309 11529 1343
rect 11563 1340 11575 1343
rect 11624 1340 11652 1380
rect 11885 1343 11943 1349
rect 11885 1340 11897 1343
rect 11563 1312 11652 1340
rect 11716 1312 11897 1340
rect 11563 1309 11575 1312
rect 11517 1303 11575 1309
rect 11054 1272 11060 1284
rect 10980 1244 11060 1272
rect 11054 1232 11060 1244
rect 11112 1232 11118 1284
rect 11716 1272 11744 1312
rect 11885 1309 11897 1312
rect 11931 1309 11943 1343
rect 11992 1340 12020 1380
rect 12066 1340 12072 1352
rect 11992 1312 12072 1340
rect 11885 1303 11943 1309
rect 12066 1300 12072 1312
rect 12124 1300 12130 1352
rect 12360 1281 12388 1448
rect 13630 1436 13636 1488
rect 13688 1476 13694 1488
rect 14844 1476 14872 1507
rect 15194 1504 15200 1556
rect 15252 1504 15258 1556
rect 16850 1504 16856 1556
rect 16908 1504 16914 1556
rect 18785 1547 18843 1553
rect 18785 1513 18797 1547
rect 18831 1544 18843 1547
rect 22094 1544 22100 1556
rect 18831 1516 22100 1544
rect 18831 1513 18843 1516
rect 18785 1507 18843 1513
rect 22094 1504 22100 1516
rect 22152 1504 22158 1556
rect 13688 1448 14872 1476
rect 13688 1436 13694 1448
rect 14918 1436 14924 1488
rect 14976 1476 14982 1488
rect 16114 1476 16120 1488
rect 14976 1448 16120 1476
rect 14976 1436 14982 1448
rect 16114 1436 16120 1448
rect 16172 1436 16178 1488
rect 12434 1368 12440 1420
rect 12492 1408 12498 1420
rect 12492 1380 13584 1408
rect 12492 1368 12498 1380
rect 12802 1300 12808 1352
rect 12860 1300 12866 1352
rect 13170 1300 13176 1352
rect 13228 1300 13234 1352
rect 13354 1300 13360 1352
rect 13412 1340 13418 1352
rect 13556 1349 13584 1380
rect 13998 1368 14004 1420
rect 14056 1408 14062 1420
rect 15102 1408 15108 1420
rect 14056 1380 15108 1408
rect 14056 1368 14062 1380
rect 15102 1368 15108 1380
rect 15160 1368 15166 1420
rect 15841 1411 15899 1417
rect 15841 1408 15853 1411
rect 15212 1380 15853 1408
rect 13541 1343 13599 1349
rect 13412 1312 13492 1340
rect 13412 1300 13418 1312
rect 11624 1244 11744 1272
rect 12345 1275 12403 1281
rect 9125 1207 9183 1213
rect 9125 1173 9137 1207
rect 9171 1173 9183 1207
rect 9125 1167 9183 1173
rect 9398 1164 9404 1216
rect 9456 1204 9462 1216
rect 9766 1204 9772 1216
rect 9456 1176 9772 1204
rect 9456 1164 9462 1176
rect 9766 1164 9772 1176
rect 9824 1164 9830 1216
rect 9858 1164 9864 1216
rect 9916 1204 9922 1216
rect 11624 1204 11652 1244
rect 12345 1241 12357 1275
rect 12391 1241 12403 1275
rect 12345 1235 12403 1241
rect 12710 1232 12716 1284
rect 12768 1272 12774 1284
rect 13464 1272 13492 1312
rect 13541 1309 13553 1343
rect 13587 1309 13599 1343
rect 13541 1303 13599 1309
rect 13814 1300 13820 1352
rect 13872 1340 13878 1352
rect 14185 1343 14243 1349
rect 14185 1340 14197 1343
rect 13872 1312 14197 1340
rect 13872 1300 13878 1312
rect 14185 1309 14197 1312
rect 14231 1309 14243 1343
rect 14185 1303 14243 1309
rect 14734 1300 14740 1352
rect 14792 1300 14798 1352
rect 15212 1272 15240 1380
rect 15841 1377 15853 1380
rect 15887 1377 15899 1411
rect 15841 1371 15899 1377
rect 15930 1368 15936 1420
rect 15988 1408 15994 1420
rect 16298 1408 16304 1420
rect 15988 1380 16304 1408
rect 15988 1368 15994 1380
rect 16298 1368 16304 1380
rect 16356 1368 16362 1420
rect 17954 1368 17960 1420
rect 18012 1408 18018 1420
rect 18506 1408 18512 1420
rect 18012 1380 18512 1408
rect 18012 1368 18018 1380
rect 18506 1368 18512 1380
rect 18564 1368 18570 1420
rect 15378 1300 15384 1352
rect 15436 1300 15442 1352
rect 15657 1343 15715 1349
rect 15657 1309 15669 1343
rect 15703 1309 15715 1343
rect 15657 1303 15715 1309
rect 12768 1244 13400 1272
rect 13464 1244 15240 1272
rect 12768 1232 12774 1244
rect 9916 1176 11652 1204
rect 9916 1164 9922 1176
rect 11698 1164 11704 1216
rect 11756 1164 11762 1216
rect 12066 1164 12072 1216
rect 12124 1164 12130 1216
rect 12526 1164 12532 1216
rect 12584 1204 12590 1216
rect 13372 1213 13400 1244
rect 12989 1207 13047 1213
rect 12989 1204 13001 1207
rect 12584 1176 13001 1204
rect 12584 1164 12590 1176
rect 12989 1173 13001 1176
rect 13035 1173 13047 1207
rect 12989 1167 13047 1173
rect 13357 1207 13415 1213
rect 13357 1173 13369 1207
rect 13403 1173 13415 1207
rect 13357 1167 13415 1173
rect 13722 1164 13728 1216
rect 13780 1164 13786 1216
rect 15672 1204 15700 1303
rect 16390 1300 16396 1352
rect 16448 1340 16454 1352
rect 16761 1343 16819 1349
rect 16761 1340 16773 1343
rect 16448 1312 16773 1340
rect 16448 1300 16454 1312
rect 16761 1309 16773 1312
rect 16807 1309 16819 1343
rect 16761 1303 16819 1309
rect 18690 1300 18696 1352
rect 18748 1340 18754 1352
rect 19337 1343 19395 1349
rect 19337 1340 19349 1343
rect 18748 1312 19349 1340
rect 18748 1300 18754 1312
rect 19337 1309 19349 1312
rect 19383 1309 19395 1343
rect 20349 1343 20407 1349
rect 20349 1340 20361 1343
rect 19337 1303 19395 1309
rect 19444 1312 20361 1340
rect 16408 1244 16988 1272
rect 16408 1204 16436 1244
rect 15672 1176 16436 1204
rect 16960 1204 16988 1244
rect 17034 1232 17040 1284
rect 17092 1272 17098 1284
rect 17313 1275 17371 1281
rect 17313 1272 17325 1275
rect 17092 1244 17325 1272
rect 17092 1232 17098 1244
rect 17313 1241 17325 1244
rect 17359 1241 17371 1275
rect 17313 1235 17371 1241
rect 17678 1232 17684 1284
rect 17736 1272 17742 1284
rect 19444 1272 19472 1312
rect 20349 1309 20361 1312
rect 20395 1309 20407 1343
rect 20349 1303 20407 1309
rect 21177 1343 21235 1349
rect 21177 1309 21189 1343
rect 21223 1340 21235 1343
rect 22738 1340 22744 1352
rect 21223 1312 22744 1340
rect 21223 1309 21235 1312
rect 21177 1303 21235 1309
rect 22738 1300 22744 1312
rect 22796 1300 22802 1352
rect 17736 1244 19472 1272
rect 20073 1275 20131 1281
rect 17736 1232 17742 1244
rect 20073 1241 20085 1275
rect 20119 1272 20131 1275
rect 22186 1272 22192 1284
rect 20119 1244 22192 1272
rect 20119 1241 20131 1244
rect 20073 1235 20131 1241
rect 22186 1232 22192 1244
rect 22244 1232 22250 1284
rect 17402 1204 17408 1216
rect 16960 1176 17408 1204
rect 17402 1164 17408 1176
rect 17460 1164 17466 1216
rect 18138 1164 18144 1216
rect 18196 1204 18202 1216
rect 18598 1204 18604 1216
rect 18196 1176 18604 1204
rect 18196 1164 18202 1176
rect 18598 1164 18604 1176
rect 18656 1164 18662 1216
rect 1104 1114 22056 1136
rect 1104 1062 6148 1114
rect 6200 1062 6212 1114
rect 6264 1062 6276 1114
rect 6328 1062 6340 1114
rect 6392 1062 6404 1114
rect 6456 1062 11346 1114
rect 11398 1062 11410 1114
rect 11462 1062 11474 1114
rect 11526 1062 11538 1114
rect 11590 1062 11602 1114
rect 11654 1062 16544 1114
rect 16596 1062 16608 1114
rect 16660 1062 16672 1114
rect 16724 1062 16736 1114
rect 16788 1062 16800 1114
rect 16852 1062 21742 1114
rect 21794 1062 21806 1114
rect 21858 1062 21870 1114
rect 21922 1062 21934 1114
rect 21986 1062 21998 1114
rect 22050 1062 22056 1114
rect 1104 1040 22056 1062
rect 2498 960 2504 1012
rect 2556 1000 2562 1012
rect 4338 1000 4344 1012
rect 2556 972 4344 1000
rect 2556 960 2562 972
rect 4338 960 4344 972
rect 4396 960 4402 1012
rect 6454 960 6460 1012
rect 6512 1000 6518 1012
rect 6730 1000 6736 1012
rect 6512 972 6736 1000
rect 6512 960 6518 972
rect 6730 960 6736 972
rect 6788 960 6794 1012
rect 6914 960 6920 1012
rect 6972 1000 6978 1012
rect 9858 1000 9864 1012
rect 6972 972 9864 1000
rect 6972 960 6978 972
rect 9858 960 9864 972
rect 9916 960 9922 1012
rect 14458 960 14464 1012
rect 14516 1000 14522 1012
rect 17494 1000 17500 1012
rect 14516 972 17500 1000
rect 14516 960 14522 972
rect 17494 960 17500 972
rect 17552 960 17558 1012
rect 22922 960 22928 1012
rect 22980 960 22986 1012
rect 842 892 848 944
rect 900 932 906 944
rect 4706 932 4712 944
rect 900 904 4712 932
rect 900 892 906 904
rect 4706 892 4712 904
rect 4764 892 4770 944
rect 8386 892 8392 944
rect 8444 932 8450 944
rect 9398 932 9404 944
rect 8444 904 9404 932
rect 8444 892 8450 904
rect 9398 892 9404 904
rect 9456 892 9462 944
rect 11790 892 11796 944
rect 11848 932 11854 944
rect 22940 932 22968 960
rect 11848 904 22968 932
rect 11848 892 11854 904
rect 11514 756 11520 808
rect 11572 796 11578 808
rect 11882 796 11888 808
rect 11572 768 11888 796
rect 11572 756 11578 768
rect 11882 756 11888 768
rect 11940 756 11946 808
rect 2774 688 2780 740
rect 2832 728 2838 740
rect 3326 728 3332 740
rect 2832 700 3332 728
rect 2832 688 2838 700
rect 3326 688 3332 700
rect 3384 688 3390 740
rect 4522 688 4528 740
rect 4580 728 4586 740
rect 5718 728 5724 740
rect 4580 700 5724 728
rect 4580 688 4586 700
rect 5718 688 5724 700
rect 5776 688 5782 740
rect 5442 620 5448 672
rect 5500 660 5506 672
rect 6178 660 6184 672
rect 5500 632 6184 660
rect 5500 620 5506 632
rect 6178 620 6184 632
rect 6236 620 6242 672
rect 9950 620 9956 672
rect 10008 660 10014 672
rect 10410 660 10416 672
rect 10008 632 10416 660
rect 10008 620 10014 632
rect 10410 620 10416 632
rect 10468 620 10474 672
rect 12894 620 12900 672
rect 12952 660 12958 672
rect 13722 660 13728 672
rect 12952 632 13728 660
rect 12952 620 12958 632
rect 13722 620 13728 632
rect 13780 620 13786 672
<< via1 >>
rect 13360 43868 13412 43920
rect 15200 43868 15252 43920
rect 16948 43868 17000 43920
rect 17408 43868 17460 43920
rect 5080 43800 5132 43852
rect 6276 43800 6328 43852
rect 16764 43800 16816 43852
rect 17776 43800 17828 43852
rect 1400 43732 1452 43784
rect 12164 43732 12216 43784
rect 12348 43732 12400 43784
rect 12440 43596 12492 43648
rect 18972 43596 19024 43648
rect 20812 43596 20864 43648
rect 6148 43494 6200 43546
rect 6212 43494 6264 43546
rect 6276 43494 6328 43546
rect 6340 43494 6392 43546
rect 6404 43494 6456 43546
rect 11346 43494 11398 43546
rect 11410 43494 11462 43546
rect 11474 43494 11526 43546
rect 11538 43494 11590 43546
rect 11602 43494 11654 43546
rect 16544 43494 16596 43546
rect 16608 43494 16660 43546
rect 16672 43494 16724 43546
rect 16736 43494 16788 43546
rect 16800 43494 16852 43546
rect 21742 43494 21794 43546
rect 21806 43494 21858 43546
rect 21870 43494 21922 43546
rect 21934 43494 21986 43546
rect 21998 43494 22050 43546
rect 2228 43435 2280 43444
rect 2228 43401 2237 43435
rect 2237 43401 2271 43435
rect 2271 43401 2280 43435
rect 2228 43392 2280 43401
rect 3148 43435 3200 43444
rect 3148 43401 3157 43435
rect 3157 43401 3191 43435
rect 3191 43401 3200 43435
rect 3148 43392 3200 43401
rect 3332 43392 3384 43444
rect 5172 43392 5224 43444
rect 5264 43435 5316 43444
rect 5264 43401 5273 43435
rect 5273 43401 5307 43435
rect 5307 43401 5316 43435
rect 5264 43392 5316 43401
rect 5448 43392 5500 43444
rect 5816 43435 5868 43444
rect 5816 43401 5825 43435
rect 5825 43401 5859 43435
rect 5859 43401 5868 43435
rect 5816 43392 5868 43401
rect 7380 43392 7432 43444
rect 8576 43392 8628 43444
rect 9036 43392 9088 43444
rect 9404 43392 9456 43444
rect 10048 43392 10100 43444
rect 12440 43435 12492 43444
rect 12440 43401 12449 43435
rect 12449 43401 12483 43435
rect 12483 43401 12492 43435
rect 12440 43392 12492 43401
rect 13728 43392 13780 43444
rect 8392 43324 8444 43376
rect 9772 43367 9824 43376
rect 9772 43333 9781 43367
rect 9781 43333 9815 43367
rect 9815 43333 9824 43367
rect 9772 43324 9824 43333
rect 10324 43367 10376 43376
rect 10324 43333 10333 43367
rect 10333 43333 10367 43367
rect 10367 43333 10376 43367
rect 10324 43324 10376 43333
rect 10876 43367 10928 43376
rect 10876 43333 10885 43367
rect 10885 43333 10919 43367
rect 10919 43333 10928 43367
rect 10876 43324 10928 43333
rect 12348 43367 12400 43376
rect 12348 43333 12357 43367
rect 12357 43333 12391 43367
rect 12391 43333 12400 43367
rect 12348 43324 12400 43333
rect 12900 43367 12952 43376
rect 12900 43333 12909 43367
rect 12909 43333 12943 43367
rect 12943 43333 12952 43367
rect 12900 43324 12952 43333
rect 13084 43324 13136 43376
rect 13912 43435 13964 43444
rect 13912 43401 13921 43435
rect 13921 43401 13955 43435
rect 13955 43401 13964 43435
rect 13912 43392 13964 43401
rect 14280 43392 14332 43444
rect 2044 43299 2096 43308
rect 2044 43265 2053 43299
rect 2053 43265 2087 43299
rect 2087 43265 2096 43299
rect 2044 43256 2096 43265
rect 2504 43299 2556 43308
rect 2504 43265 2513 43299
rect 2513 43265 2547 43299
rect 2547 43265 2556 43299
rect 2504 43256 2556 43265
rect 3056 43299 3108 43308
rect 3056 43265 3065 43299
rect 3065 43265 3099 43299
rect 3099 43265 3108 43299
rect 3056 43256 3108 43265
rect 3976 43256 4028 43308
rect 4344 43256 4396 43308
rect 2596 43188 2648 43240
rect 2964 43120 3016 43172
rect 4160 43120 4212 43172
rect 4712 43256 4764 43308
rect 5540 43256 5592 43308
rect 5080 43188 5132 43240
rect 7380 43256 7432 43308
rect 7656 43256 7708 43308
rect 7472 43120 7524 43172
rect 8944 43299 8996 43308
rect 8944 43265 8953 43299
rect 8953 43265 8987 43299
rect 8987 43265 8996 43299
rect 8944 43256 8996 43265
rect 9680 43256 9732 43308
rect 11612 43256 11664 43308
rect 11888 43256 11940 43308
rect 12072 43256 12124 43308
rect 13360 43256 13412 43308
rect 10600 43188 10652 43240
rect 13268 43188 13320 43240
rect 14740 43256 14792 43308
rect 15292 43299 15344 43308
rect 15292 43265 15301 43299
rect 15301 43265 15335 43299
rect 15335 43265 15344 43299
rect 15292 43256 15344 43265
rect 15568 43299 15620 43308
rect 15568 43265 15577 43299
rect 15577 43265 15611 43299
rect 15611 43265 15620 43299
rect 15568 43256 15620 43265
rect 15660 43256 15712 43308
rect 16120 43299 16172 43308
rect 16120 43265 16129 43299
rect 16129 43265 16163 43299
rect 16163 43265 16172 43299
rect 16120 43256 16172 43265
rect 16580 43392 16632 43444
rect 16948 43392 17000 43444
rect 17776 43435 17828 43444
rect 17776 43401 17785 43435
rect 17785 43401 17819 43435
rect 17819 43401 17828 43435
rect 17776 43392 17828 43401
rect 17316 43324 17368 43376
rect 18420 43392 18472 43444
rect 14280 43188 14332 43240
rect 14648 43188 14700 43240
rect 16304 43188 16356 43240
rect 17776 43256 17828 43308
rect 18420 43256 18472 43308
rect 18604 43299 18656 43308
rect 18604 43265 18613 43299
rect 18613 43265 18647 43299
rect 18647 43265 18656 43299
rect 18604 43256 18656 43265
rect 20720 43324 20772 43376
rect 20812 43367 20864 43376
rect 20812 43333 20821 43367
rect 20821 43333 20855 43367
rect 20855 43333 20864 43367
rect 20812 43324 20864 43333
rect 17316 43188 17368 43240
rect 18512 43188 18564 43240
rect 20996 43299 21048 43308
rect 20996 43265 21005 43299
rect 21005 43265 21039 43299
rect 21039 43265 21048 43299
rect 20996 43256 21048 43265
rect 21640 43188 21692 43240
rect 8484 43120 8536 43172
rect 8576 43120 8628 43172
rect 8116 43052 8168 43104
rect 8208 43052 8260 43104
rect 10232 43120 10284 43172
rect 13084 43163 13136 43172
rect 13084 43129 13093 43163
rect 13093 43129 13127 43163
rect 13127 43129 13136 43163
rect 13084 43120 13136 43129
rect 13452 43163 13504 43172
rect 13452 43129 13461 43163
rect 13461 43129 13495 43163
rect 13495 43129 13504 43163
rect 13452 43120 13504 43129
rect 13544 43120 13596 43172
rect 17684 43120 17736 43172
rect 10784 43052 10836 43104
rect 11152 43095 11204 43104
rect 11152 43061 11161 43095
rect 11161 43061 11195 43095
rect 11195 43061 11204 43095
rect 11152 43052 11204 43061
rect 11704 43052 11756 43104
rect 13360 43052 13412 43104
rect 14648 43095 14700 43104
rect 14648 43061 14657 43095
rect 14657 43061 14691 43095
rect 14691 43061 14700 43095
rect 14648 43052 14700 43061
rect 14832 43095 14884 43104
rect 14832 43061 14841 43095
rect 14841 43061 14875 43095
rect 14875 43061 14884 43095
rect 14832 43052 14884 43061
rect 15292 43052 15344 43104
rect 15384 43095 15436 43104
rect 15384 43061 15393 43095
rect 15393 43061 15427 43095
rect 15427 43061 15436 43095
rect 15384 43052 15436 43061
rect 15660 43095 15712 43104
rect 15660 43061 15669 43095
rect 15669 43061 15703 43095
rect 15703 43061 15712 43095
rect 15660 43052 15712 43061
rect 15936 43095 15988 43104
rect 15936 43061 15945 43095
rect 15945 43061 15979 43095
rect 15979 43061 15988 43095
rect 15936 43052 15988 43061
rect 19432 43120 19484 43172
rect 18788 43052 18840 43104
rect 3549 42950 3601 43002
rect 3613 42950 3665 43002
rect 3677 42950 3729 43002
rect 3741 42950 3793 43002
rect 3805 42950 3857 43002
rect 8747 42950 8799 43002
rect 8811 42950 8863 43002
rect 8875 42950 8927 43002
rect 8939 42950 8991 43002
rect 9003 42950 9055 43002
rect 13945 42950 13997 43002
rect 14009 42950 14061 43002
rect 14073 42950 14125 43002
rect 14137 42950 14189 43002
rect 14201 42950 14253 43002
rect 19143 42950 19195 43002
rect 19207 42950 19259 43002
rect 19271 42950 19323 43002
rect 19335 42950 19387 43002
rect 19399 42950 19451 43002
rect 6000 42848 6052 42900
rect 1952 42687 2004 42696
rect 1952 42653 1961 42687
rect 1961 42653 1995 42687
rect 1995 42653 2004 42687
rect 1952 42644 2004 42653
rect 2872 42712 2924 42764
rect 4436 42780 4488 42832
rect 7656 42848 7708 42900
rect 9680 42848 9732 42900
rect 8576 42780 8628 42832
rect 3148 42712 3200 42764
rect 3424 42712 3476 42764
rect 4620 42712 4672 42764
rect 4988 42712 5040 42764
rect 6828 42712 6880 42764
rect 7012 42755 7064 42764
rect 7012 42721 7021 42755
rect 7021 42721 7055 42755
rect 7055 42721 7064 42755
rect 7012 42712 7064 42721
rect 7564 42755 7616 42764
rect 7564 42721 7573 42755
rect 7573 42721 7607 42755
rect 7607 42721 7616 42755
rect 7564 42712 7616 42721
rect 8208 42712 8260 42764
rect 8668 42755 8720 42764
rect 8668 42721 8677 42755
rect 8677 42721 8711 42755
rect 8711 42721 8720 42755
rect 8668 42712 8720 42721
rect 8760 42712 8812 42764
rect 9220 42712 9272 42764
rect 12164 42848 12216 42900
rect 14648 42848 14700 42900
rect 15660 42848 15712 42900
rect 16028 42848 16080 42900
rect 16396 42848 16448 42900
rect 17224 42891 17276 42900
rect 17224 42857 17233 42891
rect 17233 42857 17267 42891
rect 17267 42857 17276 42891
rect 17224 42848 17276 42857
rect 17500 42848 17552 42900
rect 11336 42780 11388 42832
rect 388 42576 440 42628
rect 1400 42576 1452 42628
rect 2136 42619 2188 42628
rect 2136 42585 2145 42619
rect 2145 42585 2179 42619
rect 2179 42585 2188 42619
rect 2136 42576 2188 42585
rect 2964 42644 3016 42696
rect 6552 42644 6604 42696
rect 9128 42687 9180 42696
rect 9128 42653 9137 42687
rect 9137 42653 9171 42687
rect 9171 42653 9180 42687
rect 9128 42644 9180 42653
rect 9588 42644 9640 42696
rect 10416 42644 10468 42696
rect 10692 42644 10744 42696
rect 10968 42644 11020 42696
rect 11152 42644 11204 42696
rect 11428 42644 11480 42696
rect 11888 42687 11940 42696
rect 11888 42653 11897 42687
rect 11897 42653 11931 42687
rect 11931 42653 11940 42687
rect 11888 42644 11940 42653
rect 12256 42712 12308 42764
rect 15752 42780 15804 42832
rect 18788 42848 18840 42900
rect 19708 42848 19760 42900
rect 18236 42780 18288 42832
rect 12624 42687 12676 42696
rect 12624 42653 12633 42687
rect 12633 42653 12667 42687
rect 12667 42653 12676 42687
rect 12624 42644 12676 42653
rect 2688 42619 2740 42628
rect 2688 42585 2697 42619
rect 2697 42585 2731 42619
rect 2731 42585 2740 42619
rect 2688 42576 2740 42585
rect 2780 42576 2832 42628
rect 4896 42576 4948 42628
rect 5080 42619 5132 42628
rect 5080 42585 5089 42619
rect 5089 42585 5123 42619
rect 5123 42585 5132 42619
rect 5080 42576 5132 42585
rect 5816 42576 5868 42628
rect 5908 42576 5960 42628
rect 6736 42619 6788 42628
rect 6736 42585 6745 42619
rect 6745 42585 6779 42619
rect 6779 42585 6788 42619
rect 6736 42576 6788 42585
rect 3056 42508 3108 42560
rect 6000 42508 6052 42560
rect 7840 42619 7892 42628
rect 7840 42585 7849 42619
rect 7849 42585 7883 42619
rect 7883 42585 7892 42619
rect 7840 42576 7892 42585
rect 8392 42619 8444 42628
rect 8392 42585 8401 42619
rect 8401 42585 8435 42619
rect 8435 42585 8444 42619
rect 8392 42576 8444 42585
rect 8024 42508 8076 42560
rect 8760 42576 8812 42628
rect 9312 42576 9364 42628
rect 9496 42576 9548 42628
rect 13176 42687 13228 42696
rect 13176 42653 13185 42687
rect 13185 42653 13219 42687
rect 13219 42653 13228 42687
rect 13176 42644 13228 42653
rect 13544 42644 13596 42696
rect 13636 42687 13688 42696
rect 13636 42653 13645 42687
rect 13645 42653 13679 42687
rect 13679 42653 13688 42687
rect 13636 42644 13688 42653
rect 8668 42508 8720 42560
rect 9220 42508 9272 42560
rect 9864 42508 9916 42560
rect 10048 42551 10100 42560
rect 10048 42517 10057 42551
rect 10057 42517 10091 42551
rect 10091 42517 10100 42551
rect 10048 42508 10100 42517
rect 10508 42508 10560 42560
rect 10692 42508 10744 42560
rect 11152 42551 11204 42560
rect 11152 42517 11161 42551
rect 11161 42517 11195 42551
rect 11195 42517 11204 42551
rect 11152 42508 11204 42517
rect 11244 42508 11296 42560
rect 12072 42551 12124 42560
rect 12072 42517 12081 42551
rect 12081 42517 12115 42551
rect 12115 42517 12124 42551
rect 12072 42508 12124 42517
rect 12348 42551 12400 42560
rect 12348 42517 12357 42551
rect 12357 42517 12391 42551
rect 12391 42517 12400 42551
rect 12348 42508 12400 42517
rect 12900 42551 12952 42560
rect 12900 42517 12909 42551
rect 12909 42517 12943 42551
rect 12943 42517 12952 42551
rect 12900 42508 12952 42517
rect 12992 42508 13044 42560
rect 13820 42644 13872 42696
rect 15476 42712 15528 42764
rect 17132 42712 17184 42764
rect 18052 42712 18104 42764
rect 19984 42712 20036 42764
rect 14096 42576 14148 42628
rect 18328 42644 18380 42696
rect 19064 42644 19116 42696
rect 15108 42619 15160 42628
rect 15108 42585 15117 42619
rect 15117 42585 15151 42619
rect 15151 42585 15160 42619
rect 15108 42576 15160 42585
rect 15476 42576 15528 42628
rect 13820 42508 13872 42560
rect 14464 42551 14516 42560
rect 14464 42517 14473 42551
rect 14473 42517 14507 42551
rect 14507 42517 14516 42551
rect 14464 42508 14516 42517
rect 14740 42551 14792 42560
rect 14740 42517 14749 42551
rect 14749 42517 14783 42551
rect 14783 42517 14792 42551
rect 14740 42508 14792 42517
rect 17040 42576 17092 42628
rect 17500 42576 17552 42628
rect 17592 42576 17644 42628
rect 18052 42576 18104 42628
rect 19340 42619 19392 42628
rect 19340 42585 19349 42619
rect 19349 42585 19383 42619
rect 19383 42585 19392 42619
rect 19340 42576 19392 42585
rect 19616 42576 19668 42628
rect 20444 42619 20496 42628
rect 20444 42585 20453 42619
rect 20453 42585 20487 42619
rect 20487 42585 20496 42619
rect 20444 42576 20496 42585
rect 21364 42576 21416 42628
rect 6148 42406 6200 42458
rect 6212 42406 6264 42458
rect 6276 42406 6328 42458
rect 6340 42406 6392 42458
rect 6404 42406 6456 42458
rect 11346 42406 11398 42458
rect 11410 42406 11462 42458
rect 11474 42406 11526 42458
rect 11538 42406 11590 42458
rect 11602 42406 11654 42458
rect 16544 42406 16596 42458
rect 16608 42406 16660 42458
rect 16672 42406 16724 42458
rect 16736 42406 16788 42458
rect 16800 42406 16852 42458
rect 21742 42406 21794 42458
rect 21806 42406 21858 42458
rect 21870 42406 21922 42458
rect 21934 42406 21986 42458
rect 21998 42406 22050 42458
rect 2044 42304 2096 42356
rect 2780 42347 2832 42356
rect 2780 42313 2789 42347
rect 2789 42313 2823 42347
rect 2823 42313 2832 42347
rect 2780 42304 2832 42313
rect 4068 42304 4120 42356
rect 4252 42304 4304 42356
rect 4528 42347 4580 42356
rect 4528 42313 4537 42347
rect 4537 42313 4571 42347
rect 4571 42313 4580 42347
rect 4528 42304 4580 42313
rect 4804 42304 4856 42356
rect 5632 42347 5684 42356
rect 5632 42313 5641 42347
rect 5641 42313 5675 42347
rect 5675 42313 5684 42347
rect 5632 42304 5684 42313
rect 6000 42347 6052 42356
rect 6000 42313 6009 42347
rect 6009 42313 6043 42347
rect 6043 42313 6052 42347
rect 6000 42304 6052 42313
rect 6644 42304 6696 42356
rect 7196 42304 7248 42356
rect 10600 42347 10652 42356
rect 10600 42313 10609 42347
rect 10609 42313 10643 42347
rect 10643 42313 10652 42347
rect 10600 42304 10652 42313
rect 12900 42304 12952 42356
rect 1860 42168 1912 42220
rect 664 42100 716 42152
rect 3240 42211 3292 42220
rect 3240 42177 3249 42211
rect 3249 42177 3283 42211
rect 3283 42177 3292 42211
rect 3240 42168 3292 42177
rect 3332 42211 3384 42220
rect 3332 42177 3341 42211
rect 3341 42177 3375 42211
rect 3375 42177 3384 42211
rect 3332 42168 3384 42177
rect 3884 42211 3936 42220
rect 3884 42177 3893 42211
rect 3893 42177 3927 42211
rect 3927 42177 3936 42211
rect 3884 42168 3936 42177
rect 5264 42168 5316 42220
rect 9864 42236 9916 42288
rect 6184 42211 6236 42220
rect 6184 42177 6193 42211
rect 6193 42177 6227 42211
rect 6227 42177 6236 42211
rect 6184 42168 6236 42177
rect 5724 42100 5776 42152
rect 7288 42168 7340 42220
rect 9404 42211 9456 42220
rect 9404 42177 9413 42211
rect 9413 42177 9447 42211
rect 9447 42177 9456 42211
rect 9404 42168 9456 42177
rect 10692 42236 10744 42288
rect 11244 42236 11296 42288
rect 6000 42032 6052 42084
rect 7748 42100 7800 42152
rect 8944 42075 8996 42084
rect 8944 42041 8953 42075
rect 8953 42041 8987 42075
rect 8987 42041 8996 42075
rect 8944 42032 8996 42041
rect 9036 42032 9088 42084
rect 1032 41964 1084 42016
rect 7748 41964 7800 42016
rect 8576 42007 8628 42016
rect 8576 41973 8585 42007
rect 8585 41973 8619 42007
rect 8619 41973 8628 42007
rect 8576 41964 8628 41973
rect 10140 42100 10192 42152
rect 14464 42304 14516 42356
rect 14740 42304 14792 42356
rect 17316 42304 17368 42356
rect 17408 42304 17460 42356
rect 18144 42304 18196 42356
rect 14832 42236 14884 42288
rect 15200 42236 15252 42288
rect 19156 42304 19208 42356
rect 22192 42304 22244 42356
rect 22376 42304 22428 42356
rect 13728 42168 13780 42220
rect 14096 42168 14148 42220
rect 15292 42168 15344 42220
rect 15936 42168 15988 42220
rect 16028 42168 16080 42220
rect 16764 42211 16816 42220
rect 16764 42177 16773 42211
rect 16773 42177 16807 42211
rect 16807 42177 16816 42211
rect 16764 42168 16816 42177
rect 15660 42100 15712 42152
rect 16304 42100 16356 42152
rect 10692 42032 10744 42084
rect 11704 42032 11756 42084
rect 11980 42032 12032 42084
rect 13820 42032 13872 42084
rect 9588 41964 9640 42016
rect 9864 41964 9916 42016
rect 9956 42007 10008 42016
rect 9956 41973 9965 42007
rect 9965 41973 9999 42007
rect 9999 41973 10008 42007
rect 9956 41964 10008 41973
rect 13544 41964 13596 42016
rect 14004 41964 14056 42016
rect 14464 41964 14516 42016
rect 14924 41964 14976 42016
rect 15200 42007 15252 42016
rect 15200 41973 15209 42007
rect 15209 41973 15243 42007
rect 15243 41973 15252 42007
rect 15200 41964 15252 41973
rect 15752 41964 15804 42016
rect 15936 42007 15988 42016
rect 15936 41973 15945 42007
rect 15945 41973 15979 42007
rect 15979 41973 15988 42007
rect 15936 41964 15988 41973
rect 16856 42007 16908 42016
rect 16856 41973 16865 42007
rect 16865 41973 16899 42007
rect 16899 41973 16908 42007
rect 16856 41964 16908 41973
rect 16948 41964 17000 42016
rect 19064 42236 19116 42288
rect 17500 42211 17552 42220
rect 17500 42177 17509 42211
rect 17509 42177 17543 42211
rect 17543 42177 17552 42211
rect 17500 42168 17552 42177
rect 17776 42211 17828 42220
rect 17776 42177 17785 42211
rect 17785 42177 17819 42211
rect 17819 42177 17828 42211
rect 17776 42168 17828 42177
rect 18604 42168 18656 42220
rect 18880 42211 18932 42220
rect 18880 42177 18889 42211
rect 18889 42177 18923 42211
rect 18923 42177 18932 42211
rect 18880 42168 18932 42177
rect 18972 42168 19024 42220
rect 19524 42211 19576 42220
rect 19524 42177 19533 42211
rect 19533 42177 19567 42211
rect 19567 42177 19576 42211
rect 19524 42168 19576 42177
rect 17408 42100 17460 42152
rect 18328 42100 18380 42152
rect 19708 42236 19760 42288
rect 19984 42211 20036 42220
rect 19984 42177 19993 42211
rect 19993 42177 20027 42211
rect 20027 42177 20036 42211
rect 19984 42168 20036 42177
rect 20444 42211 20496 42220
rect 20444 42177 20453 42211
rect 20453 42177 20487 42211
rect 20487 42177 20496 42211
rect 20444 42168 20496 42177
rect 20904 42168 20956 42220
rect 21548 42100 21600 42152
rect 18880 42032 18932 42084
rect 20812 42032 20864 42084
rect 17776 41964 17828 42016
rect 19708 41964 19760 42016
rect 3549 41862 3601 41914
rect 3613 41862 3665 41914
rect 3677 41862 3729 41914
rect 3741 41862 3793 41914
rect 3805 41862 3857 41914
rect 8747 41862 8799 41914
rect 8811 41862 8863 41914
rect 8875 41862 8927 41914
rect 8939 41862 8991 41914
rect 9003 41862 9055 41914
rect 13945 41862 13997 41914
rect 14009 41862 14061 41914
rect 14073 41862 14125 41914
rect 14137 41862 14189 41914
rect 14201 41862 14253 41914
rect 19143 41862 19195 41914
rect 19207 41862 19259 41914
rect 19271 41862 19323 41914
rect 19335 41862 19387 41914
rect 19399 41862 19451 41914
rect 2688 41760 2740 41812
rect 3332 41760 3384 41812
rect 3884 41760 3936 41812
rect 3976 41760 4028 41812
rect 4712 41760 4764 41812
rect 5264 41760 5316 41812
rect 4068 41735 4120 41744
rect 4068 41701 4077 41735
rect 4077 41701 4111 41735
rect 4111 41701 4120 41735
rect 4068 41692 4120 41701
rect 5540 41692 5592 41744
rect 5724 41803 5776 41812
rect 5724 41769 5733 41803
rect 5733 41769 5767 41803
rect 5767 41769 5776 41803
rect 5724 41760 5776 41769
rect 5908 41760 5960 41812
rect 6184 41760 6236 41812
rect 6460 41803 6512 41812
rect 6460 41769 6469 41803
rect 6469 41769 6503 41803
rect 6503 41769 6512 41803
rect 6460 41760 6512 41769
rect 756 41556 808 41608
rect 2964 41556 3016 41608
rect 1492 41488 1544 41540
rect 2228 41531 2280 41540
rect 2228 41497 2237 41531
rect 2237 41497 2271 41531
rect 2271 41497 2280 41531
rect 2228 41488 2280 41497
rect 3608 41599 3660 41608
rect 3608 41565 3617 41599
rect 3617 41565 3651 41599
rect 3651 41565 3660 41599
rect 3608 41556 3660 41565
rect 3976 41599 4028 41608
rect 3976 41565 3985 41599
rect 3985 41565 4019 41599
rect 4019 41565 4028 41599
rect 3976 41556 4028 41565
rect 4252 41599 4304 41608
rect 4252 41565 4261 41599
rect 4261 41565 4295 41599
rect 4295 41565 4304 41599
rect 4252 41556 4304 41565
rect 4528 41599 4580 41608
rect 4528 41565 4537 41599
rect 4537 41565 4571 41599
rect 4571 41565 4580 41599
rect 4528 41556 4580 41565
rect 4804 41599 4856 41608
rect 4804 41565 4813 41599
rect 4813 41565 4847 41599
rect 4847 41565 4856 41599
rect 4804 41556 4856 41565
rect 5172 41556 5224 41608
rect 5356 41599 5408 41608
rect 5356 41565 5365 41599
rect 5365 41565 5399 41599
rect 5399 41565 5408 41599
rect 5356 41556 5408 41565
rect 5908 41599 5960 41608
rect 5908 41565 5917 41599
rect 5917 41565 5951 41599
rect 5951 41565 5960 41599
rect 5908 41556 5960 41565
rect 4160 41488 4212 41540
rect 5264 41488 5316 41540
rect 4988 41420 5040 41472
rect 7380 41760 7432 41812
rect 7840 41760 7892 41812
rect 12256 41760 12308 41812
rect 13728 41760 13780 41812
rect 7380 41599 7432 41608
rect 7380 41565 7389 41599
rect 7389 41565 7423 41599
rect 7423 41565 7432 41599
rect 7380 41556 7432 41565
rect 7748 41624 7800 41676
rect 9128 41692 9180 41744
rect 8484 41488 8536 41540
rect 8668 41556 8720 41608
rect 9312 41624 9364 41676
rect 9588 41624 9640 41676
rect 9404 41599 9456 41608
rect 9404 41565 9421 41599
rect 9421 41565 9455 41599
rect 9455 41565 9456 41599
rect 9404 41556 9456 41565
rect 9680 41599 9732 41608
rect 9680 41565 9689 41599
rect 9689 41565 9723 41599
rect 9723 41565 9732 41599
rect 9680 41556 9732 41565
rect 7932 41420 7984 41472
rect 13912 41624 13964 41676
rect 14372 41599 14424 41608
rect 14372 41565 14381 41599
rect 14381 41565 14415 41599
rect 14415 41565 14424 41599
rect 14372 41556 14424 41565
rect 15384 41760 15436 41812
rect 16028 41760 16080 41812
rect 16764 41760 16816 41812
rect 16948 41760 17000 41812
rect 17132 41692 17184 41744
rect 15384 41624 15436 41676
rect 15476 41624 15528 41676
rect 16304 41556 16356 41608
rect 17316 41624 17368 41676
rect 17408 41624 17460 41676
rect 17592 41735 17644 41744
rect 17592 41701 17601 41735
rect 17601 41701 17635 41735
rect 17635 41701 17644 41735
rect 17592 41692 17644 41701
rect 17868 41735 17920 41744
rect 17868 41701 17877 41735
rect 17877 41701 17911 41735
rect 17911 41701 17920 41735
rect 17868 41692 17920 41701
rect 18420 41760 18472 41812
rect 18880 41692 18932 41744
rect 16672 41599 16724 41608
rect 16672 41565 16681 41599
rect 16681 41565 16715 41599
rect 16715 41565 16724 41599
rect 16672 41556 16724 41565
rect 16948 41599 17000 41608
rect 16948 41565 16957 41599
rect 16957 41565 16991 41599
rect 16991 41565 17000 41599
rect 16948 41556 17000 41565
rect 17224 41599 17276 41608
rect 17224 41565 17233 41599
rect 17233 41565 17267 41599
rect 17267 41565 17276 41599
rect 17224 41556 17276 41565
rect 18420 41624 18472 41676
rect 19340 41692 19392 41744
rect 20536 41803 20588 41812
rect 20536 41769 20545 41803
rect 20545 41769 20579 41803
rect 20579 41769 20588 41803
rect 20536 41760 20588 41769
rect 21916 41760 21968 41812
rect 21456 41692 21508 41744
rect 9864 41420 9916 41472
rect 12532 41420 12584 41472
rect 14188 41420 14240 41472
rect 14832 41420 14884 41472
rect 15200 41420 15252 41472
rect 15384 41463 15436 41472
rect 15384 41429 15393 41463
rect 15393 41429 15427 41463
rect 15427 41429 15436 41463
rect 15384 41420 15436 41429
rect 15476 41420 15528 41472
rect 16856 41420 16908 41472
rect 17040 41420 17092 41472
rect 17408 41488 17460 41540
rect 17776 41599 17828 41608
rect 17776 41565 17785 41599
rect 17785 41565 17819 41599
rect 17819 41565 17828 41599
rect 17776 41556 17828 41565
rect 18328 41599 18380 41608
rect 18328 41565 18337 41599
rect 18337 41565 18371 41599
rect 18371 41565 18380 41599
rect 18328 41556 18380 41565
rect 22652 41624 22704 41676
rect 19800 41556 19852 41608
rect 18236 41420 18288 41472
rect 18420 41463 18472 41472
rect 18420 41429 18429 41463
rect 18429 41429 18463 41463
rect 18463 41429 18472 41463
rect 18420 41420 18472 41429
rect 20352 41599 20404 41608
rect 20352 41565 20361 41599
rect 20361 41565 20395 41599
rect 20395 41565 20404 41599
rect 20352 41556 20404 41565
rect 21088 41556 21140 41608
rect 21180 41531 21232 41540
rect 21180 41497 21189 41531
rect 21189 41497 21223 41531
rect 21223 41497 21232 41531
rect 21180 41488 21232 41497
rect 22284 41488 22336 41540
rect 22560 41420 22612 41472
rect 6148 41318 6200 41370
rect 6212 41318 6264 41370
rect 6276 41318 6328 41370
rect 6340 41318 6392 41370
rect 6404 41318 6456 41370
rect 11346 41318 11398 41370
rect 11410 41318 11462 41370
rect 11474 41318 11526 41370
rect 11538 41318 11590 41370
rect 11602 41318 11654 41370
rect 16544 41318 16596 41370
rect 16608 41318 16660 41370
rect 16672 41318 16724 41370
rect 16736 41318 16788 41370
rect 16800 41318 16852 41370
rect 21742 41318 21794 41370
rect 21806 41318 21858 41370
rect 21870 41318 21922 41370
rect 21934 41318 21986 41370
rect 21998 41318 22050 41370
rect 2504 41216 2556 41268
rect 4896 41216 4948 41268
rect 4712 41148 4764 41200
rect 5080 41148 5132 41200
rect 6000 41259 6052 41268
rect 6000 41225 6009 41259
rect 6009 41225 6043 41259
rect 6043 41225 6052 41259
rect 6000 41216 6052 41225
rect 6736 41216 6788 41268
rect 8392 41259 8444 41268
rect 8392 41225 8401 41259
rect 8401 41225 8435 41259
rect 8435 41225 8444 41259
rect 8392 41216 8444 41225
rect 14648 41259 14700 41268
rect 14648 41225 14657 41259
rect 14657 41225 14691 41259
rect 14691 41225 14700 41259
rect 14648 41216 14700 41225
rect 15016 41216 15068 41268
rect 15568 41216 15620 41268
rect 17316 41216 17368 41268
rect 1216 41080 1268 41132
rect 1584 41055 1636 41064
rect 1584 41021 1593 41055
rect 1593 41021 1627 41055
rect 1627 41021 1636 41055
rect 1584 41012 1636 41021
rect 2780 41080 2832 41132
rect 4160 41123 4212 41132
rect 4160 41089 4169 41123
rect 4169 41089 4203 41123
rect 4203 41089 4212 41123
rect 4160 41080 4212 41089
rect 5264 41080 5316 41132
rect 4068 41012 4120 41064
rect 5724 41080 5776 41132
rect 7656 41148 7708 41200
rect 14280 41148 14332 41200
rect 6552 41123 6604 41132
rect 6552 41089 6561 41123
rect 6561 41089 6595 41123
rect 6595 41089 6604 41123
rect 6552 41080 6604 41089
rect 7288 41080 7340 41132
rect 8576 41123 8628 41132
rect 8576 41089 8585 41123
rect 8585 41089 8619 41123
rect 8619 41089 8628 41123
rect 8576 41080 8628 41089
rect 11152 41080 11204 41132
rect 14556 41080 14608 41132
rect 15476 41148 15528 41200
rect 15200 41080 15252 41132
rect 2872 40944 2924 40996
rect 5908 40944 5960 40996
rect 7748 41012 7800 41064
rect 14740 41012 14792 41064
rect 15844 41080 15896 41132
rect 16396 41148 16448 41200
rect 16856 41123 16908 41132
rect 16856 41089 16865 41123
rect 16865 41089 16899 41123
rect 16899 41089 16908 41123
rect 16856 41080 16908 41089
rect 17316 41080 17368 41132
rect 16580 41012 16632 41064
rect 17592 41216 17644 41268
rect 17868 41216 17920 41268
rect 17960 41216 18012 41268
rect 18696 41216 18748 41268
rect 18788 41216 18840 41268
rect 19064 41216 19116 41268
rect 17592 41080 17644 41132
rect 18236 41080 18288 41132
rect 17500 41012 17552 41064
rect 17684 41012 17736 41064
rect 19708 41216 19760 41268
rect 21548 41216 21600 41268
rect 19064 41123 19116 41132
rect 19064 41089 19073 41123
rect 19073 41089 19107 41123
rect 19107 41089 19116 41123
rect 19064 41080 19116 41089
rect 19524 41080 19576 41132
rect 19892 41123 19944 41132
rect 19892 41089 19901 41123
rect 19901 41089 19935 41123
rect 19935 41089 19944 41123
rect 19892 41080 19944 41089
rect 20168 41123 20220 41132
rect 20168 41089 20177 41123
rect 20177 41089 20211 41123
rect 20211 41089 20220 41123
rect 20168 41080 20220 41089
rect 20444 41123 20496 41132
rect 20444 41089 20453 41123
rect 20453 41089 20487 41123
rect 20487 41089 20496 41123
rect 20444 41080 20496 41089
rect 7380 40944 7432 40996
rect 11060 40944 11112 40996
rect 16120 40944 16172 40996
rect 17224 40944 17276 40996
rect 7748 40919 7800 40928
rect 7748 40885 7757 40919
rect 7757 40885 7791 40919
rect 7791 40885 7800 40919
rect 7748 40876 7800 40885
rect 16764 40876 16816 40928
rect 17868 40944 17920 40996
rect 18696 40944 18748 40996
rect 18788 40876 18840 40928
rect 18880 40919 18932 40928
rect 18880 40885 18889 40919
rect 18889 40885 18923 40919
rect 18923 40885 18932 40919
rect 18880 40876 18932 40885
rect 19340 40944 19392 40996
rect 19984 41012 20036 41064
rect 20812 41080 20864 41132
rect 21272 41123 21324 41132
rect 21272 41089 21281 41123
rect 21281 41089 21315 41123
rect 21315 41089 21324 41123
rect 21272 41080 21324 41089
rect 21640 41012 21692 41064
rect 20904 40944 20956 40996
rect 20996 40944 21048 40996
rect 22192 40876 22244 40928
rect 3549 40774 3601 40826
rect 3613 40774 3665 40826
rect 3677 40774 3729 40826
rect 3741 40774 3793 40826
rect 3805 40774 3857 40826
rect 8747 40774 8799 40826
rect 8811 40774 8863 40826
rect 8875 40774 8927 40826
rect 8939 40774 8991 40826
rect 9003 40774 9055 40826
rect 13945 40774 13997 40826
rect 14009 40774 14061 40826
rect 14073 40774 14125 40826
rect 14137 40774 14189 40826
rect 14201 40774 14253 40826
rect 19143 40774 19195 40826
rect 19207 40774 19259 40826
rect 19271 40774 19323 40826
rect 19335 40774 19387 40826
rect 19399 40774 19451 40826
rect 5448 40715 5500 40724
rect 5448 40681 5457 40715
rect 5457 40681 5491 40715
rect 5491 40681 5500 40715
rect 5448 40672 5500 40681
rect 8576 40672 8628 40724
rect 16212 40672 16264 40724
rect 1952 40604 2004 40656
rect 4344 40604 4396 40656
rect 7472 40604 7524 40656
rect 7748 40604 7800 40656
rect 17132 40604 17184 40656
rect 17500 40647 17552 40656
rect 17500 40613 17509 40647
rect 17509 40613 17543 40647
rect 17543 40613 17552 40647
rect 17500 40604 17552 40613
rect 17868 40604 17920 40656
rect 19432 40604 19484 40656
rect 7380 40536 7432 40588
rect 8208 40536 8260 40588
rect 20444 40672 20496 40724
rect 20720 40672 20772 40724
rect 21272 40672 21324 40724
rect 19800 40604 19852 40656
rect 296 40468 348 40520
rect 1952 40511 2004 40520
rect 1952 40477 1961 40511
rect 1961 40477 1995 40511
rect 1995 40477 2004 40511
rect 1952 40468 2004 40477
rect 2044 40468 2096 40520
rect 5632 40511 5684 40520
rect 5632 40477 5641 40511
rect 5641 40477 5675 40511
rect 5675 40477 5684 40511
rect 5632 40468 5684 40477
rect 1676 40443 1728 40452
rect 1676 40409 1685 40443
rect 1685 40409 1719 40443
rect 1719 40409 1728 40443
rect 1676 40400 1728 40409
rect 2228 40443 2280 40452
rect 2228 40409 2237 40443
rect 2237 40409 2271 40443
rect 2271 40409 2280 40443
rect 2228 40400 2280 40409
rect 6552 40400 6604 40452
rect 17684 40511 17736 40520
rect 17684 40477 17693 40511
rect 17693 40477 17727 40511
rect 17727 40477 17736 40511
rect 17684 40468 17736 40477
rect 17960 40511 18012 40520
rect 17960 40477 17969 40511
rect 17969 40477 18003 40511
rect 18003 40477 18012 40511
rect 17960 40468 18012 40477
rect 18236 40511 18288 40520
rect 18236 40477 18245 40511
rect 18245 40477 18279 40511
rect 18279 40477 18288 40511
rect 18236 40468 18288 40477
rect 18328 40468 18380 40520
rect 18788 40511 18840 40520
rect 18788 40477 18797 40511
rect 18797 40477 18831 40511
rect 18831 40477 18840 40511
rect 18788 40468 18840 40477
rect 21180 40604 21232 40656
rect 19616 40511 19668 40520
rect 19616 40477 19625 40511
rect 19625 40477 19659 40511
rect 19659 40477 19668 40511
rect 19616 40468 19668 40477
rect 20076 40468 20128 40520
rect 19156 40400 19208 40452
rect 20720 40511 20772 40520
rect 20720 40477 20729 40511
rect 20729 40477 20763 40511
rect 20763 40477 20772 40511
rect 20720 40468 20772 40477
rect 20812 40468 20864 40520
rect 21272 40511 21324 40520
rect 21272 40477 21281 40511
rect 21281 40477 21315 40511
rect 21315 40477 21324 40511
rect 21272 40468 21324 40477
rect 8208 40332 8260 40384
rect 17224 40375 17276 40384
rect 17224 40341 17233 40375
rect 17233 40341 17267 40375
rect 17267 40341 17276 40375
rect 17224 40332 17276 40341
rect 18512 40332 18564 40384
rect 18604 40375 18656 40384
rect 18604 40341 18613 40375
rect 18613 40341 18647 40375
rect 18647 40341 18656 40375
rect 18604 40332 18656 40341
rect 19432 40375 19484 40384
rect 19432 40341 19441 40375
rect 19441 40341 19475 40375
rect 19475 40341 19484 40375
rect 19432 40332 19484 40341
rect 20260 40375 20312 40384
rect 20260 40341 20269 40375
rect 20269 40341 20303 40375
rect 20303 40341 20312 40375
rect 20260 40332 20312 40341
rect 20536 40375 20588 40384
rect 20536 40341 20545 40375
rect 20545 40341 20579 40375
rect 20579 40341 20588 40375
rect 20536 40332 20588 40341
rect 22192 40332 22244 40384
rect 6148 40230 6200 40282
rect 6212 40230 6264 40282
rect 6276 40230 6328 40282
rect 6340 40230 6392 40282
rect 6404 40230 6456 40282
rect 11346 40230 11398 40282
rect 11410 40230 11462 40282
rect 11474 40230 11526 40282
rect 11538 40230 11590 40282
rect 11602 40230 11654 40282
rect 16544 40230 16596 40282
rect 16608 40230 16660 40282
rect 16672 40230 16724 40282
rect 16736 40230 16788 40282
rect 16800 40230 16852 40282
rect 21742 40230 21794 40282
rect 21806 40230 21858 40282
rect 21870 40230 21922 40282
rect 21934 40230 21986 40282
rect 21998 40230 22050 40282
rect 2136 40128 2188 40180
rect 9220 40128 9272 40180
rect 15660 40128 15712 40180
rect 17592 40128 17644 40180
rect 17684 40128 17736 40180
rect 17776 40171 17828 40180
rect 17776 40137 17785 40171
rect 17785 40137 17819 40171
rect 17819 40137 17828 40171
rect 17776 40128 17828 40137
rect 18052 40171 18104 40180
rect 18052 40137 18061 40171
rect 18061 40137 18095 40171
rect 18095 40137 18104 40171
rect 18052 40128 18104 40137
rect 18420 40128 18472 40180
rect 18788 40128 18840 40180
rect 18880 40128 18932 40180
rect 18972 40128 19024 40180
rect 19156 40171 19208 40180
rect 19156 40137 19165 40171
rect 19165 40137 19199 40171
rect 19199 40137 19208 40171
rect 19156 40128 19208 40137
rect 3148 40060 3200 40112
rect 1768 40035 1820 40044
rect 1768 40001 1777 40035
rect 1777 40001 1811 40035
rect 1811 40001 1820 40035
rect 1768 39992 1820 40001
rect 2688 39992 2740 40044
rect 2596 39967 2648 39976
rect 2596 39933 2605 39967
rect 2605 39933 2639 39967
rect 2639 39933 2648 39967
rect 2596 39924 2648 39933
rect 1124 39856 1176 39908
rect 16304 40035 16356 40044
rect 16304 40001 16313 40035
rect 16313 40001 16347 40035
rect 16347 40001 16356 40035
rect 16304 39992 16356 40001
rect 17684 40035 17736 40044
rect 17684 40001 17693 40035
rect 17693 40001 17727 40035
rect 17727 40001 17736 40035
rect 17684 39992 17736 40001
rect 3424 39924 3476 39976
rect 4712 39856 4764 39908
rect 5540 39856 5592 39908
rect 4068 39788 4120 39840
rect 6828 39788 6880 39840
rect 13544 39856 13596 39908
rect 15936 39856 15988 39908
rect 18144 40060 18196 40112
rect 20260 40128 20312 40180
rect 20352 40128 20404 40180
rect 18696 39992 18748 40044
rect 18788 40035 18840 40044
rect 18788 40001 18797 40035
rect 18797 40001 18831 40035
rect 18831 40001 18840 40035
rect 18788 39992 18840 40001
rect 18972 39992 19024 40044
rect 18052 39924 18104 39976
rect 19708 39992 19760 40044
rect 19432 39924 19484 39976
rect 16212 39788 16264 39840
rect 19892 39856 19944 39908
rect 20904 40060 20956 40112
rect 21088 39992 21140 40044
rect 21364 39924 21416 39976
rect 20996 39856 21048 39908
rect 22468 39856 22520 39908
rect 21456 39831 21508 39840
rect 21456 39797 21465 39831
rect 21465 39797 21499 39831
rect 21499 39797 21508 39831
rect 21456 39788 21508 39797
rect 3549 39686 3601 39738
rect 3613 39686 3665 39738
rect 3677 39686 3729 39738
rect 3741 39686 3793 39738
rect 3805 39686 3857 39738
rect 8747 39686 8799 39738
rect 8811 39686 8863 39738
rect 8875 39686 8927 39738
rect 8939 39686 8991 39738
rect 9003 39686 9055 39738
rect 13945 39686 13997 39738
rect 14009 39686 14061 39738
rect 14073 39686 14125 39738
rect 14137 39686 14189 39738
rect 14201 39686 14253 39738
rect 19143 39686 19195 39738
rect 19207 39686 19259 39738
rect 19271 39686 19323 39738
rect 19335 39686 19387 39738
rect 19399 39686 19451 39738
rect 5816 39584 5868 39636
rect 10140 39584 10192 39636
rect 16304 39584 16356 39636
rect 17684 39584 17736 39636
rect 18052 39627 18104 39636
rect 18052 39593 18061 39627
rect 18061 39593 18095 39627
rect 18095 39593 18104 39627
rect 18052 39584 18104 39593
rect 19616 39584 19668 39636
rect 20720 39584 20772 39636
rect 21272 39584 21324 39636
rect 8116 39516 8168 39568
rect 1676 39380 1728 39432
rect 1860 39380 1912 39432
rect 3056 39448 3108 39500
rect 3700 39448 3752 39500
rect 18972 39516 19024 39568
rect 19340 39516 19392 39568
rect 1308 39312 1360 39364
rect 5724 39380 5776 39432
rect 16120 39423 16172 39432
rect 16120 39389 16129 39423
rect 16129 39389 16163 39423
rect 16163 39389 16172 39423
rect 16120 39380 16172 39389
rect 17500 39380 17552 39432
rect 17684 39380 17736 39432
rect 3976 39312 4028 39364
rect 2504 39287 2556 39296
rect 2504 39253 2513 39287
rect 2513 39253 2547 39287
rect 2547 39253 2556 39287
rect 2504 39244 2556 39253
rect 4160 39244 4212 39296
rect 8392 39244 8444 39296
rect 17040 39244 17092 39296
rect 19616 39448 19668 39500
rect 18880 39380 18932 39432
rect 19524 39380 19576 39432
rect 19708 39423 19760 39432
rect 19708 39389 19717 39423
rect 19717 39389 19751 39423
rect 19751 39389 19760 39423
rect 19708 39380 19760 39389
rect 19800 39380 19852 39432
rect 18788 39312 18840 39364
rect 20352 39380 20404 39432
rect 20444 39312 20496 39364
rect 20812 39380 20864 39432
rect 20996 39423 21048 39432
rect 20996 39389 21005 39423
rect 21005 39389 21039 39423
rect 21039 39389 21048 39423
rect 20996 39380 21048 39389
rect 20720 39312 20772 39364
rect 20812 39287 20864 39296
rect 20812 39253 20821 39287
rect 20821 39253 20855 39287
rect 20855 39253 20864 39287
rect 20812 39244 20864 39253
rect 22192 39244 22244 39296
rect 6148 39142 6200 39194
rect 6212 39142 6264 39194
rect 6276 39142 6328 39194
rect 6340 39142 6392 39194
rect 6404 39142 6456 39194
rect 11346 39142 11398 39194
rect 11410 39142 11462 39194
rect 11474 39142 11526 39194
rect 11538 39142 11590 39194
rect 11602 39142 11654 39194
rect 16544 39142 16596 39194
rect 16608 39142 16660 39194
rect 16672 39142 16724 39194
rect 16736 39142 16788 39194
rect 16800 39142 16852 39194
rect 21742 39142 21794 39194
rect 21806 39142 21858 39194
rect 21870 39142 21922 39194
rect 21934 39142 21986 39194
rect 21998 39142 22050 39194
rect 1584 39040 1636 39092
rect 5080 39040 5132 39092
rect 6000 39083 6052 39092
rect 6000 39049 6009 39083
rect 6009 39049 6043 39083
rect 6043 39049 6052 39083
rect 6000 39040 6052 39049
rect 16120 39040 16172 39092
rect 18788 39083 18840 39092
rect 18788 39049 18797 39083
rect 18797 39049 18831 39083
rect 18831 39049 18840 39083
rect 18788 39040 18840 39049
rect 1860 38972 1912 39024
rect 2964 38972 3016 39024
rect 3148 38972 3200 39024
rect 3332 38972 3384 39024
rect 2596 38904 2648 38956
rect 3700 38904 3752 38956
rect 8300 38972 8352 39024
rect 20168 39040 20220 39092
rect 20352 39040 20404 39092
rect 20720 39040 20772 39092
rect 20812 39040 20864 39092
rect 6000 38904 6052 38956
rect 1676 38836 1728 38888
rect 1492 38700 1544 38752
rect 1676 38700 1728 38752
rect 2964 38836 3016 38888
rect 3424 38836 3476 38888
rect 5264 38768 5316 38820
rect 6552 38904 6604 38956
rect 6736 38904 6788 38956
rect 15844 38947 15896 38956
rect 15844 38913 15853 38947
rect 15853 38913 15887 38947
rect 15887 38913 15896 38947
rect 15844 38904 15896 38913
rect 17040 38904 17092 38956
rect 18972 38947 19024 38956
rect 18972 38913 18981 38947
rect 18981 38913 19015 38947
rect 19015 38913 19024 38947
rect 18972 38904 19024 38913
rect 19800 38904 19852 38956
rect 16212 38836 16264 38888
rect 20260 38947 20312 38956
rect 20260 38913 20269 38947
rect 20269 38913 20303 38947
rect 20303 38913 20312 38947
rect 20260 38904 20312 38913
rect 20720 38947 20772 38956
rect 20720 38913 20729 38947
rect 20729 38913 20763 38947
rect 20763 38913 20772 38947
rect 20720 38904 20772 38913
rect 20904 38904 20956 38956
rect 2320 38700 2372 38752
rect 3148 38700 3200 38752
rect 3884 38700 3936 38752
rect 4528 38700 4580 38752
rect 5172 38700 5224 38752
rect 5908 38700 5960 38752
rect 11888 38768 11940 38820
rect 12256 38768 12308 38820
rect 6644 38700 6696 38752
rect 7380 38743 7432 38752
rect 7380 38709 7389 38743
rect 7389 38709 7423 38743
rect 7423 38709 7432 38743
rect 7380 38700 7432 38709
rect 7564 38700 7616 38752
rect 12624 38700 12676 38752
rect 15752 38700 15804 38752
rect 16212 38700 16264 38752
rect 21180 38700 21232 38752
rect 21456 38743 21508 38752
rect 21456 38709 21465 38743
rect 21465 38709 21499 38743
rect 21499 38709 21508 38743
rect 21456 38700 21508 38709
rect 3549 38598 3601 38650
rect 3613 38598 3665 38650
rect 3677 38598 3729 38650
rect 3741 38598 3793 38650
rect 3805 38598 3857 38650
rect 8747 38598 8799 38650
rect 8811 38598 8863 38650
rect 8875 38598 8927 38650
rect 8939 38598 8991 38650
rect 9003 38598 9055 38650
rect 13945 38598 13997 38650
rect 14009 38598 14061 38650
rect 14073 38598 14125 38650
rect 14137 38598 14189 38650
rect 14201 38598 14253 38650
rect 19143 38598 19195 38650
rect 19207 38598 19259 38650
rect 19271 38598 19323 38650
rect 19335 38598 19387 38650
rect 19399 38598 19451 38650
rect 1124 38360 1176 38412
rect 6828 38496 6880 38548
rect 9680 38496 9732 38548
rect 13176 38496 13228 38548
rect 16028 38496 16080 38548
rect 17684 38496 17736 38548
rect 18972 38496 19024 38548
rect 20720 38496 20772 38548
rect 20996 38496 21048 38548
rect 19984 38471 20036 38480
rect 19984 38437 19993 38471
rect 19993 38437 20027 38471
rect 20027 38437 20036 38471
rect 19984 38428 20036 38437
rect 3884 38403 3936 38412
rect 3884 38369 3893 38403
rect 3893 38369 3927 38403
rect 3927 38369 3936 38403
rect 3884 38360 3936 38369
rect 5264 38360 5316 38412
rect 7564 38360 7616 38412
rect 12716 38360 12768 38412
rect 14556 38360 14608 38412
rect 16028 38360 16080 38412
rect 1860 38292 1912 38344
rect 1308 38224 1360 38276
rect 4068 38292 4120 38344
rect 4896 38292 4948 38344
rect 3424 38267 3476 38276
rect 3424 38233 3433 38267
rect 3433 38233 3467 38267
rect 3467 38233 3476 38267
rect 3424 38224 3476 38233
rect 5540 38292 5592 38344
rect 6644 38292 6696 38344
rect 6920 38292 6972 38344
rect 9128 38292 9180 38344
rect 13544 38292 13596 38344
rect 7840 38224 7892 38276
rect 11704 38224 11756 38276
rect 18604 38292 18656 38344
rect 20168 38335 20220 38344
rect 20168 38301 20177 38335
rect 20177 38301 20211 38335
rect 20211 38301 20220 38335
rect 20168 38292 20220 38301
rect 20444 38335 20496 38344
rect 20444 38301 20453 38335
rect 20453 38301 20487 38335
rect 20487 38301 20496 38335
rect 20444 38292 20496 38301
rect 20720 38335 20772 38344
rect 20720 38301 20729 38335
rect 20729 38301 20763 38335
rect 20763 38301 20772 38335
rect 20720 38292 20772 38301
rect 20812 38292 20864 38344
rect 2688 38199 2740 38208
rect 2688 38165 2697 38199
rect 2697 38165 2731 38199
rect 2731 38165 2740 38199
rect 2688 38156 2740 38165
rect 4988 38156 5040 38208
rect 5264 38156 5316 38208
rect 6552 38156 6604 38208
rect 7196 38156 7248 38208
rect 7748 38199 7800 38208
rect 7748 38165 7757 38199
rect 7757 38165 7791 38199
rect 7791 38165 7800 38199
rect 7748 38156 7800 38165
rect 8208 38156 8260 38208
rect 14832 38156 14884 38208
rect 15200 38156 15252 38208
rect 21088 38156 21140 38208
rect 22192 38156 22244 38208
rect 6148 38054 6200 38106
rect 6212 38054 6264 38106
rect 6276 38054 6328 38106
rect 6340 38054 6392 38106
rect 6404 38054 6456 38106
rect 11346 38054 11398 38106
rect 11410 38054 11462 38106
rect 11474 38054 11526 38106
rect 11538 38054 11590 38106
rect 11602 38054 11654 38106
rect 16544 38054 16596 38106
rect 16608 38054 16660 38106
rect 16672 38054 16724 38106
rect 16736 38054 16788 38106
rect 16800 38054 16852 38106
rect 21742 38054 21794 38106
rect 21806 38054 21858 38106
rect 21870 38054 21922 38106
rect 21934 38054 21986 38106
rect 21998 38054 22050 38106
rect 3240 37952 3292 38004
rect 6000 37995 6052 38004
rect 6000 37961 6009 37995
rect 6009 37961 6043 37995
rect 6043 37961 6052 37995
rect 6000 37952 6052 37961
rect 1492 37816 1544 37868
rect 3148 37859 3200 37868
rect 3148 37825 3157 37859
rect 3157 37825 3191 37859
rect 3191 37825 3200 37859
rect 3148 37816 3200 37825
rect 3884 37816 3936 37868
rect 4896 37859 4948 37868
rect 4896 37825 4903 37859
rect 4903 37825 4937 37859
rect 4937 37825 4948 37859
rect 4896 37816 4948 37825
rect 7104 37927 7156 37936
rect 7104 37893 7113 37927
rect 7113 37893 7147 37927
rect 7147 37893 7156 37927
rect 7104 37884 7156 37893
rect 6276 37816 6328 37868
rect 7288 37816 7340 37868
rect 7656 37816 7708 37868
rect 7840 37859 7892 37868
rect 7840 37825 7849 37859
rect 7849 37825 7883 37859
rect 7883 37825 7892 37859
rect 7840 37816 7892 37825
rect 8300 37816 8352 37868
rect 10048 37952 10100 38004
rect 15844 37952 15896 38004
rect 18604 37995 18656 38004
rect 18604 37961 18613 37995
rect 18613 37961 18647 37995
rect 18647 37961 18656 37995
rect 18604 37952 18656 37961
rect 20168 37952 20220 38004
rect 20720 37952 20772 38004
rect 11244 37816 11296 37868
rect 12256 37816 12308 37868
rect 13544 37884 13596 37936
rect 14188 37884 14240 37936
rect 13176 37816 13228 37868
rect 1860 37748 1912 37800
rect 2504 37748 2556 37800
rect 2872 37791 2924 37800
rect 2872 37757 2881 37791
rect 2881 37757 2915 37791
rect 2915 37757 2924 37791
rect 2872 37748 2924 37757
rect 2412 37680 2464 37732
rect 4160 37748 4212 37800
rect 7748 37748 7800 37800
rect 3148 37612 3200 37664
rect 4528 37655 4580 37664
rect 4528 37621 4537 37655
rect 4537 37621 4571 37655
rect 4571 37621 4580 37655
rect 4528 37612 4580 37621
rect 5540 37612 5592 37664
rect 6644 37655 6696 37664
rect 6644 37621 6653 37655
rect 6653 37621 6687 37655
rect 6687 37621 6696 37655
rect 6644 37612 6696 37621
rect 6920 37612 6972 37664
rect 8484 37612 8536 37664
rect 9220 37612 9272 37664
rect 10692 37655 10744 37664
rect 10692 37621 10701 37655
rect 10701 37621 10735 37655
rect 10735 37621 10744 37655
rect 10692 37612 10744 37621
rect 11152 37612 11204 37664
rect 12072 37612 12124 37664
rect 14280 37612 14332 37664
rect 15200 37816 15252 37868
rect 18788 37859 18840 37868
rect 18788 37825 18797 37859
rect 18797 37825 18831 37859
rect 18831 37825 18840 37859
rect 18788 37816 18840 37825
rect 20076 37859 20128 37868
rect 20076 37825 20085 37859
rect 20085 37825 20119 37859
rect 20119 37825 20128 37859
rect 20076 37816 20128 37825
rect 20168 37816 20220 37868
rect 20720 37859 20772 37868
rect 20720 37825 20729 37859
rect 20729 37825 20763 37859
rect 20763 37825 20772 37859
rect 20720 37816 20772 37825
rect 20996 37859 21048 37868
rect 20996 37825 21005 37859
rect 21005 37825 21039 37859
rect 21039 37825 21048 37859
rect 20996 37816 21048 37825
rect 21180 37816 21232 37868
rect 14556 37791 14608 37800
rect 14556 37757 14565 37791
rect 14565 37757 14599 37791
rect 14599 37757 14608 37791
rect 14556 37748 14608 37757
rect 19708 37748 19760 37800
rect 20812 37748 20864 37800
rect 18328 37680 18380 37732
rect 20904 37680 20956 37732
rect 15568 37655 15620 37664
rect 15568 37621 15577 37655
rect 15577 37621 15611 37655
rect 15611 37621 15620 37655
rect 15568 37612 15620 37621
rect 20812 37655 20864 37664
rect 20812 37621 20821 37655
rect 20821 37621 20855 37655
rect 20855 37621 20864 37655
rect 20812 37612 20864 37621
rect 21456 37655 21508 37664
rect 21456 37621 21465 37655
rect 21465 37621 21499 37655
rect 21499 37621 21508 37655
rect 21456 37612 21508 37621
rect 3549 37510 3601 37562
rect 3613 37510 3665 37562
rect 3677 37510 3729 37562
rect 3741 37510 3793 37562
rect 3805 37510 3857 37562
rect 8747 37510 8799 37562
rect 8811 37510 8863 37562
rect 8875 37510 8927 37562
rect 8939 37510 8991 37562
rect 9003 37510 9055 37562
rect 13945 37510 13997 37562
rect 14009 37510 14061 37562
rect 14073 37510 14125 37562
rect 14137 37510 14189 37562
rect 14201 37510 14253 37562
rect 19143 37510 19195 37562
rect 19207 37510 19259 37562
rect 19271 37510 19323 37562
rect 19335 37510 19387 37562
rect 19399 37510 19451 37562
rect 1860 37408 1912 37460
rect 4252 37408 4304 37460
rect 2320 37340 2372 37392
rect 2872 37340 2924 37392
rect 5448 37408 5500 37460
rect 5724 37451 5776 37460
rect 5724 37417 5733 37451
rect 5733 37417 5767 37451
rect 5767 37417 5776 37451
rect 5724 37408 5776 37417
rect 14004 37408 14056 37460
rect 19708 37451 19760 37460
rect 19708 37417 19717 37451
rect 19717 37417 19751 37451
rect 19751 37417 19760 37451
rect 19708 37408 19760 37417
rect 20168 37408 20220 37460
rect 20444 37408 20496 37460
rect 20720 37408 20772 37460
rect 4436 37383 4488 37392
rect 4436 37349 4445 37383
rect 4445 37349 4479 37383
rect 4479 37349 4488 37383
rect 4436 37340 4488 37349
rect 4528 37340 4580 37392
rect 15660 37340 15712 37392
rect 16948 37340 17000 37392
rect 4068 37272 4120 37324
rect 4988 37315 5040 37324
rect 4988 37281 4997 37315
rect 4997 37281 5031 37315
rect 5031 37281 5040 37315
rect 4988 37272 5040 37281
rect 3056 37247 3108 37256
rect 3056 37213 3065 37247
rect 3065 37213 3099 37247
rect 3099 37213 3108 37247
rect 3056 37204 3108 37213
rect 3148 37204 3200 37256
rect 3240 37136 3292 37188
rect 3976 37247 4028 37256
rect 3976 37213 3985 37247
rect 3985 37213 4019 37247
rect 4019 37213 4028 37247
rect 3976 37204 4028 37213
rect 4896 37204 4948 37256
rect 1860 37068 1912 37120
rect 2964 37068 3016 37120
rect 3884 37068 3936 37120
rect 6552 37272 6604 37324
rect 7380 37272 7432 37324
rect 6368 37204 6420 37256
rect 6644 37204 6696 37256
rect 4712 37068 4764 37120
rect 5448 37068 5500 37120
rect 6276 37068 6328 37120
rect 6920 37179 6972 37188
rect 6920 37145 6929 37179
rect 6929 37145 6963 37179
rect 6963 37145 6972 37179
rect 6920 37136 6972 37145
rect 9956 37272 10008 37324
rect 10692 37272 10744 37324
rect 12256 37272 12308 37324
rect 13084 37272 13136 37324
rect 10876 37204 10928 37256
rect 11704 37247 11756 37256
rect 11704 37213 11713 37247
rect 11713 37213 11747 37247
rect 11747 37213 11756 37247
rect 11704 37204 11756 37213
rect 10416 37136 10468 37188
rect 10968 37179 11020 37188
rect 10968 37145 10977 37179
rect 10977 37145 11011 37179
rect 11011 37145 11020 37179
rect 10968 37136 11020 37145
rect 12624 37183 12649 37188
rect 12649 37183 12676 37188
rect 12624 37136 12676 37183
rect 15568 37272 15620 37324
rect 15108 37204 15160 37256
rect 15752 37247 15804 37256
rect 15752 37213 15761 37247
rect 15761 37213 15795 37247
rect 15795 37213 15804 37247
rect 15752 37204 15804 37213
rect 14556 37179 14608 37188
rect 7104 37068 7156 37120
rect 7748 37068 7800 37120
rect 8576 37068 8628 37120
rect 8852 37068 8904 37120
rect 9772 37111 9824 37120
rect 9772 37077 9781 37111
rect 9781 37077 9815 37111
rect 9815 37077 9824 37111
rect 9772 37068 9824 37077
rect 10232 37111 10284 37120
rect 10232 37077 10241 37111
rect 10241 37077 10275 37111
rect 10275 37077 10284 37111
rect 10232 37068 10284 37077
rect 11336 37111 11388 37120
rect 11336 37077 11345 37111
rect 11345 37077 11379 37111
rect 11379 37077 11388 37111
rect 11336 37068 11388 37077
rect 12072 37068 12124 37120
rect 13452 37068 13504 37120
rect 14556 37145 14568 37179
rect 14568 37145 14608 37179
rect 14556 37136 14608 37145
rect 13912 37068 13964 37120
rect 14004 37068 14056 37120
rect 14372 37068 14424 37120
rect 15844 37111 15896 37120
rect 15844 37077 15853 37111
rect 15853 37077 15887 37111
rect 15887 37077 15896 37111
rect 15844 37068 15896 37077
rect 16120 37111 16172 37120
rect 16120 37077 16129 37111
rect 16129 37077 16163 37111
rect 16163 37077 16172 37111
rect 16120 37068 16172 37077
rect 17224 37247 17276 37256
rect 17224 37213 17233 37247
rect 17233 37213 17267 37247
rect 17267 37213 17276 37247
rect 17224 37204 17276 37213
rect 17868 37247 17920 37256
rect 17868 37213 17877 37247
rect 17877 37213 17911 37247
rect 17911 37213 17920 37247
rect 17868 37204 17920 37213
rect 18052 37204 18104 37256
rect 18236 37204 18288 37256
rect 19708 37204 19760 37256
rect 20444 37247 20496 37256
rect 20444 37213 20453 37247
rect 20453 37213 20487 37247
rect 20487 37213 20496 37247
rect 20444 37204 20496 37213
rect 20536 37204 20588 37256
rect 20904 37204 20956 37256
rect 21088 37204 21140 37256
rect 17316 37111 17368 37120
rect 17316 37077 17325 37111
rect 17325 37077 17359 37111
rect 17359 37077 17368 37111
rect 17316 37068 17368 37077
rect 18144 37111 18196 37120
rect 18144 37077 18153 37111
rect 18153 37077 18187 37111
rect 18187 37077 18196 37111
rect 18144 37068 18196 37077
rect 22284 37136 22336 37188
rect 21088 37068 21140 37120
rect 6148 36966 6200 37018
rect 6212 36966 6264 37018
rect 6276 36966 6328 37018
rect 6340 36966 6392 37018
rect 6404 36966 6456 37018
rect 11346 36966 11398 37018
rect 11410 36966 11462 37018
rect 11474 36966 11526 37018
rect 11538 36966 11590 37018
rect 11602 36966 11654 37018
rect 16544 36966 16596 37018
rect 16608 36966 16660 37018
rect 16672 36966 16724 37018
rect 16736 36966 16788 37018
rect 16800 36966 16852 37018
rect 21742 36966 21794 37018
rect 21806 36966 21858 37018
rect 21870 36966 21922 37018
rect 21934 36966 21986 37018
rect 21998 36966 22050 37018
rect 3792 36864 3844 36916
rect 5632 36864 5684 36916
rect 8300 36907 8352 36916
rect 8300 36873 8309 36907
rect 8309 36873 8343 36907
rect 8343 36873 8352 36907
rect 8300 36864 8352 36873
rect 572 36728 624 36780
rect 1676 36728 1728 36780
rect 2504 36728 2556 36780
rect 3332 36728 3384 36780
rect 4344 36771 4396 36780
rect 4344 36737 4351 36771
rect 4351 36737 4385 36771
rect 4385 36737 4396 36771
rect 4344 36728 4396 36737
rect 4896 36728 4948 36780
rect 5448 36728 5500 36780
rect 6000 36728 6052 36780
rect 6368 36771 6420 36780
rect 6368 36737 6377 36771
rect 6377 36737 6411 36771
rect 6411 36737 6420 36771
rect 6368 36728 6420 36737
rect 7564 36771 7616 36780
rect 7564 36737 7573 36771
rect 7573 36737 7616 36771
rect 7564 36728 7616 36737
rect 7656 36728 7708 36780
rect 9956 36864 10008 36916
rect 10232 36864 10284 36916
rect 9128 36796 9180 36848
rect 10416 36864 10468 36916
rect 14556 36864 14608 36916
rect 15752 36864 15804 36916
rect 15844 36864 15896 36916
rect 16120 36864 16172 36916
rect 16396 36864 16448 36916
rect 16580 36864 16632 36916
rect 17224 36864 17276 36916
rect 17316 36864 17368 36916
rect 17868 36864 17920 36916
rect 18144 36864 18196 36916
rect 8852 36728 8904 36780
rect 9404 36728 9456 36780
rect 1860 36660 1912 36712
rect 2412 36660 2464 36712
rect 3424 36660 3476 36712
rect 4068 36703 4120 36712
rect 4068 36669 4077 36703
rect 4077 36669 4111 36703
rect 4111 36669 4120 36703
rect 4068 36660 4120 36669
rect 2412 36524 2464 36576
rect 6828 36660 6880 36712
rect 7196 36660 7248 36712
rect 5448 36592 5500 36644
rect 6920 36592 6972 36644
rect 4988 36524 5040 36576
rect 5724 36524 5776 36576
rect 9588 36524 9640 36576
rect 9864 36524 9916 36576
rect 12992 36796 13044 36848
rect 10048 36771 10100 36780
rect 10048 36737 10057 36771
rect 10057 36737 10091 36771
rect 10091 36737 10100 36771
rect 10048 36728 10100 36737
rect 10232 36728 10284 36780
rect 11704 36728 11756 36780
rect 14004 36728 14056 36780
rect 15108 36728 15160 36780
rect 11796 36635 11848 36644
rect 11796 36601 11805 36635
rect 11805 36601 11839 36635
rect 11839 36601 11848 36635
rect 11796 36592 11848 36601
rect 13176 36660 13228 36712
rect 13452 36660 13504 36712
rect 13636 36660 13688 36712
rect 13820 36703 13872 36712
rect 13820 36669 13829 36703
rect 13829 36669 13863 36703
rect 13863 36669 13872 36703
rect 13820 36660 13872 36669
rect 14280 36660 14332 36712
rect 16304 36728 16356 36780
rect 16396 36771 16448 36780
rect 16396 36737 16405 36771
rect 16405 36737 16439 36771
rect 16439 36737 16448 36771
rect 16396 36728 16448 36737
rect 16488 36728 16540 36780
rect 20812 36864 20864 36916
rect 20996 36864 21048 36916
rect 19616 36771 19668 36780
rect 19616 36737 19625 36771
rect 19625 36737 19659 36771
rect 19659 36737 19668 36771
rect 19616 36728 19668 36737
rect 20352 36771 20404 36780
rect 20352 36737 20361 36771
rect 20361 36737 20395 36771
rect 20395 36737 20404 36771
rect 20352 36728 20404 36737
rect 15568 36592 15620 36644
rect 14556 36524 14608 36576
rect 16488 36524 16540 36576
rect 18512 36660 18564 36712
rect 20444 36660 20496 36712
rect 19800 36592 19852 36644
rect 20812 36771 20864 36780
rect 20812 36737 20821 36771
rect 20821 36737 20855 36771
rect 20855 36737 20864 36771
rect 20812 36728 20864 36737
rect 17960 36524 18012 36576
rect 18144 36524 18196 36576
rect 19708 36524 19760 36576
rect 19984 36524 20036 36576
rect 20904 36524 20956 36576
rect 21456 36567 21508 36576
rect 21456 36533 21465 36567
rect 21465 36533 21499 36567
rect 21499 36533 21508 36567
rect 21456 36524 21508 36533
rect 3549 36422 3601 36474
rect 3613 36422 3665 36474
rect 3677 36422 3729 36474
rect 3741 36422 3793 36474
rect 3805 36422 3857 36474
rect 8747 36422 8799 36474
rect 8811 36422 8863 36474
rect 8875 36422 8927 36474
rect 8939 36422 8991 36474
rect 9003 36422 9055 36474
rect 13945 36422 13997 36474
rect 14009 36422 14061 36474
rect 14073 36422 14125 36474
rect 14137 36422 14189 36474
rect 14201 36422 14253 36474
rect 19143 36422 19195 36474
rect 19207 36422 19259 36474
rect 19271 36422 19323 36474
rect 19335 36422 19387 36474
rect 19399 36422 19451 36474
rect 1216 36320 1268 36372
rect 1584 36320 1636 36372
rect 4804 36320 4856 36372
rect 5632 36320 5684 36372
rect 5816 36320 5868 36372
rect 1124 36116 1176 36168
rect 1400 36159 1452 36168
rect 1400 36125 1409 36159
rect 1409 36125 1443 36159
rect 1443 36125 1452 36159
rect 1400 36116 1452 36125
rect 2596 36116 2648 36168
rect 5448 36184 5500 36236
rect 6920 36184 6972 36236
rect 7196 36184 7248 36236
rect 9772 36320 9824 36372
rect 10968 36320 11020 36372
rect 13820 36320 13872 36372
rect 14740 36320 14792 36372
rect 15016 36320 15068 36372
rect 16396 36320 16448 36372
rect 16580 36363 16632 36372
rect 16580 36329 16589 36363
rect 16589 36329 16623 36363
rect 16623 36329 16632 36363
rect 16580 36320 16632 36329
rect 10048 36252 10100 36304
rect 12256 36295 12308 36304
rect 12256 36261 12265 36295
rect 12265 36261 12299 36295
rect 12299 36261 12308 36295
rect 12256 36252 12308 36261
rect 14556 36252 14608 36304
rect 18144 36320 18196 36372
rect 21180 36320 21232 36372
rect 19708 36252 19760 36304
rect 4068 36048 4120 36100
rect 1584 35980 1636 36032
rect 2228 35980 2280 36032
rect 2596 35980 2648 36032
rect 3332 35980 3384 36032
rect 6092 36159 6144 36168
rect 6092 36125 6101 36159
rect 6101 36125 6135 36159
rect 6135 36125 6144 36159
rect 6092 36116 6144 36125
rect 7288 36116 7340 36168
rect 7656 36116 7708 36168
rect 7748 36159 7800 36168
rect 7748 36125 7755 36159
rect 7755 36125 7789 36159
rect 7789 36125 7800 36159
rect 7748 36116 7800 36125
rect 10600 36116 10652 36168
rect 5724 35980 5776 36032
rect 6184 35980 6236 36032
rect 8024 36048 8076 36100
rect 8300 36048 8352 36100
rect 6920 36023 6972 36032
rect 6920 35989 6929 36023
rect 6929 35989 6963 36023
rect 6963 35989 6972 36023
rect 6920 35980 6972 35989
rect 7840 35980 7892 36032
rect 8760 35980 8812 36032
rect 9128 35980 9180 36032
rect 9312 35980 9364 36032
rect 9772 35980 9824 36032
rect 11428 36116 11480 36168
rect 12164 36116 12216 36168
rect 13820 35980 13872 36032
rect 16028 36184 16080 36236
rect 16212 36184 16264 36236
rect 18052 36184 18104 36236
rect 19340 36184 19392 36236
rect 19892 36252 19944 36304
rect 20996 36252 21048 36304
rect 16488 36116 16540 36168
rect 18328 36116 18380 36168
rect 18972 36116 19024 36168
rect 19708 36155 19760 36168
rect 19708 36121 19717 36155
rect 19717 36121 19751 36155
rect 19751 36121 19760 36155
rect 19708 36116 19760 36121
rect 20444 36116 20496 36168
rect 21364 36116 21416 36168
rect 14740 36048 14792 36100
rect 18420 36048 18472 36100
rect 15844 35980 15896 36032
rect 18512 35980 18564 36032
rect 19064 35980 19116 36032
rect 22284 36048 22336 36100
rect 20444 36023 20496 36032
rect 20444 35989 20453 36023
rect 20453 35989 20487 36023
rect 20487 35989 20496 36023
rect 20444 35980 20496 35989
rect 20812 36023 20864 36032
rect 20812 35989 20821 36023
rect 20821 35989 20855 36023
rect 20855 35989 20864 36023
rect 20812 35980 20864 35989
rect 6148 35878 6200 35930
rect 6212 35878 6264 35930
rect 6276 35878 6328 35930
rect 6340 35878 6392 35930
rect 6404 35878 6456 35930
rect 11346 35878 11398 35930
rect 11410 35878 11462 35930
rect 11474 35878 11526 35930
rect 11538 35878 11590 35930
rect 11602 35878 11654 35930
rect 16544 35878 16596 35930
rect 16608 35878 16660 35930
rect 16672 35878 16724 35930
rect 16736 35878 16788 35930
rect 16800 35878 16852 35930
rect 21742 35878 21794 35930
rect 21806 35878 21858 35930
rect 21870 35878 21922 35930
rect 21934 35878 21986 35930
rect 21998 35878 22050 35930
rect 2872 35776 2924 35828
rect 4620 35776 4672 35828
rect 3516 35708 3568 35760
rect 5816 35776 5868 35828
rect 1768 35615 1820 35624
rect 1768 35581 1777 35615
rect 1777 35581 1811 35615
rect 1811 35581 1820 35615
rect 1768 35572 1820 35581
rect 2964 35683 3016 35692
rect 2964 35649 2973 35683
rect 2973 35649 3007 35683
rect 3007 35649 3016 35683
rect 2964 35640 3016 35649
rect 2136 35572 2188 35624
rect 2412 35615 2464 35624
rect 2412 35581 2421 35615
rect 2421 35581 2455 35615
rect 2455 35581 2464 35615
rect 2412 35572 2464 35581
rect 2228 35504 2280 35556
rect 2780 35615 2832 35624
rect 2780 35581 2814 35615
rect 2814 35581 2832 35615
rect 2780 35572 2832 35581
rect 3148 35572 3200 35624
rect 4252 35683 4304 35692
rect 4252 35649 4261 35683
rect 4261 35649 4295 35683
rect 4295 35649 4304 35683
rect 4252 35640 4304 35649
rect 4344 35640 4396 35692
rect 7564 35708 7616 35760
rect 13084 35776 13136 35828
rect 14556 35776 14608 35828
rect 8576 35708 8628 35760
rect 18972 35751 19024 35760
rect 7748 35640 7800 35692
rect 9312 35683 9364 35692
rect 9312 35649 9321 35683
rect 9321 35649 9355 35683
rect 9355 35649 9364 35683
rect 9312 35640 9364 35649
rect 11704 35640 11756 35692
rect 13452 35640 13504 35692
rect 1308 35436 1360 35488
rect 3976 35436 4028 35488
rect 4528 35615 4580 35624
rect 4528 35581 4537 35615
rect 4537 35581 4571 35615
rect 4571 35581 4580 35615
rect 4528 35572 4580 35581
rect 4896 35615 4948 35624
rect 4896 35581 4905 35615
rect 4905 35581 4939 35615
rect 4939 35581 4948 35615
rect 4896 35572 4948 35581
rect 6828 35572 6880 35624
rect 5724 35504 5776 35556
rect 6644 35504 6696 35556
rect 8576 35615 8628 35624
rect 8576 35581 8585 35615
rect 8585 35581 8619 35615
rect 8619 35581 8628 35615
rect 8576 35572 8628 35581
rect 8760 35572 8812 35624
rect 9429 35615 9481 35624
rect 9429 35581 9438 35615
rect 9438 35581 9472 35615
rect 9472 35581 9481 35615
rect 9429 35572 9481 35581
rect 9588 35615 9640 35624
rect 9588 35581 9597 35615
rect 9597 35581 9631 35615
rect 9631 35581 9640 35615
rect 9588 35572 9640 35581
rect 10968 35572 11020 35624
rect 11152 35572 11204 35624
rect 15200 35640 15252 35692
rect 16028 35640 16080 35692
rect 4896 35436 4948 35488
rect 8024 35479 8076 35488
rect 8024 35445 8033 35479
rect 8033 35445 8067 35479
rect 8067 35445 8076 35479
rect 8024 35436 8076 35445
rect 17040 35615 17092 35624
rect 17040 35581 17049 35615
rect 17049 35581 17083 35615
rect 17083 35581 17092 35615
rect 17040 35572 17092 35581
rect 12532 35504 12584 35556
rect 14280 35504 14332 35556
rect 17500 35504 17552 35556
rect 12164 35436 12216 35488
rect 12808 35479 12860 35488
rect 12808 35445 12817 35479
rect 12817 35445 12851 35479
rect 12851 35445 12860 35479
rect 12808 35436 12860 35445
rect 15292 35479 15344 35488
rect 15292 35445 15301 35479
rect 15301 35445 15335 35479
rect 15335 35445 15344 35479
rect 15292 35436 15344 35445
rect 17592 35436 17644 35488
rect 17776 35504 17828 35556
rect 18972 35717 18984 35751
rect 18984 35717 19024 35751
rect 18972 35708 19024 35717
rect 19708 35776 19760 35828
rect 21272 35776 21324 35828
rect 17960 35640 18012 35692
rect 18236 35640 18288 35692
rect 18328 35640 18380 35692
rect 18512 35640 18564 35692
rect 19524 35640 19576 35692
rect 20444 35640 20496 35692
rect 20996 35683 21048 35692
rect 20996 35649 21005 35683
rect 21005 35649 21039 35683
rect 21039 35649 21048 35683
rect 20996 35640 21048 35649
rect 21088 35640 21140 35692
rect 17960 35504 18012 35556
rect 18420 35547 18472 35556
rect 18420 35513 18429 35547
rect 18429 35513 18463 35547
rect 18463 35513 18472 35547
rect 18420 35504 18472 35513
rect 22836 35572 22888 35624
rect 22928 35572 22980 35624
rect 20720 35504 20772 35556
rect 20996 35436 21048 35488
rect 21456 35479 21508 35488
rect 21456 35445 21465 35479
rect 21465 35445 21499 35479
rect 21499 35445 21508 35479
rect 21456 35436 21508 35445
rect 3549 35334 3601 35386
rect 3613 35334 3665 35386
rect 3677 35334 3729 35386
rect 3741 35334 3793 35386
rect 3805 35334 3857 35386
rect 8747 35334 8799 35386
rect 8811 35334 8863 35386
rect 8875 35334 8927 35386
rect 8939 35334 8991 35386
rect 9003 35334 9055 35386
rect 13945 35334 13997 35386
rect 14009 35334 14061 35386
rect 14073 35334 14125 35386
rect 14137 35334 14189 35386
rect 14201 35334 14253 35386
rect 19143 35334 19195 35386
rect 19207 35334 19259 35386
rect 19271 35334 19323 35386
rect 19335 35334 19387 35386
rect 19399 35334 19451 35386
rect 3516 35232 3568 35284
rect 4160 35232 4212 35284
rect 4804 35232 4856 35284
rect 5356 35232 5408 35284
rect 5816 35232 5868 35284
rect 1768 35164 1820 35216
rect 1768 35028 1820 35080
rect 1676 35003 1728 35012
rect 1676 34969 1685 35003
rect 1685 34969 1719 35003
rect 1719 34969 1728 35003
rect 1676 34960 1728 34969
rect 4344 35164 4396 35216
rect 2688 35096 2740 35148
rect 4528 35096 4580 35148
rect 6644 35232 6696 35284
rect 7196 35232 7248 35284
rect 7288 35275 7340 35284
rect 7288 35241 7297 35275
rect 7297 35241 7331 35275
rect 7331 35241 7340 35275
rect 7288 35232 7340 35241
rect 11796 35232 11848 35284
rect 14556 35232 14608 35284
rect 7012 35164 7064 35216
rect 8300 35164 8352 35216
rect 12256 35207 12308 35216
rect 12256 35173 12265 35207
rect 12265 35173 12299 35207
rect 12299 35173 12308 35207
rect 12256 35164 12308 35173
rect 2136 35028 2188 35080
rect 2596 35071 2648 35080
rect 2596 35037 2605 35071
rect 2605 35037 2639 35071
rect 2639 35037 2648 35071
rect 2596 35028 2648 35037
rect 8024 35096 8076 35148
rect 12532 35139 12584 35148
rect 12532 35105 12541 35139
rect 12541 35105 12575 35139
rect 12575 35105 12584 35139
rect 12532 35096 12584 35105
rect 12808 35139 12860 35148
rect 12808 35105 12817 35139
rect 12817 35105 12851 35139
rect 12851 35105 12860 35139
rect 12808 35096 12860 35105
rect 15108 35232 15160 35284
rect 17040 35232 17092 35284
rect 16212 35096 16264 35148
rect 3608 34960 3660 35012
rect 3884 35003 3936 35012
rect 3884 34969 3893 35003
rect 3893 34969 3927 35003
rect 3927 34969 3936 35003
rect 3884 34960 3936 34969
rect 4068 34960 4120 35012
rect 1308 34892 1360 34944
rect 1860 34892 1912 34944
rect 2320 34892 2372 34944
rect 2872 34892 2924 34944
rect 3056 34892 3108 34944
rect 3516 34935 3568 34944
rect 3516 34901 3525 34935
rect 3525 34901 3559 34935
rect 3559 34901 3568 34935
rect 3516 34892 3568 34901
rect 4528 34935 4580 34944
rect 4528 34901 4537 34935
rect 4537 34901 4571 34935
rect 4571 34901 4580 34935
rect 4528 34892 4580 34901
rect 7288 35028 7340 35080
rect 8668 35028 8720 35080
rect 9496 35071 9548 35080
rect 9496 35037 9505 35071
rect 9505 35037 9539 35071
rect 9539 35037 9548 35071
rect 9496 35028 9548 35037
rect 6644 34960 6696 35012
rect 10600 35028 10652 35080
rect 11612 35071 11664 35080
rect 11612 35037 11621 35071
rect 11621 35037 11655 35071
rect 11655 35037 11664 35071
rect 11612 35028 11664 35037
rect 9864 35003 9916 35012
rect 9864 34969 9873 35003
rect 9873 34969 9907 35003
rect 9907 34969 9916 35003
rect 9864 34960 9916 34969
rect 10232 35003 10284 35012
rect 10232 34969 10241 35003
rect 10241 34969 10275 35003
rect 10275 34969 10284 35003
rect 10232 34960 10284 34969
rect 10876 34960 10928 35012
rect 11244 35003 11296 35012
rect 11244 34969 11253 35003
rect 11253 34969 11287 35003
rect 11287 34969 11296 35003
rect 11244 34960 11296 34969
rect 5816 34892 5868 34944
rect 6000 34892 6052 34944
rect 8024 34892 8076 34944
rect 9220 34892 9272 34944
rect 9496 34892 9548 34944
rect 9956 34892 10008 34944
rect 10508 34892 10560 34944
rect 11796 35071 11848 35080
rect 11796 35037 11805 35071
rect 11805 35037 11839 35071
rect 11839 35037 11848 35071
rect 11796 35028 11848 35037
rect 12624 35071 12676 35080
rect 12624 35037 12658 35071
rect 12658 35037 12676 35071
rect 12624 35028 12676 35037
rect 15200 34960 15252 35012
rect 12256 34892 12308 34944
rect 16212 34935 16264 34944
rect 16212 34901 16221 34935
rect 16221 34901 16255 34935
rect 16255 34901 16264 34935
rect 16212 34892 16264 34901
rect 16948 35028 17000 35080
rect 17500 35232 17552 35284
rect 17776 35275 17828 35284
rect 17776 35241 17785 35275
rect 17785 35241 17819 35275
rect 17819 35241 17828 35275
rect 17776 35232 17828 35241
rect 19708 35232 19760 35284
rect 20352 35232 20404 35284
rect 21180 35232 21232 35284
rect 16396 34960 16448 35012
rect 17040 34892 17092 34944
rect 19064 35028 19116 35080
rect 20536 35028 20588 35080
rect 18328 34892 18380 34944
rect 19616 34892 19668 34944
rect 20904 35028 20956 35080
rect 22008 34960 22060 35012
rect 22192 34892 22244 34944
rect 6148 34790 6200 34842
rect 6212 34790 6264 34842
rect 6276 34790 6328 34842
rect 6340 34790 6392 34842
rect 6404 34790 6456 34842
rect 11346 34790 11398 34842
rect 11410 34790 11462 34842
rect 11474 34790 11526 34842
rect 11538 34790 11590 34842
rect 11602 34790 11654 34842
rect 16544 34790 16596 34842
rect 16608 34790 16660 34842
rect 16672 34790 16724 34842
rect 16736 34790 16788 34842
rect 16800 34790 16852 34842
rect 21742 34790 21794 34842
rect 21806 34790 21858 34842
rect 21870 34790 21922 34842
rect 21934 34790 21986 34842
rect 21998 34790 22050 34842
rect 2136 34688 2188 34740
rect 4896 34688 4948 34740
rect 6000 34688 6052 34740
rect 6460 34688 6512 34740
rect 6828 34688 6880 34740
rect 7104 34688 7156 34740
rect 10416 34688 10468 34740
rect 2320 34620 2372 34672
rect 4528 34620 4580 34672
rect 4804 34663 4856 34672
rect 4804 34629 4813 34663
rect 4813 34629 4847 34663
rect 4847 34629 4856 34663
rect 4804 34620 4856 34629
rect 5080 34663 5132 34672
rect 5080 34629 5089 34663
rect 5089 34629 5123 34663
rect 5123 34629 5132 34663
rect 5080 34620 5132 34629
rect 5816 34620 5868 34672
rect 6092 34620 6144 34672
rect 9404 34620 9456 34672
rect 9680 34620 9732 34672
rect 10876 34731 10928 34740
rect 10876 34697 10885 34731
rect 10885 34697 10919 34731
rect 10919 34697 10928 34731
rect 10876 34688 10928 34697
rect 11336 34620 11388 34672
rect 2044 34552 2096 34604
rect 2596 34552 2648 34604
rect 4896 34552 4948 34604
rect 6000 34552 6052 34604
rect 2964 34484 3016 34536
rect 4988 34484 5040 34536
rect 5908 34484 5960 34536
rect 7196 34552 7248 34604
rect 7932 34595 7984 34604
rect 388 34348 440 34400
rect 2872 34391 2924 34400
rect 2872 34357 2881 34391
rect 2881 34357 2915 34391
rect 2915 34357 2924 34391
rect 2872 34348 2924 34357
rect 6828 34416 6880 34468
rect 4252 34391 4304 34400
rect 4252 34357 4261 34391
rect 4261 34357 4295 34391
rect 4295 34357 4304 34391
rect 4252 34348 4304 34357
rect 4620 34348 4672 34400
rect 7932 34561 7939 34595
rect 7939 34561 7973 34595
rect 7973 34561 7984 34595
rect 7932 34552 7984 34561
rect 9588 34595 9640 34604
rect 9588 34561 9597 34595
rect 9597 34561 9631 34595
rect 9631 34561 9640 34595
rect 9588 34552 9640 34561
rect 9956 34595 10008 34604
rect 9956 34561 9965 34595
rect 9965 34561 9999 34595
rect 9999 34561 10008 34595
rect 9956 34552 10008 34561
rect 10048 34552 10100 34604
rect 10692 34552 10744 34604
rect 12624 34552 12676 34604
rect 13084 34620 13136 34672
rect 15292 34688 15344 34740
rect 16028 34731 16080 34740
rect 16028 34697 16037 34731
rect 16037 34697 16071 34731
rect 16071 34697 16080 34731
rect 16028 34688 16080 34697
rect 16212 34688 16264 34740
rect 16396 34688 16448 34740
rect 18052 34688 18104 34740
rect 18788 34688 18840 34740
rect 19524 34688 19576 34740
rect 19892 34688 19944 34740
rect 13820 34620 13872 34672
rect 14280 34552 14332 34604
rect 16948 34595 17000 34604
rect 16948 34561 16957 34595
rect 16957 34561 16991 34595
rect 16991 34561 17000 34595
rect 16948 34552 17000 34561
rect 17040 34552 17092 34604
rect 17960 34552 18012 34604
rect 20168 34688 20220 34740
rect 20444 34688 20496 34740
rect 20720 34688 20772 34740
rect 20812 34620 20864 34672
rect 10600 34416 10652 34468
rect 20168 34595 20220 34604
rect 20168 34561 20177 34595
rect 20177 34561 20211 34595
rect 20211 34561 20220 34595
rect 20168 34552 20220 34561
rect 20444 34595 20496 34604
rect 20444 34561 20453 34595
rect 20453 34561 20487 34595
rect 20487 34561 20496 34595
rect 20444 34552 20496 34561
rect 20904 34552 20956 34604
rect 22284 34552 22336 34604
rect 21364 34484 21416 34536
rect 8484 34348 8536 34400
rect 11060 34348 11112 34400
rect 13820 34348 13872 34400
rect 15384 34391 15436 34400
rect 15384 34357 15393 34391
rect 15393 34357 15427 34391
rect 15427 34357 15436 34391
rect 15384 34348 15436 34357
rect 16212 34348 16264 34400
rect 17960 34348 18012 34400
rect 18604 34348 18656 34400
rect 21088 34348 21140 34400
rect 21456 34391 21508 34400
rect 21456 34357 21465 34391
rect 21465 34357 21499 34391
rect 21499 34357 21508 34391
rect 21456 34348 21508 34357
rect 3549 34246 3601 34298
rect 3613 34246 3665 34298
rect 3677 34246 3729 34298
rect 3741 34246 3793 34298
rect 3805 34246 3857 34298
rect 8747 34246 8799 34298
rect 8811 34246 8863 34298
rect 8875 34246 8927 34298
rect 8939 34246 8991 34298
rect 9003 34246 9055 34298
rect 13945 34246 13997 34298
rect 14009 34246 14061 34298
rect 14073 34246 14125 34298
rect 14137 34246 14189 34298
rect 14201 34246 14253 34298
rect 19143 34246 19195 34298
rect 19207 34246 19259 34298
rect 19271 34246 19323 34298
rect 19335 34246 19387 34298
rect 19399 34246 19451 34298
rect 4252 34144 4304 34196
rect 2780 34076 2832 34128
rect 4528 34076 4580 34128
rect 2688 34008 2740 34060
rect 3976 34008 4028 34060
rect 8116 34144 8168 34196
rect 9588 34144 9640 34196
rect 7564 34076 7616 34128
rect 8760 34076 8812 34128
rect 11060 34144 11112 34196
rect 12164 34144 12216 34196
rect 13912 34144 13964 34196
rect 15200 34144 15252 34196
rect 7380 34008 7432 34060
rect 8116 34008 8168 34060
rect 9036 34008 9088 34060
rect 2964 33983 3016 33992
rect 2964 33949 2973 33983
rect 2973 33949 3007 33983
rect 3007 33949 3016 33983
rect 2964 33940 3016 33949
rect 1860 33919 1885 33924
rect 1885 33919 1912 33924
rect 1860 33872 1912 33919
rect 2412 33804 2464 33856
rect 2596 33847 2648 33856
rect 2596 33813 2605 33847
rect 2605 33813 2639 33847
rect 2639 33813 2648 33847
rect 2596 33804 2648 33813
rect 3332 33940 3384 33992
rect 5080 33940 5132 33992
rect 5448 33940 5500 33992
rect 6000 33940 6052 33992
rect 6552 33940 6604 33992
rect 7012 33940 7064 33992
rect 7104 33940 7156 33992
rect 18236 34144 18288 34196
rect 20444 34144 20496 34196
rect 21180 34144 21232 34196
rect 10692 34051 10744 34060
rect 10692 34017 10701 34051
rect 10701 34017 10735 34051
rect 10735 34017 10744 34051
rect 10692 34008 10744 34017
rect 13176 34008 13228 34060
rect 14280 34008 14332 34060
rect 16304 34051 16356 34060
rect 16304 34017 16313 34051
rect 16313 34017 16347 34051
rect 16347 34017 16356 34051
rect 16304 34008 16356 34017
rect 4344 33872 4396 33924
rect 4804 33872 4856 33924
rect 10416 33940 10468 33992
rect 4988 33804 5040 33856
rect 5172 33804 5224 33856
rect 5264 33804 5316 33856
rect 6092 33804 6144 33856
rect 8024 33872 8076 33924
rect 12900 33872 12952 33924
rect 14556 33940 14608 33992
rect 14740 33940 14792 33992
rect 15292 33872 15344 33924
rect 16948 33872 17000 33924
rect 18052 34008 18104 34060
rect 18604 34008 18656 34060
rect 17960 33940 18012 33992
rect 6644 33804 6696 33856
rect 6920 33804 6972 33856
rect 9312 33804 9364 33856
rect 9588 33804 9640 33856
rect 10968 33804 11020 33856
rect 13544 33804 13596 33856
rect 15936 33847 15988 33856
rect 15936 33813 15945 33847
rect 15945 33813 15979 33847
rect 15979 33813 15988 33847
rect 15936 33804 15988 33813
rect 19432 33983 19484 33992
rect 19432 33949 19441 33983
rect 19441 33949 19475 33983
rect 19475 33949 19484 33983
rect 19432 33940 19484 33949
rect 19892 33983 19944 33992
rect 19892 33949 19901 33983
rect 19901 33949 19935 33983
rect 19935 33949 19944 33983
rect 19892 33940 19944 33949
rect 19156 33872 19208 33924
rect 20352 33983 20404 33992
rect 20352 33949 20361 33983
rect 20361 33949 20395 33983
rect 20395 33949 20404 33983
rect 20352 33940 20404 33949
rect 20628 33983 20680 33992
rect 20628 33949 20637 33983
rect 20637 33949 20671 33983
rect 20671 33949 20680 33983
rect 20628 33940 20680 33949
rect 20720 33940 20772 33992
rect 21456 34008 21508 34060
rect 21272 33983 21324 33992
rect 21272 33949 21281 33983
rect 21281 33949 21315 33983
rect 21315 33949 21324 33983
rect 21272 33940 21324 33949
rect 20260 33872 20312 33924
rect 20536 33872 20588 33924
rect 19708 33847 19760 33856
rect 19708 33813 19717 33847
rect 19717 33813 19751 33847
rect 19751 33813 19760 33847
rect 19708 33804 19760 33813
rect 20720 33804 20772 33856
rect 20812 33847 20864 33856
rect 20812 33813 20821 33847
rect 20821 33813 20855 33847
rect 20855 33813 20864 33847
rect 20812 33804 20864 33813
rect 21272 33804 21324 33856
rect 22192 33804 22244 33856
rect 6148 33702 6200 33754
rect 6212 33702 6264 33754
rect 6276 33702 6328 33754
rect 6340 33702 6392 33754
rect 6404 33702 6456 33754
rect 11346 33702 11398 33754
rect 11410 33702 11462 33754
rect 11474 33702 11526 33754
rect 11538 33702 11590 33754
rect 11602 33702 11654 33754
rect 16544 33702 16596 33754
rect 16608 33702 16660 33754
rect 16672 33702 16724 33754
rect 16736 33702 16788 33754
rect 16800 33702 16852 33754
rect 21742 33702 21794 33754
rect 21806 33702 21858 33754
rect 21870 33702 21922 33754
rect 21934 33702 21986 33754
rect 21998 33702 22050 33754
rect 2780 33532 2832 33584
rect 3884 33532 3936 33584
rect 1400 33507 1452 33516
rect 1400 33473 1409 33507
rect 1409 33473 1443 33507
rect 1443 33473 1452 33507
rect 1400 33464 1452 33473
rect 1952 33507 2004 33516
rect 1952 33473 1961 33507
rect 1961 33473 1995 33507
rect 1995 33473 2004 33507
rect 1952 33464 2004 33473
rect 3240 33507 3292 33516
rect 3240 33473 3249 33507
rect 3249 33473 3283 33507
rect 3283 33473 3292 33507
rect 3240 33464 3292 33473
rect 4804 33464 4856 33516
rect 5080 33532 5132 33584
rect 5540 33532 5592 33584
rect 6736 33532 6788 33584
rect 5908 33464 5960 33516
rect 8024 33464 8076 33516
rect 9680 33532 9732 33584
rect 10876 33532 10928 33584
rect 11060 33532 11112 33584
rect 12072 33532 12124 33584
rect 13084 33532 13136 33584
rect 10416 33464 10468 33516
rect 10784 33464 10836 33516
rect 13360 33532 13412 33584
rect 15384 33600 15436 33652
rect 13728 33532 13780 33584
rect 14280 33575 14332 33584
rect 14280 33541 14289 33575
rect 14289 33541 14323 33575
rect 14323 33541 14332 33575
rect 14280 33532 14332 33541
rect 14556 33532 14608 33584
rect 15016 33532 15068 33584
rect 16580 33532 16632 33584
rect 17132 33600 17184 33652
rect 19156 33643 19208 33652
rect 19156 33609 19165 33643
rect 19165 33609 19199 33643
rect 19199 33609 19208 33643
rect 19156 33600 19208 33609
rect 19708 33600 19760 33652
rect 19892 33600 19944 33652
rect 2044 33396 2096 33448
rect 2228 33439 2280 33448
rect 2228 33405 2237 33439
rect 2237 33405 2271 33439
rect 2271 33405 2280 33439
rect 2228 33396 2280 33405
rect 2872 33396 2924 33448
rect 3976 33396 4028 33448
rect 4252 33396 4304 33448
rect 5356 33396 5408 33448
rect 6736 33396 6788 33448
rect 8484 33396 8536 33448
rect 9036 33439 9088 33448
rect 9036 33405 9045 33439
rect 9045 33405 9079 33439
rect 9079 33405 9088 33439
rect 9036 33396 9088 33405
rect 9772 33396 9824 33448
rect 9956 33396 10008 33448
rect 11152 33396 11204 33448
rect 11428 33396 11480 33448
rect 13820 33396 13872 33448
rect 14464 33396 14516 33448
rect 7012 33328 7064 33380
rect 5632 33303 5684 33312
rect 5632 33269 5641 33303
rect 5641 33269 5675 33303
rect 5675 33269 5684 33303
rect 5632 33260 5684 33269
rect 5816 33260 5868 33312
rect 6920 33260 6972 33312
rect 7104 33260 7156 33312
rect 9772 33260 9824 33312
rect 10784 33303 10836 33312
rect 10784 33269 10793 33303
rect 10793 33269 10827 33303
rect 10827 33269 10836 33303
rect 10784 33260 10836 33269
rect 11244 33260 11296 33312
rect 12624 33260 12676 33312
rect 12808 33260 12860 33312
rect 12992 33260 13044 33312
rect 15844 33464 15896 33516
rect 16764 33396 16816 33448
rect 17224 33507 17276 33516
rect 17224 33473 17233 33507
rect 17233 33473 17267 33507
rect 17267 33473 17276 33507
rect 17224 33464 17276 33473
rect 20996 33575 21048 33584
rect 20996 33541 21005 33575
rect 21005 33541 21039 33575
rect 21039 33541 21048 33575
rect 20996 33532 21048 33541
rect 19340 33507 19392 33516
rect 19340 33473 19349 33507
rect 19349 33473 19383 33507
rect 19383 33473 19392 33507
rect 19340 33464 19392 33473
rect 19708 33464 19760 33516
rect 18880 33396 18932 33448
rect 20352 33464 20404 33516
rect 16580 33328 16632 33380
rect 17132 33328 17184 33380
rect 15660 33303 15712 33312
rect 15660 33269 15669 33303
rect 15669 33269 15703 33303
rect 15703 33269 15712 33303
rect 15660 33260 15712 33269
rect 18052 33260 18104 33312
rect 19892 33260 19944 33312
rect 20444 33260 20496 33312
rect 21180 33260 21232 33312
rect 21272 33303 21324 33312
rect 21272 33269 21281 33303
rect 21281 33269 21315 33303
rect 21315 33269 21324 33303
rect 21272 33260 21324 33269
rect 3549 33158 3601 33210
rect 3613 33158 3665 33210
rect 3677 33158 3729 33210
rect 3741 33158 3793 33210
rect 3805 33158 3857 33210
rect 8747 33158 8799 33210
rect 8811 33158 8863 33210
rect 8875 33158 8927 33210
rect 8939 33158 8991 33210
rect 9003 33158 9055 33210
rect 13945 33158 13997 33210
rect 14009 33158 14061 33210
rect 14073 33158 14125 33210
rect 14137 33158 14189 33210
rect 14201 33158 14253 33210
rect 19143 33158 19195 33210
rect 19207 33158 19259 33210
rect 19271 33158 19323 33210
rect 19335 33158 19387 33210
rect 19399 33158 19451 33210
rect 2412 33056 2464 33108
rect 3240 33056 3292 33108
rect 4896 33056 4948 33108
rect 5080 33056 5132 33108
rect 6644 33056 6696 33108
rect 7380 33056 7432 33108
rect 1124 32920 1176 32972
rect 1584 32920 1636 32972
rect 2136 32920 2188 32972
rect 5356 32988 5408 33040
rect 5632 32920 5684 32972
rect 1492 32827 1544 32836
rect 1492 32793 1501 32827
rect 1501 32793 1535 32827
rect 1535 32793 1544 32827
rect 1492 32784 1544 32793
rect 1768 32784 1820 32836
rect 3792 32784 3844 32836
rect 5540 32852 5592 32904
rect 5172 32784 5224 32836
rect 5356 32784 5408 32836
rect 5816 32895 5868 32904
rect 5816 32861 5825 32895
rect 5825 32861 5859 32895
rect 5859 32861 5868 32895
rect 5816 32852 5868 32861
rect 388 32716 440 32768
rect 3148 32716 3200 32768
rect 4068 32716 4120 32768
rect 4896 32716 4948 32768
rect 5448 32759 5500 32768
rect 5448 32725 5457 32759
rect 5457 32725 5491 32759
rect 5491 32725 5500 32759
rect 5448 32716 5500 32725
rect 6920 32895 6972 32904
rect 6920 32861 6929 32895
rect 6929 32861 6963 32895
rect 6963 32861 6972 32895
rect 6920 32852 6972 32861
rect 6000 32784 6052 32836
rect 6552 32759 6604 32768
rect 6552 32725 6561 32759
rect 6561 32725 6595 32759
rect 6595 32725 6604 32759
rect 6552 32716 6604 32725
rect 6736 32716 6788 32768
rect 8392 33056 8444 33108
rect 8484 32920 8536 32972
rect 8852 32920 8904 32972
rect 7104 32852 7156 32904
rect 7380 32895 7432 32904
rect 7380 32861 7389 32895
rect 7389 32861 7423 32895
rect 7423 32861 7432 32895
rect 7380 32852 7432 32861
rect 8392 32852 8444 32904
rect 7564 32784 7616 32836
rect 9312 32831 9337 32836
rect 9337 32831 9364 32836
rect 9312 32784 9364 32831
rect 10968 32920 11020 32972
rect 14556 32988 14608 33040
rect 15660 33056 15712 33108
rect 15752 33056 15804 33108
rect 17500 33056 17552 33108
rect 17960 33056 18012 33108
rect 18052 33099 18104 33108
rect 18052 33065 18061 33099
rect 18061 33065 18095 33099
rect 18095 33065 18104 33099
rect 18052 33056 18104 33065
rect 18144 33056 18196 33108
rect 18328 32988 18380 33040
rect 12624 32963 12676 32972
rect 12624 32929 12633 32963
rect 12633 32929 12667 32963
rect 12667 32929 12676 32963
rect 12624 32920 12676 32929
rect 10876 32895 10928 32904
rect 10876 32861 10885 32895
rect 10885 32861 10919 32895
rect 10919 32861 10928 32895
rect 10876 32852 10928 32861
rect 11244 32852 11296 32904
rect 11704 32895 11756 32904
rect 11704 32861 11727 32895
rect 11727 32861 11756 32895
rect 11704 32852 11756 32861
rect 12532 32852 12584 32904
rect 15936 32920 15988 32972
rect 16304 32920 16356 32972
rect 7104 32716 7156 32768
rect 7932 32716 7984 32768
rect 8484 32759 8536 32768
rect 8484 32725 8493 32759
rect 8493 32725 8527 32759
rect 8527 32725 8536 32759
rect 8484 32716 8536 32725
rect 10048 32759 10100 32768
rect 10048 32725 10057 32759
rect 10057 32725 10091 32759
rect 10091 32725 10100 32759
rect 10048 32716 10100 32725
rect 10784 32716 10836 32768
rect 12532 32716 12584 32768
rect 12624 32716 12676 32768
rect 14372 32852 14424 32904
rect 14280 32784 14332 32836
rect 15476 32895 15528 32904
rect 15476 32861 15485 32895
rect 15485 32861 15519 32895
rect 15519 32861 15528 32895
rect 15476 32852 15528 32861
rect 18144 32920 18196 32972
rect 18880 33099 18932 33108
rect 18880 33065 18889 33099
rect 18889 33065 18923 33099
rect 18923 33065 18932 33099
rect 18880 33056 18932 33065
rect 20812 33056 20864 33108
rect 20628 32988 20680 33040
rect 16764 32827 16816 32836
rect 16764 32793 16798 32827
rect 16798 32793 16816 32827
rect 16764 32784 16816 32793
rect 18328 32852 18380 32904
rect 13360 32716 13412 32768
rect 17868 32716 17920 32768
rect 18236 32759 18288 32768
rect 18236 32725 18245 32759
rect 18245 32725 18279 32759
rect 18279 32725 18288 32759
rect 18236 32716 18288 32725
rect 18880 32852 18932 32904
rect 19156 32852 19208 32904
rect 21640 32988 21692 33040
rect 22836 32920 22888 32972
rect 20812 32895 20864 32904
rect 20812 32861 20821 32895
rect 20821 32861 20855 32895
rect 20855 32861 20864 32895
rect 20812 32852 20864 32861
rect 20904 32852 20956 32904
rect 21180 32852 21232 32904
rect 21548 32895 21600 32904
rect 21548 32861 21557 32895
rect 21557 32861 21591 32895
rect 21591 32861 21600 32895
rect 21548 32852 21600 32861
rect 19708 32784 19760 32836
rect 18788 32716 18840 32768
rect 19984 32716 20036 32768
rect 22836 32784 22888 32836
rect 21364 32759 21416 32768
rect 21364 32725 21373 32759
rect 21373 32725 21407 32759
rect 21407 32725 21416 32759
rect 21364 32716 21416 32725
rect 6148 32614 6200 32666
rect 6212 32614 6264 32666
rect 6276 32614 6328 32666
rect 6340 32614 6392 32666
rect 6404 32614 6456 32666
rect 11346 32614 11398 32666
rect 11410 32614 11462 32666
rect 11474 32614 11526 32666
rect 11538 32614 11590 32666
rect 11602 32614 11654 32666
rect 16544 32614 16596 32666
rect 16608 32614 16660 32666
rect 16672 32614 16724 32666
rect 16736 32614 16788 32666
rect 16800 32614 16852 32666
rect 21742 32614 21794 32666
rect 21806 32614 21858 32666
rect 21870 32614 21922 32666
rect 21934 32614 21986 32666
rect 21998 32614 22050 32666
rect 2780 32512 2832 32564
rect 3148 32512 3200 32564
rect 4160 32512 4212 32564
rect 4712 32512 4764 32564
rect 5816 32512 5868 32564
rect 6920 32512 6972 32564
rect 7380 32512 7432 32564
rect 756 32444 808 32496
rect 2320 32376 2372 32428
rect 3240 32487 3292 32496
rect 3240 32453 3249 32487
rect 3249 32453 3283 32487
rect 3283 32453 3292 32487
rect 3240 32444 3292 32453
rect 3884 32444 3936 32496
rect 6736 32444 6788 32496
rect 7196 32419 7248 32428
rect 7196 32385 7205 32419
rect 7205 32385 7239 32419
rect 7239 32385 7248 32419
rect 7196 32376 7248 32385
rect 7380 32386 7432 32438
rect 8944 32512 8996 32564
rect 9036 32444 9088 32496
rect 9312 32512 9364 32564
rect 10968 32512 11020 32564
rect 11796 32512 11848 32564
rect 12532 32512 12584 32564
rect 13084 32512 13136 32564
rect 13452 32512 13504 32564
rect 13912 32512 13964 32564
rect 15936 32512 15988 32564
rect 17868 32555 17920 32564
rect 17868 32521 17877 32555
rect 17877 32521 17911 32555
rect 17911 32521 17920 32555
rect 17868 32512 17920 32521
rect 1400 32308 1452 32360
rect 2596 32308 2648 32360
rect 3332 32308 3384 32360
rect 4252 32240 4304 32292
rect 1584 32172 1636 32224
rect 2964 32172 3016 32224
rect 4712 32308 4764 32360
rect 4896 32351 4948 32360
rect 4896 32317 4905 32351
rect 4905 32317 4939 32351
rect 4939 32317 4948 32351
rect 4896 32308 4948 32317
rect 6184 32308 6236 32360
rect 7012 32308 7064 32360
rect 7564 32419 7616 32428
rect 7564 32385 7571 32419
rect 7571 32385 7605 32419
rect 7605 32385 7616 32419
rect 9772 32444 9824 32496
rect 10232 32487 10284 32496
rect 10232 32453 10241 32487
rect 10241 32453 10275 32487
rect 10275 32453 10284 32487
rect 10232 32444 10284 32453
rect 10416 32444 10468 32496
rect 7564 32376 7616 32385
rect 9680 32376 9732 32428
rect 10692 32376 10744 32428
rect 11060 32419 11112 32428
rect 11060 32385 11069 32419
rect 11069 32385 11103 32419
rect 11103 32385 11112 32419
rect 11060 32376 11112 32385
rect 11336 32376 11388 32428
rect 12808 32376 12860 32428
rect 13636 32376 13688 32428
rect 13820 32376 13872 32428
rect 15476 32376 15528 32428
rect 17684 32444 17736 32496
rect 17960 32444 18012 32496
rect 18972 32376 19024 32428
rect 19984 32444 20036 32496
rect 20076 32444 20128 32496
rect 20628 32555 20680 32564
rect 20628 32521 20637 32555
rect 20637 32521 20671 32555
rect 20671 32521 20680 32555
rect 20628 32512 20680 32521
rect 20812 32512 20864 32564
rect 21180 32512 21232 32564
rect 19432 32419 19484 32428
rect 19432 32385 19441 32419
rect 19441 32385 19475 32419
rect 19475 32385 19484 32419
rect 19432 32376 19484 32385
rect 19524 32376 19576 32428
rect 19616 32419 19668 32428
rect 19616 32385 19625 32419
rect 19625 32385 19659 32419
rect 19659 32385 19668 32419
rect 19616 32376 19668 32385
rect 21180 32419 21232 32428
rect 21180 32385 21189 32419
rect 21189 32385 21223 32419
rect 21223 32385 21232 32419
rect 21180 32376 21232 32385
rect 22284 32444 22336 32496
rect 8484 32308 8536 32360
rect 13544 32308 13596 32360
rect 13912 32308 13964 32360
rect 5908 32240 5960 32292
rect 8852 32240 8904 32292
rect 10416 32283 10468 32292
rect 10416 32249 10425 32283
rect 10425 32249 10459 32283
rect 10459 32249 10468 32283
rect 10416 32240 10468 32249
rect 6000 32172 6052 32224
rect 6644 32172 6696 32224
rect 8024 32172 8076 32224
rect 8576 32172 8628 32224
rect 10324 32172 10376 32224
rect 10692 32172 10744 32224
rect 11244 32240 11296 32292
rect 11796 32240 11848 32292
rect 13636 32215 13688 32224
rect 13636 32181 13645 32215
rect 13645 32181 13679 32215
rect 13679 32181 13688 32215
rect 13636 32172 13688 32181
rect 15660 32240 15712 32292
rect 18788 32308 18840 32360
rect 14372 32172 14424 32224
rect 15016 32215 15068 32224
rect 15016 32181 15025 32215
rect 15025 32181 15059 32215
rect 15059 32181 15068 32215
rect 15016 32172 15068 32181
rect 15752 32172 15804 32224
rect 16212 32172 16264 32224
rect 16488 32172 16540 32224
rect 16856 32172 16908 32224
rect 17132 32172 17184 32224
rect 17960 32172 18012 32224
rect 19708 32172 19760 32224
rect 19892 32172 19944 32224
rect 21456 32308 21508 32360
rect 22284 32308 22336 32360
rect 22744 32308 22796 32360
rect 22836 32240 22888 32292
rect 20904 32172 20956 32224
rect 20996 32215 21048 32224
rect 20996 32181 21005 32215
rect 21005 32181 21039 32215
rect 21039 32181 21048 32215
rect 20996 32172 21048 32181
rect 21456 32215 21508 32224
rect 21456 32181 21465 32215
rect 21465 32181 21499 32215
rect 21499 32181 21508 32215
rect 21456 32172 21508 32181
rect 3549 32070 3601 32122
rect 3613 32070 3665 32122
rect 3677 32070 3729 32122
rect 3741 32070 3793 32122
rect 3805 32070 3857 32122
rect 8747 32070 8799 32122
rect 8811 32070 8863 32122
rect 8875 32070 8927 32122
rect 8939 32070 8991 32122
rect 9003 32070 9055 32122
rect 13945 32070 13997 32122
rect 14009 32070 14061 32122
rect 14073 32070 14125 32122
rect 14137 32070 14189 32122
rect 14201 32070 14253 32122
rect 19143 32070 19195 32122
rect 19207 32070 19259 32122
rect 19271 32070 19323 32122
rect 19335 32070 19387 32122
rect 19399 32070 19451 32122
rect 22836 32036 22888 32088
rect 2412 31968 2464 32020
rect 3332 31968 3384 32020
rect 5172 31968 5224 32020
rect 5540 31968 5592 32020
rect 7196 31968 7248 32020
rect 1400 31807 1452 31816
rect 1400 31773 1409 31807
rect 1409 31773 1443 31807
rect 1443 31773 1452 31807
rect 1400 31764 1452 31773
rect 1768 31807 1820 31816
rect 1768 31773 1777 31807
rect 1777 31773 1811 31807
rect 1811 31773 1820 31807
rect 1768 31764 1820 31773
rect 1860 31764 1912 31816
rect 2412 31875 2464 31884
rect 2412 31841 2421 31875
rect 2421 31841 2455 31875
rect 2455 31841 2464 31875
rect 2412 31832 2464 31841
rect 2780 31875 2832 31884
rect 2780 31841 2814 31875
rect 2814 31841 2832 31875
rect 2780 31832 2832 31841
rect 2964 31807 3016 31816
rect 2964 31773 2973 31807
rect 2973 31773 3007 31807
rect 3007 31773 3016 31807
rect 2964 31764 3016 31773
rect 3792 31807 3844 31816
rect 3792 31773 3801 31807
rect 3801 31773 3835 31807
rect 3835 31773 3844 31807
rect 3792 31764 3844 31773
rect 4068 31807 4120 31816
rect 4068 31773 4077 31807
rect 4077 31773 4111 31807
rect 4111 31773 4120 31807
rect 4068 31764 4120 31773
rect 4896 31832 4948 31884
rect 5264 31832 5316 31884
rect 5724 31832 5776 31884
rect 6000 31875 6052 31884
rect 6000 31841 6034 31875
rect 6034 31841 6052 31875
rect 6000 31832 6052 31841
rect 7380 31832 7432 31884
rect 10048 31968 10100 32020
rect 10876 31968 10928 32020
rect 4436 31764 4488 31816
rect 4528 31764 4580 31816
rect 4712 31807 4764 31816
rect 4712 31773 4721 31807
rect 4721 31773 4755 31807
rect 4755 31773 4764 31807
rect 4712 31764 4764 31773
rect 6184 31807 6236 31816
rect 6184 31773 6193 31807
rect 6193 31773 6227 31807
rect 6227 31773 6236 31807
rect 6184 31764 6236 31773
rect 9588 31832 9640 31884
rect 10324 31832 10376 31884
rect 10692 31875 10744 31884
rect 10692 31841 10701 31875
rect 10701 31841 10735 31875
rect 10735 31841 10744 31875
rect 10692 31832 10744 31841
rect 11152 31832 11204 31884
rect 8484 31764 8536 31816
rect 9956 31807 10008 31816
rect 9956 31773 9965 31807
rect 9965 31773 9999 31807
rect 9999 31773 10008 31807
rect 9956 31764 10008 31773
rect 10968 31807 11020 31816
rect 10968 31773 10977 31807
rect 10977 31773 11011 31807
rect 11011 31773 11020 31807
rect 10968 31764 11020 31773
rect 13912 31900 13964 31952
rect 15016 31968 15068 32020
rect 16488 31968 16540 32020
rect 15936 31900 15988 31952
rect 13360 31832 13412 31884
rect 13636 31832 13688 31884
rect 14280 31875 14332 31884
rect 12624 31764 12676 31816
rect 7656 31696 7708 31748
rect 7932 31696 7984 31748
rect 9312 31696 9364 31748
rect 1860 31628 1912 31680
rect 4160 31628 4212 31680
rect 4252 31628 4304 31680
rect 4712 31628 4764 31680
rect 4896 31628 4948 31680
rect 5356 31628 5408 31680
rect 6000 31628 6052 31680
rect 6276 31628 6328 31680
rect 7288 31628 7340 31680
rect 8208 31628 8260 31680
rect 8484 31671 8536 31680
rect 8484 31637 8493 31671
rect 8493 31637 8527 31671
rect 8527 31637 8536 31671
rect 8484 31628 8536 31637
rect 8576 31628 8628 31680
rect 9680 31628 9732 31680
rect 13360 31696 13412 31748
rect 13544 31696 13596 31748
rect 14280 31841 14289 31875
rect 14289 31841 14323 31875
rect 14323 31841 14332 31875
rect 14280 31832 14332 31841
rect 14096 31807 14148 31816
rect 14096 31773 14105 31807
rect 14105 31773 14139 31807
rect 14139 31773 14148 31807
rect 14096 31764 14148 31773
rect 15660 31832 15712 31884
rect 17224 31832 17276 31884
rect 18880 31968 18932 32020
rect 19892 31968 19944 32020
rect 19984 32011 20036 32020
rect 19984 31977 19993 32011
rect 19993 31977 20027 32011
rect 20027 31977 20036 32011
rect 19984 31968 20036 31977
rect 21548 31968 21600 32020
rect 10232 31628 10284 31680
rect 10784 31628 10836 31680
rect 12164 31628 12216 31680
rect 15108 31807 15160 31816
rect 15108 31773 15142 31807
rect 15142 31773 15160 31807
rect 15108 31764 15160 31773
rect 16212 31764 16264 31816
rect 16948 31764 17000 31816
rect 18328 31807 18380 31816
rect 18328 31773 18337 31807
rect 18337 31773 18371 31807
rect 18371 31773 18380 31807
rect 18328 31764 18380 31773
rect 20904 31900 20956 31952
rect 18972 31764 19024 31816
rect 19708 31832 19760 31884
rect 19800 31807 19852 31816
rect 19800 31773 19809 31807
rect 19809 31773 19843 31807
rect 19843 31773 19852 31807
rect 19800 31764 19852 31773
rect 20720 31875 20772 31884
rect 20720 31841 20729 31875
rect 20729 31841 20763 31875
rect 20763 31841 20772 31875
rect 20720 31832 20772 31841
rect 20444 31807 20496 31816
rect 20444 31773 20453 31807
rect 20453 31773 20487 31807
rect 20487 31773 20496 31807
rect 20444 31764 20496 31773
rect 19708 31696 19760 31748
rect 21088 31764 21140 31816
rect 22560 31714 22612 31766
rect 22928 31764 22980 31816
rect 14832 31628 14884 31680
rect 15568 31628 15620 31680
rect 18144 31628 18196 31680
rect 18512 31671 18564 31680
rect 18512 31637 18521 31671
rect 18521 31637 18555 31671
rect 18555 31637 18564 31671
rect 18512 31628 18564 31637
rect 20076 31628 20128 31680
rect 22192 31628 22244 31680
rect 6148 31526 6200 31578
rect 6212 31526 6264 31578
rect 6276 31526 6328 31578
rect 6340 31526 6392 31578
rect 6404 31526 6456 31578
rect 11346 31526 11398 31578
rect 11410 31526 11462 31578
rect 11474 31526 11526 31578
rect 11538 31526 11590 31578
rect 11602 31526 11654 31578
rect 16544 31526 16596 31578
rect 16608 31526 16660 31578
rect 16672 31526 16724 31578
rect 16736 31526 16788 31578
rect 16800 31526 16852 31578
rect 21742 31526 21794 31578
rect 21806 31526 21858 31578
rect 21870 31526 21922 31578
rect 21934 31526 21986 31578
rect 21998 31526 22050 31578
rect 2412 31467 2464 31476
rect 2412 31433 2421 31467
rect 2421 31433 2455 31467
rect 2455 31433 2464 31467
rect 2412 31424 2464 31433
rect 2780 31424 2832 31476
rect 1308 31356 1360 31408
rect 1492 31356 1544 31408
rect 2136 31356 2188 31408
rect 2596 31356 2648 31408
rect 2044 31288 2096 31340
rect 2504 31288 2556 31340
rect 2688 31288 2740 31340
rect 2780 31288 2832 31340
rect 3332 31424 3384 31476
rect 6460 31424 6512 31476
rect 7380 31424 7432 31476
rect 6736 31356 6788 31408
rect 10416 31356 10468 31408
rect 10968 31424 11020 31476
rect 2872 31263 2924 31272
rect 2872 31229 2881 31263
rect 2881 31229 2915 31263
rect 2915 31229 2924 31263
rect 2872 31220 2924 31229
rect 4436 31263 4488 31272
rect 4436 31229 4445 31263
rect 4445 31229 4479 31263
rect 4479 31229 4488 31263
rect 4436 31220 4488 31229
rect 5264 31288 5316 31340
rect 5724 31288 5776 31340
rect 5908 31288 5960 31340
rect 6460 31288 6512 31340
rect 7012 31288 7064 31340
rect 7196 31288 7248 31340
rect 8484 31331 8536 31340
rect 8484 31297 8493 31331
rect 8493 31297 8527 31331
rect 8527 31297 8536 31331
rect 8484 31288 8536 31297
rect 10048 31331 10100 31340
rect 6828 31220 6880 31272
rect 7932 31263 7984 31272
rect 7932 31229 7941 31263
rect 7941 31229 7975 31263
rect 7975 31229 7984 31263
rect 7932 31220 7984 31229
rect 8208 31263 8260 31272
rect 8208 31229 8217 31263
rect 8217 31229 8251 31263
rect 8251 31229 8260 31263
rect 8208 31220 8260 31229
rect 1492 31084 1544 31136
rect 3884 31127 3936 31136
rect 3884 31093 3893 31127
rect 3893 31093 3927 31127
rect 3927 31093 3936 31127
rect 3884 31084 3936 31093
rect 4068 31084 4120 31136
rect 5908 31127 5960 31136
rect 5908 31093 5917 31127
rect 5917 31093 5951 31127
rect 5951 31093 5960 31127
rect 5908 31084 5960 31093
rect 6092 31084 6144 31136
rect 7564 31152 7616 31204
rect 8024 31084 8076 31136
rect 8484 31084 8536 31136
rect 9680 31220 9732 31272
rect 10048 31297 10055 31331
rect 10055 31297 10089 31331
rect 10089 31297 10100 31331
rect 10048 31288 10100 31297
rect 11244 31288 11296 31340
rect 16120 31424 16172 31476
rect 17224 31424 17276 31476
rect 18328 31424 18380 31476
rect 10876 31220 10928 31272
rect 11888 31084 11940 31136
rect 13084 31331 13136 31340
rect 13084 31297 13093 31331
rect 13093 31297 13127 31331
rect 13127 31297 13136 31331
rect 13084 31288 13136 31297
rect 13544 31288 13596 31340
rect 12256 31220 12308 31272
rect 15292 31356 15344 31408
rect 18604 31356 18656 31408
rect 19708 31424 19760 31476
rect 20444 31424 20496 31476
rect 21180 31424 21232 31476
rect 15200 31220 15252 31272
rect 16304 31288 16356 31340
rect 17224 31288 17276 31340
rect 17960 31288 18012 31340
rect 18880 31288 18932 31340
rect 19708 31288 19760 31340
rect 18972 31220 19024 31272
rect 20628 31288 20680 31340
rect 12992 31127 13044 31136
rect 12992 31093 13001 31127
rect 13001 31093 13035 31127
rect 13035 31093 13044 31127
rect 12992 31084 13044 31093
rect 14740 31084 14792 31136
rect 18144 31152 18196 31204
rect 21272 31331 21324 31340
rect 21272 31297 21281 31331
rect 21281 31297 21315 31331
rect 21315 31297 21324 31331
rect 21272 31288 21324 31297
rect 15476 31127 15528 31136
rect 15476 31093 15485 31127
rect 15485 31093 15519 31127
rect 15519 31093 15528 31127
rect 15476 31084 15528 31093
rect 21088 31084 21140 31136
rect 21456 31127 21508 31136
rect 21456 31093 21465 31127
rect 21465 31093 21499 31127
rect 21499 31093 21508 31127
rect 21456 31084 21508 31093
rect 3549 30982 3601 31034
rect 3613 30982 3665 31034
rect 3677 30982 3729 31034
rect 3741 30982 3793 31034
rect 3805 30982 3857 31034
rect 8747 30982 8799 31034
rect 8811 30982 8863 31034
rect 8875 30982 8927 31034
rect 8939 30982 8991 31034
rect 9003 30982 9055 31034
rect 13945 30982 13997 31034
rect 14009 30982 14061 31034
rect 14073 30982 14125 31034
rect 14137 30982 14189 31034
rect 14201 30982 14253 31034
rect 19143 30982 19195 31034
rect 19207 30982 19259 31034
rect 19271 30982 19323 31034
rect 19335 30982 19387 31034
rect 19399 30982 19451 31034
rect 1492 30880 1544 30932
rect 2412 30880 2464 30932
rect 5356 30880 5408 30932
rect 8208 30880 8260 30932
rect 10048 30880 10100 30932
rect 11060 30880 11112 30932
rect 2964 30812 3016 30864
rect 3424 30812 3476 30864
rect 3884 30812 3936 30864
rect 12256 30812 12308 30864
rect 3240 30744 3292 30796
rect 4160 30744 4212 30796
rect 5356 30744 5408 30796
rect 5908 30744 5960 30796
rect 8024 30744 8076 30796
rect 9404 30744 9456 30796
rect 1124 30676 1176 30728
rect 2136 30676 2188 30728
rect 2780 30719 2832 30728
rect 2780 30685 2789 30719
rect 2789 30685 2823 30719
rect 2823 30685 2832 30719
rect 2780 30676 2832 30685
rect 2872 30676 2924 30728
rect 3424 30676 3476 30728
rect 3792 30719 3844 30728
rect 3792 30685 3801 30719
rect 3801 30685 3835 30719
rect 3835 30685 3844 30719
rect 3792 30676 3844 30685
rect 4712 30719 4764 30728
rect 4712 30685 4721 30719
rect 4721 30685 4755 30719
rect 4755 30685 4764 30719
rect 4712 30676 4764 30685
rect 4988 30719 5040 30728
rect 4988 30685 4997 30719
rect 4997 30685 5031 30719
rect 5031 30685 5040 30719
rect 4988 30676 5040 30685
rect 6644 30676 6696 30728
rect 2320 30540 2372 30592
rect 2688 30540 2740 30592
rect 2872 30540 2924 30592
rect 4252 30540 4304 30592
rect 4896 30540 4948 30592
rect 5264 30540 5316 30592
rect 6368 30651 6420 30660
rect 6368 30617 6377 30651
rect 6377 30617 6411 30651
rect 6411 30617 6420 30651
rect 6368 30608 6420 30617
rect 7380 30676 7432 30728
rect 11888 30744 11940 30796
rect 12992 30880 13044 30932
rect 13084 30880 13136 30932
rect 13268 30880 13320 30932
rect 15108 30880 15160 30932
rect 16028 30880 16080 30932
rect 18328 30880 18380 30932
rect 18512 30880 18564 30932
rect 13452 30744 13504 30796
rect 6828 30651 6880 30660
rect 6828 30617 6837 30651
rect 6837 30617 6871 30651
rect 6871 30617 6880 30651
rect 6828 30608 6880 30617
rect 12624 30719 12676 30728
rect 12624 30685 12633 30719
rect 12633 30685 12667 30719
rect 12667 30685 12676 30719
rect 12624 30676 12676 30685
rect 12900 30719 12952 30728
rect 12900 30685 12909 30719
rect 12909 30685 12943 30719
rect 12943 30685 12952 30719
rect 12900 30676 12952 30685
rect 15292 30676 15344 30728
rect 16304 30676 16356 30728
rect 7196 30583 7248 30592
rect 7196 30549 7205 30583
rect 7205 30549 7239 30583
rect 7239 30549 7248 30583
rect 7196 30540 7248 30549
rect 7932 30540 7984 30592
rect 14188 30608 14240 30660
rect 16212 30608 16264 30660
rect 17224 30608 17276 30660
rect 18144 30719 18196 30728
rect 18144 30685 18153 30719
rect 18153 30685 18187 30719
rect 18187 30685 18196 30719
rect 18144 30676 18196 30685
rect 20812 30880 20864 30932
rect 21364 30812 21416 30864
rect 22284 30744 22336 30796
rect 22560 30744 22612 30796
rect 13544 30540 13596 30592
rect 14464 30540 14516 30592
rect 16028 30540 16080 30592
rect 18880 30676 18932 30728
rect 19156 30676 19208 30728
rect 19800 30676 19852 30728
rect 20904 30676 20956 30728
rect 21180 30719 21232 30728
rect 21180 30685 21189 30719
rect 21189 30685 21223 30719
rect 21223 30685 21232 30719
rect 21180 30676 21232 30685
rect 18788 30608 18840 30660
rect 19064 30608 19116 30660
rect 19708 30608 19760 30660
rect 22284 30608 22336 30660
rect 20812 30583 20864 30592
rect 20812 30549 20821 30583
rect 20821 30549 20855 30583
rect 20855 30549 20864 30583
rect 20812 30540 20864 30549
rect 6148 30438 6200 30490
rect 6212 30438 6264 30490
rect 6276 30438 6328 30490
rect 6340 30438 6392 30490
rect 6404 30438 6456 30490
rect 11346 30438 11398 30490
rect 11410 30438 11462 30490
rect 11474 30438 11526 30490
rect 11538 30438 11590 30490
rect 11602 30438 11654 30490
rect 16544 30438 16596 30490
rect 16608 30438 16660 30490
rect 16672 30438 16724 30490
rect 16736 30438 16788 30490
rect 16800 30438 16852 30490
rect 21742 30438 21794 30490
rect 21806 30438 21858 30490
rect 21870 30438 21922 30490
rect 21934 30438 21986 30490
rect 21998 30438 22050 30490
rect 1768 30336 1820 30388
rect 3976 30336 4028 30388
rect 4988 30336 5040 30388
rect 5908 30336 5960 30388
rect 6092 30336 6144 30388
rect 7196 30336 7248 30388
rect 7380 30379 7432 30388
rect 7380 30345 7389 30379
rect 7389 30345 7423 30379
rect 7423 30345 7432 30379
rect 7380 30336 7432 30345
rect 7656 30336 7708 30388
rect 10048 30336 10100 30388
rect 12624 30336 12676 30388
rect 13820 30336 13872 30388
rect 14648 30336 14700 30388
rect 1952 30273 2004 30320
rect 1400 30243 1452 30252
rect 1400 30209 1409 30243
rect 1409 30209 1443 30243
rect 1443 30209 1452 30243
rect 1400 30200 1452 30209
rect 1492 30200 1544 30252
rect 1952 30268 1977 30273
rect 1977 30268 2004 30273
rect 2412 30268 2464 30320
rect 3884 30268 3936 30320
rect 3240 30200 3292 30252
rect 3608 30243 3660 30252
rect 3608 30209 3615 30243
rect 3615 30209 3649 30243
rect 3649 30209 3660 30243
rect 3608 30200 3660 30209
rect 4160 30200 4212 30252
rect 5816 30268 5868 30320
rect 5172 30243 5224 30252
rect 5172 30209 5179 30243
rect 5179 30209 5213 30243
rect 5213 30209 5224 30243
rect 5172 30200 5224 30209
rect 9036 30268 9088 30320
rect 10692 30268 10744 30320
rect 7104 30200 7156 30252
rect 9220 30200 9272 30252
rect 11612 30200 11664 30252
rect 12440 30243 12492 30252
rect 12440 30209 12449 30243
rect 12449 30209 12483 30243
rect 12483 30209 12492 30243
rect 12440 30200 12492 30209
rect 13452 30243 13504 30252
rect 13452 30209 13461 30243
rect 13461 30209 13495 30243
rect 13495 30209 13504 30243
rect 13452 30200 13504 30209
rect 13636 30200 13688 30252
rect 15844 30336 15896 30388
rect 15200 30268 15252 30320
rect 16028 30268 16080 30320
rect 17592 30336 17644 30388
rect 18788 30336 18840 30388
rect 18972 30336 19024 30388
rect 20444 30336 20496 30388
rect 22652 30336 22704 30388
rect 2872 30132 2924 30184
rect 4896 30175 4948 30184
rect 4896 30141 4905 30175
rect 4905 30141 4939 30175
rect 4939 30141 4948 30175
rect 4896 30132 4948 30141
rect 6368 30175 6420 30184
rect 6368 30141 6377 30175
rect 6377 30141 6411 30175
rect 6411 30141 6420 30175
rect 6368 30132 6420 30141
rect 11244 30132 11296 30184
rect 11704 30175 11756 30184
rect 11704 30141 11713 30175
rect 11713 30141 11747 30175
rect 11747 30141 11756 30175
rect 11704 30132 11756 30141
rect 11888 30132 11940 30184
rect 2688 30039 2740 30048
rect 2688 30005 2697 30039
rect 2697 30005 2731 30039
rect 2731 30005 2740 30039
rect 2688 29996 2740 30005
rect 3056 29996 3108 30048
rect 3332 29996 3384 30048
rect 5908 30039 5960 30048
rect 5908 30005 5917 30039
rect 5917 30005 5951 30039
rect 5951 30005 5960 30039
rect 5908 29996 5960 30005
rect 9404 30064 9456 30116
rect 7840 29996 7892 30048
rect 8576 29996 8628 30048
rect 11612 30064 11664 30116
rect 12716 30175 12768 30184
rect 12716 30141 12725 30175
rect 12725 30141 12759 30175
rect 12759 30141 12768 30175
rect 12716 30132 12768 30141
rect 13084 30132 13136 30184
rect 14740 30132 14792 30184
rect 16856 30200 16908 30252
rect 17500 30200 17552 30252
rect 19524 30243 19576 30252
rect 19524 30209 19533 30243
rect 19533 30209 19567 30243
rect 19567 30209 19576 30243
rect 19524 30200 19576 30209
rect 19800 30243 19852 30252
rect 19800 30209 19807 30243
rect 19807 30209 19841 30243
rect 19841 30209 19852 30243
rect 19800 30200 19852 30209
rect 20996 30268 21048 30320
rect 21640 30200 21692 30252
rect 13360 29996 13412 30048
rect 13820 29996 13872 30048
rect 15844 30039 15896 30048
rect 15844 30005 15853 30039
rect 15853 30005 15887 30039
rect 15887 30005 15896 30039
rect 15844 29996 15896 30005
rect 16396 30039 16448 30048
rect 16396 30005 16405 30039
rect 16405 30005 16439 30039
rect 16439 30005 16448 30039
rect 16396 29996 16448 30005
rect 16764 29996 16816 30048
rect 19064 30039 19116 30048
rect 19064 30005 19073 30039
rect 19073 30005 19107 30039
rect 19107 30005 19116 30039
rect 19064 29996 19116 30005
rect 20996 29996 21048 30048
rect 21456 30039 21508 30048
rect 21456 30005 21465 30039
rect 21465 30005 21499 30039
rect 21499 30005 21508 30039
rect 21456 29996 21508 30005
rect 3549 29894 3601 29946
rect 3613 29894 3665 29946
rect 3677 29894 3729 29946
rect 3741 29894 3793 29946
rect 3805 29894 3857 29946
rect 8747 29894 8799 29946
rect 8811 29894 8863 29946
rect 8875 29894 8927 29946
rect 8939 29894 8991 29946
rect 9003 29894 9055 29946
rect 13945 29894 13997 29946
rect 14009 29894 14061 29946
rect 14073 29894 14125 29946
rect 14137 29894 14189 29946
rect 14201 29894 14253 29946
rect 19143 29894 19195 29946
rect 19207 29894 19259 29946
rect 19271 29894 19323 29946
rect 19335 29894 19387 29946
rect 19399 29894 19451 29946
rect 4160 29792 4212 29844
rect 5172 29792 5224 29844
rect 7840 29792 7892 29844
rect 9220 29792 9272 29844
rect 4620 29724 4672 29776
rect 6736 29724 6788 29776
rect 7472 29724 7524 29776
rect 10968 29792 11020 29844
rect 12256 29792 12308 29844
rect 2320 29656 2372 29708
rect 756 29588 808 29640
rect 2688 29588 2740 29640
rect 2964 29588 3016 29640
rect 1676 29563 1728 29572
rect 1676 29529 1685 29563
rect 1685 29529 1719 29563
rect 1719 29529 1728 29563
rect 1676 29520 1728 29529
rect 1860 29520 1912 29572
rect 2504 29520 2556 29572
rect 3516 29588 3568 29640
rect 5908 29656 5960 29708
rect 7104 29656 7156 29708
rect 11612 29724 11664 29776
rect 12900 29792 12952 29844
rect 15844 29792 15896 29844
rect 16396 29792 16448 29844
rect 18328 29792 18380 29844
rect 18512 29792 18564 29844
rect 19064 29792 19116 29844
rect 20628 29792 20680 29844
rect 20720 29792 20772 29844
rect 7380 29588 7432 29640
rect 7840 29588 7892 29640
rect 9036 29656 9088 29708
rect 9496 29656 9548 29708
rect 10600 29656 10652 29708
rect 8300 29588 8352 29640
rect 9220 29588 9272 29640
rect 1768 29452 1820 29504
rect 3240 29452 3292 29504
rect 4160 29520 4212 29572
rect 5448 29520 5500 29572
rect 5632 29563 5684 29572
rect 5632 29529 5641 29563
rect 5641 29529 5675 29563
rect 5675 29529 5684 29563
rect 5632 29520 5684 29529
rect 5724 29563 5776 29572
rect 5724 29529 5733 29563
rect 5733 29529 5767 29563
rect 5767 29529 5776 29563
rect 5724 29520 5776 29529
rect 6000 29520 6052 29572
rect 6552 29520 6604 29572
rect 6828 29520 6880 29572
rect 7196 29520 7248 29572
rect 7564 29520 7616 29572
rect 10140 29588 10192 29640
rect 10876 29588 10928 29640
rect 11336 29699 11388 29708
rect 11336 29665 11345 29699
rect 11345 29665 11379 29699
rect 11379 29665 11388 29699
rect 11336 29656 11388 29665
rect 12164 29656 12216 29708
rect 12716 29656 12768 29708
rect 12900 29656 12952 29708
rect 13912 29656 13964 29708
rect 14188 29656 14240 29708
rect 5908 29452 5960 29504
rect 6460 29495 6512 29504
rect 6460 29461 6469 29495
rect 6469 29461 6503 29495
rect 6503 29461 6512 29495
rect 6460 29452 6512 29461
rect 6644 29495 6696 29504
rect 6644 29461 6653 29495
rect 6653 29461 6687 29495
rect 6687 29461 6696 29495
rect 6644 29452 6696 29461
rect 7380 29452 7432 29504
rect 8116 29452 8168 29504
rect 10048 29452 10100 29504
rect 13268 29588 13320 29640
rect 15476 29656 15528 29708
rect 15108 29631 15160 29640
rect 15108 29597 15142 29631
rect 15142 29597 15160 29631
rect 15108 29588 15160 29597
rect 14004 29452 14056 29504
rect 14188 29452 14240 29504
rect 15016 29452 15068 29504
rect 16212 29631 16264 29640
rect 16212 29597 16221 29631
rect 16221 29597 16255 29631
rect 16255 29597 16264 29631
rect 16212 29588 16264 29597
rect 18052 29656 18104 29708
rect 18328 29656 18380 29708
rect 20904 29724 20956 29776
rect 16764 29588 16816 29640
rect 18144 29631 18196 29640
rect 18144 29597 18153 29631
rect 18153 29597 18187 29631
rect 18187 29597 18196 29631
rect 18144 29588 18196 29597
rect 19984 29631 20036 29640
rect 19984 29597 19993 29631
rect 19993 29597 20027 29631
rect 20027 29597 20036 29631
rect 19984 29588 20036 29597
rect 17040 29452 17092 29504
rect 19708 29520 19760 29572
rect 20536 29631 20588 29640
rect 20536 29597 20545 29631
rect 20545 29597 20579 29631
rect 20579 29597 20588 29631
rect 20536 29588 20588 29597
rect 17224 29495 17276 29504
rect 17224 29461 17233 29495
rect 17233 29461 17267 29495
rect 17267 29461 17276 29495
rect 17224 29452 17276 29461
rect 17960 29495 18012 29504
rect 17960 29461 17969 29495
rect 17969 29461 18003 29495
rect 18003 29461 18012 29495
rect 17960 29452 18012 29461
rect 20444 29520 20496 29572
rect 20996 29588 21048 29640
rect 21088 29588 21140 29640
rect 20996 29452 21048 29504
rect 21180 29495 21232 29504
rect 21180 29461 21189 29495
rect 21189 29461 21223 29495
rect 21223 29461 21232 29495
rect 21180 29452 21232 29461
rect 22192 29452 22244 29504
rect 6148 29350 6200 29402
rect 6212 29350 6264 29402
rect 6276 29350 6328 29402
rect 6340 29350 6392 29402
rect 6404 29350 6456 29402
rect 11346 29350 11398 29402
rect 11410 29350 11462 29402
rect 11474 29350 11526 29402
rect 11538 29350 11590 29402
rect 11602 29350 11654 29402
rect 16544 29350 16596 29402
rect 16608 29350 16660 29402
rect 16672 29350 16724 29402
rect 16736 29350 16788 29402
rect 16800 29350 16852 29402
rect 21742 29350 21794 29402
rect 21806 29350 21858 29402
rect 21870 29350 21922 29402
rect 21934 29350 21986 29402
rect 21998 29350 22050 29402
rect 20 29248 72 29300
rect 2596 29248 2648 29300
rect 3148 29291 3200 29300
rect 3148 29257 3157 29291
rect 3157 29257 3191 29291
rect 3191 29257 3200 29291
rect 3148 29248 3200 29257
rect 5724 29248 5776 29300
rect 2044 29180 2096 29232
rect 2412 29180 2464 29232
rect 2872 29180 2924 29232
rect 1308 29044 1360 29096
rect 2964 29155 3016 29164
rect 2964 29121 2973 29155
rect 2973 29121 3007 29155
rect 3007 29121 3016 29155
rect 2964 29112 3016 29121
rect 9220 29223 9272 29232
rect 9220 29189 9229 29223
rect 9229 29189 9263 29223
rect 9263 29189 9272 29223
rect 9220 29180 9272 29189
rect 9429 29223 9481 29232
rect 9429 29189 9459 29223
rect 9459 29189 9481 29223
rect 9429 29180 9481 29189
rect 4620 29112 4672 29164
rect 4896 29155 4948 29164
rect 4896 29121 4905 29155
rect 4905 29121 4939 29155
rect 4939 29121 4948 29155
rect 4896 29112 4948 29121
rect 5172 29155 5224 29164
rect 5172 29121 5179 29155
rect 5179 29121 5213 29155
rect 5213 29121 5224 29155
rect 5172 29112 5224 29121
rect 7380 29155 7432 29164
rect 7380 29121 7389 29155
rect 7389 29121 7423 29155
rect 7423 29121 7432 29155
rect 7380 29112 7432 29121
rect 8484 29112 8536 29164
rect 8576 29155 8628 29164
rect 8576 29121 8585 29155
rect 8585 29121 8619 29155
rect 8619 29121 8628 29155
rect 8576 29112 8628 29121
rect 2320 28976 2372 29028
rect 3148 28976 3200 29028
rect 4068 28976 4120 29028
rect 8116 29044 8168 29096
rect 10140 29112 10192 29164
rect 10232 29155 10284 29164
rect 10232 29121 10241 29155
rect 10241 29121 10275 29155
rect 10275 29121 10284 29155
rect 10232 29112 10284 29121
rect 10968 29180 11020 29232
rect 10876 29112 10928 29164
rect 11888 29248 11940 29300
rect 12348 29248 12400 29300
rect 12716 29248 12768 29300
rect 13268 29248 13320 29300
rect 14280 29248 14332 29300
rect 14740 29248 14792 29300
rect 16212 29248 16264 29300
rect 17040 29248 17092 29300
rect 18144 29248 18196 29300
rect 18512 29248 18564 29300
rect 9404 29044 9456 29096
rect 10600 29044 10652 29096
rect 7840 28976 7892 29028
rect 9036 28976 9088 29028
rect 9220 28976 9272 29028
rect 10784 29019 10836 29028
rect 10784 28985 10793 29019
rect 10793 28985 10827 29019
rect 10827 28985 10836 29019
rect 10784 28976 10836 28985
rect 12256 29044 12308 29096
rect 13268 29087 13320 29096
rect 13268 29053 13277 29087
rect 13277 29053 13311 29087
rect 13311 29053 13320 29087
rect 13268 29044 13320 29053
rect 14280 29155 14332 29164
rect 14280 29121 14314 29155
rect 14314 29121 14332 29155
rect 14280 29112 14332 29121
rect 14464 29155 14516 29164
rect 14464 29121 14473 29155
rect 14473 29121 14507 29155
rect 14507 29121 14516 29155
rect 14464 29112 14516 29121
rect 16028 29180 16080 29232
rect 15936 29112 15988 29164
rect 16304 29112 16356 29164
rect 16672 29155 16724 29164
rect 16672 29121 16681 29155
rect 16681 29121 16715 29155
rect 16715 29121 16724 29155
rect 16672 29112 16724 29121
rect 18972 29180 19024 29232
rect 17500 29112 17552 29164
rect 18052 29112 18104 29164
rect 18512 29112 18564 29164
rect 20444 29291 20496 29300
rect 20444 29257 20453 29291
rect 20453 29257 20487 29291
rect 20487 29257 20496 29291
rect 20444 29248 20496 29257
rect 20536 29248 20588 29300
rect 19984 29112 20036 29164
rect 20168 29155 20220 29164
rect 20168 29121 20177 29155
rect 20177 29121 20211 29155
rect 20211 29121 20220 29155
rect 20168 29112 20220 29121
rect 20812 29180 20864 29232
rect 21272 29112 21324 29164
rect 13912 29087 13964 29096
rect 13912 29053 13921 29087
rect 13921 29053 13955 29087
rect 13955 29053 13964 29087
rect 13912 29044 13964 29053
rect 14004 29044 14056 29096
rect 1860 28908 1912 28960
rect 2412 28908 2464 28960
rect 2688 28908 2740 28960
rect 3332 28908 3384 28960
rect 8484 28908 8536 28960
rect 10692 28908 10744 28960
rect 11520 28908 11572 28960
rect 12440 28908 12492 28960
rect 13452 28908 13504 28960
rect 16212 28951 16264 28960
rect 16212 28917 16221 28951
rect 16221 28917 16255 28951
rect 16255 28917 16264 28951
rect 16212 28908 16264 28917
rect 19524 29044 19576 29096
rect 19708 29044 19760 29096
rect 22192 29044 22244 29096
rect 19524 28908 19576 28960
rect 21456 28951 21508 28960
rect 21456 28917 21465 28951
rect 21465 28917 21499 28951
rect 21499 28917 21508 28951
rect 21456 28908 21508 28917
rect 3549 28806 3601 28858
rect 3613 28806 3665 28858
rect 3677 28806 3729 28858
rect 3741 28806 3793 28858
rect 3805 28806 3857 28858
rect 8747 28806 8799 28858
rect 8811 28806 8863 28858
rect 8875 28806 8927 28858
rect 8939 28806 8991 28858
rect 9003 28806 9055 28858
rect 13945 28806 13997 28858
rect 14009 28806 14061 28858
rect 14073 28806 14125 28858
rect 14137 28806 14189 28858
rect 14201 28806 14253 28858
rect 19143 28806 19195 28858
rect 19207 28806 19259 28858
rect 19271 28806 19323 28858
rect 19335 28806 19387 28858
rect 19399 28806 19451 28858
rect 3332 28704 3384 28756
rect 3792 28704 3844 28756
rect 1860 28636 1912 28688
rect 756 28500 808 28552
rect 1584 28500 1636 28552
rect 1768 28543 1820 28552
rect 1768 28509 1777 28543
rect 1777 28509 1811 28543
rect 1811 28509 1820 28543
rect 1768 28500 1820 28509
rect 3148 28568 3200 28620
rect 2504 28543 2556 28552
rect 2504 28509 2513 28543
rect 2513 28509 2556 28543
rect 2504 28500 2556 28509
rect 2872 28500 2924 28552
rect 5172 28636 5224 28688
rect 5172 28500 5224 28552
rect 7840 28636 7892 28688
rect 8116 28679 8168 28688
rect 8116 28645 8125 28679
rect 8125 28645 8159 28679
rect 8159 28645 8168 28679
rect 8116 28636 8168 28645
rect 10416 28704 10468 28756
rect 15200 28704 15252 28756
rect 15292 28704 15344 28756
rect 12164 28636 12216 28688
rect 12532 28636 12584 28688
rect 14372 28636 14424 28688
rect 5540 28611 5592 28620
rect 5540 28577 5549 28611
rect 5549 28577 5583 28611
rect 5583 28577 5592 28611
rect 5540 28568 5592 28577
rect 9036 28568 9088 28620
rect 7104 28543 7156 28552
rect 7104 28509 7113 28543
rect 7113 28509 7147 28543
rect 7147 28509 7156 28543
rect 7104 28500 7156 28509
rect 7288 28500 7340 28552
rect 7840 28500 7892 28552
rect 8852 28500 8904 28552
rect 13452 28568 13504 28620
rect 14740 28611 14792 28620
rect 14740 28577 14749 28611
rect 14749 28577 14783 28611
rect 14783 28577 14792 28611
rect 14740 28568 14792 28577
rect 16948 28636 17000 28688
rect 18052 28704 18104 28756
rect 15844 28568 15896 28620
rect 19800 28636 19852 28688
rect 20168 28636 20220 28688
rect 1860 28432 1912 28484
rect 1584 28364 1636 28416
rect 9312 28432 9364 28484
rect 11060 28500 11112 28552
rect 11612 28500 11664 28552
rect 14004 28500 14056 28552
rect 10140 28432 10192 28484
rect 13268 28432 13320 28484
rect 15016 28543 15068 28552
rect 15016 28509 15025 28543
rect 15025 28509 15059 28543
rect 15059 28509 15068 28543
rect 15016 28500 15068 28509
rect 15292 28543 15344 28552
rect 15292 28509 15301 28543
rect 15301 28509 15335 28543
rect 15335 28509 15344 28543
rect 15292 28500 15344 28509
rect 16028 28543 16080 28552
rect 16028 28509 16037 28543
rect 16037 28509 16071 28543
rect 16071 28509 16080 28543
rect 16028 28500 16080 28509
rect 16212 28500 16264 28552
rect 17224 28500 17276 28552
rect 2504 28364 2556 28416
rect 3700 28364 3752 28416
rect 3976 28364 4028 28416
rect 4252 28364 4304 28416
rect 4620 28364 4672 28416
rect 4896 28407 4948 28416
rect 4896 28373 4905 28407
rect 4905 28373 4939 28407
rect 4939 28373 4948 28407
rect 4896 28364 4948 28373
rect 5540 28364 5592 28416
rect 8484 28364 8536 28416
rect 8668 28364 8720 28416
rect 10416 28364 10468 28416
rect 11244 28364 11296 28416
rect 12256 28364 12308 28416
rect 12624 28364 12676 28416
rect 15844 28364 15896 28416
rect 19340 28543 19392 28552
rect 19340 28509 19349 28543
rect 19349 28509 19383 28543
rect 19383 28509 19392 28543
rect 19340 28500 19392 28509
rect 20536 28568 20588 28620
rect 19432 28432 19484 28484
rect 17500 28407 17552 28416
rect 17500 28373 17509 28407
rect 17509 28373 17543 28407
rect 17543 28373 17552 28407
rect 17500 28364 17552 28373
rect 19524 28407 19576 28416
rect 19524 28373 19533 28407
rect 19533 28373 19567 28407
rect 19567 28373 19576 28407
rect 19524 28364 19576 28373
rect 19616 28407 19668 28416
rect 19616 28373 19625 28407
rect 19625 28373 19659 28407
rect 19659 28373 19668 28407
rect 19616 28364 19668 28373
rect 20628 28543 20680 28552
rect 20628 28509 20637 28543
rect 20637 28509 20671 28543
rect 20671 28509 20680 28543
rect 20628 28500 20680 28509
rect 20996 28500 21048 28552
rect 20720 28407 20772 28416
rect 20720 28373 20729 28407
rect 20729 28373 20763 28407
rect 20763 28373 20772 28407
rect 20720 28364 20772 28373
rect 20996 28407 21048 28416
rect 20996 28373 21005 28407
rect 21005 28373 21039 28407
rect 21039 28373 21048 28407
rect 20996 28364 21048 28373
rect 22192 28364 22244 28416
rect 6148 28262 6200 28314
rect 6212 28262 6264 28314
rect 6276 28262 6328 28314
rect 6340 28262 6392 28314
rect 6404 28262 6456 28314
rect 11346 28262 11398 28314
rect 11410 28262 11462 28314
rect 11474 28262 11526 28314
rect 11538 28262 11590 28314
rect 11602 28262 11654 28314
rect 16544 28262 16596 28314
rect 16608 28262 16660 28314
rect 16672 28262 16724 28314
rect 16736 28262 16788 28314
rect 16800 28262 16852 28314
rect 21742 28262 21794 28314
rect 21806 28262 21858 28314
rect 21870 28262 21922 28314
rect 21934 28262 21986 28314
rect 21998 28262 22050 28314
rect 3332 28160 3384 28212
rect 5172 28160 5224 28212
rect 8944 28160 8996 28212
rect 9036 28160 9088 28212
rect 2504 28092 2556 28144
rect 756 28024 808 28076
rect 1676 28024 1728 28076
rect 1952 28067 2004 28076
rect 1952 28033 1961 28067
rect 1961 28033 1995 28067
rect 1995 28033 2004 28067
rect 1952 28024 2004 28033
rect 2872 28024 2924 28076
rect 3884 28092 3936 28144
rect 3608 28024 3660 28076
rect 3700 28024 3752 28076
rect 4896 28092 4948 28144
rect 7656 28092 7708 28144
rect 4068 28024 4120 28076
rect 4528 28024 4580 28076
rect 4804 28024 4856 28076
rect 5172 28024 5224 28076
rect 8576 28092 8628 28144
rect 8852 28024 8904 28076
rect 9588 28160 9640 28212
rect 10324 28160 10376 28212
rect 10968 28160 11020 28212
rect 9496 28092 9548 28144
rect 13912 28160 13964 28212
rect 15660 28160 15712 28212
rect 15844 28092 15896 28144
rect 15936 28092 15988 28144
rect 10140 28024 10192 28076
rect 13912 28024 13964 28076
rect 14188 28024 14240 28076
rect 14648 28024 14700 28076
rect 17040 28203 17092 28212
rect 17040 28169 17049 28203
rect 17049 28169 17083 28203
rect 17083 28169 17092 28203
rect 17040 28160 17092 28169
rect 17500 28160 17552 28212
rect 17960 28160 18012 28212
rect 19340 28160 19392 28212
rect 19616 28160 19668 28212
rect 20536 28160 20588 28212
rect 20628 28160 20680 28212
rect 20720 28160 20772 28212
rect 2688 27956 2740 28008
rect 1676 27931 1728 27940
rect 1676 27897 1685 27931
rect 1685 27897 1719 27931
rect 1719 27897 1728 27931
rect 1676 27888 1728 27897
rect 7288 27956 7340 28008
rect 8668 27956 8720 28008
rect 9772 27956 9824 28008
rect 11060 27956 11112 28008
rect 8484 27888 8536 27940
rect 2320 27820 2372 27872
rect 3884 27820 3936 27872
rect 5264 27820 5316 27872
rect 6000 27820 6052 27872
rect 7748 27820 7800 27872
rect 11244 27820 11296 27872
rect 11888 27820 11940 27872
rect 16212 27956 16264 28008
rect 17040 27956 17092 28008
rect 15200 27888 15252 27940
rect 19616 28067 19668 28076
rect 19616 28033 19625 28067
rect 19625 28033 19659 28067
rect 19659 28033 19668 28067
rect 19616 28024 19668 28033
rect 20168 28067 20220 28076
rect 20168 28033 20177 28067
rect 20177 28033 20211 28067
rect 20211 28033 20220 28067
rect 20168 28024 20220 28033
rect 14372 27820 14424 27872
rect 15292 27820 15344 27872
rect 16396 27820 16448 27872
rect 19064 27888 19116 27940
rect 20812 28067 20864 28076
rect 20812 28033 20821 28067
rect 20821 28033 20855 28067
rect 20855 28033 20864 28067
rect 20812 28024 20864 28033
rect 21272 28067 21324 28076
rect 21272 28033 21281 28067
rect 21281 28033 21315 28067
rect 21315 28033 21324 28067
rect 21272 28024 21324 28033
rect 19616 27820 19668 27872
rect 19800 27820 19852 27872
rect 20904 27820 20956 27872
rect 21088 27863 21140 27872
rect 21088 27829 21097 27863
rect 21097 27829 21131 27863
rect 21131 27829 21140 27863
rect 21088 27820 21140 27829
rect 21456 27863 21508 27872
rect 21456 27829 21465 27863
rect 21465 27829 21499 27863
rect 21499 27829 21508 27863
rect 21456 27820 21508 27829
rect 756 27684 808 27736
rect 3549 27718 3601 27770
rect 3613 27718 3665 27770
rect 3677 27718 3729 27770
rect 3741 27718 3793 27770
rect 3805 27718 3857 27770
rect 8747 27718 8799 27770
rect 8811 27718 8863 27770
rect 8875 27718 8927 27770
rect 8939 27718 8991 27770
rect 9003 27718 9055 27770
rect 13945 27718 13997 27770
rect 14009 27718 14061 27770
rect 14073 27718 14125 27770
rect 14137 27718 14189 27770
rect 14201 27718 14253 27770
rect 19143 27718 19195 27770
rect 19207 27718 19259 27770
rect 19271 27718 19323 27770
rect 19335 27718 19387 27770
rect 19399 27718 19451 27770
rect 1676 27616 1728 27668
rect 2872 27616 2924 27668
rect 3148 27548 3200 27600
rect 4252 27548 4304 27600
rect 9128 27616 9180 27668
rect 9496 27616 9548 27668
rect 5172 27548 5224 27600
rect 1584 27455 1636 27464
rect 1584 27421 1593 27455
rect 1593 27421 1627 27455
rect 1627 27421 1636 27455
rect 1584 27412 1636 27421
rect 1860 27455 1912 27464
rect 1860 27421 1867 27455
rect 1867 27421 1901 27455
rect 1901 27421 1912 27455
rect 1860 27412 1912 27421
rect 1308 27344 1360 27396
rect 2412 27412 2464 27464
rect 8116 27480 8168 27532
rect 2504 27344 2556 27396
rect 4160 27412 4212 27464
rect 3700 27344 3752 27396
rect 4068 27344 4120 27396
rect 5540 27412 5592 27464
rect 6000 27412 6052 27464
rect 4896 27344 4948 27396
rect 7288 27412 7340 27464
rect 7472 27412 7524 27464
rect 2596 27319 2648 27328
rect 2596 27285 2605 27319
rect 2605 27285 2639 27319
rect 2639 27285 2648 27319
rect 2596 27276 2648 27285
rect 3148 27319 3200 27328
rect 3148 27285 3157 27319
rect 3157 27285 3191 27319
rect 3191 27285 3200 27319
rect 3148 27276 3200 27285
rect 3332 27276 3384 27328
rect 4804 27276 4856 27328
rect 6000 27276 6052 27328
rect 7564 27344 7616 27396
rect 7656 27387 7708 27396
rect 7656 27353 7665 27387
rect 7665 27353 7699 27387
rect 7699 27353 7708 27387
rect 7656 27344 7708 27353
rect 7748 27387 7800 27396
rect 7748 27353 7757 27387
rect 7757 27353 7791 27387
rect 7791 27353 7800 27387
rect 7748 27344 7800 27353
rect 8024 27412 8076 27464
rect 9772 27480 9824 27532
rect 14372 27616 14424 27668
rect 14556 27616 14608 27668
rect 16212 27616 16264 27668
rect 17040 27616 17092 27668
rect 17500 27616 17552 27668
rect 18052 27616 18104 27668
rect 18144 27616 18196 27668
rect 19524 27616 19576 27668
rect 20720 27616 20772 27668
rect 20812 27616 20864 27668
rect 17776 27548 17828 27600
rect 11612 27412 11664 27464
rect 9220 27344 9272 27396
rect 9588 27344 9640 27396
rect 9956 27344 10008 27396
rect 10600 27344 10652 27396
rect 7104 27276 7156 27328
rect 8392 27276 8444 27328
rect 8484 27319 8536 27328
rect 8484 27285 8493 27319
rect 8493 27285 8527 27319
rect 8527 27285 8536 27319
rect 8484 27276 8536 27285
rect 9404 27276 9456 27328
rect 10784 27276 10836 27328
rect 11152 27276 11204 27328
rect 11888 27387 11940 27396
rect 11888 27353 11897 27387
rect 11897 27353 11931 27387
rect 11931 27353 11940 27387
rect 11888 27344 11940 27353
rect 11980 27344 12032 27396
rect 12256 27387 12308 27396
rect 12256 27353 12265 27387
rect 12265 27353 12299 27387
rect 12299 27353 12308 27387
rect 12256 27344 12308 27353
rect 12992 27412 13044 27464
rect 13084 27412 13136 27464
rect 13268 27412 13320 27464
rect 18144 27480 18196 27532
rect 19064 27480 19116 27532
rect 20260 27480 20312 27532
rect 21640 27480 21692 27532
rect 17316 27455 17368 27464
rect 17316 27421 17325 27455
rect 17325 27421 17359 27455
rect 17359 27421 17368 27455
rect 17316 27412 17368 27421
rect 17408 27455 17460 27464
rect 17408 27421 17417 27455
rect 17417 27421 17451 27455
rect 17451 27421 17460 27455
rect 17408 27412 17460 27421
rect 15936 27344 15988 27396
rect 20996 27455 21048 27464
rect 20996 27421 21005 27455
rect 21005 27421 21039 27455
rect 21039 27421 21048 27455
rect 20996 27412 21048 27421
rect 12716 27276 12768 27328
rect 14464 27276 14516 27328
rect 15476 27276 15528 27328
rect 19616 27344 19668 27396
rect 20720 27276 20772 27328
rect 22192 27344 22244 27396
rect 20996 27276 21048 27328
rect 6148 27174 6200 27226
rect 6212 27174 6264 27226
rect 6276 27174 6328 27226
rect 6340 27174 6392 27226
rect 6404 27174 6456 27226
rect 11346 27174 11398 27226
rect 11410 27174 11462 27226
rect 11474 27174 11526 27226
rect 11538 27174 11590 27226
rect 11602 27174 11654 27226
rect 16544 27174 16596 27226
rect 16608 27174 16660 27226
rect 16672 27174 16724 27226
rect 16736 27174 16788 27226
rect 16800 27174 16852 27226
rect 21742 27174 21794 27226
rect 21806 27174 21858 27226
rect 21870 27174 21922 27226
rect 21934 27174 21986 27226
rect 21998 27174 22050 27226
rect 1216 27072 1268 27124
rect 2412 27072 2464 27124
rect 2504 27072 2556 27124
rect 2596 27072 2648 27124
rect 2688 27072 2740 27124
rect 3332 27072 3384 27124
rect 3700 27072 3752 27124
rect 3976 27072 4028 27124
rect 4252 27072 4304 27124
rect 1308 27004 1360 27056
rect 1400 26979 1452 26988
rect 1400 26945 1409 26979
rect 1409 26945 1443 26979
rect 1443 26945 1452 26979
rect 1400 26936 1452 26945
rect 1492 26936 1544 26988
rect 480 26868 532 26920
rect 1032 26868 1084 26920
rect 2044 26868 2096 26920
rect 2688 26936 2740 26988
rect 2964 26936 3016 26988
rect 3148 26979 3200 26988
rect 3148 26945 3157 26979
rect 3157 26945 3191 26979
rect 3191 26945 3200 26979
rect 3148 26936 3200 26945
rect 3792 27004 3844 27056
rect 4160 27004 4212 27056
rect 5540 27072 5592 27124
rect 10692 27072 10744 27124
rect 11152 27072 11204 27124
rect 3976 26936 4028 26988
rect 5264 27004 5316 27056
rect 5356 27004 5408 27056
rect 6000 27004 6052 27056
rect 8116 27004 8168 27056
rect 9312 27004 9364 27056
rect 2320 26732 2372 26784
rect 4068 26868 4120 26920
rect 4620 26868 4672 26920
rect 2504 26843 2556 26852
rect 2504 26809 2513 26843
rect 2513 26809 2547 26843
rect 2547 26809 2556 26843
rect 2504 26800 2556 26809
rect 2596 26732 2648 26784
rect 4068 26775 4120 26784
rect 4068 26741 4077 26775
rect 4077 26741 4111 26775
rect 4111 26741 4120 26775
rect 4068 26732 4120 26741
rect 4436 26775 4488 26784
rect 4436 26741 4445 26775
rect 4445 26741 4479 26775
rect 4479 26741 4488 26775
rect 4436 26732 4488 26741
rect 5632 26868 5684 26920
rect 6552 26911 6604 26920
rect 6552 26877 6561 26911
rect 6561 26877 6595 26911
rect 6595 26877 6604 26911
rect 6552 26868 6604 26877
rect 7380 26979 7432 26988
rect 7380 26945 7414 26979
rect 7414 26945 7432 26979
rect 7380 26936 7432 26945
rect 7564 26979 7616 26988
rect 7564 26945 7573 26979
rect 7573 26945 7607 26979
rect 7607 26945 7616 26979
rect 7564 26936 7616 26945
rect 8668 26936 8720 26988
rect 7104 26868 7156 26920
rect 8116 26868 8168 26920
rect 6000 26732 6052 26784
rect 9772 26936 9824 26988
rect 10140 27004 10192 27056
rect 10784 27004 10836 27056
rect 11796 27004 11848 27056
rect 11980 27047 12032 27056
rect 11980 27013 11989 27047
rect 11989 27013 12023 27047
rect 12023 27013 12032 27047
rect 11980 27004 12032 27013
rect 12164 27004 12216 27056
rect 12256 27004 12308 27056
rect 12624 27004 12676 27056
rect 12992 27004 13044 27056
rect 9404 26868 9456 26920
rect 10692 26936 10744 26988
rect 14832 27072 14884 27124
rect 16120 27072 16172 27124
rect 16856 27072 16908 27124
rect 17316 27072 17368 27124
rect 18052 27072 18104 27124
rect 18144 27115 18196 27124
rect 18144 27081 18153 27115
rect 18153 27081 18187 27115
rect 18187 27081 18196 27115
rect 18144 27072 18196 27081
rect 20260 27072 20312 27124
rect 21272 27072 21324 27124
rect 15660 27004 15712 27056
rect 16304 27004 16356 27056
rect 14648 26979 14700 26988
rect 14648 26945 14657 26979
rect 14657 26945 14691 26979
rect 14691 26945 14700 26979
rect 14648 26936 14700 26945
rect 16120 26979 16172 26988
rect 16120 26945 16129 26979
rect 16129 26945 16163 26979
rect 16163 26945 16172 26979
rect 16120 26936 16172 26945
rect 13360 26868 13412 26920
rect 13636 26868 13688 26920
rect 14464 26868 14516 26920
rect 14740 26911 14792 26920
rect 14740 26877 14774 26911
rect 14774 26877 14792 26911
rect 14740 26868 14792 26877
rect 15292 26868 15344 26920
rect 16856 26936 16908 26988
rect 19892 27009 19944 27056
rect 8760 26732 8812 26784
rect 9312 26775 9364 26784
rect 9312 26741 9321 26775
rect 9321 26741 9355 26775
rect 9355 26741 9364 26775
rect 9312 26732 9364 26741
rect 9772 26775 9824 26784
rect 9772 26741 9781 26775
rect 9781 26741 9815 26775
rect 9815 26741 9824 26775
rect 9772 26732 9824 26741
rect 12992 26775 13044 26784
rect 12992 26741 13001 26775
rect 13001 26741 13035 26775
rect 13035 26741 13044 26775
rect 12992 26732 13044 26741
rect 13636 26732 13688 26784
rect 14740 26732 14792 26784
rect 15660 26775 15712 26784
rect 15660 26741 15669 26775
rect 15669 26741 15703 26775
rect 15703 26741 15712 26775
rect 15660 26732 15712 26741
rect 15752 26732 15804 26784
rect 19892 27004 19917 27009
rect 19917 27004 19944 27009
rect 20076 27004 20128 27056
rect 18144 26868 18196 26920
rect 17040 26732 17092 26784
rect 18880 26732 18932 26784
rect 21272 26911 21324 26920
rect 21272 26877 21281 26911
rect 21281 26877 21315 26911
rect 21315 26877 21324 26911
rect 21272 26868 21324 26877
rect 20628 26843 20680 26852
rect 20628 26809 20637 26843
rect 20637 26809 20671 26843
rect 20671 26809 20680 26843
rect 20628 26800 20680 26809
rect 20444 26732 20496 26784
rect 22652 26732 22704 26784
rect 3549 26630 3601 26682
rect 3613 26630 3665 26682
rect 3677 26630 3729 26682
rect 3741 26630 3793 26682
rect 3805 26630 3857 26682
rect 8747 26630 8799 26682
rect 8811 26630 8863 26682
rect 8875 26630 8927 26682
rect 8939 26630 8991 26682
rect 9003 26630 9055 26682
rect 13945 26630 13997 26682
rect 14009 26630 14061 26682
rect 14073 26630 14125 26682
rect 14137 26630 14189 26682
rect 14201 26630 14253 26682
rect 19143 26630 19195 26682
rect 19207 26630 19259 26682
rect 19271 26630 19323 26682
rect 19335 26630 19387 26682
rect 19399 26630 19451 26682
rect 2964 26571 3016 26580
rect 2964 26537 2973 26571
rect 2973 26537 3007 26571
rect 3007 26537 3016 26571
rect 2964 26528 3016 26537
rect 3148 26528 3200 26580
rect 1400 26435 1452 26444
rect 1400 26401 1409 26435
rect 1409 26401 1443 26435
rect 1443 26401 1452 26435
rect 1400 26392 1452 26401
rect 2044 26324 2096 26376
rect 2504 26460 2556 26512
rect 3332 26460 3384 26512
rect 3424 26460 3476 26512
rect 4620 26460 4672 26512
rect 1584 26256 1636 26308
rect 3056 26367 3108 26376
rect 3056 26333 3065 26367
rect 3065 26333 3099 26367
rect 3099 26333 3108 26367
rect 3056 26324 3108 26333
rect 3332 26367 3384 26376
rect 3332 26333 3341 26367
rect 3341 26333 3375 26367
rect 3375 26333 3384 26367
rect 3332 26324 3384 26333
rect 2412 26231 2464 26240
rect 2412 26197 2421 26231
rect 2421 26197 2455 26231
rect 2455 26197 2464 26231
rect 2412 26188 2464 26197
rect 2780 26188 2832 26240
rect 5172 26324 5224 26376
rect 5356 26367 5408 26376
rect 5356 26333 5365 26367
rect 5365 26333 5399 26367
rect 5399 26333 5408 26367
rect 5356 26324 5408 26333
rect 6000 26435 6052 26444
rect 6000 26401 6009 26435
rect 6009 26401 6043 26435
rect 6043 26401 6052 26435
rect 6000 26392 6052 26401
rect 6920 26392 6972 26444
rect 6276 26367 6328 26376
rect 6276 26333 6285 26367
rect 6285 26333 6319 26367
rect 6319 26333 6328 26367
rect 6276 26324 6328 26333
rect 6644 26188 6696 26240
rect 7196 26231 7248 26240
rect 7196 26197 7205 26231
rect 7205 26197 7239 26231
rect 7239 26197 7248 26231
rect 7196 26188 7248 26197
rect 8484 26528 8536 26580
rect 9128 26528 9180 26580
rect 9772 26528 9824 26580
rect 12532 26528 12584 26580
rect 13636 26528 13688 26580
rect 14464 26528 14516 26580
rect 9312 26435 9364 26444
rect 9312 26401 9321 26435
rect 9321 26401 9355 26435
rect 9355 26401 9364 26435
rect 9312 26392 9364 26401
rect 7840 26324 7892 26376
rect 8116 26324 8168 26376
rect 9772 26367 9824 26376
rect 9772 26333 9781 26367
rect 9781 26333 9815 26367
rect 9815 26333 9824 26367
rect 9772 26324 9824 26333
rect 9956 26324 10008 26376
rect 12716 26392 12768 26444
rect 15016 26528 15068 26580
rect 16120 26528 16172 26580
rect 17408 26528 17460 26580
rect 18236 26528 18288 26580
rect 15200 26392 15252 26444
rect 15292 26435 15344 26444
rect 15292 26401 15301 26435
rect 15301 26401 15335 26435
rect 15335 26401 15344 26435
rect 15292 26392 15344 26401
rect 20076 26571 20128 26580
rect 20076 26537 20085 26571
rect 20085 26537 20119 26571
rect 20119 26537 20128 26571
rect 20076 26528 20128 26537
rect 20444 26571 20496 26580
rect 20444 26537 20453 26571
rect 20453 26537 20487 26571
rect 20487 26537 20496 26571
rect 20444 26528 20496 26537
rect 20628 26528 20680 26580
rect 20720 26528 20772 26580
rect 21272 26528 21324 26580
rect 10784 26324 10836 26376
rect 10876 26324 10928 26376
rect 13912 26324 13964 26376
rect 14188 26324 14240 26376
rect 9220 26256 9272 26308
rect 11980 26256 12032 26308
rect 12256 26256 12308 26308
rect 12624 26256 12676 26308
rect 12992 26256 13044 26308
rect 16120 26256 16172 26308
rect 16396 26324 16448 26376
rect 16304 26303 16329 26308
rect 16329 26303 16356 26308
rect 16304 26256 16356 26303
rect 19524 26324 19576 26376
rect 19156 26256 19208 26308
rect 19800 26324 19852 26376
rect 20260 26367 20312 26376
rect 20260 26333 20269 26367
rect 20269 26333 20303 26367
rect 20303 26333 20312 26367
rect 20260 26324 20312 26333
rect 20904 26324 20956 26376
rect 21272 26256 21324 26308
rect 22284 26256 22336 26308
rect 7840 26188 7892 26240
rect 8484 26231 8536 26240
rect 8484 26197 8493 26231
rect 8493 26197 8527 26231
rect 8527 26197 8536 26231
rect 8484 26188 8536 26197
rect 9312 26188 9364 26240
rect 10508 26188 10560 26240
rect 11152 26188 11204 26240
rect 12164 26188 12216 26240
rect 13544 26188 13596 26240
rect 16212 26188 16264 26240
rect 18512 26188 18564 26240
rect 19800 26188 19852 26240
rect 6148 26086 6200 26138
rect 6212 26086 6264 26138
rect 6276 26086 6328 26138
rect 6340 26086 6392 26138
rect 6404 26086 6456 26138
rect 11346 26086 11398 26138
rect 11410 26086 11462 26138
rect 11474 26086 11526 26138
rect 11538 26086 11590 26138
rect 11602 26086 11654 26138
rect 16544 26086 16596 26138
rect 16608 26086 16660 26138
rect 16672 26086 16724 26138
rect 16736 26086 16788 26138
rect 16800 26086 16852 26138
rect 21742 26086 21794 26138
rect 21806 26086 21858 26138
rect 21870 26086 21922 26138
rect 21934 26086 21986 26138
rect 21998 26086 22050 26138
rect 3884 25984 3936 26036
rect 5356 25984 5408 26036
rect 7196 25984 7248 26036
rect 7288 25984 7340 26036
rect 8208 26027 8260 26036
rect 8208 25993 8217 26027
rect 8217 25993 8251 26027
rect 8251 25993 8260 26027
rect 8208 25984 8260 25993
rect 1584 25891 1636 25900
rect 1584 25857 1593 25891
rect 1593 25857 1627 25891
rect 1627 25857 1636 25891
rect 1584 25848 1636 25857
rect 2228 25916 2280 25968
rect 2320 25916 2372 25968
rect 3332 25916 3384 25968
rect 3976 25959 4028 25968
rect 3976 25925 3985 25959
rect 3985 25925 4019 25959
rect 4019 25925 4028 25959
rect 3976 25916 4028 25925
rect 2044 25848 2096 25900
rect 3516 25891 3568 25900
rect 3516 25857 3525 25891
rect 3525 25857 3559 25891
rect 3559 25857 3568 25891
rect 3516 25848 3568 25857
rect 8392 25916 8444 25968
rect 10876 25984 10928 26036
rect 8668 25916 8720 25968
rect 7748 25848 7800 25900
rect 7840 25848 7892 25900
rect 13268 25916 13320 25968
rect 13912 26027 13964 26036
rect 13912 25993 13921 26027
rect 13921 25993 13955 26027
rect 13955 25993 13964 26027
rect 13912 25984 13964 25993
rect 14648 25984 14700 26036
rect 15660 25984 15712 26036
rect 9864 25848 9916 25900
rect 10600 25848 10652 25900
rect 11060 25848 11112 25900
rect 11244 25848 11296 25900
rect 12164 25848 12216 25900
rect 13636 25848 13688 25900
rect 14924 25848 14976 25900
rect 15292 25848 15344 25900
rect 15752 25848 15804 25900
rect 16212 25891 16264 25900
rect 16212 25857 16221 25891
rect 16221 25857 16255 25891
rect 16255 25857 16264 25891
rect 16212 25848 16264 25857
rect 17040 25984 17092 26036
rect 18604 25984 18656 26036
rect 19156 26027 19208 26036
rect 19156 25993 19165 26027
rect 19165 25993 19199 26027
rect 19199 25993 19208 26027
rect 19156 25984 19208 25993
rect 19708 25984 19760 26036
rect 17776 25891 17828 25900
rect 17776 25857 17785 25891
rect 17785 25857 17819 25891
rect 17819 25857 17828 25891
rect 17776 25848 17828 25857
rect 6644 25823 6696 25832
rect 6644 25789 6653 25823
rect 6653 25789 6687 25823
rect 6687 25789 6696 25823
rect 6644 25780 6696 25789
rect 4528 25755 4580 25764
rect 4528 25721 4537 25755
rect 4537 25721 4571 25755
rect 4571 25721 4580 25755
rect 4528 25712 4580 25721
rect 12900 25823 12952 25832
rect 12900 25789 12909 25823
rect 12909 25789 12943 25823
rect 12943 25789 12952 25823
rect 12900 25780 12952 25789
rect 18512 25848 18564 25900
rect 19616 25916 19668 25968
rect 20904 25891 20956 25900
rect 20904 25857 20913 25891
rect 20913 25857 20947 25891
rect 20947 25857 20956 25891
rect 20904 25848 20956 25857
rect 18880 25780 18932 25832
rect 20076 25780 20128 25832
rect 7104 25644 7156 25696
rect 9588 25644 9640 25696
rect 10784 25644 10836 25696
rect 12808 25712 12860 25764
rect 12532 25687 12584 25696
rect 12532 25653 12541 25687
rect 12541 25653 12575 25687
rect 12575 25653 12584 25687
rect 12532 25644 12584 25653
rect 13268 25644 13320 25696
rect 15936 25687 15988 25696
rect 15936 25653 15945 25687
rect 15945 25653 15979 25687
rect 15979 25653 15988 25687
rect 15936 25644 15988 25653
rect 17684 25644 17736 25696
rect 18696 25644 18748 25696
rect 19708 25644 19760 25696
rect 20720 25687 20772 25696
rect 20720 25653 20729 25687
rect 20729 25653 20763 25687
rect 20763 25653 20772 25687
rect 20720 25644 20772 25653
rect 21088 25687 21140 25696
rect 21088 25653 21097 25687
rect 21097 25653 21131 25687
rect 21131 25653 21140 25687
rect 21088 25644 21140 25653
rect 21456 25687 21508 25696
rect 21456 25653 21465 25687
rect 21465 25653 21499 25687
rect 21499 25653 21508 25687
rect 21456 25644 21508 25653
rect 3549 25542 3601 25594
rect 3613 25542 3665 25594
rect 3677 25542 3729 25594
rect 3741 25542 3793 25594
rect 3805 25542 3857 25594
rect 8747 25542 8799 25594
rect 8811 25542 8863 25594
rect 8875 25542 8927 25594
rect 8939 25542 8991 25594
rect 9003 25542 9055 25594
rect 13945 25542 13997 25594
rect 14009 25542 14061 25594
rect 14073 25542 14125 25594
rect 14137 25542 14189 25594
rect 14201 25542 14253 25594
rect 19143 25542 19195 25594
rect 19207 25542 19259 25594
rect 19271 25542 19323 25594
rect 19335 25542 19387 25594
rect 19399 25542 19451 25594
rect 2136 25440 2188 25492
rect 3332 25483 3384 25492
rect 3332 25449 3341 25483
rect 3341 25449 3375 25483
rect 3375 25449 3384 25483
rect 3332 25440 3384 25449
rect 1676 25347 1728 25356
rect 1676 25313 1685 25347
rect 1685 25313 1719 25347
rect 1719 25313 1728 25347
rect 1676 25304 1728 25313
rect 1400 25279 1452 25288
rect 1400 25245 1409 25279
rect 1409 25245 1443 25279
rect 1443 25245 1452 25279
rect 1400 25236 1452 25245
rect 6736 25440 6788 25492
rect 7104 25440 7156 25492
rect 6000 25372 6052 25424
rect 2228 25304 2280 25356
rect 5908 25347 5960 25356
rect 5908 25313 5917 25347
rect 5917 25313 5951 25347
rect 5951 25313 5960 25347
rect 5908 25304 5960 25313
rect 6092 25304 6144 25356
rect 2504 25236 2556 25288
rect 3240 25236 3292 25288
rect 4528 25168 4580 25220
rect 5356 25236 5408 25288
rect 5632 25236 5684 25288
rect 6920 25279 6972 25288
rect 6920 25245 6929 25279
rect 6929 25245 6963 25279
rect 6963 25245 6972 25279
rect 6920 25236 6972 25245
rect 8116 25483 8168 25492
rect 8116 25449 8125 25483
rect 8125 25449 8159 25483
rect 8159 25449 8168 25483
rect 8116 25440 8168 25449
rect 8484 25440 8536 25492
rect 9128 25440 9180 25492
rect 8208 25304 8260 25356
rect 8668 25304 8720 25356
rect 10784 25483 10836 25492
rect 10784 25449 10793 25483
rect 10793 25449 10827 25483
rect 10827 25449 10836 25483
rect 10784 25440 10836 25449
rect 12808 25440 12860 25492
rect 12532 25304 12584 25356
rect 9864 25279 9916 25288
rect 9864 25245 9873 25279
rect 9873 25245 9907 25279
rect 9907 25245 9916 25279
rect 9864 25236 9916 25245
rect 10140 25279 10192 25288
rect 10140 25245 10149 25279
rect 10149 25245 10183 25279
rect 10183 25245 10192 25279
rect 10140 25236 10192 25245
rect 11980 25236 12032 25288
rect 12348 25236 12400 25288
rect 12808 25236 12860 25288
rect 14832 25236 14884 25288
rect 15016 25236 15068 25288
rect 15384 25279 15436 25288
rect 8392 25168 8444 25220
rect 8668 25168 8720 25220
rect 11888 25211 11940 25220
rect 11888 25177 11897 25211
rect 11897 25177 11931 25211
rect 11931 25177 11940 25211
rect 11888 25168 11940 25177
rect 12256 25211 12308 25220
rect 12256 25177 12265 25211
rect 12265 25177 12299 25211
rect 12299 25177 12308 25211
rect 12256 25168 12308 25177
rect 15384 25245 15391 25279
rect 15391 25245 15425 25279
rect 15425 25245 15436 25279
rect 15384 25236 15436 25245
rect 16028 25168 16080 25220
rect 6920 25100 6972 25152
rect 9404 25100 9456 25152
rect 11152 25100 11204 25152
rect 12348 25100 12400 25152
rect 12624 25143 12676 25152
rect 12624 25109 12633 25143
rect 12633 25109 12667 25143
rect 12667 25109 12676 25143
rect 12624 25100 12676 25109
rect 13360 25100 13412 25152
rect 14280 25100 14332 25152
rect 14924 25100 14976 25152
rect 15844 25100 15896 25152
rect 16120 25143 16172 25152
rect 16120 25109 16129 25143
rect 16129 25109 16163 25143
rect 16163 25109 16172 25143
rect 16120 25100 16172 25109
rect 18512 25236 18564 25288
rect 18880 25279 18932 25288
rect 18880 25245 18889 25279
rect 18889 25245 18923 25279
rect 18923 25245 18932 25279
rect 18880 25236 18932 25245
rect 19524 25483 19576 25492
rect 19524 25449 19533 25483
rect 19533 25449 19567 25483
rect 19567 25449 19576 25483
rect 19524 25440 19576 25449
rect 19616 25483 19668 25492
rect 19616 25449 19625 25483
rect 19625 25449 19659 25483
rect 19659 25449 19668 25483
rect 19616 25440 19668 25449
rect 19708 25440 19760 25492
rect 19800 25440 19852 25492
rect 20076 25483 20128 25492
rect 20076 25449 20085 25483
rect 20085 25449 20119 25483
rect 20119 25449 20128 25483
rect 20076 25440 20128 25449
rect 20720 25440 20772 25492
rect 17040 25100 17092 25152
rect 17408 25100 17460 25152
rect 17500 25143 17552 25152
rect 17500 25109 17509 25143
rect 17509 25109 17543 25143
rect 17543 25109 17552 25143
rect 17500 25100 17552 25109
rect 18972 25168 19024 25220
rect 19892 25168 19944 25220
rect 18604 25143 18656 25152
rect 18604 25109 18613 25143
rect 18613 25109 18647 25143
rect 18647 25109 18656 25143
rect 18604 25100 18656 25109
rect 19708 25100 19760 25152
rect 20536 25304 20588 25356
rect 20444 25279 20496 25288
rect 20444 25245 20453 25279
rect 20453 25245 20487 25279
rect 20487 25245 20496 25279
rect 20444 25236 20496 25245
rect 20536 25168 20588 25220
rect 21272 25236 21324 25288
rect 22284 25168 22336 25220
rect 20628 25143 20680 25152
rect 20628 25109 20637 25143
rect 20637 25109 20671 25143
rect 20671 25109 20680 25143
rect 20628 25100 20680 25109
rect 20720 25143 20772 25152
rect 20720 25109 20729 25143
rect 20729 25109 20763 25143
rect 20763 25109 20772 25143
rect 20720 25100 20772 25109
rect 20 25032 72 25084
rect 296 25032 348 25084
rect 6148 24998 6200 25050
rect 6212 24998 6264 25050
rect 6276 24998 6328 25050
rect 6340 24998 6392 25050
rect 6404 24998 6456 25050
rect 11346 24998 11398 25050
rect 11410 24998 11462 25050
rect 11474 24998 11526 25050
rect 11538 24998 11590 25050
rect 11602 24998 11654 25050
rect 16544 24998 16596 25050
rect 16608 24998 16660 25050
rect 16672 24998 16724 25050
rect 16736 24998 16788 25050
rect 16800 24998 16852 25050
rect 21742 24998 21794 25050
rect 21806 24998 21858 25050
rect 21870 24998 21922 25050
rect 21934 24998 21986 25050
rect 21998 24998 22050 25050
rect 2872 24896 2924 24948
rect 4068 24896 4120 24948
rect 4988 24896 5040 24948
rect 5448 24896 5500 24948
rect 6000 24896 6052 24948
rect 1860 24871 1912 24880
rect 1860 24837 1869 24871
rect 1869 24837 1903 24871
rect 1903 24837 1912 24871
rect 1860 24828 1912 24837
rect 2136 24871 2188 24880
rect 2136 24837 2145 24871
rect 2145 24837 2179 24871
rect 2179 24837 2188 24871
rect 2136 24828 2188 24837
rect 3332 24828 3384 24880
rect 4528 24828 4580 24880
rect 5908 24828 5960 24880
rect 8116 24896 8168 24948
rect 9864 24896 9916 24948
rect 10140 24896 10192 24948
rect 11888 24896 11940 24948
rect 6552 24828 6604 24880
rect 9496 24828 9548 24880
rect 10784 24828 10836 24880
rect 12440 24828 12492 24880
rect 848 24760 900 24812
rect 2504 24760 2556 24812
rect 3424 24760 3476 24812
rect 6828 24760 6880 24812
rect 7288 24760 7340 24812
rect 8760 24760 8812 24812
rect 14372 24896 14424 24948
rect 13820 24828 13872 24880
rect 10508 24760 10560 24812
rect 11244 24760 11296 24812
rect 12532 24760 12584 24812
rect 12992 24760 13044 24812
rect 13452 24779 13459 24812
rect 13459 24779 13493 24812
rect 13493 24779 13504 24812
rect 13452 24760 13504 24779
rect 2412 24692 2464 24744
rect 3884 24692 3936 24744
rect 3608 24556 3660 24608
rect 4344 24556 4396 24608
rect 5724 24624 5776 24676
rect 7380 24692 7432 24744
rect 7840 24735 7892 24744
rect 7840 24701 7849 24735
rect 7849 24701 7883 24735
rect 7883 24701 7892 24735
rect 7840 24692 7892 24701
rect 7104 24624 7156 24676
rect 9036 24692 9088 24744
rect 9220 24692 9272 24744
rect 8300 24667 8352 24676
rect 8300 24633 8309 24667
rect 8309 24633 8343 24667
rect 8343 24633 8352 24667
rect 8300 24624 8352 24633
rect 5632 24556 5684 24608
rect 8392 24556 8444 24608
rect 9404 24624 9456 24676
rect 9496 24599 9548 24608
rect 9496 24565 9505 24599
rect 9505 24565 9539 24599
rect 9539 24565 9548 24599
rect 9496 24556 9548 24565
rect 14740 24803 14792 24812
rect 14740 24769 14749 24803
rect 14749 24769 14783 24803
rect 14783 24769 14792 24803
rect 14740 24760 14792 24769
rect 14924 24760 14976 24812
rect 18144 24896 18196 24948
rect 18880 24896 18932 24948
rect 19524 24896 19576 24948
rect 20720 24896 20772 24948
rect 20904 24896 20956 24948
rect 22008 24896 22060 24948
rect 22192 24896 22244 24948
rect 17776 24828 17828 24880
rect 19892 24871 19944 24880
rect 17408 24760 17460 24812
rect 18604 24760 18656 24812
rect 18696 24760 18748 24812
rect 18880 24760 18932 24812
rect 18972 24760 19024 24812
rect 19892 24837 19926 24871
rect 19926 24837 19944 24871
rect 19892 24828 19944 24837
rect 20076 24828 20128 24880
rect 19340 24692 19392 24744
rect 14372 24624 14424 24676
rect 13176 24556 13228 24608
rect 14648 24599 14700 24608
rect 14648 24565 14657 24599
rect 14657 24565 14691 24599
rect 14691 24565 14700 24599
rect 14648 24556 14700 24565
rect 15016 24556 15068 24608
rect 16028 24599 16080 24608
rect 16028 24565 16037 24599
rect 16037 24565 16071 24599
rect 16071 24565 16080 24599
rect 16028 24556 16080 24565
rect 21456 24599 21508 24608
rect 21456 24565 21465 24599
rect 21465 24565 21499 24599
rect 21499 24565 21508 24599
rect 21456 24556 21508 24565
rect 3549 24454 3601 24506
rect 3613 24454 3665 24506
rect 3677 24454 3729 24506
rect 3741 24454 3793 24506
rect 3805 24454 3857 24506
rect 8747 24454 8799 24506
rect 8811 24454 8863 24506
rect 8875 24454 8927 24506
rect 8939 24454 8991 24506
rect 9003 24454 9055 24506
rect 13945 24454 13997 24506
rect 14009 24454 14061 24506
rect 14073 24454 14125 24506
rect 14137 24454 14189 24506
rect 14201 24454 14253 24506
rect 19143 24454 19195 24506
rect 19207 24454 19259 24506
rect 19271 24454 19323 24506
rect 19335 24454 19387 24506
rect 19399 24454 19451 24506
rect 1768 24352 1820 24404
rect 2504 24352 2556 24404
rect 3240 24352 3292 24404
rect 4252 24352 4304 24404
rect 1400 24284 1452 24336
rect 4988 24284 5040 24336
rect 5632 24352 5684 24404
rect 5724 24352 5776 24404
rect 756 24148 808 24200
rect 1492 24148 1544 24200
rect 2596 24148 2648 24200
rect 4344 24080 4396 24132
rect 4528 24148 4580 24200
rect 4804 24148 4856 24200
rect 4896 24191 4948 24200
rect 4896 24157 4905 24191
rect 4905 24157 4939 24191
rect 4939 24157 4948 24191
rect 4896 24148 4948 24157
rect 6092 24216 6144 24268
rect 8300 24352 8352 24404
rect 9496 24352 9548 24404
rect 10048 24352 10100 24404
rect 5908 24191 5960 24200
rect 5908 24157 5917 24191
rect 5917 24157 5951 24191
rect 5951 24157 5960 24191
rect 5908 24148 5960 24157
rect 6828 24148 6880 24200
rect 7564 24148 7616 24200
rect 7932 24148 7984 24200
rect 10048 24191 10100 24200
rect 10048 24157 10057 24191
rect 10057 24157 10091 24191
rect 10091 24157 10100 24191
rect 10048 24148 10100 24157
rect 10324 24148 10376 24200
rect 6552 24055 6604 24064
rect 6552 24021 6561 24055
rect 6561 24021 6595 24055
rect 6595 24021 6604 24055
rect 6552 24012 6604 24021
rect 7748 24012 7800 24064
rect 11244 24080 11296 24132
rect 12440 24352 12492 24404
rect 13176 24352 13228 24404
rect 14372 24352 14424 24404
rect 14648 24352 14700 24404
rect 14832 24352 14884 24404
rect 15476 24352 15528 24404
rect 16948 24352 17000 24404
rect 17408 24352 17460 24404
rect 13820 24148 13872 24200
rect 14280 24191 14332 24200
rect 14280 24157 14289 24191
rect 14289 24157 14323 24191
rect 14323 24157 14332 24191
rect 14280 24148 14332 24157
rect 16120 24284 16172 24336
rect 17500 24216 17552 24268
rect 18696 24352 18748 24404
rect 18880 24352 18932 24404
rect 20536 24352 20588 24404
rect 20628 24352 20680 24404
rect 21088 24352 21140 24404
rect 18972 24216 19024 24268
rect 19064 24216 19116 24268
rect 14924 24191 14976 24200
rect 14924 24157 14933 24191
rect 14933 24157 14967 24191
rect 14967 24157 14976 24191
rect 14924 24148 14976 24157
rect 15200 24148 15252 24200
rect 15292 24148 15344 24200
rect 16304 24191 16356 24200
rect 16304 24157 16313 24191
rect 16313 24157 16347 24191
rect 16347 24157 16356 24191
rect 16304 24148 16356 24157
rect 16396 24191 16448 24200
rect 16396 24157 16430 24191
rect 16430 24157 16448 24191
rect 16396 24148 16448 24157
rect 14372 24080 14424 24132
rect 14832 24080 14884 24132
rect 17500 24080 17552 24132
rect 17684 24080 17736 24132
rect 18880 24148 18932 24200
rect 17868 24127 17893 24132
rect 17893 24127 17920 24132
rect 17868 24080 17920 24127
rect 18052 24080 18104 24132
rect 19340 24080 19392 24132
rect 19708 24080 19760 24132
rect 19892 24080 19944 24132
rect 9864 24055 9916 24064
rect 9864 24021 9873 24055
rect 9873 24021 9907 24055
rect 9907 24021 9916 24055
rect 9864 24012 9916 24021
rect 10140 24012 10192 24064
rect 10876 24012 10928 24064
rect 11152 24055 11204 24064
rect 11152 24021 11161 24055
rect 11161 24021 11195 24055
rect 11195 24021 11204 24055
rect 11152 24012 11204 24021
rect 11704 24055 11756 24064
rect 11704 24021 11713 24055
rect 11713 24021 11747 24055
rect 11747 24021 11756 24055
rect 11704 24012 11756 24021
rect 13452 24055 13504 24064
rect 13452 24021 13461 24055
rect 13461 24021 13495 24055
rect 13495 24021 13504 24055
rect 13452 24012 13504 24021
rect 13820 24012 13872 24064
rect 14648 24012 14700 24064
rect 16304 24012 16356 24064
rect 17316 24012 17368 24064
rect 20168 24012 20220 24064
rect 20628 24148 20680 24200
rect 20904 24148 20956 24200
rect 21088 24080 21140 24132
rect 21548 24080 21600 24132
rect 20996 24055 21048 24064
rect 20996 24021 21005 24055
rect 21005 24021 21039 24055
rect 21039 24021 21048 24055
rect 20996 24012 21048 24021
rect 22192 24012 22244 24064
rect 6148 23910 6200 23962
rect 6212 23910 6264 23962
rect 6276 23910 6328 23962
rect 6340 23910 6392 23962
rect 6404 23910 6456 23962
rect 11346 23910 11398 23962
rect 11410 23910 11462 23962
rect 11474 23910 11526 23962
rect 11538 23910 11590 23962
rect 11602 23910 11654 23962
rect 16544 23910 16596 23962
rect 16608 23910 16660 23962
rect 16672 23910 16724 23962
rect 16736 23910 16788 23962
rect 16800 23910 16852 23962
rect 21742 23910 21794 23962
rect 21806 23910 21858 23962
rect 21870 23910 21922 23962
rect 21934 23910 21986 23962
rect 21998 23910 22050 23962
rect 5356 23740 5408 23792
rect 1400 23715 1452 23724
rect 1400 23681 1409 23715
rect 1409 23681 1443 23715
rect 1443 23681 1452 23715
rect 1400 23672 1452 23681
rect 1768 23672 1820 23724
rect 3884 23672 3936 23724
rect 5172 23715 5224 23724
rect 5172 23681 5179 23715
rect 5179 23681 5213 23715
rect 5213 23681 5224 23715
rect 5172 23672 5224 23681
rect 6552 23672 6604 23724
rect 2780 23647 2832 23656
rect 2780 23613 2789 23647
rect 2789 23613 2823 23647
rect 2823 23613 2832 23647
rect 2780 23604 2832 23613
rect 3976 23604 4028 23656
rect 7472 23672 7524 23724
rect 7564 23672 7616 23724
rect 8116 23672 8168 23724
rect 664 23468 716 23520
rect 4436 23536 4488 23588
rect 8024 23604 8076 23656
rect 8300 23604 8352 23656
rect 8760 23647 8812 23656
rect 8760 23613 8794 23647
rect 8794 23613 8812 23647
rect 8760 23604 8812 23613
rect 9128 23604 9180 23656
rect 9864 23808 9916 23860
rect 10968 23808 11020 23860
rect 11612 23808 11664 23860
rect 11704 23808 11756 23860
rect 11888 23808 11940 23860
rect 12808 23808 12860 23860
rect 11244 23672 11296 23724
rect 11704 23672 11756 23724
rect 11980 23672 12032 23724
rect 12716 23740 12768 23792
rect 12900 23740 12952 23792
rect 14924 23808 14976 23860
rect 15200 23740 15252 23792
rect 20628 23851 20680 23860
rect 20628 23817 20637 23851
rect 20637 23817 20671 23851
rect 20671 23817 20680 23851
rect 20628 23808 20680 23817
rect 12624 23672 12676 23724
rect 12900 23647 12952 23656
rect 12900 23613 12909 23647
rect 12909 23613 12943 23647
rect 12943 23613 12952 23647
rect 12900 23604 12952 23613
rect 2320 23468 2372 23520
rect 5908 23511 5960 23520
rect 5908 23477 5917 23511
rect 5917 23477 5951 23511
rect 5951 23477 5960 23511
rect 5908 23468 5960 23477
rect 6460 23468 6512 23520
rect 6552 23468 6604 23520
rect 9588 23536 9640 23588
rect 10508 23536 10560 23588
rect 10968 23536 11020 23588
rect 7472 23511 7524 23520
rect 7472 23477 7481 23511
rect 7481 23477 7515 23511
rect 7515 23477 7524 23511
rect 7472 23468 7524 23477
rect 7656 23468 7708 23520
rect 8760 23468 8812 23520
rect 11152 23468 11204 23520
rect 11428 23468 11480 23520
rect 11612 23536 11664 23588
rect 11980 23536 12032 23588
rect 12716 23536 12768 23588
rect 13084 23468 13136 23520
rect 13820 23715 13872 23724
rect 13820 23681 13829 23715
rect 13829 23681 13863 23715
rect 13863 23681 13872 23715
rect 13820 23672 13872 23681
rect 13452 23604 13504 23656
rect 13912 23647 13964 23656
rect 13912 23613 13946 23647
rect 13946 23613 13964 23647
rect 13912 23604 13964 23613
rect 14280 23604 14332 23656
rect 17316 23672 17368 23724
rect 14832 23647 14884 23656
rect 14832 23613 14841 23647
rect 14841 23613 14875 23647
rect 14875 23613 14884 23647
rect 14832 23604 14884 23613
rect 15844 23604 15896 23656
rect 16120 23604 16172 23656
rect 19248 23715 19300 23724
rect 19248 23681 19257 23715
rect 19257 23681 19291 23715
rect 19291 23681 19300 23715
rect 19248 23672 19300 23681
rect 19340 23672 19392 23724
rect 19892 23715 19944 23724
rect 19892 23681 19899 23715
rect 19899 23681 19933 23715
rect 19933 23681 19944 23715
rect 19892 23672 19944 23681
rect 20536 23672 20588 23724
rect 19524 23536 19576 23588
rect 14556 23468 14608 23520
rect 17684 23511 17736 23520
rect 17684 23477 17693 23511
rect 17693 23477 17727 23511
rect 17727 23477 17736 23511
rect 17684 23468 17736 23477
rect 18972 23468 19024 23520
rect 19616 23468 19668 23520
rect 20720 23468 20772 23520
rect 3549 23366 3601 23418
rect 3613 23366 3665 23418
rect 3677 23366 3729 23418
rect 3741 23366 3793 23418
rect 3805 23366 3857 23418
rect 8747 23366 8799 23418
rect 8811 23366 8863 23418
rect 8875 23366 8927 23418
rect 8939 23366 8991 23418
rect 9003 23366 9055 23418
rect 13945 23366 13997 23418
rect 14009 23366 14061 23418
rect 14073 23366 14125 23418
rect 14137 23366 14189 23418
rect 14201 23366 14253 23418
rect 19143 23366 19195 23418
rect 19207 23366 19259 23418
rect 19271 23366 19323 23418
rect 19335 23366 19387 23418
rect 19399 23366 19451 23418
rect 1124 23264 1176 23316
rect 3240 23239 3292 23248
rect 3240 23205 3249 23239
rect 3249 23205 3283 23239
rect 3283 23205 3292 23239
rect 3240 23196 3292 23205
rect 1492 23128 1544 23180
rect 1400 23103 1452 23112
rect 1400 23069 1409 23103
rect 1409 23069 1443 23103
rect 1443 23069 1452 23103
rect 1400 23060 1452 23069
rect 1860 23060 1912 23112
rect 2688 23060 2740 23112
rect 3424 23264 3476 23316
rect 4804 23264 4856 23316
rect 5724 23264 5776 23316
rect 5816 23264 5868 23316
rect 6276 23264 6328 23316
rect 5632 23196 5684 23248
rect 6276 23171 6328 23180
rect 6276 23137 6310 23171
rect 6310 23137 6328 23171
rect 6276 23128 6328 23137
rect 6460 23171 6512 23180
rect 6460 23137 6469 23171
rect 6469 23137 6503 23171
rect 6503 23137 6512 23171
rect 6460 23128 6512 23137
rect 6828 23128 6880 23180
rect 7748 23264 7800 23316
rect 7932 23264 7984 23316
rect 9128 23264 9180 23316
rect 1308 22992 1360 23044
rect 3424 23060 3476 23112
rect 3792 23103 3844 23112
rect 3792 23069 3801 23103
rect 3801 23069 3835 23103
rect 3835 23069 3844 23103
rect 3792 23060 3844 23069
rect 3976 23060 4028 23112
rect 4712 23060 4764 23112
rect 5264 23103 5316 23112
rect 5264 23069 5273 23103
rect 5273 23069 5307 23103
rect 5307 23069 5316 23103
rect 5264 23060 5316 23069
rect 5356 23060 5408 23112
rect 7748 23103 7800 23112
rect 4620 22992 4672 23044
rect 4988 22992 5040 23044
rect 7748 23069 7755 23103
rect 7755 23069 7789 23103
rect 7789 23069 7800 23103
rect 7748 23060 7800 23069
rect 9680 23103 9732 23112
rect 9680 23069 9689 23103
rect 9689 23069 9723 23103
rect 9723 23069 9732 23103
rect 9680 23060 9732 23069
rect 10048 23060 10100 23112
rect 1584 22967 1636 22976
rect 1584 22933 1593 22967
rect 1593 22933 1627 22967
rect 1627 22933 1636 22967
rect 1584 22924 1636 22933
rect 2504 22924 2556 22976
rect 4068 22924 4120 22976
rect 4344 22924 4396 22976
rect 4804 22967 4856 22976
rect 4804 22933 4813 22967
rect 4813 22933 4847 22967
rect 4847 22933 4856 22967
rect 4804 22924 4856 22933
rect 5448 22924 5500 22976
rect 6552 22924 6604 22976
rect 9772 22992 9824 23044
rect 10324 22992 10376 23044
rect 10692 23264 10744 23316
rect 11520 23264 11572 23316
rect 11244 23060 11296 23112
rect 12164 23264 12216 23316
rect 14280 23264 14332 23316
rect 14556 23264 14608 23316
rect 14740 23264 14792 23316
rect 13820 23196 13872 23248
rect 16396 23264 16448 23316
rect 16028 23239 16080 23248
rect 16028 23205 16037 23239
rect 16037 23205 16071 23239
rect 16071 23205 16080 23239
rect 16028 23196 16080 23205
rect 19524 23264 19576 23316
rect 19616 23264 19668 23316
rect 19892 23264 19944 23316
rect 20536 23307 20588 23316
rect 20536 23273 20545 23307
rect 20545 23273 20579 23307
rect 20579 23273 20588 23307
rect 20536 23264 20588 23273
rect 21548 23264 21600 23316
rect 17960 23196 18012 23248
rect 18512 23196 18564 23248
rect 12164 23128 12216 23180
rect 12348 23128 12400 23180
rect 15200 23128 15252 23180
rect 15752 23128 15804 23180
rect 17684 23128 17736 23180
rect 12624 23060 12676 23112
rect 12808 23060 12860 23112
rect 8024 22924 8076 22976
rect 8208 22924 8260 22976
rect 9864 22924 9916 22976
rect 10692 22967 10744 22976
rect 10692 22933 10701 22967
rect 10701 22933 10735 22967
rect 10735 22933 10744 22967
rect 10692 22924 10744 22933
rect 11520 22924 11572 22976
rect 14556 22992 14608 23044
rect 12624 22924 12676 22976
rect 13268 22924 13320 22976
rect 14832 23103 14884 23112
rect 14832 23069 14841 23103
rect 14841 23069 14875 23103
rect 14875 23069 14884 23103
rect 14832 23060 14884 23069
rect 15292 23060 15344 23112
rect 16396 23103 16448 23112
rect 16396 23069 16430 23103
rect 16430 23069 16448 23103
rect 16396 23060 16448 23069
rect 17500 22992 17552 23044
rect 17684 22992 17736 23044
rect 18420 23128 18472 23180
rect 20444 23196 20496 23248
rect 21180 23196 21232 23248
rect 19340 23060 19392 23112
rect 19892 23060 19944 23112
rect 20996 23060 21048 23112
rect 18144 22924 18196 22976
rect 18328 22967 18380 22976
rect 18328 22933 18337 22967
rect 18337 22933 18371 22967
rect 18371 22933 18380 22967
rect 18328 22924 18380 22933
rect 19064 22967 19116 22976
rect 19064 22933 19073 22967
rect 19073 22933 19107 22967
rect 19107 22933 19116 22967
rect 19064 22924 19116 22933
rect 19156 22924 19208 22976
rect 19294 22924 19346 22976
rect 19432 22924 19484 22976
rect 6148 22822 6200 22874
rect 6212 22822 6264 22874
rect 6276 22822 6328 22874
rect 6340 22822 6392 22874
rect 6404 22822 6456 22874
rect 11346 22822 11398 22874
rect 11410 22822 11462 22874
rect 11474 22822 11526 22874
rect 11538 22822 11590 22874
rect 11602 22822 11654 22874
rect 16544 22822 16596 22874
rect 16608 22822 16660 22874
rect 16672 22822 16724 22874
rect 16736 22822 16788 22874
rect 16800 22822 16852 22874
rect 21742 22822 21794 22874
rect 21806 22822 21858 22874
rect 21870 22822 21922 22874
rect 21934 22822 21986 22874
rect 21998 22822 22050 22874
rect 1676 22763 1728 22772
rect 1676 22729 1685 22763
rect 1685 22729 1719 22763
rect 1719 22729 1728 22763
rect 1676 22720 1728 22729
rect 2872 22720 2924 22772
rect 3056 22720 3108 22772
rect 2504 22652 2556 22704
rect 2780 22695 2832 22704
rect 2780 22661 2789 22695
rect 2789 22661 2823 22695
rect 2823 22661 2832 22695
rect 2780 22652 2832 22661
rect 1952 22627 2004 22636
rect 1952 22593 1961 22627
rect 1961 22593 1995 22627
rect 1995 22593 2004 22627
rect 1952 22584 2004 22593
rect 2412 22627 2464 22636
rect 2412 22593 2421 22627
rect 2421 22593 2455 22627
rect 2455 22593 2464 22627
rect 2412 22584 2464 22593
rect 3516 22652 3568 22704
rect 3608 22695 3660 22704
rect 3608 22661 3617 22695
rect 3617 22661 3651 22695
rect 3651 22661 3660 22695
rect 3608 22652 3660 22661
rect 4804 22720 4856 22772
rect 5908 22720 5960 22772
rect 7380 22720 7432 22772
rect 7932 22720 7984 22772
rect 4344 22652 4396 22704
rect 4436 22695 4488 22704
rect 4436 22661 4445 22695
rect 4445 22661 4479 22695
rect 4479 22661 4488 22695
rect 4436 22652 4488 22661
rect 10324 22720 10376 22772
rect 10508 22720 10560 22772
rect 12808 22720 12860 22772
rect 3424 22584 3476 22636
rect 6828 22627 6880 22636
rect 6828 22593 6837 22627
rect 6837 22593 6871 22627
rect 6871 22593 6880 22627
rect 6828 22584 6880 22593
rect 10048 22652 10100 22704
rect 10692 22652 10744 22704
rect 10876 22652 10928 22704
rect 10968 22695 11020 22704
rect 10968 22661 10977 22695
rect 10977 22661 11011 22695
rect 11011 22661 11020 22695
rect 10968 22652 11020 22661
rect 11796 22652 11848 22704
rect 12348 22652 12400 22704
rect 7472 22584 7524 22636
rect 8668 22584 8720 22636
rect 9496 22584 9548 22636
rect 10324 22584 10376 22636
rect 10508 22584 10560 22636
rect 11244 22584 11296 22636
rect 2320 22516 2372 22568
rect 2964 22516 3016 22568
rect 3884 22516 3936 22568
rect 5080 22516 5132 22568
rect 5448 22516 5500 22568
rect 6552 22516 6604 22568
rect 4620 22491 4672 22500
rect 4620 22457 4629 22491
rect 4629 22457 4663 22491
rect 4663 22457 4672 22491
rect 4620 22448 4672 22457
rect 7932 22448 7984 22500
rect 10048 22516 10100 22568
rect 11152 22516 11204 22568
rect 8484 22448 8536 22500
rect 7748 22380 7800 22432
rect 9128 22380 9180 22432
rect 9864 22380 9916 22432
rect 11152 22423 11204 22432
rect 11152 22389 11161 22423
rect 11161 22389 11195 22423
rect 11195 22389 11204 22423
rect 11152 22380 11204 22389
rect 12808 22584 12860 22636
rect 14832 22720 14884 22772
rect 15752 22720 15804 22772
rect 16396 22720 16448 22772
rect 18052 22720 18104 22772
rect 19064 22720 19116 22772
rect 19432 22720 19484 22772
rect 20352 22763 20404 22772
rect 20352 22729 20361 22763
rect 20361 22729 20395 22763
rect 20395 22729 20404 22763
rect 20352 22720 20404 22729
rect 22192 22720 22244 22772
rect 13084 22627 13136 22636
rect 13084 22593 13093 22627
rect 13093 22593 13127 22627
rect 13127 22593 13136 22627
rect 13084 22584 13136 22593
rect 13452 22516 13504 22568
rect 13084 22448 13136 22500
rect 13912 22559 13964 22568
rect 13912 22525 13946 22559
rect 13946 22525 13964 22559
rect 13912 22516 13964 22525
rect 14280 22516 14332 22568
rect 14740 22516 14792 22568
rect 15016 22380 15068 22432
rect 16396 22584 16448 22636
rect 16948 22584 17000 22636
rect 17776 22584 17828 22636
rect 18144 22627 18196 22636
rect 18144 22593 18178 22627
rect 18178 22593 18196 22627
rect 18144 22584 18196 22593
rect 19340 22652 19392 22704
rect 19156 22584 19208 22636
rect 19493 22594 19545 22646
rect 20168 22584 20220 22636
rect 20812 22584 20864 22636
rect 21916 22652 21968 22704
rect 22744 22652 22796 22704
rect 21732 22584 21784 22636
rect 22376 22584 22428 22636
rect 21548 22559 21600 22568
rect 21548 22525 21557 22559
rect 21557 22525 21591 22559
rect 21591 22525 21600 22559
rect 21548 22516 21600 22525
rect 21272 22448 21324 22500
rect 15936 22423 15988 22432
rect 15936 22389 15945 22423
rect 15945 22389 15979 22423
rect 15979 22389 15988 22423
rect 15936 22380 15988 22389
rect 17776 22380 17828 22432
rect 18972 22380 19024 22432
rect 21364 22423 21416 22432
rect 21364 22389 21373 22423
rect 21373 22389 21407 22423
rect 21407 22389 21416 22423
rect 21364 22380 21416 22389
rect 3549 22278 3601 22330
rect 3613 22278 3665 22330
rect 3677 22278 3729 22330
rect 3741 22278 3793 22330
rect 3805 22278 3857 22330
rect 8747 22278 8799 22330
rect 8811 22278 8863 22330
rect 8875 22278 8927 22330
rect 8939 22278 8991 22330
rect 9003 22278 9055 22330
rect 13945 22278 13997 22330
rect 14009 22278 14061 22330
rect 14073 22278 14125 22330
rect 14137 22278 14189 22330
rect 14201 22278 14253 22330
rect 19143 22278 19195 22330
rect 19207 22278 19259 22330
rect 19271 22278 19323 22330
rect 19335 22278 19387 22330
rect 19399 22278 19451 22330
rect 4160 22176 4212 22228
rect 4620 22176 4672 22228
rect 7380 22176 7432 22228
rect 8208 22176 8260 22228
rect 1952 22108 2004 22160
rect 2412 22108 2464 22160
rect 480 22040 532 22092
rect 664 22040 716 22092
rect 1400 22083 1452 22092
rect 1400 22049 1409 22083
rect 1409 22049 1443 22083
rect 1443 22049 1452 22083
rect 1400 22040 1452 22049
rect 3332 22108 3384 22160
rect 4252 22108 4304 22160
rect 4804 22108 4856 22160
rect 6368 22151 6420 22160
rect 6368 22117 6377 22151
rect 6377 22117 6411 22151
rect 6411 22117 6420 22151
rect 6368 22108 6420 22117
rect 7288 22108 7340 22160
rect 8576 22108 8628 22160
rect 1216 21972 1268 22024
rect 1676 22015 1728 22024
rect 1676 21981 1685 22015
rect 1685 21981 1719 22015
rect 1719 21981 1728 22015
rect 1676 21972 1728 21981
rect 2320 22015 2372 22024
rect 2320 21981 2329 22015
rect 2329 21981 2363 22015
rect 2363 21981 2372 22015
rect 2320 21972 2372 21981
rect 4620 21972 4672 22024
rect 4896 22040 4948 22092
rect 6460 22040 6512 22092
rect 8668 22040 8720 22092
rect 10048 22176 10100 22228
rect 9864 22108 9916 22160
rect 10876 22176 10928 22228
rect 11060 22176 11112 22228
rect 12072 22176 12124 22228
rect 12624 22108 12676 22160
rect 10600 22083 10652 22092
rect 10600 22049 10609 22083
rect 10609 22049 10643 22083
rect 10643 22049 10652 22083
rect 10600 22040 10652 22049
rect 11704 22040 11756 22092
rect 13820 22176 13872 22228
rect 14188 22176 14240 22228
rect 14372 22176 14424 22228
rect 14740 22176 14792 22228
rect 15200 22176 15252 22228
rect 15568 22108 15620 22160
rect 15936 22108 15988 22160
rect 13268 22083 13320 22092
rect 13268 22049 13277 22083
rect 13277 22049 13311 22083
rect 13311 22049 13320 22083
rect 13268 22040 13320 22049
rect 13820 22040 13872 22092
rect 15384 22083 15436 22092
rect 15384 22049 15393 22083
rect 15393 22049 15427 22083
rect 15427 22049 15436 22083
rect 15384 22040 15436 22049
rect 17408 22176 17460 22228
rect 19432 22176 19484 22228
rect 20352 22176 20404 22228
rect 21456 22219 21508 22228
rect 21456 22185 21465 22219
rect 21465 22185 21499 22219
rect 21499 22185 21508 22219
rect 21456 22176 21508 22185
rect 22928 22176 22980 22228
rect 4988 21972 5040 22024
rect 5356 22015 5408 22024
rect 5356 21981 5365 22015
rect 5365 21981 5399 22015
rect 5399 21981 5408 22015
rect 5356 21972 5408 21981
rect 756 21904 808 21956
rect 2688 21836 2740 21888
rect 2872 21836 2924 21888
rect 3240 21836 3292 21888
rect 4988 21836 5040 21888
rect 5356 21836 5408 21888
rect 7748 21972 7800 22024
rect 7932 22015 7984 22024
rect 7932 21981 7941 22015
rect 7941 21981 7975 22015
rect 7975 21981 7984 22015
rect 7932 21972 7984 21981
rect 8300 21972 8352 22024
rect 8392 21972 8444 22024
rect 9772 21972 9824 22024
rect 10324 21972 10376 22024
rect 12256 22015 12308 22024
rect 12256 21981 12265 22015
rect 12265 21981 12299 22015
rect 12299 21981 12308 22015
rect 12256 21972 12308 21981
rect 13084 22015 13136 22024
rect 13084 21981 13118 22015
rect 13118 21981 13136 22015
rect 13084 21972 13136 21981
rect 5632 21836 5684 21888
rect 6736 21904 6788 21956
rect 8024 21904 8076 21956
rect 8668 21904 8720 21956
rect 15200 21972 15252 22024
rect 11704 21836 11756 21888
rect 16304 22015 16356 22024
rect 16304 21981 16313 22015
rect 16313 21981 16347 22015
rect 16347 21981 16356 22015
rect 16304 21972 16356 21981
rect 14372 21836 14424 21888
rect 17040 21836 17092 21888
rect 18328 21972 18380 22024
rect 18972 21972 19024 22024
rect 21456 22040 21508 22092
rect 21272 22015 21324 22024
rect 21272 21981 21281 22015
rect 21281 21981 21315 22015
rect 21315 21981 21324 22015
rect 21272 21972 21324 21981
rect 21364 21972 21416 22024
rect 21548 21972 21600 22024
rect 22192 21972 22244 22024
rect 17684 21904 17736 21956
rect 20076 21904 20128 21956
rect 20996 21836 21048 21888
rect 22192 21836 22244 21888
rect 6148 21734 6200 21786
rect 6212 21734 6264 21786
rect 6276 21734 6328 21786
rect 6340 21734 6392 21786
rect 6404 21734 6456 21786
rect 11346 21734 11398 21786
rect 11410 21734 11462 21786
rect 11474 21734 11526 21786
rect 11538 21734 11590 21786
rect 11602 21734 11654 21786
rect 16544 21734 16596 21786
rect 16608 21734 16660 21786
rect 16672 21734 16724 21786
rect 16736 21734 16788 21786
rect 16800 21734 16852 21786
rect 21742 21734 21794 21786
rect 21806 21734 21858 21786
rect 21870 21734 21922 21786
rect 21934 21734 21986 21786
rect 21998 21734 22050 21786
rect 1676 21496 1728 21548
rect 3424 21632 3476 21684
rect 3884 21675 3936 21684
rect 3884 21641 3893 21675
rect 3893 21641 3927 21675
rect 3927 21641 3936 21675
rect 3884 21632 3936 21641
rect 4528 21632 4580 21684
rect 5632 21632 5684 21684
rect 5724 21632 5776 21684
rect 7748 21632 7800 21684
rect 9496 21632 9548 21684
rect 9956 21632 10008 21684
rect 10232 21675 10284 21684
rect 10232 21641 10241 21675
rect 10241 21641 10275 21675
rect 10275 21641 10284 21675
rect 10232 21632 10284 21641
rect 12624 21632 12676 21684
rect 12716 21632 12768 21684
rect 12900 21632 12952 21684
rect 13084 21632 13136 21684
rect 15200 21632 15252 21684
rect 3056 21496 3108 21548
rect 4068 21496 4120 21548
rect 1216 21428 1268 21480
rect 4344 21564 4396 21616
rect 9036 21564 9088 21616
rect 9128 21607 9180 21616
rect 9128 21573 9137 21607
rect 9137 21573 9171 21607
rect 9171 21573 9180 21607
rect 9128 21564 9180 21573
rect 9772 21564 9824 21616
rect 11060 21564 11112 21616
rect 4896 21496 4948 21548
rect 7380 21496 7432 21548
rect 9404 21539 9456 21548
rect 9404 21505 9413 21539
rect 9413 21505 9447 21539
rect 9447 21505 9456 21539
rect 9404 21496 9456 21505
rect 11244 21496 11296 21548
rect 12072 21539 12124 21548
rect 12072 21505 12081 21539
rect 12081 21505 12115 21539
rect 12115 21505 12124 21539
rect 12072 21496 12124 21505
rect 13636 21564 13688 21616
rect 13452 21496 13504 21548
rect 15200 21496 15252 21548
rect 20076 21564 20128 21616
rect 20628 21564 20680 21616
rect 17592 21539 17644 21548
rect 17592 21505 17601 21539
rect 17601 21505 17635 21539
rect 17635 21505 17644 21539
rect 17592 21496 17644 21505
rect 19432 21496 19484 21548
rect 20904 21496 20956 21548
rect 204 21292 256 21344
rect 2412 21292 2464 21344
rect 3884 21292 3936 21344
rect 4252 21292 4304 21344
rect 6920 21428 6972 21480
rect 7564 21471 7616 21480
rect 7564 21437 7573 21471
rect 7573 21437 7607 21471
rect 7607 21437 7616 21471
rect 7564 21428 7616 21437
rect 5632 21292 5684 21344
rect 5908 21292 5960 21344
rect 6184 21292 6236 21344
rect 6736 21292 6788 21344
rect 11612 21428 11664 21480
rect 13268 21360 13320 21412
rect 13452 21360 13504 21412
rect 16212 21428 16264 21480
rect 16856 21471 16908 21480
rect 16856 21437 16865 21471
rect 16865 21437 16899 21471
rect 16899 21437 16908 21471
rect 16856 21428 16908 21437
rect 14464 21360 14516 21412
rect 15384 21360 15436 21412
rect 17868 21471 17920 21480
rect 17868 21437 17877 21471
rect 17877 21437 17911 21471
rect 17911 21437 17920 21471
rect 17868 21428 17920 21437
rect 19524 21428 19576 21480
rect 17408 21360 17460 21412
rect 21364 21428 21416 21480
rect 7932 21292 7984 21344
rect 10324 21292 10376 21344
rect 12992 21335 13044 21344
rect 12992 21301 13001 21335
rect 13001 21301 13035 21335
rect 13035 21301 13044 21335
rect 12992 21292 13044 21301
rect 13728 21292 13780 21344
rect 14280 21292 14332 21344
rect 15752 21292 15804 21344
rect 17592 21292 17644 21344
rect 19064 21292 19116 21344
rect 20076 21292 20128 21344
rect 20352 21292 20404 21344
rect 20536 21292 20588 21344
rect 21180 21335 21232 21344
rect 21180 21301 21189 21335
rect 21189 21301 21223 21335
rect 21223 21301 21232 21335
rect 21180 21292 21232 21301
rect 21272 21292 21324 21344
rect 3549 21190 3601 21242
rect 3613 21190 3665 21242
rect 3677 21190 3729 21242
rect 3741 21190 3793 21242
rect 3805 21190 3857 21242
rect 8747 21190 8799 21242
rect 8811 21190 8863 21242
rect 8875 21190 8927 21242
rect 8939 21190 8991 21242
rect 9003 21190 9055 21242
rect 13945 21190 13997 21242
rect 14009 21190 14061 21242
rect 14073 21190 14125 21242
rect 14137 21190 14189 21242
rect 14201 21190 14253 21242
rect 19143 21190 19195 21242
rect 19207 21190 19259 21242
rect 19271 21190 19323 21242
rect 19335 21190 19387 21242
rect 19399 21190 19451 21242
rect 2044 21088 2096 21140
rect 756 20952 808 21004
rect 2228 21020 2280 21072
rect 3148 21088 3200 21140
rect 4528 21088 4580 21140
rect 6184 21088 6236 21140
rect 8116 21088 8168 21140
rect 9036 21088 9088 21140
rect 9220 21088 9272 21140
rect 9772 21088 9824 21140
rect 11244 21088 11296 21140
rect 12072 21088 12124 21140
rect 12624 21088 12676 21140
rect 5448 20952 5500 21004
rect 15016 21020 15068 21072
rect 15568 21020 15620 21072
rect 16120 21020 16172 21072
rect 17408 21088 17460 21140
rect 20536 21088 20588 21140
rect 20812 21088 20864 21140
rect 18788 21020 18840 21072
rect 1952 20884 2004 20936
rect 2504 20884 2556 20936
rect 1308 20816 1360 20868
rect 4252 20884 4304 20936
rect 5724 20884 5776 20936
rect 2964 20816 3016 20868
rect 4436 20816 4488 20868
rect 5908 20884 5960 20936
rect 6736 20884 6788 20936
rect 7748 20952 7800 21004
rect 10048 20952 10100 21004
rect 10508 20952 10560 21004
rect 13360 20952 13412 21004
rect 13820 20952 13872 21004
rect 14096 20995 14148 21004
rect 14096 20961 14105 20995
rect 14105 20961 14139 20995
rect 14139 20961 14148 20995
rect 14096 20952 14148 20961
rect 7932 20884 7984 20936
rect 2136 20748 2188 20800
rect 2504 20748 2556 20800
rect 2688 20748 2740 20800
rect 3424 20748 3476 20800
rect 4528 20748 4580 20800
rect 4896 20748 4948 20800
rect 5172 20748 5224 20800
rect 6184 20791 6236 20800
rect 6184 20757 6193 20791
rect 6193 20757 6227 20791
rect 6227 20757 6236 20791
rect 6184 20748 6236 20757
rect 6828 20816 6880 20868
rect 9128 20884 9180 20936
rect 9588 20884 9640 20936
rect 10600 20884 10652 20936
rect 7104 20748 7156 20800
rect 9496 20748 9548 20800
rect 10324 20748 10376 20800
rect 11428 20884 11480 20936
rect 12624 20884 12676 20936
rect 11796 20816 11848 20868
rect 16028 20927 16080 20936
rect 16028 20893 16037 20927
rect 16037 20893 16071 20927
rect 16071 20893 16080 20927
rect 16028 20884 16080 20893
rect 13912 20748 13964 20800
rect 16212 20884 16264 20936
rect 14924 20748 14976 20800
rect 15844 20791 15896 20800
rect 15844 20757 15853 20791
rect 15853 20757 15887 20791
rect 15887 20757 15896 20791
rect 15844 20748 15896 20757
rect 16120 20748 16172 20800
rect 16304 20791 16356 20800
rect 16304 20757 16313 20791
rect 16313 20757 16347 20791
rect 16347 20757 16356 20791
rect 16304 20748 16356 20757
rect 18604 20952 18656 21004
rect 20352 20952 20404 21004
rect 22652 20952 22704 21004
rect 17040 20884 17092 20936
rect 17960 20884 18012 20936
rect 21272 20884 21324 20936
rect 17224 20816 17276 20868
rect 18880 20816 18932 20868
rect 20628 20816 20680 20868
rect 17592 20748 17644 20800
rect 22192 20816 22244 20868
rect 21456 20748 21508 20800
rect 6148 20646 6200 20698
rect 6212 20646 6264 20698
rect 6276 20646 6328 20698
rect 6340 20646 6392 20698
rect 6404 20646 6456 20698
rect 11346 20646 11398 20698
rect 11410 20646 11462 20698
rect 11474 20646 11526 20698
rect 11538 20646 11590 20698
rect 11602 20646 11654 20698
rect 16544 20646 16596 20698
rect 16608 20646 16660 20698
rect 16672 20646 16724 20698
rect 16736 20646 16788 20698
rect 16800 20646 16852 20698
rect 21742 20646 21794 20698
rect 21806 20646 21858 20698
rect 21870 20646 21922 20698
rect 21934 20646 21986 20698
rect 21998 20646 22050 20698
rect 22928 20612 22980 20664
rect 940 20544 992 20596
rect 1308 20544 1360 20596
rect 2320 20587 2372 20596
rect 2320 20553 2329 20587
rect 2329 20553 2363 20587
rect 2363 20553 2372 20587
rect 2320 20544 2372 20553
rect 1492 20408 1544 20460
rect 2504 20476 2556 20528
rect 3148 20476 3200 20528
rect 3332 20476 3384 20528
rect 4160 20544 4212 20596
rect 4344 20544 4396 20596
rect 4528 20544 4580 20596
rect 6828 20544 6880 20596
rect 6460 20476 6512 20528
rect 6552 20476 6604 20528
rect 6736 20476 6788 20528
rect 2688 20451 2740 20460
rect 2688 20417 2697 20451
rect 2697 20417 2731 20451
rect 2731 20417 2740 20451
rect 2688 20408 2740 20417
rect 2872 20408 2924 20460
rect 4436 20408 4488 20460
rect 4528 20408 4580 20460
rect 5448 20408 5500 20460
rect 7932 20544 7984 20596
rect 8024 20544 8076 20596
rect 7656 20476 7708 20528
rect 7840 20519 7892 20528
rect 7840 20485 7849 20519
rect 7849 20485 7883 20519
rect 7883 20485 7892 20519
rect 7840 20476 7892 20485
rect 8300 20519 8352 20528
rect 8300 20485 8309 20519
rect 8309 20485 8343 20519
rect 8343 20485 8352 20519
rect 8300 20476 8352 20485
rect 8576 20544 8628 20596
rect 9404 20544 9456 20596
rect 9220 20476 9272 20528
rect 7932 20451 7984 20460
rect 7932 20417 7941 20451
rect 7941 20417 7975 20451
rect 7975 20417 7984 20451
rect 7932 20408 7984 20417
rect 12900 20544 12952 20596
rect 13084 20544 13136 20596
rect 13176 20544 13228 20596
rect 14096 20544 14148 20596
rect 10324 20451 10376 20460
rect 10324 20417 10331 20451
rect 10331 20417 10365 20451
rect 10365 20417 10376 20451
rect 10324 20408 10376 20417
rect 11428 20408 11480 20460
rect 12808 20408 12860 20460
rect 12900 20408 12952 20460
rect 15568 20544 15620 20596
rect 15660 20476 15712 20528
rect 15200 20408 15252 20460
rect 17868 20544 17920 20596
rect 20812 20544 20864 20596
rect 21180 20544 21232 20596
rect 15936 20476 15988 20528
rect 2504 20340 2556 20392
rect 3884 20340 3936 20392
rect 5356 20340 5408 20392
rect 6920 20340 6972 20392
rect 7012 20340 7064 20392
rect 7104 20340 7156 20392
rect 11520 20383 11572 20392
rect 1584 20315 1636 20324
rect 1584 20281 1593 20315
rect 1593 20281 1627 20315
rect 1627 20281 1636 20315
rect 1584 20272 1636 20281
rect 5724 20272 5776 20324
rect 6460 20272 6512 20324
rect 6552 20272 6604 20324
rect 3516 20204 3568 20256
rect 5264 20247 5316 20256
rect 5264 20213 5273 20247
rect 5273 20213 5307 20247
rect 5307 20213 5316 20247
rect 5264 20204 5316 20213
rect 6644 20247 6696 20256
rect 6644 20213 6653 20247
rect 6653 20213 6687 20247
rect 6687 20213 6696 20247
rect 6644 20204 6696 20213
rect 9128 20204 9180 20256
rect 9864 20204 9916 20256
rect 11520 20349 11529 20383
rect 11529 20349 11563 20383
rect 11563 20349 11572 20383
rect 11520 20340 11572 20349
rect 13176 20340 13228 20392
rect 10968 20272 11020 20324
rect 11336 20272 11388 20324
rect 14142 20383 14194 20392
rect 14142 20349 14151 20383
rect 14151 20349 14185 20383
rect 14185 20349 14194 20383
rect 14142 20340 14194 20349
rect 14924 20340 14976 20392
rect 11060 20247 11112 20256
rect 11060 20213 11069 20247
rect 11069 20213 11103 20247
rect 11103 20213 11112 20247
rect 11060 20204 11112 20213
rect 11244 20204 11296 20256
rect 13728 20315 13780 20324
rect 13728 20281 13737 20315
rect 13737 20281 13771 20315
rect 13771 20281 13780 20315
rect 13728 20272 13780 20281
rect 12624 20204 12676 20256
rect 15384 20204 15436 20256
rect 16120 20204 16172 20256
rect 17592 20340 17644 20392
rect 20168 20408 20220 20460
rect 20996 20408 21048 20460
rect 19524 20383 19576 20392
rect 19524 20349 19533 20383
rect 19533 20349 19567 20383
rect 19567 20349 19576 20383
rect 19524 20340 19576 20349
rect 19984 20204 20036 20256
rect 20536 20247 20588 20256
rect 20536 20213 20545 20247
rect 20545 20213 20579 20247
rect 20579 20213 20588 20247
rect 20536 20204 20588 20213
rect 21180 20204 21232 20256
rect 21456 20247 21508 20256
rect 21456 20213 21465 20247
rect 21465 20213 21499 20247
rect 21499 20213 21508 20247
rect 21456 20204 21508 20213
rect 3549 20102 3601 20154
rect 3613 20102 3665 20154
rect 3677 20102 3729 20154
rect 3741 20102 3793 20154
rect 3805 20102 3857 20154
rect 8747 20102 8799 20154
rect 8811 20102 8863 20154
rect 8875 20102 8927 20154
rect 8939 20102 8991 20154
rect 9003 20102 9055 20154
rect 13945 20102 13997 20154
rect 14009 20102 14061 20154
rect 14073 20102 14125 20154
rect 14137 20102 14189 20154
rect 14201 20102 14253 20154
rect 19143 20102 19195 20154
rect 19207 20102 19259 20154
rect 19271 20102 19323 20154
rect 19335 20102 19387 20154
rect 19399 20102 19451 20154
rect 756 20000 808 20052
rect 1768 20000 1820 20052
rect 2780 20000 2832 20052
rect 2044 19975 2096 19984
rect 2044 19941 2053 19975
rect 2053 19941 2087 19975
rect 2087 19941 2096 19975
rect 2044 19932 2096 19941
rect 4436 20000 4488 20052
rect 5356 20000 5408 20052
rect 5724 20000 5776 20052
rect 6092 20000 6144 20052
rect 8208 20000 8260 20052
rect 8668 20000 8720 20052
rect 11152 20000 11204 20052
rect 11336 20000 11388 20052
rect 11520 20000 11572 20052
rect 1216 19864 1268 19916
rect 2320 19907 2372 19916
rect 2320 19873 2329 19907
rect 2329 19873 2363 19907
rect 2363 19873 2372 19907
rect 2320 19864 2372 19873
rect 3240 19864 3292 19916
rect 4528 19907 4580 19916
rect 4528 19873 4537 19907
rect 4537 19873 4571 19907
rect 4571 19873 4580 19907
rect 4528 19864 4580 19873
rect 10416 19864 10468 19916
rect 11060 19864 11112 19916
rect 756 19796 808 19848
rect 1768 19796 1820 19848
rect 1860 19771 1912 19780
rect 1860 19737 1869 19771
rect 1869 19737 1903 19771
rect 1903 19737 1912 19771
rect 1860 19728 1912 19737
rect 2320 19728 2372 19780
rect 2780 19728 2832 19780
rect 4436 19796 4488 19848
rect 6644 19796 6696 19848
rect 6920 19796 6972 19848
rect 10140 19796 10192 19848
rect 13360 20000 13412 20052
rect 15384 20000 15436 20052
rect 13728 19932 13780 19984
rect 14464 19864 14516 19916
rect 14648 19864 14700 19916
rect 14832 19864 14884 19916
rect 15108 19907 15160 19916
rect 15108 19873 15142 19907
rect 15142 19873 15160 19907
rect 15108 19864 15160 19873
rect 16028 20000 16080 20052
rect 19984 20000 20036 20052
rect 16948 19864 17000 19916
rect 17316 19864 17368 19916
rect 20352 19864 20404 19916
rect 12072 19796 12124 19848
rect 756 19660 808 19712
rect 3056 19660 3108 19712
rect 3148 19660 3200 19712
rect 6184 19728 6236 19780
rect 4988 19660 5040 19712
rect 9680 19660 9732 19712
rect 10692 19771 10744 19780
rect 10692 19737 10701 19771
rect 10701 19737 10735 19771
rect 10735 19737 10744 19771
rect 10692 19728 10744 19737
rect 11704 19771 11756 19780
rect 11704 19737 11713 19771
rect 11713 19737 11747 19771
rect 11747 19737 11756 19771
rect 11704 19728 11756 19737
rect 14280 19839 14332 19848
rect 14280 19805 14289 19839
rect 14289 19805 14323 19839
rect 14323 19805 14332 19839
rect 14280 19796 14332 19805
rect 16764 19796 16816 19848
rect 13084 19728 13136 19780
rect 13728 19728 13780 19780
rect 11060 19703 11112 19712
rect 11060 19669 11069 19703
rect 11069 19669 11103 19703
rect 11103 19669 11112 19703
rect 11060 19660 11112 19669
rect 11152 19660 11204 19712
rect 11796 19660 11848 19712
rect 12440 19660 12492 19712
rect 12716 19660 12768 19712
rect 16028 19728 16080 19780
rect 17132 19796 17184 19848
rect 18420 19796 18472 19848
rect 18972 19796 19024 19848
rect 19064 19839 19116 19848
rect 19064 19805 19073 19839
rect 19073 19805 19107 19839
rect 19107 19805 19116 19839
rect 19064 19796 19116 19805
rect 20904 19839 20956 19848
rect 20904 19805 20913 19839
rect 20913 19805 20947 19839
rect 20947 19805 20956 19839
rect 20904 19796 20956 19805
rect 21180 19796 21232 19848
rect 21364 19796 21416 19848
rect 17316 19771 17368 19780
rect 15752 19660 15804 19712
rect 17316 19737 17325 19771
rect 17325 19737 17359 19771
rect 17359 19737 17368 19771
rect 17316 19728 17368 19737
rect 17132 19660 17184 19712
rect 19616 19728 19668 19780
rect 20168 19728 20220 19780
rect 20444 19728 20496 19780
rect 18880 19703 18932 19712
rect 18880 19669 18889 19703
rect 18889 19669 18923 19703
rect 18923 19669 18932 19703
rect 18880 19660 18932 19669
rect 22192 19660 22244 19712
rect 664 19524 716 19576
rect 6148 19558 6200 19610
rect 6212 19558 6264 19610
rect 6276 19558 6328 19610
rect 6340 19558 6392 19610
rect 6404 19558 6456 19610
rect 11346 19558 11398 19610
rect 11410 19558 11462 19610
rect 11474 19558 11526 19610
rect 11538 19558 11590 19610
rect 11602 19558 11654 19610
rect 16544 19558 16596 19610
rect 16608 19558 16660 19610
rect 16672 19558 16724 19610
rect 16736 19558 16788 19610
rect 16800 19558 16852 19610
rect 21742 19558 21794 19610
rect 21806 19558 21858 19610
rect 21870 19558 21922 19610
rect 21934 19558 21986 19610
rect 21998 19558 22050 19610
rect 2504 19499 2556 19508
rect 2504 19465 2513 19499
rect 2513 19465 2547 19499
rect 2547 19465 2556 19499
rect 2504 19456 2556 19465
rect 1952 19388 2004 19440
rect 2596 19320 2648 19372
rect 2688 19320 2740 19372
rect 2872 19363 2924 19372
rect 2872 19329 2881 19363
rect 2881 19329 2915 19363
rect 2915 19329 2924 19363
rect 2872 19320 2924 19329
rect 3332 19320 3384 19372
rect 4436 19388 4488 19440
rect 4252 19320 4304 19372
rect 5356 19388 5408 19440
rect 5908 19499 5960 19508
rect 5908 19465 5917 19499
rect 5917 19465 5951 19499
rect 5951 19465 5960 19499
rect 5908 19456 5960 19465
rect 6552 19456 6604 19508
rect 7012 19456 7064 19508
rect 7932 19456 7984 19508
rect 9680 19456 9732 19508
rect 9772 19388 9824 19440
rect 11428 19456 11480 19508
rect 11888 19456 11940 19508
rect 12440 19456 12492 19508
rect 11060 19388 11112 19440
rect 5540 19320 5592 19372
rect 8208 19320 8260 19372
rect 9864 19320 9916 19372
rect 10692 19320 10744 19372
rect 4344 19184 4396 19236
rect 4804 19184 4856 19236
rect 11888 19320 11940 19372
rect 12072 19320 12124 19372
rect 13544 19320 13596 19372
rect 15936 19456 15988 19508
rect 16856 19456 16908 19508
rect 17132 19456 17184 19508
rect 14648 19363 14700 19372
rect 14648 19329 14655 19363
rect 14655 19329 14689 19363
rect 14689 19329 14700 19363
rect 14648 19320 14700 19329
rect 15384 19320 15436 19372
rect 16120 19363 16172 19372
rect 16120 19329 16129 19363
rect 16129 19329 16163 19363
rect 16163 19329 16172 19363
rect 16120 19320 16172 19329
rect 16304 19431 16356 19440
rect 16304 19397 16313 19431
rect 16313 19397 16347 19431
rect 16347 19397 16356 19431
rect 16304 19388 16356 19397
rect 17592 19388 17644 19440
rect 18420 19388 18472 19440
rect 13360 19295 13412 19304
rect 13360 19261 13369 19295
rect 13369 19261 13403 19295
rect 13403 19261 13412 19295
rect 13360 19252 13412 19261
rect 4620 19116 4672 19168
rect 8300 19184 8352 19236
rect 9772 19184 9824 19236
rect 5356 19116 5408 19168
rect 6920 19116 6972 19168
rect 7564 19116 7616 19168
rect 8668 19116 8720 19168
rect 9588 19116 9640 19168
rect 11796 19184 11848 19236
rect 12072 19184 12124 19236
rect 13084 19227 13136 19236
rect 13084 19193 13093 19227
rect 13093 19193 13127 19227
rect 13127 19193 13136 19227
rect 13084 19184 13136 19193
rect 15200 19252 15252 19304
rect 16856 19320 16908 19372
rect 12440 19116 12492 19168
rect 14280 19159 14332 19168
rect 14280 19125 14289 19159
rect 14289 19125 14323 19159
rect 14323 19125 14332 19159
rect 14280 19116 14332 19125
rect 15108 19184 15160 19236
rect 15844 19184 15896 19236
rect 16304 19116 16356 19168
rect 18604 19320 18656 19372
rect 18880 19320 18932 19372
rect 20628 19320 20680 19372
rect 21180 19363 21232 19372
rect 21180 19329 21189 19363
rect 21189 19329 21223 19363
rect 21223 19329 21232 19363
rect 21180 19320 21232 19329
rect 18972 19252 19024 19304
rect 20444 19159 20496 19168
rect 20444 19125 20453 19159
rect 20453 19125 20487 19159
rect 20487 19125 20496 19159
rect 20444 19116 20496 19125
rect 20720 19159 20772 19168
rect 20720 19125 20729 19159
rect 20729 19125 20763 19159
rect 20763 19125 20772 19159
rect 20720 19116 20772 19125
rect 20996 19116 21048 19168
rect 21456 19159 21508 19168
rect 21456 19125 21465 19159
rect 21465 19125 21499 19159
rect 21499 19125 21508 19159
rect 21456 19116 21508 19125
rect 3549 19014 3601 19066
rect 3613 19014 3665 19066
rect 3677 19014 3729 19066
rect 3741 19014 3793 19066
rect 3805 19014 3857 19066
rect 8747 19014 8799 19066
rect 8811 19014 8863 19066
rect 8875 19014 8927 19066
rect 8939 19014 8991 19066
rect 9003 19014 9055 19066
rect 13945 19014 13997 19066
rect 14009 19014 14061 19066
rect 14073 19014 14125 19066
rect 14137 19014 14189 19066
rect 14201 19014 14253 19066
rect 19143 19014 19195 19066
rect 19207 19014 19259 19066
rect 19271 19014 19323 19066
rect 19335 19014 19387 19066
rect 19399 19014 19451 19066
rect 1032 18912 1084 18964
rect 4528 18912 4580 18964
rect 1492 18776 1544 18828
rect 1676 18819 1728 18828
rect 1676 18785 1685 18819
rect 1685 18785 1719 18819
rect 1719 18785 1728 18819
rect 1676 18776 1728 18785
rect 2320 18819 2372 18828
rect 2320 18785 2329 18819
rect 2329 18785 2363 18819
rect 2363 18785 2372 18819
rect 2320 18776 2372 18785
rect 3240 18776 3292 18828
rect 4068 18819 4120 18828
rect 4068 18785 4077 18819
rect 4077 18785 4111 18819
rect 4111 18785 4120 18819
rect 4068 18776 4120 18785
rect 5448 18912 5500 18964
rect 5724 18955 5776 18964
rect 5724 18921 5733 18955
rect 5733 18921 5767 18955
rect 5767 18921 5776 18955
rect 5724 18912 5776 18921
rect 7104 18955 7156 18964
rect 7104 18921 7113 18955
rect 7113 18921 7147 18955
rect 7147 18921 7156 18955
rect 7104 18912 7156 18921
rect 9772 18912 9824 18964
rect 10416 18955 10468 18964
rect 10416 18921 10425 18955
rect 10425 18921 10459 18955
rect 10459 18921 10468 18955
rect 10416 18912 10468 18921
rect 7288 18844 7340 18896
rect 12624 18912 12676 18964
rect 12808 18912 12860 18964
rect 13360 18912 13412 18964
rect 15200 18912 15252 18964
rect 15384 18955 15436 18964
rect 15384 18921 15393 18955
rect 15393 18921 15427 18955
rect 15427 18921 15436 18955
rect 15384 18912 15436 18921
rect 16120 18912 16172 18964
rect 14648 18844 14700 18896
rect 16948 18912 17000 18964
rect 5540 18776 5592 18828
rect 2228 18708 2280 18760
rect 2596 18751 2648 18760
rect 2596 18717 2605 18751
rect 2605 18717 2648 18751
rect 2596 18708 2648 18717
rect 4620 18640 4672 18692
rect 4804 18640 4856 18692
rect 5264 18640 5316 18692
rect 7104 18640 7156 18692
rect 7564 18640 7616 18692
rect 7840 18640 7892 18692
rect 3332 18615 3384 18624
rect 3332 18581 3341 18615
rect 3341 18581 3375 18615
rect 3375 18581 3384 18615
rect 3332 18572 3384 18581
rect 4896 18572 4948 18624
rect 5356 18572 5408 18624
rect 5448 18572 5500 18624
rect 8852 18708 8904 18760
rect 8300 18640 8352 18692
rect 8208 18572 8260 18624
rect 8392 18572 8444 18624
rect 9404 18819 9456 18828
rect 9404 18785 9413 18819
rect 9413 18785 9447 18819
rect 9447 18785 9456 18819
rect 9404 18776 9456 18785
rect 10140 18776 10192 18828
rect 11060 18819 11112 18828
rect 11060 18785 11069 18819
rect 11069 18785 11103 18819
rect 11103 18785 11112 18819
rect 11060 18776 11112 18785
rect 11612 18776 11664 18828
rect 12072 18819 12124 18828
rect 12072 18785 12106 18819
rect 12106 18785 12124 18819
rect 12072 18776 12124 18785
rect 12440 18776 12492 18828
rect 15108 18776 15160 18828
rect 9956 18640 10008 18692
rect 11428 18708 11480 18760
rect 15200 18708 15252 18760
rect 16948 18708 17000 18760
rect 17408 18819 17460 18828
rect 17408 18785 17417 18819
rect 17417 18785 17451 18819
rect 17451 18785 17460 18819
rect 17408 18776 17460 18785
rect 19524 18912 19576 18964
rect 19708 18912 19760 18964
rect 20536 18912 20588 18964
rect 21180 18912 21232 18964
rect 20352 18844 20404 18896
rect 17776 18708 17828 18760
rect 11152 18572 11204 18624
rect 17960 18640 18012 18692
rect 19616 18708 19668 18760
rect 20536 18640 20588 18692
rect 22744 18708 22796 18760
rect 22652 18640 22704 18692
rect 14280 18572 14332 18624
rect 19524 18572 19576 18624
rect 20628 18572 20680 18624
rect 22192 18572 22244 18624
rect 6148 18470 6200 18522
rect 6212 18470 6264 18522
rect 6276 18470 6328 18522
rect 6340 18470 6392 18522
rect 6404 18470 6456 18522
rect 11346 18470 11398 18522
rect 11410 18470 11462 18522
rect 11474 18470 11526 18522
rect 11538 18470 11590 18522
rect 11602 18470 11654 18522
rect 16544 18470 16596 18522
rect 16608 18470 16660 18522
rect 16672 18470 16724 18522
rect 16736 18470 16788 18522
rect 16800 18470 16852 18522
rect 21742 18470 21794 18522
rect 21806 18470 21858 18522
rect 21870 18470 21922 18522
rect 21934 18470 21986 18522
rect 21998 18470 22050 18522
rect 22652 18436 22704 18488
rect 3148 18368 3200 18420
rect 6736 18368 6788 18420
rect 6920 18368 6972 18420
rect 7564 18368 7616 18420
rect 7932 18368 7984 18420
rect 8300 18368 8352 18420
rect 940 18300 992 18352
rect 2964 18300 3016 18352
rect 8116 18300 8168 18352
rect 8852 18300 8904 18352
rect 9220 18368 9272 18420
rect 10600 18368 10652 18420
rect 12716 18368 12768 18420
rect 13084 18411 13136 18420
rect 13084 18377 13093 18411
rect 13093 18377 13127 18411
rect 13127 18377 13136 18411
rect 13084 18368 13136 18377
rect 13728 18368 13780 18420
rect 10692 18300 10744 18352
rect 10876 18300 10928 18352
rect 1952 18232 2004 18284
rect 2688 18275 2740 18284
rect 2688 18241 2697 18275
rect 2697 18241 2740 18275
rect 2688 18232 2740 18241
rect 4988 18275 5040 18284
rect 4988 18241 4997 18275
rect 4997 18241 5031 18275
rect 5031 18241 5040 18275
rect 4988 18232 5040 18241
rect 7104 18275 7156 18284
rect 7104 18241 7111 18275
rect 7111 18241 7145 18275
rect 7145 18241 7156 18275
rect 7104 18232 7156 18241
rect 7472 18232 7524 18284
rect 7932 18232 7984 18284
rect 9956 18232 10008 18284
rect 10232 18232 10284 18284
rect 15660 18300 15712 18352
rect 16212 18368 16264 18420
rect 20076 18368 20128 18420
rect 20352 18368 20404 18420
rect 20444 18368 20496 18420
rect 20536 18411 20588 18420
rect 20536 18377 20545 18411
rect 20545 18377 20579 18411
rect 20579 18377 20588 18411
rect 20536 18368 20588 18377
rect 20720 18368 20772 18420
rect 13820 18232 13872 18284
rect 16396 18232 16448 18284
rect 17960 18300 18012 18352
rect 19064 18300 19116 18352
rect 2320 18164 2372 18216
rect 3424 18164 3476 18216
rect 4068 18164 4120 18216
rect 4160 18164 4212 18216
rect 3884 18096 3936 18148
rect 1584 18071 1636 18080
rect 1584 18037 1593 18071
rect 1593 18037 1627 18071
rect 1627 18037 1636 18071
rect 1584 18028 1636 18037
rect 2228 18028 2280 18080
rect 3976 18028 4028 18080
rect 4804 18207 4856 18216
rect 4804 18173 4838 18207
rect 4838 18173 4856 18207
rect 4804 18164 4856 18173
rect 5356 18164 5408 18216
rect 5540 18164 5592 18216
rect 8392 18164 8444 18216
rect 10048 18207 10100 18216
rect 10048 18173 10057 18207
rect 10057 18173 10091 18207
rect 10091 18173 10100 18207
rect 10048 18164 10100 18173
rect 11796 18164 11848 18216
rect 4804 18028 4856 18080
rect 13084 18164 13136 18216
rect 7288 18028 7340 18080
rect 7840 18071 7892 18080
rect 7840 18037 7849 18071
rect 7849 18037 7883 18071
rect 7883 18037 7892 18071
rect 7840 18028 7892 18037
rect 11060 18071 11112 18080
rect 11060 18037 11069 18071
rect 11069 18037 11103 18071
rect 11103 18037 11112 18071
rect 11060 18028 11112 18037
rect 11152 18028 11204 18080
rect 12808 18028 12860 18080
rect 15384 18164 15436 18216
rect 16672 18207 16724 18216
rect 16672 18173 16681 18207
rect 16681 18173 16715 18207
rect 16715 18173 16724 18207
rect 16672 18164 16724 18173
rect 15200 18096 15252 18148
rect 16396 18096 16448 18148
rect 14740 18028 14792 18080
rect 15292 18028 15344 18080
rect 15752 18028 15804 18080
rect 16212 18028 16264 18080
rect 16580 18028 16632 18080
rect 18972 18028 19024 18080
rect 20720 18028 20772 18080
rect 21456 18071 21508 18080
rect 21456 18037 21465 18071
rect 21465 18037 21499 18071
rect 21499 18037 21508 18071
rect 21456 18028 21508 18037
rect 3549 17926 3601 17978
rect 3613 17926 3665 17978
rect 3677 17926 3729 17978
rect 3741 17926 3793 17978
rect 3805 17926 3857 17978
rect 8747 17926 8799 17978
rect 8811 17926 8863 17978
rect 8875 17926 8927 17978
rect 8939 17926 8991 17978
rect 9003 17926 9055 17978
rect 13945 17926 13997 17978
rect 14009 17926 14061 17978
rect 14073 17926 14125 17978
rect 14137 17926 14189 17978
rect 14201 17926 14253 17978
rect 19143 17926 19195 17978
rect 19207 17926 19259 17978
rect 19271 17926 19323 17978
rect 19335 17926 19387 17978
rect 19399 17926 19451 17978
rect 1768 17824 1820 17876
rect 6092 17824 6144 17876
rect 6184 17824 6236 17876
rect 2504 17756 2556 17808
rect 6736 17799 6788 17808
rect 6736 17765 6745 17799
rect 6745 17765 6779 17799
rect 6779 17765 6788 17799
rect 6736 17756 6788 17765
rect 2044 17688 2096 17740
rect 2412 17731 2464 17740
rect 2412 17697 2421 17731
rect 2421 17697 2455 17731
rect 2455 17697 2464 17731
rect 2412 17688 2464 17697
rect 2688 17731 2740 17740
rect 2688 17697 2697 17731
rect 2697 17697 2731 17731
rect 2731 17697 2740 17731
rect 2688 17688 2740 17697
rect 4068 17688 4120 17740
rect 5724 17731 5776 17740
rect 1676 17620 1728 17672
rect 2136 17620 2188 17672
rect 2964 17663 3016 17672
rect 2964 17629 2973 17663
rect 2973 17629 3007 17663
rect 3007 17629 3016 17663
rect 2964 17620 3016 17629
rect 3700 17620 3752 17672
rect 5724 17697 5733 17731
rect 5733 17697 5767 17731
rect 5767 17697 5776 17731
rect 5724 17688 5776 17697
rect 7012 17688 7064 17740
rect 4252 17620 4304 17672
rect 4712 17620 4764 17672
rect 5908 17620 5960 17672
rect 8576 17824 8628 17876
rect 9956 17867 10008 17876
rect 9956 17833 9965 17867
rect 9965 17833 9999 17867
rect 9999 17833 10008 17867
rect 9956 17824 10008 17833
rect 10048 17824 10100 17876
rect 12072 17824 12124 17876
rect 12900 17824 12952 17876
rect 7196 17688 7248 17740
rect 7472 17620 7524 17672
rect 7564 17620 7616 17672
rect 7840 17620 7892 17672
rect 8116 17663 8168 17672
rect 8116 17629 8125 17663
rect 8125 17629 8159 17663
rect 8159 17629 8168 17663
rect 8116 17620 8168 17629
rect 8300 17620 8352 17672
rect 11796 17688 11848 17740
rect 11980 17688 12032 17740
rect 12624 17731 12676 17740
rect 12624 17697 12633 17731
rect 12633 17697 12667 17731
rect 12667 17697 12676 17731
rect 12624 17688 12676 17697
rect 15936 17824 15988 17876
rect 16120 17824 16172 17876
rect 20904 17824 20956 17876
rect 20996 17867 21048 17876
rect 20996 17833 21005 17867
rect 21005 17833 21039 17867
rect 21039 17833 21048 17867
rect 20996 17824 21048 17833
rect 20812 17756 20864 17808
rect 15292 17731 15344 17740
rect 15292 17697 15301 17731
rect 15301 17697 15335 17731
rect 15335 17697 15344 17731
rect 15292 17688 15344 17697
rect 16212 17688 16264 17740
rect 20628 17731 20680 17740
rect 20628 17697 20637 17731
rect 20637 17697 20671 17731
rect 20671 17697 20680 17731
rect 20628 17688 20680 17697
rect 8944 17663 8996 17672
rect 8944 17629 8953 17663
rect 8953 17629 8987 17663
rect 8987 17629 8996 17663
rect 8944 17620 8996 17629
rect 9220 17663 9272 17672
rect 9220 17629 9227 17663
rect 9227 17629 9261 17663
rect 9261 17629 9272 17663
rect 9220 17620 9272 17629
rect 6828 17552 6880 17604
rect 7012 17552 7064 17604
rect 10600 17620 10652 17672
rect 10692 17663 10744 17672
rect 10692 17629 10701 17663
rect 10701 17629 10735 17663
rect 10735 17629 10744 17663
rect 10692 17620 10744 17629
rect 1676 17484 1728 17536
rect 2596 17484 2648 17536
rect 3056 17484 3108 17536
rect 4620 17527 4672 17536
rect 4620 17493 4629 17527
rect 4629 17493 4663 17527
rect 4663 17493 4672 17527
rect 4620 17484 4672 17493
rect 4988 17484 5040 17536
rect 5908 17484 5960 17536
rect 6092 17484 6144 17536
rect 10416 17552 10468 17604
rect 8116 17484 8168 17536
rect 8760 17484 8812 17536
rect 13360 17620 13412 17672
rect 12624 17552 12676 17604
rect 13084 17552 13136 17604
rect 11704 17527 11756 17536
rect 11704 17493 11713 17527
rect 11713 17493 11747 17527
rect 11747 17493 11756 17527
rect 11704 17484 11756 17493
rect 11888 17484 11940 17536
rect 12072 17484 12124 17536
rect 12440 17484 12492 17536
rect 14464 17620 14516 17672
rect 15108 17663 15160 17672
rect 15108 17629 15142 17663
rect 15142 17629 15160 17663
rect 15108 17620 15160 17629
rect 17040 17620 17092 17672
rect 17960 17663 18012 17672
rect 17960 17629 17967 17663
rect 17967 17629 18001 17663
rect 18001 17629 18012 17663
rect 17960 17620 18012 17629
rect 19064 17620 19116 17672
rect 19524 17620 19576 17672
rect 16028 17552 16080 17604
rect 16580 17595 16632 17604
rect 16580 17561 16589 17595
rect 16589 17561 16623 17595
rect 16623 17561 16632 17595
rect 16580 17552 16632 17561
rect 17776 17552 17828 17604
rect 14832 17484 14884 17536
rect 15292 17484 15344 17536
rect 16120 17484 16172 17536
rect 16672 17484 16724 17536
rect 17224 17484 17276 17536
rect 17316 17527 17368 17536
rect 17316 17493 17325 17527
rect 17325 17493 17359 17527
rect 17359 17493 17368 17527
rect 17316 17484 17368 17493
rect 17500 17527 17552 17536
rect 17500 17493 17509 17527
rect 17509 17493 17543 17527
rect 17543 17493 17552 17527
rect 17500 17484 17552 17493
rect 17868 17484 17920 17536
rect 20536 17620 20588 17672
rect 21272 17663 21324 17672
rect 21272 17629 21281 17663
rect 21281 17629 21315 17663
rect 21315 17629 21324 17663
rect 21272 17620 21324 17629
rect 20352 17484 20404 17536
rect 20904 17484 20956 17536
rect 22192 17484 22244 17536
rect 6148 17382 6200 17434
rect 6212 17382 6264 17434
rect 6276 17382 6328 17434
rect 6340 17382 6392 17434
rect 6404 17382 6456 17434
rect 11346 17382 11398 17434
rect 11410 17382 11462 17434
rect 11474 17382 11526 17434
rect 11538 17382 11590 17434
rect 11602 17382 11654 17434
rect 16544 17382 16596 17434
rect 16608 17382 16660 17434
rect 16672 17382 16724 17434
rect 16736 17382 16788 17434
rect 16800 17382 16852 17434
rect 21742 17382 21794 17434
rect 21806 17382 21858 17434
rect 21870 17382 21922 17434
rect 21934 17382 21986 17434
rect 21998 17382 22050 17434
rect 1768 17280 1820 17332
rect 1584 17255 1636 17264
rect 1584 17221 1593 17255
rect 1593 17221 1627 17255
rect 1627 17221 1636 17255
rect 1584 17212 1636 17221
rect 2688 17280 2740 17332
rect 3884 17280 3936 17332
rect 3976 17280 4028 17332
rect 4988 17280 5040 17332
rect 7472 17280 7524 17332
rect 3700 17212 3752 17264
rect 7012 17212 7064 17264
rect 7564 17255 7616 17264
rect 7564 17221 7573 17255
rect 7573 17221 7607 17255
rect 7607 17221 7616 17255
rect 7564 17212 7616 17221
rect 7840 17280 7892 17332
rect 10232 17280 10284 17332
rect 8116 17212 8168 17264
rect 8576 17212 8628 17264
rect 9772 17212 9824 17264
rect 2596 17144 2648 17196
rect 2780 17144 2832 17196
rect 3332 17076 3384 17128
rect 4988 17187 5040 17196
rect 4988 17153 4997 17187
rect 4997 17153 5031 17187
rect 5031 17153 5040 17187
rect 4988 17144 5040 17153
rect 4712 17119 4764 17128
rect 1860 17008 1912 17060
rect 2320 17008 2372 17060
rect 1216 16940 1268 16992
rect 3792 17008 3844 17060
rect 4344 17008 4396 17060
rect 4712 17085 4721 17119
rect 4721 17085 4755 17119
rect 4755 17085 4764 17119
rect 4712 17076 4764 17085
rect 5540 17076 5592 17128
rect 7472 17187 7524 17196
rect 7472 17153 7481 17187
rect 7481 17153 7515 17187
rect 7515 17153 7524 17187
rect 10968 17212 11020 17264
rect 12992 17280 13044 17332
rect 15016 17323 15068 17332
rect 15016 17289 15025 17323
rect 15025 17289 15059 17323
rect 15059 17289 15068 17323
rect 15016 17280 15068 17289
rect 15292 17280 15344 17332
rect 16212 17323 16264 17332
rect 16212 17289 16221 17323
rect 16221 17289 16255 17323
rect 16255 17289 16264 17323
rect 16212 17280 16264 17289
rect 16856 17280 16908 17332
rect 17316 17280 17368 17332
rect 17684 17280 17736 17332
rect 7472 17144 7524 17153
rect 10600 17144 10652 17196
rect 11244 17144 11296 17196
rect 15660 17212 15712 17264
rect 6000 17076 6052 17128
rect 6552 17076 6604 17128
rect 9864 17076 9916 17128
rect 5448 17008 5500 17060
rect 3424 16940 3476 16992
rect 3976 16940 4028 16992
rect 4068 16940 4120 16992
rect 8944 16940 8996 16992
rect 9496 16940 9548 16992
rect 10876 17076 10928 17128
rect 12808 17051 12860 17060
rect 12808 17017 12817 17051
rect 12817 17017 12851 17051
rect 12851 17017 12860 17051
rect 12808 17008 12860 17017
rect 10416 16940 10468 16992
rect 10692 16940 10744 16992
rect 10968 16983 11020 16992
rect 10968 16949 10977 16983
rect 10977 16949 11011 16983
rect 11011 16949 11020 16983
rect 10968 16940 11020 16949
rect 11152 16940 11204 16992
rect 12440 16940 12492 16992
rect 12624 16940 12676 16992
rect 13268 17076 13320 17128
rect 13360 17119 13412 17128
rect 13360 17085 13369 17119
rect 13369 17085 13403 17119
rect 13403 17085 13412 17119
rect 13360 17076 13412 17085
rect 14740 17076 14792 17128
rect 17592 17187 17644 17196
rect 17592 17153 17601 17187
rect 17601 17153 17635 17187
rect 17635 17153 17644 17187
rect 17592 17144 17644 17153
rect 16856 17119 16908 17128
rect 16856 17085 16865 17119
rect 16865 17085 16899 17119
rect 16899 17085 16908 17119
rect 16856 17076 16908 17085
rect 17684 17119 17736 17128
rect 17684 17085 17718 17119
rect 17718 17085 17736 17119
rect 17684 17076 17736 17085
rect 17866 17119 17918 17128
rect 17866 17085 17875 17119
rect 17875 17085 17909 17119
rect 17909 17085 17918 17119
rect 17866 17076 17918 17085
rect 20904 17280 20956 17332
rect 19524 17187 19576 17196
rect 19524 17153 19558 17187
rect 19558 17153 19576 17187
rect 19524 17144 19576 17153
rect 20720 17144 20772 17196
rect 18972 17076 19024 17128
rect 17316 17051 17368 17060
rect 17316 17017 17325 17051
rect 17325 17017 17359 17051
rect 17359 17017 17368 17051
rect 17316 17008 17368 17017
rect 20352 17008 20404 17060
rect 13544 16940 13596 16992
rect 14280 16940 14332 16992
rect 15292 16940 15344 16992
rect 16212 16940 16264 16992
rect 17040 16940 17092 16992
rect 18512 16983 18564 16992
rect 18512 16949 18521 16983
rect 18521 16949 18555 16983
rect 18555 16949 18564 16983
rect 18512 16940 18564 16949
rect 19524 16940 19576 16992
rect 20168 16940 20220 16992
rect 20536 16940 20588 16992
rect 20628 16940 20680 16992
rect 21456 16983 21508 16992
rect 21456 16949 21465 16983
rect 21465 16949 21499 16983
rect 21499 16949 21508 16983
rect 21456 16940 21508 16949
rect 3549 16838 3601 16890
rect 3613 16838 3665 16890
rect 3677 16838 3729 16890
rect 3741 16838 3793 16890
rect 3805 16838 3857 16890
rect 8747 16838 8799 16890
rect 8811 16838 8863 16890
rect 8875 16838 8927 16890
rect 8939 16838 8991 16890
rect 9003 16838 9055 16890
rect 13945 16838 13997 16890
rect 14009 16838 14061 16890
rect 14073 16838 14125 16890
rect 14137 16838 14189 16890
rect 14201 16838 14253 16890
rect 19143 16838 19195 16890
rect 19207 16838 19259 16890
rect 19271 16838 19323 16890
rect 19335 16838 19387 16890
rect 19399 16838 19451 16890
rect 1952 16736 2004 16788
rect 2964 16736 3016 16788
rect 3608 16736 3660 16788
rect 6736 16736 6788 16788
rect 6828 16779 6880 16788
rect 6828 16745 6837 16779
rect 6837 16745 6871 16779
rect 6871 16745 6880 16779
rect 6828 16736 6880 16745
rect 7564 16736 7616 16788
rect 3976 16600 4028 16652
rect 4896 16600 4948 16652
rect 2228 16532 2280 16584
rect 2596 16532 2648 16584
rect 2780 16532 2832 16584
rect 4344 16532 4396 16584
rect 5632 16643 5684 16652
rect 5632 16609 5641 16643
rect 5641 16609 5675 16643
rect 5675 16609 5684 16643
rect 5632 16600 5684 16609
rect 5908 16643 5960 16652
rect 5908 16609 5917 16643
rect 5917 16609 5951 16643
rect 5951 16609 5960 16643
rect 5908 16600 5960 16609
rect 480 16464 532 16516
rect 3240 16464 3292 16516
rect 3332 16464 3384 16516
rect 1492 16396 1544 16448
rect 3976 16439 4028 16448
rect 3976 16405 3985 16439
rect 3985 16405 4019 16439
rect 4019 16405 4028 16439
rect 3976 16396 4028 16405
rect 6092 16532 6144 16584
rect 4528 16464 4580 16516
rect 4712 16464 4764 16516
rect 6736 16464 6788 16516
rect 7012 16668 7064 16720
rect 8668 16600 8720 16652
rect 12164 16736 12216 16788
rect 12716 16736 12768 16788
rect 10692 16668 10744 16720
rect 13360 16736 13412 16788
rect 15200 16736 15252 16788
rect 7012 16532 7064 16584
rect 6920 16464 6972 16516
rect 9312 16532 9364 16584
rect 10140 16532 10192 16584
rect 10876 16600 10928 16652
rect 11704 16600 11756 16652
rect 10508 16575 10560 16584
rect 10508 16541 10517 16575
rect 10517 16541 10551 16575
rect 10551 16541 10560 16575
rect 10508 16532 10560 16541
rect 11336 16575 11388 16584
rect 11336 16541 11370 16575
rect 11370 16541 11388 16575
rect 11336 16532 11388 16541
rect 12440 16575 12492 16584
rect 12440 16541 12449 16575
rect 12449 16541 12483 16575
rect 12483 16541 12492 16575
rect 12440 16532 12492 16541
rect 12624 16532 12676 16584
rect 15292 16668 15344 16720
rect 15936 16736 15988 16788
rect 16028 16736 16080 16788
rect 16764 16779 16816 16788
rect 16764 16745 16773 16779
rect 16773 16745 16807 16779
rect 16807 16745 16816 16779
rect 16764 16736 16816 16745
rect 14648 16600 14700 16652
rect 14740 16600 14792 16652
rect 14280 16532 14332 16584
rect 15200 16600 15252 16652
rect 20352 16779 20404 16788
rect 20352 16745 20361 16779
rect 20361 16745 20395 16779
rect 20395 16745 20404 16779
rect 20352 16736 20404 16745
rect 20904 16600 20956 16652
rect 21456 16643 21508 16652
rect 21456 16609 21465 16643
rect 21465 16609 21499 16643
rect 21499 16609 21508 16643
rect 21456 16600 21508 16609
rect 15844 16575 15896 16584
rect 15844 16541 15853 16575
rect 15853 16541 15887 16575
rect 15887 16541 15896 16575
rect 15844 16532 15896 16541
rect 5448 16396 5500 16448
rect 5540 16396 5592 16448
rect 6092 16396 6144 16448
rect 7564 16396 7616 16448
rect 10048 16396 10100 16448
rect 11060 16396 11112 16448
rect 11336 16396 11388 16448
rect 12164 16439 12216 16448
rect 12164 16405 12173 16439
rect 12173 16405 12207 16439
rect 12207 16405 12216 16439
rect 12164 16396 12216 16405
rect 15292 16396 15344 16448
rect 15384 16396 15436 16448
rect 17592 16532 17644 16584
rect 17040 16396 17092 16448
rect 20168 16532 20220 16584
rect 20720 16575 20772 16584
rect 20720 16541 20729 16575
rect 20729 16541 20763 16575
rect 20763 16541 20772 16575
rect 20720 16532 20772 16541
rect 21088 16532 21140 16584
rect 19984 16464 20036 16516
rect 19616 16396 19668 16448
rect 20996 16439 21048 16448
rect 20996 16405 21005 16439
rect 21005 16405 21039 16439
rect 21039 16405 21048 16439
rect 20996 16396 21048 16405
rect 6148 16294 6200 16346
rect 6212 16294 6264 16346
rect 6276 16294 6328 16346
rect 6340 16294 6392 16346
rect 6404 16294 6456 16346
rect 11346 16294 11398 16346
rect 11410 16294 11462 16346
rect 11474 16294 11526 16346
rect 11538 16294 11590 16346
rect 11602 16294 11654 16346
rect 16544 16294 16596 16346
rect 16608 16294 16660 16346
rect 16672 16294 16724 16346
rect 16736 16294 16788 16346
rect 16800 16294 16852 16346
rect 21742 16294 21794 16346
rect 21806 16294 21858 16346
rect 21870 16294 21922 16346
rect 21934 16294 21986 16346
rect 21998 16294 22050 16346
rect 1308 16192 1360 16244
rect 2780 16192 2832 16244
rect 5264 16192 5316 16244
rect 1492 16167 1544 16176
rect 1492 16133 1501 16167
rect 1501 16133 1535 16167
rect 1535 16133 1544 16167
rect 1492 16124 1544 16133
rect 2320 16056 2372 16108
rect 3424 16099 3476 16108
rect 3424 16065 3433 16099
rect 3433 16065 3467 16099
rect 3467 16065 3476 16099
rect 3424 16056 3476 16065
rect 4252 16099 4304 16108
rect 4252 16065 4261 16099
rect 4261 16065 4295 16099
rect 4295 16065 4304 16099
rect 4252 16056 4304 16065
rect 2044 15988 2096 16040
rect 2596 15988 2648 16040
rect 2964 15988 3016 16040
rect 4896 16124 4948 16176
rect 4988 16124 5040 16176
rect 7196 16192 7248 16244
rect 7288 16192 7340 16244
rect 6000 16124 6052 16176
rect 9220 16124 9272 16176
rect 6920 16056 6972 16108
rect 7012 16056 7064 16108
rect 7288 16056 7340 16108
rect 8300 16056 8352 16108
rect 9956 16192 10008 16244
rect 11244 16192 11296 16244
rect 12808 16192 12860 16244
rect 13452 16192 13504 16244
rect 9680 16124 9732 16176
rect 10600 16056 10652 16108
rect 12440 16124 12492 16176
rect 13636 16124 13688 16176
rect 15936 16192 15988 16244
rect 12072 16056 12124 16108
rect 2504 15920 2556 15972
rect 3792 15852 3844 15904
rect 3884 15852 3936 15904
rect 4988 15852 5040 15904
rect 5356 15852 5408 15904
rect 9680 16031 9732 16040
rect 9680 15997 9689 16031
rect 9689 15997 9723 16031
rect 9723 15997 9732 16031
rect 9680 15988 9732 15997
rect 10048 15988 10100 16040
rect 10232 15988 10284 16040
rect 10416 16031 10468 16040
rect 10416 15997 10425 16031
rect 10425 15997 10459 16031
rect 10459 15997 10468 16031
rect 10416 15988 10468 15997
rect 10876 15988 10928 16040
rect 9128 15895 9180 15904
rect 9128 15861 9137 15895
rect 9137 15861 9171 15895
rect 9171 15861 9180 15895
rect 9128 15852 9180 15861
rect 10692 15852 10744 15904
rect 13084 16056 13136 16108
rect 15384 16124 15436 16176
rect 16120 16124 16172 16176
rect 17316 16192 17368 16244
rect 17960 16192 18012 16244
rect 18328 16192 18380 16244
rect 20720 16192 20772 16244
rect 20812 16192 20864 16244
rect 20996 16192 21048 16244
rect 21088 16235 21140 16244
rect 21088 16201 21097 16235
rect 21097 16201 21131 16235
rect 21131 16201 21140 16235
rect 21088 16192 21140 16201
rect 15844 16056 15896 16108
rect 16856 16056 16908 16108
rect 13268 16031 13320 16040
rect 13268 15997 13277 16031
rect 13277 15997 13311 16031
rect 13311 15997 13320 16031
rect 13268 15988 13320 15997
rect 14648 16031 14700 16040
rect 14648 15997 14657 16031
rect 14657 15997 14691 16031
rect 14691 15997 14700 16031
rect 14648 15988 14700 15997
rect 15752 15988 15804 16040
rect 14280 15895 14332 15904
rect 14280 15861 14289 15895
rect 14289 15861 14323 15895
rect 14323 15861 14332 15895
rect 14280 15852 14332 15861
rect 16212 15920 16264 15972
rect 18328 16099 18380 16108
rect 18328 16065 18337 16099
rect 18337 16065 18371 16099
rect 18371 16065 18380 16099
rect 18328 16056 18380 16065
rect 18696 16056 18748 16108
rect 17408 15988 17460 16040
rect 17868 15988 17920 16040
rect 18880 15988 18932 16040
rect 19248 15920 19300 15972
rect 19616 16031 19668 16040
rect 19616 15997 19625 16031
rect 19625 15997 19659 16031
rect 19659 15997 19668 16031
rect 19616 15988 19668 15997
rect 16120 15852 16172 15904
rect 16304 15852 16356 15904
rect 17408 15852 17460 15904
rect 18420 15895 18472 15904
rect 18420 15861 18429 15895
rect 18429 15861 18463 15895
rect 18463 15861 18472 15895
rect 18420 15852 18472 15861
rect 19064 15852 19116 15904
rect 21456 15895 21508 15904
rect 21456 15861 21465 15895
rect 21465 15861 21499 15895
rect 21499 15861 21508 15895
rect 21456 15852 21508 15861
rect 3549 15750 3601 15802
rect 3613 15750 3665 15802
rect 3677 15750 3729 15802
rect 3741 15750 3793 15802
rect 3805 15750 3857 15802
rect 8747 15750 8799 15802
rect 8811 15750 8863 15802
rect 8875 15750 8927 15802
rect 8939 15750 8991 15802
rect 9003 15750 9055 15802
rect 13945 15750 13997 15802
rect 14009 15750 14061 15802
rect 14073 15750 14125 15802
rect 14137 15750 14189 15802
rect 14201 15750 14253 15802
rect 19143 15750 19195 15802
rect 19207 15750 19259 15802
rect 19271 15750 19323 15802
rect 19335 15750 19387 15802
rect 19399 15750 19451 15802
rect 2412 15691 2464 15700
rect 2412 15657 2421 15691
rect 2421 15657 2455 15691
rect 2455 15657 2464 15691
rect 2412 15648 2464 15657
rect 4252 15648 4304 15700
rect 4344 15648 4396 15700
rect 9128 15648 9180 15700
rect 9220 15648 9272 15700
rect 14280 15648 14332 15700
rect 18328 15648 18380 15700
rect 18420 15648 18472 15700
rect 19064 15648 19116 15700
rect 19524 15648 19576 15700
rect 3148 15580 3200 15632
rect 3976 15580 4028 15632
rect 4528 15580 4580 15632
rect 1676 15487 1728 15496
rect 1676 15453 1683 15487
rect 1683 15453 1717 15487
rect 1717 15453 1728 15487
rect 1676 15444 1728 15453
rect 2044 15444 2096 15496
rect 4160 15512 4212 15564
rect 4344 15512 4396 15564
rect 5080 15555 5132 15564
rect 5080 15521 5114 15555
rect 5114 15521 5132 15555
rect 5080 15512 5132 15521
rect 5448 15512 5500 15564
rect 10784 15580 10836 15632
rect 12624 15512 12676 15564
rect 12716 15555 12768 15564
rect 12716 15521 12725 15555
rect 12725 15521 12759 15555
rect 12759 15521 12768 15555
rect 12716 15512 12768 15521
rect 18696 15623 18748 15632
rect 18696 15589 18705 15623
rect 18705 15589 18739 15623
rect 18739 15589 18748 15623
rect 18696 15580 18748 15589
rect 14556 15555 14608 15564
rect 14556 15521 14565 15555
rect 14565 15521 14599 15555
rect 14599 15521 14608 15555
rect 14556 15512 14608 15521
rect 15384 15512 15436 15564
rect 15568 15512 15620 15564
rect 18880 15512 18932 15564
rect 20904 15691 20956 15700
rect 20904 15657 20913 15691
rect 20913 15657 20947 15691
rect 20947 15657 20956 15691
rect 20904 15648 20956 15657
rect 4252 15487 4304 15496
rect 4252 15453 4261 15487
rect 4261 15453 4295 15487
rect 4295 15453 4304 15487
rect 4252 15444 4304 15453
rect 5264 15487 5316 15496
rect 5264 15453 5273 15487
rect 5273 15453 5307 15487
rect 5307 15453 5316 15487
rect 5264 15444 5316 15453
rect 5908 15444 5960 15496
rect 8024 15444 8076 15496
rect 8668 15444 8720 15496
rect 9220 15487 9272 15496
rect 9220 15453 9229 15487
rect 9229 15453 9263 15487
rect 9263 15453 9272 15487
rect 9220 15444 9272 15453
rect 11888 15444 11940 15496
rect 13176 15444 13228 15496
rect 14372 15444 14424 15496
rect 3056 15308 3108 15360
rect 4068 15308 4120 15360
rect 6736 15376 6788 15428
rect 5540 15308 5592 15360
rect 6000 15351 6052 15360
rect 6000 15317 6009 15351
rect 6009 15317 6043 15351
rect 6043 15317 6052 15351
rect 6000 15308 6052 15317
rect 7380 15419 7432 15428
rect 7380 15385 7389 15419
rect 7389 15385 7423 15419
rect 7423 15385 7432 15419
rect 7380 15376 7432 15385
rect 7472 15376 7524 15428
rect 7840 15376 7892 15428
rect 9312 15376 9364 15428
rect 15200 15444 15252 15496
rect 16212 15444 16264 15496
rect 17132 15444 17184 15496
rect 7012 15308 7064 15360
rect 7564 15308 7616 15360
rect 10232 15351 10284 15360
rect 10232 15317 10241 15351
rect 10241 15317 10275 15351
rect 10275 15317 10284 15351
rect 10232 15308 10284 15317
rect 11704 15308 11756 15360
rect 12072 15308 12124 15360
rect 19156 15444 19208 15496
rect 19800 15444 19852 15496
rect 20720 15444 20772 15496
rect 21180 15487 21232 15496
rect 21180 15453 21189 15487
rect 21189 15453 21223 15487
rect 21223 15453 21232 15487
rect 21180 15444 21232 15453
rect 18972 15376 19024 15428
rect 13820 15308 13872 15360
rect 15568 15351 15620 15360
rect 15568 15317 15577 15351
rect 15577 15317 15611 15351
rect 15611 15317 15620 15351
rect 15568 15308 15620 15317
rect 16856 15308 16908 15360
rect 18420 15308 18472 15360
rect 21088 15376 21140 15428
rect 22560 15376 22612 15428
rect 20720 15308 20772 15360
rect 6148 15206 6200 15258
rect 6212 15206 6264 15258
rect 6276 15206 6328 15258
rect 6340 15206 6392 15258
rect 6404 15206 6456 15258
rect 11346 15206 11398 15258
rect 11410 15206 11462 15258
rect 11474 15206 11526 15258
rect 11538 15206 11590 15258
rect 11602 15206 11654 15258
rect 16544 15206 16596 15258
rect 16608 15206 16660 15258
rect 16672 15206 16724 15258
rect 16736 15206 16788 15258
rect 16800 15206 16852 15258
rect 21742 15206 21794 15258
rect 21806 15206 21858 15258
rect 21870 15206 21922 15258
rect 21934 15206 21986 15258
rect 21998 15206 22050 15258
rect 22192 15172 22244 15224
rect 22560 15172 22612 15224
rect 3148 15104 3200 15156
rect 5908 15104 5960 15156
rect 5080 15036 5132 15088
rect 3976 15011 4028 15020
rect 3976 14977 4010 15011
rect 4010 14977 4028 15011
rect 3976 14968 4028 14977
rect 4160 15011 4212 15020
rect 4160 14977 4169 15011
rect 4169 14977 4203 15011
rect 4203 14977 4212 15011
rect 4160 14968 4212 14977
rect 5724 14968 5776 15020
rect 7380 15104 7432 15156
rect 8300 15104 8352 15156
rect 9496 15104 9548 15156
rect 2964 14943 3016 14952
rect 2964 14909 2973 14943
rect 2973 14909 3007 14943
rect 3007 14909 3016 14943
rect 2964 14900 3016 14909
rect 1860 14764 1912 14816
rect 3976 14764 4028 14816
rect 4252 14764 4304 14816
rect 6092 14900 6144 14952
rect 6368 14943 6420 14952
rect 6368 14909 6377 14943
rect 6377 14909 6411 14943
rect 6411 14909 6420 14943
rect 6368 14900 6420 14909
rect 8208 14968 8260 15020
rect 9220 15036 9272 15088
rect 10324 15041 10376 15088
rect 10324 15036 10349 15041
rect 10349 15036 10376 15041
rect 12440 15036 12492 15088
rect 12716 15104 12768 15156
rect 15752 15104 15804 15156
rect 16120 15104 16172 15156
rect 16396 15104 16448 15156
rect 17132 15104 17184 15156
rect 18880 15104 18932 15156
rect 19800 15104 19852 15156
rect 20720 15104 20772 15156
rect 7472 14900 7524 14952
rect 7564 14943 7616 14952
rect 7564 14909 7573 14943
rect 7573 14909 7607 14943
rect 7607 14909 7616 14943
rect 7564 14900 7616 14909
rect 7932 14900 7984 14952
rect 8668 14943 8720 14952
rect 8668 14909 8677 14943
rect 8677 14909 8711 14943
rect 8711 14909 8720 14943
rect 8668 14900 8720 14909
rect 15568 14968 15620 15020
rect 18052 15011 18104 15020
rect 18052 14977 18059 15011
rect 18059 14977 18093 15011
rect 18093 14977 18104 15011
rect 18052 14968 18104 14977
rect 12900 14900 12952 14952
rect 14280 14900 14332 14952
rect 4620 14832 4672 14884
rect 4896 14764 4948 14816
rect 5172 14764 5224 14816
rect 6552 14764 6604 14816
rect 6920 14832 6972 14884
rect 7472 14764 7524 14816
rect 8208 14807 8260 14816
rect 8208 14773 8217 14807
rect 8217 14773 8251 14807
rect 8251 14773 8260 14807
rect 8208 14764 8260 14773
rect 8392 14764 8444 14816
rect 10048 14764 10100 14816
rect 11060 14807 11112 14816
rect 11060 14773 11069 14807
rect 11069 14773 11103 14807
rect 11103 14773 11112 14807
rect 11060 14764 11112 14773
rect 12808 14832 12860 14884
rect 13544 14832 13596 14884
rect 13636 14764 13688 14816
rect 14372 14875 14424 14884
rect 14372 14841 14381 14875
rect 14381 14841 14415 14875
rect 14415 14841 14424 14875
rect 14372 14832 14424 14841
rect 14832 14900 14884 14952
rect 17684 14900 17736 14952
rect 20904 15011 20956 15020
rect 20904 14977 20913 15011
rect 20913 14977 20947 15011
rect 20947 14977 20956 15011
rect 20904 14968 20956 14977
rect 22744 14968 22796 15020
rect 14832 14764 14884 14816
rect 15568 14807 15620 14816
rect 15568 14773 15577 14807
rect 15577 14773 15611 14807
rect 15611 14773 15620 14807
rect 15568 14764 15620 14773
rect 16396 14764 16448 14816
rect 17316 14764 17368 14816
rect 20352 14807 20404 14816
rect 20352 14773 20361 14807
rect 20361 14773 20395 14807
rect 20395 14773 20404 14807
rect 20352 14764 20404 14773
rect 22744 14832 22796 14884
rect 20996 14807 21048 14816
rect 20996 14773 21005 14807
rect 21005 14773 21039 14807
rect 21039 14773 21048 14807
rect 20996 14764 21048 14773
rect 21456 14807 21508 14816
rect 21456 14773 21465 14807
rect 21465 14773 21499 14807
rect 21499 14773 21508 14807
rect 21456 14764 21508 14773
rect 3549 14662 3601 14714
rect 3613 14662 3665 14714
rect 3677 14662 3729 14714
rect 3741 14662 3793 14714
rect 3805 14662 3857 14714
rect 8747 14662 8799 14714
rect 8811 14662 8863 14714
rect 8875 14662 8927 14714
rect 8939 14662 8991 14714
rect 9003 14662 9055 14714
rect 13945 14662 13997 14714
rect 14009 14662 14061 14714
rect 14073 14662 14125 14714
rect 14137 14662 14189 14714
rect 14201 14662 14253 14714
rect 19143 14662 19195 14714
rect 19207 14662 19259 14714
rect 19271 14662 19323 14714
rect 19335 14662 19387 14714
rect 19399 14662 19451 14714
rect 1768 14603 1820 14612
rect 1768 14569 1777 14603
rect 1777 14569 1811 14603
rect 1811 14569 1820 14603
rect 1768 14560 1820 14569
rect 4344 14560 4396 14612
rect 5264 14603 5316 14612
rect 5264 14569 5273 14603
rect 5273 14569 5307 14603
rect 5307 14569 5316 14603
rect 5264 14560 5316 14569
rect 4252 14492 4304 14544
rect 3424 14424 3476 14476
rect 3608 14424 3660 14476
rect 1216 14356 1268 14408
rect 2688 14288 2740 14340
rect 4344 14288 4396 14340
rect 4620 14356 4672 14408
rect 5908 14399 5960 14408
rect 4712 14288 4764 14340
rect 5356 14288 5408 14340
rect 1216 14220 1268 14272
rect 2412 14220 2464 14272
rect 3240 14220 3292 14272
rect 5908 14365 5915 14399
rect 5915 14365 5949 14399
rect 5949 14365 5960 14399
rect 6460 14560 6512 14612
rect 7472 14560 7524 14612
rect 8024 14603 8076 14612
rect 8024 14569 8033 14603
rect 8033 14569 8067 14603
rect 8067 14569 8076 14603
rect 8024 14560 8076 14569
rect 9772 14560 9824 14612
rect 10968 14560 11020 14612
rect 11612 14560 11664 14612
rect 12900 14560 12952 14612
rect 13636 14603 13688 14612
rect 13636 14569 13645 14603
rect 13645 14569 13679 14603
rect 13679 14569 13688 14603
rect 13636 14560 13688 14569
rect 14372 14560 14424 14612
rect 15568 14560 15620 14612
rect 6368 14492 6420 14544
rect 7012 14492 7064 14544
rect 10232 14492 10284 14544
rect 6552 14424 6604 14476
rect 6736 14424 6788 14476
rect 10140 14424 10192 14476
rect 10600 14424 10652 14476
rect 11612 14424 11664 14476
rect 12440 14467 12492 14476
rect 12440 14433 12449 14467
rect 12449 14433 12483 14467
rect 12483 14433 12492 14467
rect 12440 14424 12492 14433
rect 12716 14467 12768 14476
rect 12716 14433 12725 14467
rect 12725 14433 12759 14467
rect 12759 14433 12768 14467
rect 12716 14424 12768 14433
rect 13360 14424 13412 14476
rect 13544 14424 13596 14476
rect 5908 14356 5960 14365
rect 9864 14399 9916 14408
rect 9864 14365 9873 14399
rect 9873 14365 9907 14399
rect 9907 14365 9916 14399
rect 9864 14356 9916 14365
rect 10784 14399 10836 14408
rect 10784 14365 10793 14399
rect 10793 14365 10827 14399
rect 10827 14365 10836 14399
rect 10784 14356 10836 14365
rect 11060 14399 11112 14408
rect 11060 14365 11069 14399
rect 11069 14365 11103 14399
rect 11103 14365 11112 14399
rect 11060 14356 11112 14365
rect 11888 14356 11940 14408
rect 12992 14399 13044 14408
rect 12992 14365 13001 14399
rect 13001 14365 13035 14399
rect 13035 14365 13044 14399
rect 12992 14356 13044 14365
rect 14096 14399 14148 14408
rect 14096 14365 14105 14399
rect 14105 14365 14139 14399
rect 14139 14365 14148 14399
rect 14096 14356 14148 14365
rect 7104 14288 7156 14340
rect 17684 14424 17736 14476
rect 19616 14560 19668 14612
rect 20352 14560 20404 14612
rect 20904 14560 20956 14612
rect 20996 14560 21048 14612
rect 15660 14356 15712 14408
rect 15752 14399 15804 14408
rect 15752 14365 15761 14399
rect 15761 14365 15795 14399
rect 15795 14365 15804 14399
rect 15752 14356 15804 14365
rect 16304 14356 16356 14408
rect 7288 14220 7340 14272
rect 7932 14220 7984 14272
rect 10968 14220 11020 14272
rect 11704 14263 11756 14272
rect 11704 14229 11713 14263
rect 11713 14229 11747 14263
rect 11747 14229 11756 14263
rect 11704 14220 11756 14229
rect 14556 14288 14608 14340
rect 15200 14288 15252 14340
rect 21088 14356 21140 14408
rect 14096 14220 14148 14272
rect 15936 14263 15988 14272
rect 15936 14229 15945 14263
rect 15945 14229 15979 14263
rect 15979 14229 15988 14263
rect 15936 14220 15988 14229
rect 17960 14220 18012 14272
rect 21180 14263 21232 14272
rect 21180 14229 21189 14263
rect 21189 14229 21223 14263
rect 21223 14229 21232 14263
rect 21180 14220 21232 14229
rect 22192 14220 22244 14272
rect 6148 14118 6200 14170
rect 6212 14118 6264 14170
rect 6276 14118 6328 14170
rect 6340 14118 6392 14170
rect 6404 14118 6456 14170
rect 11346 14118 11398 14170
rect 11410 14118 11462 14170
rect 11474 14118 11526 14170
rect 11538 14118 11590 14170
rect 11602 14118 11654 14170
rect 16544 14118 16596 14170
rect 16608 14118 16660 14170
rect 16672 14118 16724 14170
rect 16736 14118 16788 14170
rect 16800 14118 16852 14170
rect 21742 14118 21794 14170
rect 21806 14118 21858 14170
rect 21870 14118 21922 14170
rect 21934 14118 21986 14170
rect 21998 14118 22050 14170
rect 940 13948 992 14000
rect 4160 14016 4212 14068
rect 4436 14016 4488 14068
rect 5264 14016 5316 14068
rect 5356 14016 5408 14068
rect 5632 14016 5684 14068
rect 1768 13923 1820 13932
rect 1768 13889 1777 13923
rect 1777 13889 1811 13923
rect 1811 13889 1820 13923
rect 1768 13880 1820 13889
rect 3240 13923 3292 13932
rect 3240 13889 3249 13923
rect 3249 13889 3283 13923
rect 3283 13889 3292 13923
rect 3240 13880 3292 13889
rect 3424 13880 3476 13932
rect 4436 13880 4488 13932
rect 5080 13880 5132 13932
rect 6276 13948 6328 14000
rect 6552 13948 6604 14000
rect 7012 13991 7064 14000
rect 7012 13957 7021 13991
rect 7021 13957 7055 13991
rect 7055 13957 7064 13991
rect 7012 13948 7064 13957
rect 7104 13923 7156 13932
rect 7104 13889 7113 13923
rect 7113 13889 7147 13923
rect 7147 13889 7156 13923
rect 7104 13880 7156 13889
rect 7380 13880 7432 13932
rect 7564 13880 7616 13932
rect 7840 13923 7892 13932
rect 7840 13889 7863 13923
rect 7863 13889 7892 13923
rect 7840 13880 7892 13889
rect 1952 13812 2004 13864
rect 2872 13812 2924 13864
rect 3056 13812 3108 13864
rect 4344 13812 4396 13864
rect 6552 13812 6604 13864
rect 9956 13880 10008 13932
rect 10048 13923 10100 13932
rect 10048 13889 10057 13923
rect 10057 13889 10091 13923
rect 10091 13889 10100 13923
rect 10048 13880 10100 13889
rect 10876 13880 10928 13932
rect 9220 13812 9272 13864
rect 10232 13812 10284 13864
rect 11060 14016 11112 14068
rect 11704 14016 11756 14068
rect 12072 14016 12124 14068
rect 11980 13948 12032 14000
rect 12992 14016 13044 14068
rect 13176 14016 13228 14068
rect 13544 14016 13596 14068
rect 14464 14016 14516 14068
rect 14740 14016 14792 14068
rect 14280 13948 14332 14000
rect 15200 13948 15252 14000
rect 16580 14016 16632 14068
rect 21088 14016 21140 14068
rect 21180 14016 21232 14068
rect 16120 13948 16172 14000
rect 16212 13991 16264 14000
rect 16212 13957 16221 13991
rect 16221 13957 16255 13991
rect 16255 13957 16264 13991
rect 16212 13948 16264 13957
rect 19800 13948 19852 14000
rect 20076 13948 20128 14000
rect 12900 13880 12952 13932
rect 13176 13880 13228 13932
rect 15844 13923 15896 13932
rect 15844 13889 15853 13923
rect 15853 13889 15887 13923
rect 15887 13889 15896 13923
rect 15844 13880 15896 13889
rect 16948 13923 17000 13932
rect 16948 13889 16955 13923
rect 16955 13889 16989 13923
rect 16989 13889 17000 13923
rect 16948 13880 17000 13889
rect 18972 13923 19024 13932
rect 18972 13889 18981 13923
rect 18981 13889 19015 13923
rect 19015 13889 19024 13923
rect 18972 13880 19024 13889
rect 19524 13880 19576 13932
rect 20720 13880 20772 13932
rect 11152 13812 11204 13864
rect 572 13744 624 13796
rect 1400 13787 1452 13796
rect 1400 13753 1409 13787
rect 1409 13753 1443 13787
rect 1443 13753 1452 13787
rect 1400 13744 1452 13753
rect 2412 13676 2464 13728
rect 2872 13719 2924 13728
rect 2872 13685 2881 13719
rect 2881 13685 2915 13719
rect 2915 13685 2924 13719
rect 2872 13676 2924 13685
rect 3240 13676 3292 13728
rect 4252 13744 4304 13796
rect 4620 13744 4672 13796
rect 9496 13787 9548 13796
rect 9496 13753 9505 13787
rect 9505 13753 9539 13787
rect 9539 13753 9548 13787
rect 9496 13744 9548 13753
rect 5908 13676 5960 13728
rect 9772 13676 9824 13728
rect 11336 13676 11388 13728
rect 13360 13676 13412 13728
rect 16396 13787 16448 13796
rect 16396 13753 16405 13787
rect 16405 13753 16439 13787
rect 16439 13753 16448 13787
rect 16396 13744 16448 13753
rect 18880 13676 18932 13728
rect 21272 13676 21324 13728
rect 21456 13719 21508 13728
rect 21456 13685 21465 13719
rect 21465 13685 21499 13719
rect 21499 13685 21508 13719
rect 21456 13676 21508 13685
rect 572 13540 624 13592
rect 3549 13574 3601 13626
rect 3613 13574 3665 13626
rect 3677 13574 3729 13626
rect 3741 13574 3793 13626
rect 3805 13574 3857 13626
rect 8747 13574 8799 13626
rect 8811 13574 8863 13626
rect 8875 13574 8927 13626
rect 8939 13574 8991 13626
rect 9003 13574 9055 13626
rect 13945 13574 13997 13626
rect 14009 13574 14061 13626
rect 14073 13574 14125 13626
rect 14137 13574 14189 13626
rect 14201 13574 14253 13626
rect 19143 13574 19195 13626
rect 19207 13574 19259 13626
rect 19271 13574 19323 13626
rect 19335 13574 19387 13626
rect 19399 13574 19451 13626
rect 940 13472 992 13524
rect 3424 13472 3476 13524
rect 4160 13472 4212 13524
rect 1400 13336 1452 13388
rect 1952 13336 2004 13388
rect 3884 13336 3936 13388
rect 4712 13379 4764 13388
rect 4712 13345 4721 13379
rect 4721 13345 4755 13379
rect 4755 13345 4764 13379
rect 4712 13336 4764 13345
rect 4896 13336 4948 13388
rect 5540 13472 5592 13524
rect 7104 13515 7156 13524
rect 7104 13481 7113 13515
rect 7113 13481 7147 13515
rect 7147 13481 7156 13515
rect 7104 13472 7156 13481
rect 9496 13472 9548 13524
rect 10048 13472 10100 13524
rect 10416 13472 10468 13524
rect 10968 13472 11020 13524
rect 7288 13404 7340 13456
rect 7472 13379 7524 13388
rect 7472 13345 7481 13379
rect 7481 13345 7515 13379
rect 7515 13345 7524 13379
rect 7472 13336 7524 13345
rect 8300 13336 8352 13388
rect 9864 13336 9916 13388
rect 10416 13379 10468 13388
rect 10416 13345 10425 13379
rect 10425 13345 10459 13379
rect 10459 13345 10468 13379
rect 10416 13336 10468 13345
rect 10692 13379 10744 13388
rect 10692 13345 10701 13379
rect 10701 13345 10735 13379
rect 10735 13345 10744 13379
rect 10692 13336 10744 13345
rect 10876 13336 10928 13388
rect 11336 13336 11388 13388
rect 2136 13268 2188 13320
rect 2596 13268 2648 13320
rect 2964 13268 3016 13320
rect 3792 13311 3844 13320
rect 3792 13277 3801 13311
rect 3801 13277 3835 13311
rect 3835 13277 3844 13311
rect 3792 13268 3844 13277
rect 3976 13311 4028 13320
rect 3976 13277 3985 13311
rect 3985 13277 4019 13311
rect 4019 13277 4028 13311
rect 3976 13268 4028 13277
rect 5724 13268 5776 13320
rect 5816 13268 5868 13320
rect 6276 13268 6328 13320
rect 7840 13268 7892 13320
rect 9220 13268 9272 13320
rect 9680 13268 9732 13320
rect 9956 13311 10008 13320
rect 9956 13277 9965 13311
rect 9965 13277 9999 13311
rect 9999 13277 10008 13311
rect 9956 13268 10008 13277
rect 10968 13311 11020 13320
rect 10968 13277 10977 13311
rect 10977 13277 11011 13311
rect 11011 13277 11020 13311
rect 10968 13268 11020 13277
rect 11980 13472 12032 13524
rect 12440 13472 12492 13524
rect 14188 13336 14240 13388
rect 14740 13447 14792 13456
rect 14740 13413 14749 13447
rect 14749 13413 14783 13447
rect 14783 13413 14792 13447
rect 14740 13404 14792 13413
rect 1308 13132 1360 13184
rect 5632 13175 5684 13184
rect 5632 13141 5641 13175
rect 5641 13141 5675 13175
rect 5675 13141 5684 13175
rect 5632 13132 5684 13141
rect 5724 13132 5776 13184
rect 6460 13132 6512 13184
rect 8576 13200 8628 13252
rect 11704 13200 11756 13252
rect 13268 13268 13320 13320
rect 15752 13472 15804 13524
rect 16580 13472 16632 13524
rect 15844 13336 15896 13388
rect 16120 13379 16172 13388
rect 16120 13345 16129 13379
rect 16129 13345 16163 13379
rect 16163 13345 16172 13379
rect 16120 13336 16172 13345
rect 15016 13311 15068 13320
rect 15016 13277 15025 13311
rect 15025 13277 15059 13311
rect 15059 13277 15068 13311
rect 15016 13268 15068 13277
rect 15292 13311 15344 13320
rect 15292 13277 15301 13311
rect 15301 13277 15335 13311
rect 15335 13277 15344 13311
rect 15292 13268 15344 13277
rect 13820 13200 13872 13252
rect 17040 13268 17092 13320
rect 18972 13472 19024 13524
rect 20812 13472 20864 13524
rect 19064 13404 19116 13456
rect 18512 13268 18564 13320
rect 19616 13311 19668 13320
rect 19616 13277 19625 13311
rect 19625 13277 19659 13311
rect 19659 13277 19668 13311
rect 19616 13268 19668 13277
rect 19984 13268 20036 13320
rect 20720 13268 20772 13320
rect 16396 13247 16421 13252
rect 16421 13247 16448 13252
rect 16396 13200 16448 13247
rect 18604 13200 18656 13252
rect 9220 13132 9272 13184
rect 12440 13132 12492 13184
rect 19064 13175 19116 13184
rect 19064 13141 19073 13175
rect 19073 13141 19107 13175
rect 19107 13141 19116 13175
rect 19064 13132 19116 13141
rect 20628 13175 20680 13184
rect 20628 13141 20637 13175
rect 20637 13141 20671 13175
rect 20671 13141 20680 13175
rect 20628 13132 20680 13141
rect 21364 13175 21416 13184
rect 21364 13141 21373 13175
rect 21373 13141 21407 13175
rect 21407 13141 21416 13175
rect 21364 13132 21416 13141
rect 6148 13030 6200 13082
rect 6212 13030 6264 13082
rect 6276 13030 6328 13082
rect 6340 13030 6392 13082
rect 6404 13030 6456 13082
rect 11346 13030 11398 13082
rect 11410 13030 11462 13082
rect 11474 13030 11526 13082
rect 11538 13030 11590 13082
rect 11602 13030 11654 13082
rect 16544 13030 16596 13082
rect 16608 13030 16660 13082
rect 16672 13030 16724 13082
rect 16736 13030 16788 13082
rect 16800 13030 16852 13082
rect 21742 13030 21794 13082
rect 21806 13030 21858 13082
rect 21870 13030 21922 13082
rect 21934 13030 21986 13082
rect 21998 13030 22050 13082
rect 13728 12928 13780 12980
rect 14740 12928 14792 12980
rect 15292 12928 15344 12980
rect 16396 12928 16448 12980
rect 18604 12928 18656 12980
rect 19064 12928 19116 12980
rect 5816 12860 5868 12912
rect 7104 12860 7156 12912
rect 7380 12903 7432 12912
rect 7380 12869 7389 12903
rect 7389 12869 7423 12903
rect 7423 12869 7432 12903
rect 7380 12860 7432 12869
rect 7564 12860 7616 12912
rect 2228 12792 2280 12844
rect 2504 12835 2556 12844
rect 2504 12801 2513 12835
rect 2513 12801 2547 12835
rect 2547 12801 2556 12835
rect 2504 12792 2556 12801
rect 3240 12835 3292 12844
rect 3240 12801 3249 12835
rect 3249 12801 3283 12835
rect 3283 12801 3292 12835
rect 3240 12792 3292 12801
rect 3516 12835 3568 12844
rect 3516 12801 3525 12835
rect 3525 12801 3559 12835
rect 3559 12801 3568 12835
rect 3516 12792 3568 12801
rect 4620 12792 4672 12844
rect 5356 12792 5408 12844
rect 5724 12792 5776 12844
rect 6276 12792 6328 12844
rect 7012 12835 7064 12844
rect 7012 12801 7021 12835
rect 7021 12801 7055 12835
rect 7055 12801 7064 12835
rect 7012 12792 7064 12801
rect 7288 12792 7340 12844
rect 8852 12792 8904 12844
rect 9312 12860 9364 12912
rect 1400 12724 1452 12776
rect 2320 12767 2372 12776
rect 2320 12733 2329 12767
rect 2329 12733 2363 12767
rect 2363 12733 2372 12767
rect 2320 12724 2372 12733
rect 3700 12724 3752 12776
rect 1492 12588 1544 12640
rect 2964 12699 3016 12708
rect 2964 12665 2973 12699
rect 2973 12665 3007 12699
rect 3007 12665 3016 12699
rect 2964 12656 3016 12665
rect 4804 12588 4856 12640
rect 6552 12724 6604 12776
rect 7748 12724 7800 12776
rect 5724 12699 5776 12708
rect 5724 12665 5733 12699
rect 5733 12665 5767 12699
rect 5767 12665 5776 12699
rect 5724 12656 5776 12665
rect 10416 12860 10468 12912
rect 11152 12860 11204 12912
rect 10324 12835 10376 12844
rect 10324 12801 10331 12835
rect 10331 12801 10365 12835
rect 10365 12801 10376 12835
rect 12532 12860 12584 12912
rect 10324 12792 10376 12801
rect 5632 12588 5684 12640
rect 6368 12588 6420 12640
rect 10048 12588 10100 12640
rect 10324 12588 10376 12640
rect 12808 12792 12860 12844
rect 10968 12724 11020 12776
rect 11152 12724 11204 12776
rect 11704 12724 11756 12776
rect 12900 12656 12952 12708
rect 13820 12792 13872 12844
rect 14556 12792 14608 12844
rect 15016 12792 15068 12844
rect 16856 12792 16908 12844
rect 17776 12835 17828 12844
rect 17776 12801 17785 12835
rect 17785 12801 17819 12835
rect 17819 12801 17828 12835
rect 17776 12792 17828 12801
rect 18512 12792 18564 12844
rect 13084 12631 13136 12640
rect 13084 12597 13093 12631
rect 13093 12597 13127 12631
rect 13127 12597 13136 12631
rect 13084 12588 13136 12597
rect 13452 12588 13504 12640
rect 17960 12767 18012 12776
rect 17960 12733 17969 12767
rect 17969 12733 18003 12767
rect 18003 12733 18012 12767
rect 17960 12724 18012 12733
rect 19524 12792 19576 12844
rect 19800 12835 19852 12844
rect 19800 12801 19809 12835
rect 19809 12801 19843 12835
rect 19843 12801 19852 12835
rect 19800 12792 19852 12801
rect 21364 12928 21416 12980
rect 20628 12860 20680 12912
rect 19064 12588 19116 12640
rect 19892 12724 19944 12776
rect 19984 12767 20036 12776
rect 19984 12733 19993 12767
rect 19993 12733 20027 12767
rect 20027 12733 20036 12767
rect 19984 12724 20036 12733
rect 20904 12724 20956 12776
rect 19616 12588 19668 12640
rect 19800 12588 19852 12640
rect 20076 12631 20128 12640
rect 20076 12597 20085 12631
rect 20085 12597 20119 12631
rect 20119 12597 20128 12631
rect 20076 12588 20128 12597
rect 20720 12588 20772 12640
rect 21088 12631 21140 12640
rect 21088 12597 21097 12631
rect 21097 12597 21131 12631
rect 21131 12597 21140 12631
rect 21088 12588 21140 12597
rect 3549 12486 3601 12538
rect 3613 12486 3665 12538
rect 3677 12486 3729 12538
rect 3741 12486 3793 12538
rect 3805 12486 3857 12538
rect 8747 12486 8799 12538
rect 8811 12486 8863 12538
rect 8875 12486 8927 12538
rect 8939 12486 8991 12538
rect 9003 12486 9055 12538
rect 13945 12486 13997 12538
rect 14009 12486 14061 12538
rect 14073 12486 14125 12538
rect 14137 12486 14189 12538
rect 14201 12486 14253 12538
rect 19143 12486 19195 12538
rect 19207 12486 19259 12538
rect 19271 12486 19323 12538
rect 19335 12486 19387 12538
rect 19399 12486 19451 12538
rect 22192 12452 22244 12504
rect 1584 12427 1636 12436
rect 1584 12393 1593 12427
rect 1593 12393 1627 12427
rect 1627 12393 1636 12427
rect 1584 12384 1636 12393
rect 2136 12316 2188 12368
rect 2228 12316 2280 12368
rect 3884 12384 3936 12436
rect 3976 12384 4028 12436
rect 4712 12384 4764 12436
rect 5172 12384 5224 12436
rect 6460 12384 6512 12436
rect 7012 12384 7064 12436
rect 7472 12384 7524 12436
rect 7748 12384 7800 12436
rect 10232 12384 10284 12436
rect 4068 12316 4120 12368
rect 4252 12316 4304 12368
rect 6828 12316 6880 12368
rect 4620 12248 4672 12300
rect 4712 12291 4764 12300
rect 4712 12257 4721 12291
rect 4721 12257 4755 12291
rect 4755 12257 4764 12291
rect 4712 12248 4764 12257
rect 7288 12248 7340 12300
rect 10140 12248 10192 12300
rect 10508 12291 10560 12300
rect 10508 12257 10517 12291
rect 10517 12257 10551 12291
rect 10551 12257 10560 12291
rect 10508 12248 10560 12257
rect 10600 12248 10652 12300
rect 12532 12384 12584 12436
rect 12900 12384 12952 12436
rect 13452 12384 13504 12436
rect 13728 12384 13780 12436
rect 14924 12384 14976 12436
rect 13636 12359 13688 12368
rect 13636 12325 13645 12359
rect 13645 12325 13679 12359
rect 13679 12325 13688 12359
rect 13636 12316 13688 12325
rect 1492 12155 1544 12164
rect 1492 12121 1501 12155
rect 1501 12121 1535 12155
rect 1535 12121 1544 12155
rect 1492 12112 1544 12121
rect 3884 12112 3936 12164
rect 5080 12180 5132 12232
rect 5632 12180 5684 12232
rect 7196 12180 7248 12232
rect 7656 12180 7708 12232
rect 9312 12180 9364 12232
rect 9680 12180 9732 12232
rect 9864 12223 9916 12232
rect 9864 12189 9873 12223
rect 9873 12189 9907 12223
rect 9907 12189 9916 12223
rect 9864 12180 9916 12189
rect 10968 12180 11020 12232
rect 12992 12180 13044 12232
rect 14740 12248 14792 12300
rect 16120 12384 16172 12436
rect 16948 12384 17000 12436
rect 17592 12384 17644 12436
rect 18788 12384 18840 12436
rect 19984 12384 20036 12436
rect 20076 12384 20128 12436
rect 20904 12384 20956 12436
rect 16396 12316 16448 12368
rect 17776 12316 17828 12368
rect 18604 12316 18656 12368
rect 18972 12316 19024 12368
rect 16856 12291 16908 12300
rect 16856 12257 16865 12291
rect 16865 12257 16899 12291
rect 16899 12257 16908 12291
rect 16856 12248 16908 12257
rect 13820 12180 13872 12232
rect 2044 12087 2096 12096
rect 2044 12053 2053 12087
rect 2053 12053 2087 12087
rect 2087 12053 2096 12087
rect 2044 12044 2096 12053
rect 3240 12044 3292 12096
rect 3424 12044 3476 12096
rect 8208 12112 8260 12164
rect 6368 12044 6420 12096
rect 6828 12044 6880 12096
rect 7288 12044 7340 12096
rect 8116 12044 8168 12096
rect 9496 12044 9548 12096
rect 11704 12087 11756 12096
rect 11704 12053 11713 12087
rect 11713 12053 11747 12087
rect 11747 12053 11756 12087
rect 11704 12044 11756 12053
rect 11980 12112 12032 12164
rect 13452 12112 13504 12164
rect 15936 12180 15988 12232
rect 17224 12180 17276 12232
rect 14648 12044 14700 12096
rect 15660 12044 15712 12096
rect 16120 12044 16172 12096
rect 17224 12044 17276 12096
rect 17592 12044 17644 12096
rect 17684 12044 17736 12096
rect 18420 12223 18472 12232
rect 18420 12189 18429 12223
rect 18429 12189 18463 12223
rect 18463 12189 18472 12223
rect 18420 12180 18472 12189
rect 19064 12180 19116 12232
rect 19432 12223 19484 12232
rect 19432 12189 19441 12223
rect 19441 12189 19475 12223
rect 19475 12189 19484 12223
rect 19432 12180 19484 12189
rect 19892 12223 19944 12232
rect 19892 12189 19901 12223
rect 19901 12189 19935 12223
rect 19935 12189 19944 12223
rect 19892 12180 19944 12189
rect 19984 12223 20036 12232
rect 19984 12189 19993 12223
rect 19993 12189 20027 12223
rect 20027 12189 20036 12223
rect 19984 12180 20036 12189
rect 20996 12316 21048 12368
rect 20628 12248 20680 12300
rect 20444 12223 20496 12232
rect 20444 12189 20453 12223
rect 20453 12189 20487 12223
rect 20487 12189 20496 12223
rect 20444 12180 20496 12189
rect 20536 12223 20588 12232
rect 20536 12189 20545 12223
rect 20545 12189 20579 12223
rect 20579 12189 20588 12223
rect 20536 12180 20588 12189
rect 20720 12180 20772 12232
rect 22836 12180 22888 12232
rect 18328 12087 18380 12096
rect 18328 12053 18337 12087
rect 18337 12053 18371 12087
rect 18371 12053 18380 12087
rect 18328 12044 18380 12053
rect 18512 12087 18564 12096
rect 18512 12053 18521 12087
rect 18521 12053 18555 12087
rect 18555 12053 18564 12087
rect 18512 12044 18564 12053
rect 18696 12044 18748 12096
rect 20628 12112 20680 12164
rect 20352 12044 20404 12096
rect 22192 12112 22244 12164
rect 21088 12087 21140 12096
rect 21088 12053 21097 12087
rect 21097 12053 21131 12087
rect 21131 12053 21140 12087
rect 21088 12044 21140 12053
rect 6148 11942 6200 11994
rect 6212 11942 6264 11994
rect 6276 11942 6328 11994
rect 6340 11942 6392 11994
rect 6404 11942 6456 11994
rect 11346 11942 11398 11994
rect 11410 11942 11462 11994
rect 11474 11942 11526 11994
rect 11538 11942 11590 11994
rect 11602 11942 11654 11994
rect 16544 11942 16596 11994
rect 16608 11942 16660 11994
rect 16672 11942 16724 11994
rect 16736 11942 16788 11994
rect 16800 11942 16852 11994
rect 21742 11942 21794 11994
rect 21806 11942 21858 11994
rect 21870 11942 21922 11994
rect 21934 11942 21986 11994
rect 21998 11942 22050 11994
rect 1584 11840 1636 11892
rect 2688 11883 2740 11892
rect 2688 11849 2697 11883
rect 2697 11849 2731 11883
rect 2731 11849 2740 11883
rect 2688 11840 2740 11849
rect 1400 11704 1452 11756
rect 1768 11772 1820 11824
rect 4528 11840 4580 11892
rect 4712 11840 4764 11892
rect 4988 11840 5040 11892
rect 5632 11840 5684 11892
rect 6552 11840 6604 11892
rect 6736 11840 6788 11892
rect 8208 11840 8260 11892
rect 2320 11704 2372 11756
rect 2872 11704 2924 11756
rect 3516 11704 3568 11756
rect 3976 11704 4028 11756
rect 4712 11747 4764 11756
rect 4712 11713 4721 11747
rect 4721 11713 4755 11747
rect 4755 11713 4764 11747
rect 4712 11704 4764 11713
rect 4988 11747 5040 11756
rect 4988 11713 4995 11747
rect 4995 11713 5029 11747
rect 5029 11713 5040 11747
rect 4988 11704 5040 11713
rect 5264 11772 5316 11824
rect 5908 11772 5960 11824
rect 6000 11772 6052 11824
rect 6276 11704 6328 11756
rect 7104 11747 7156 11756
rect 7104 11713 7113 11747
rect 7113 11713 7147 11747
rect 7147 11713 7156 11747
rect 7104 11704 7156 11713
rect 7380 11747 7432 11756
rect 7380 11713 7389 11747
rect 7389 11713 7423 11747
rect 7423 11713 7432 11747
rect 7380 11704 7432 11713
rect 8576 11747 8628 11756
rect 8576 11713 8585 11747
rect 8585 11713 8619 11747
rect 8619 11713 8628 11747
rect 8576 11704 8628 11713
rect 9588 11704 9640 11756
rect 10048 11747 10100 11756
rect 10048 11713 10057 11747
rect 10057 11713 10091 11747
rect 10091 11713 10100 11747
rect 10048 11704 10100 11713
rect 14464 11772 14516 11824
rect 14832 11772 14884 11824
rect 18512 11840 18564 11892
rect 19064 11840 19116 11892
rect 19524 11840 19576 11892
rect 19800 11840 19852 11892
rect 20352 11840 20404 11892
rect 20444 11840 20496 11892
rect 16580 11772 16632 11824
rect 3056 11636 3108 11688
rect 3240 11636 3292 11688
rect 3056 11500 3108 11552
rect 7012 11636 7064 11688
rect 7564 11679 7616 11688
rect 7564 11645 7573 11679
rect 7573 11645 7607 11679
rect 7607 11645 7616 11679
rect 7564 11636 7616 11645
rect 8300 11679 8352 11688
rect 8300 11645 8309 11679
rect 8309 11645 8343 11679
rect 8343 11645 8352 11679
rect 8300 11636 8352 11645
rect 9772 11636 9824 11688
rect 11888 11704 11940 11756
rect 13360 11747 13412 11756
rect 13360 11713 13369 11747
rect 13369 11713 13403 11747
rect 13403 11713 13412 11747
rect 13360 11704 13412 11713
rect 13544 11704 13596 11756
rect 13636 11747 13688 11756
rect 13636 11713 13645 11747
rect 13645 11713 13679 11747
rect 13679 11713 13688 11747
rect 13636 11704 13688 11713
rect 14280 11704 14332 11756
rect 15108 11704 15160 11756
rect 15752 11747 15804 11756
rect 15752 11713 15761 11747
rect 15761 11713 15795 11747
rect 15795 11713 15804 11747
rect 15752 11704 15804 11713
rect 11612 11636 11664 11688
rect 12532 11636 12584 11688
rect 16212 11704 16264 11756
rect 17040 11704 17092 11756
rect 17316 11704 17368 11756
rect 18696 11704 18748 11756
rect 19800 11704 19852 11756
rect 21180 11704 21232 11756
rect 12992 11568 13044 11620
rect 13084 11611 13136 11620
rect 13084 11577 13093 11611
rect 13093 11577 13127 11611
rect 13127 11577 13136 11611
rect 13084 11568 13136 11577
rect 18512 11636 18564 11688
rect 19984 11636 20036 11688
rect 16396 11568 16448 11620
rect 20996 11611 21048 11620
rect 20996 11577 21005 11611
rect 21005 11577 21039 11611
rect 21039 11577 21048 11611
rect 20996 11568 21048 11577
rect 5724 11500 5776 11552
rect 6644 11500 6696 11552
rect 7288 11500 7340 11552
rect 7932 11500 7984 11552
rect 8116 11500 8168 11552
rect 12348 11500 12400 11552
rect 13360 11500 13412 11552
rect 13636 11500 13688 11552
rect 16488 11500 16540 11552
rect 17868 11500 17920 11552
rect 18788 11500 18840 11552
rect 3549 11398 3601 11450
rect 3613 11398 3665 11450
rect 3677 11398 3729 11450
rect 3741 11398 3793 11450
rect 3805 11398 3857 11450
rect 8747 11398 8799 11450
rect 8811 11398 8863 11450
rect 8875 11398 8927 11450
rect 8939 11398 8991 11450
rect 9003 11398 9055 11450
rect 13945 11398 13997 11450
rect 14009 11398 14061 11450
rect 14073 11398 14125 11450
rect 14137 11398 14189 11450
rect 14201 11398 14253 11450
rect 19143 11398 19195 11450
rect 19207 11398 19259 11450
rect 19271 11398 19323 11450
rect 19335 11398 19387 11450
rect 19399 11398 19451 11450
rect 2228 11296 2280 11348
rect 940 11228 992 11280
rect 1584 11092 1636 11144
rect 3424 11296 3476 11348
rect 3608 11296 3660 11348
rect 3976 11296 4028 11348
rect 4068 11296 4120 11348
rect 4988 11228 5040 11280
rect 7104 11296 7156 11348
rect 8208 11296 8260 11348
rect 9036 11296 9088 11348
rect 9680 11296 9732 11348
rect 4252 11160 4304 11212
rect 5448 11160 5500 11212
rect 5540 11203 5592 11212
rect 5540 11169 5549 11203
rect 5549 11169 5583 11203
rect 5583 11169 5592 11203
rect 5540 11160 5592 11169
rect 6000 11160 6052 11212
rect 6460 11160 6512 11212
rect 940 11024 992 11076
rect 2412 11024 2464 11076
rect 4436 11092 4488 11144
rect 3056 11024 3108 11076
rect 3792 11024 3844 11076
rect 4160 11024 4212 11076
rect 4252 11067 4304 11076
rect 4252 11033 4261 11067
rect 4261 11033 4295 11067
rect 4295 11033 4304 11067
rect 4252 11024 4304 11033
rect 4804 11024 4856 11076
rect 6092 11135 6144 11144
rect 6092 11101 6101 11135
rect 6101 11101 6135 11135
rect 6135 11101 6144 11135
rect 6092 11092 6144 11101
rect 6828 11092 6880 11144
rect 7288 11160 7340 11212
rect 7748 11135 7800 11144
rect 7748 11101 7755 11135
rect 7755 11101 7789 11135
rect 7789 11101 7800 11135
rect 7748 11092 7800 11101
rect 9036 11092 9088 11144
rect 9772 11160 9824 11212
rect 10784 11296 10836 11348
rect 10876 11228 10928 11280
rect 11796 11271 11848 11280
rect 11796 11237 11805 11271
rect 11805 11237 11839 11271
rect 11839 11237 11848 11271
rect 11796 11228 11848 11237
rect 11336 11203 11388 11212
rect 11336 11169 11345 11203
rect 11345 11169 11379 11203
rect 11379 11169 11388 11203
rect 11336 11160 11388 11169
rect 12072 11296 12124 11348
rect 13360 11296 13412 11348
rect 12072 11203 12124 11212
rect 12072 11169 12081 11203
rect 12081 11169 12115 11203
rect 12115 11169 12124 11203
rect 12072 11160 12124 11169
rect 13544 11228 13596 11280
rect 10416 11135 10468 11144
rect 10416 11101 10425 11135
rect 10425 11101 10459 11135
rect 10459 11101 10468 11135
rect 10416 11092 10468 11101
rect 11244 11092 11296 11144
rect 13452 11160 13504 11212
rect 14096 11203 14148 11212
rect 14096 11169 14105 11203
rect 14105 11169 14139 11203
rect 14139 11169 14148 11203
rect 14096 11160 14148 11169
rect 12348 11135 12400 11144
rect 12348 11101 12357 11135
rect 12357 11101 12391 11135
rect 12391 11101 12400 11135
rect 12348 11092 12400 11101
rect 12992 11092 13044 11144
rect 11060 11067 11112 11076
rect 11060 11033 11069 11067
rect 11069 11033 11103 11067
rect 11103 11033 11112 11067
rect 11060 11024 11112 11033
rect 2872 10956 2924 11008
rect 6644 10956 6696 11008
rect 7012 10956 7064 11008
rect 10968 10956 11020 11008
rect 12072 10956 12124 11008
rect 13544 11024 13596 11076
rect 15292 11296 15344 11348
rect 15568 11203 15620 11212
rect 15568 11169 15577 11203
rect 15577 11169 15611 11203
rect 15611 11169 15620 11203
rect 15568 11160 15620 11169
rect 14924 11024 14976 11076
rect 15936 11092 15988 11144
rect 16580 11339 16632 11348
rect 16580 11305 16589 11339
rect 16589 11305 16623 11339
rect 16623 11305 16632 11339
rect 16580 11296 16632 11305
rect 17684 11296 17736 11348
rect 18420 11296 18472 11348
rect 19800 11339 19852 11348
rect 19800 11305 19809 11339
rect 19809 11305 19843 11339
rect 19843 11305 19852 11339
rect 19800 11296 19852 11305
rect 19340 11228 19392 11280
rect 19708 11228 19760 11280
rect 17776 11092 17828 11144
rect 17868 11135 17920 11144
rect 17868 11101 17877 11135
rect 17877 11101 17911 11135
rect 17911 11101 17920 11135
rect 17868 11092 17920 11101
rect 18328 11135 18380 11144
rect 18328 11101 18337 11135
rect 18337 11101 18371 11135
rect 18371 11101 18380 11135
rect 18328 11092 18380 11101
rect 18788 11092 18840 11144
rect 16304 11024 16356 11076
rect 13452 10956 13504 11008
rect 18144 10956 18196 11008
rect 19708 11135 19760 11144
rect 19708 11101 19717 11135
rect 19717 11101 19751 11135
rect 19751 11101 19760 11135
rect 19708 11092 19760 11101
rect 19708 10956 19760 11008
rect 21364 10999 21416 11008
rect 21364 10965 21373 10999
rect 21373 10965 21407 10999
rect 21407 10965 21416 10999
rect 21364 10956 21416 10965
rect 6148 10854 6200 10906
rect 6212 10854 6264 10906
rect 6276 10854 6328 10906
rect 6340 10854 6392 10906
rect 6404 10854 6456 10906
rect 11346 10854 11398 10906
rect 11410 10854 11462 10906
rect 11474 10854 11526 10906
rect 11538 10854 11590 10906
rect 11602 10854 11654 10906
rect 16544 10854 16596 10906
rect 16608 10854 16660 10906
rect 16672 10854 16724 10906
rect 16736 10854 16788 10906
rect 16800 10854 16852 10906
rect 21742 10854 21794 10906
rect 21806 10854 21858 10906
rect 21870 10854 21922 10906
rect 21934 10854 21986 10906
rect 21998 10854 22050 10906
rect 3792 10752 3844 10804
rect 6368 10752 6420 10804
rect 7656 10752 7708 10804
rect 8576 10752 8628 10804
rect 10416 10752 10468 10804
rect 11888 10752 11940 10804
rect 1216 10684 1268 10736
rect 3516 10659 3568 10668
rect 3516 10625 3525 10659
rect 3525 10625 3559 10659
rect 3559 10625 3568 10659
rect 3516 10616 3568 10625
rect 2412 10548 2464 10600
rect 2688 10548 2740 10600
rect 2872 10548 2924 10600
rect 3884 10548 3936 10600
rect 4436 10684 4488 10736
rect 9128 10684 9180 10736
rect 4712 10616 4764 10668
rect 5356 10659 5408 10668
rect 5356 10625 5390 10659
rect 5390 10625 5408 10659
rect 5356 10616 5408 10625
rect 5540 10659 5592 10668
rect 5540 10625 5549 10659
rect 5549 10625 5583 10659
rect 5583 10625 5592 10659
rect 5540 10616 5592 10625
rect 6828 10616 6880 10668
rect 1216 10480 1268 10532
rect 1768 10455 1820 10464
rect 1768 10421 1777 10455
rect 1777 10421 1811 10455
rect 1811 10421 1820 10455
rect 1768 10412 1820 10421
rect 3056 10480 3108 10532
rect 4988 10523 5040 10532
rect 4988 10489 4997 10523
rect 4997 10489 5031 10523
rect 5031 10489 5040 10523
rect 4988 10480 5040 10489
rect 9588 10616 9640 10668
rect 9680 10616 9732 10668
rect 10048 10659 10100 10668
rect 10048 10625 10057 10659
rect 10057 10625 10091 10659
rect 10091 10625 10100 10659
rect 10048 10616 10100 10625
rect 10232 10616 10284 10668
rect 10324 10659 10376 10668
rect 10324 10625 10331 10659
rect 10331 10625 10365 10659
rect 10365 10625 10376 10659
rect 13268 10752 13320 10804
rect 13452 10752 13504 10804
rect 14096 10752 14148 10804
rect 10324 10616 10376 10625
rect 13544 10659 13596 10668
rect 13544 10625 13553 10659
rect 13553 10625 13587 10659
rect 13587 10625 13596 10659
rect 13544 10616 13596 10625
rect 13636 10659 13688 10668
rect 14648 10752 14700 10804
rect 17040 10752 17092 10804
rect 17316 10752 17368 10804
rect 17776 10752 17828 10804
rect 19340 10752 19392 10804
rect 19800 10752 19852 10804
rect 19892 10752 19944 10804
rect 22192 10752 22244 10804
rect 13636 10625 13670 10659
rect 13670 10625 13688 10659
rect 13636 10616 13688 10625
rect 14740 10616 14792 10668
rect 19432 10659 19484 10668
rect 19432 10625 19441 10659
rect 19441 10625 19475 10659
rect 19475 10625 19484 10659
rect 19432 10616 19484 10625
rect 20720 10684 20772 10736
rect 7288 10591 7340 10600
rect 7288 10557 7297 10591
rect 7297 10557 7331 10591
rect 7331 10557 7340 10591
rect 7288 10548 7340 10557
rect 3608 10412 3660 10464
rect 4160 10455 4212 10464
rect 4160 10421 4169 10455
rect 4169 10421 4203 10455
rect 4203 10421 4212 10455
rect 4160 10412 4212 10421
rect 5724 10412 5776 10464
rect 5908 10412 5960 10464
rect 6460 10455 6512 10464
rect 6460 10421 6469 10455
rect 6469 10421 6503 10455
rect 6503 10421 6512 10455
rect 6460 10412 6512 10421
rect 6920 10455 6972 10464
rect 6920 10421 6929 10455
rect 6929 10421 6963 10455
rect 6963 10421 6972 10455
rect 6920 10412 6972 10421
rect 7564 10412 7616 10464
rect 11888 10548 11940 10600
rect 12532 10548 12584 10600
rect 13360 10548 13412 10600
rect 17224 10548 17276 10600
rect 9036 10412 9088 10464
rect 10324 10412 10376 10464
rect 13084 10412 13136 10464
rect 13728 10412 13780 10464
rect 15292 10480 15344 10532
rect 15752 10480 15804 10532
rect 18420 10548 18472 10600
rect 19524 10591 19576 10600
rect 19524 10557 19533 10591
rect 19533 10557 19567 10591
rect 19567 10557 19576 10591
rect 19524 10548 19576 10557
rect 18328 10455 18380 10464
rect 18328 10421 18337 10455
rect 18337 10421 18371 10455
rect 18371 10421 18380 10455
rect 18328 10412 18380 10421
rect 20352 10412 20404 10464
rect 3549 10310 3601 10362
rect 3613 10310 3665 10362
rect 3677 10310 3729 10362
rect 3741 10310 3793 10362
rect 3805 10310 3857 10362
rect 8747 10310 8799 10362
rect 8811 10310 8863 10362
rect 8875 10310 8927 10362
rect 8939 10310 8991 10362
rect 9003 10310 9055 10362
rect 13945 10310 13997 10362
rect 14009 10310 14061 10362
rect 14073 10310 14125 10362
rect 14137 10310 14189 10362
rect 14201 10310 14253 10362
rect 19143 10310 19195 10362
rect 19207 10310 19259 10362
rect 19271 10310 19323 10362
rect 19335 10310 19387 10362
rect 19399 10310 19451 10362
rect 1492 10208 1544 10260
rect 1676 10251 1728 10260
rect 1676 10217 1685 10251
rect 1685 10217 1719 10251
rect 1719 10217 1728 10251
rect 1676 10208 1728 10217
rect 2780 10208 2832 10260
rect 3332 10251 3384 10260
rect 3332 10217 3341 10251
rect 3341 10217 3375 10251
rect 3375 10217 3384 10251
rect 3332 10208 3384 10217
rect 3976 10251 4028 10260
rect 3976 10217 3985 10251
rect 3985 10217 4019 10251
rect 4019 10217 4028 10251
rect 3976 10208 4028 10217
rect 3056 10140 3108 10192
rect 6000 10208 6052 10260
rect 1400 10072 1452 10124
rect 2136 10004 2188 10056
rect 3056 10004 3108 10056
rect 4068 10072 4120 10124
rect 6644 10115 6696 10124
rect 6644 10081 6653 10115
rect 6653 10081 6687 10115
rect 6687 10081 6696 10115
rect 6644 10072 6696 10081
rect 4528 10004 4580 10056
rect 6368 10004 6420 10056
rect 6460 10004 6512 10056
rect 3884 9979 3936 9988
rect 3884 9945 3893 9979
rect 3893 9945 3927 9979
rect 3927 9945 3936 9979
rect 3884 9936 3936 9945
rect 2136 9868 2188 9920
rect 2872 9868 2924 9920
rect 4620 9868 4672 9920
rect 7012 10072 7064 10124
rect 7288 10115 7340 10124
rect 7288 10081 7297 10115
rect 7297 10081 7331 10115
rect 7331 10081 7340 10115
rect 7288 10072 7340 10081
rect 8300 10140 8352 10192
rect 10508 10208 10560 10260
rect 14556 10208 14608 10260
rect 15936 10208 15988 10260
rect 18052 10208 18104 10260
rect 18604 10208 18656 10260
rect 20260 10208 20312 10260
rect 20352 10208 20404 10260
rect 20904 10251 20956 10260
rect 20904 10217 20913 10251
rect 20913 10217 20947 10251
rect 20947 10217 20956 10251
rect 20904 10208 20956 10217
rect 7656 10115 7708 10124
rect 7656 10081 7690 10115
rect 7690 10081 7708 10115
rect 7656 10072 7708 10081
rect 10416 10072 10468 10124
rect 12072 10140 12124 10192
rect 11888 10115 11940 10124
rect 11888 10081 11897 10115
rect 11897 10081 11931 10115
rect 11931 10081 11940 10115
rect 11888 10072 11940 10081
rect 12348 10115 12400 10124
rect 12348 10081 12357 10115
rect 12357 10081 12391 10115
rect 12391 10081 12400 10115
rect 12348 10072 12400 10081
rect 18144 10183 18196 10192
rect 18144 10149 18153 10183
rect 18153 10149 18187 10183
rect 18187 10149 18196 10183
rect 18144 10140 18196 10149
rect 18420 10140 18472 10192
rect 12716 10072 12768 10124
rect 7840 10047 7892 10056
rect 7840 10013 7849 10047
rect 7849 10013 7883 10047
rect 7883 10013 7892 10047
rect 7840 10004 7892 10013
rect 8760 10047 8812 10056
rect 8760 10013 8769 10047
rect 8769 10013 8803 10047
rect 8803 10013 8812 10047
rect 8760 10004 8812 10013
rect 9680 10047 9732 10056
rect 9680 10013 9687 10047
rect 9687 10013 9721 10047
rect 9721 10013 9732 10047
rect 9680 10004 9732 10013
rect 10692 10004 10744 10056
rect 11704 10047 11756 10056
rect 11704 10013 11713 10047
rect 11713 10013 11747 10047
rect 11747 10013 11756 10047
rect 11704 10004 11756 10013
rect 11796 9936 11848 9988
rect 8484 9911 8536 9920
rect 8484 9877 8493 9911
rect 8493 9877 8527 9911
rect 8527 9877 8536 9911
rect 8484 9868 8536 9877
rect 9128 9868 9180 9920
rect 12900 10047 12952 10056
rect 12900 10013 12909 10047
rect 12909 10013 12943 10047
rect 12943 10013 12952 10047
rect 12900 10004 12952 10013
rect 13544 10115 13596 10124
rect 13544 10081 13553 10115
rect 13553 10081 13587 10115
rect 13587 10081 13596 10115
rect 13544 10072 13596 10081
rect 15108 10072 15160 10124
rect 16764 10072 16816 10124
rect 14372 9936 14424 9988
rect 14280 9868 14332 9920
rect 15016 9936 15068 9988
rect 15292 9979 15344 9988
rect 15292 9945 15301 9979
rect 15301 9945 15335 9979
rect 15335 9945 15344 9979
rect 15292 9936 15344 9945
rect 16028 10047 16080 10056
rect 16028 10013 16037 10047
rect 16037 10013 16071 10047
rect 16071 10013 16080 10047
rect 16028 10004 16080 10013
rect 16396 10004 16448 10056
rect 18144 10047 18196 10056
rect 18144 10013 18153 10047
rect 18153 10013 18187 10047
rect 18187 10013 18196 10047
rect 18144 10004 18196 10013
rect 18328 10004 18380 10056
rect 18788 10047 18840 10056
rect 18788 10013 18797 10047
rect 18797 10013 18831 10047
rect 18831 10013 18840 10047
rect 18788 10004 18840 10013
rect 15752 9868 15804 9920
rect 17684 9868 17736 9920
rect 19064 10047 19116 10056
rect 19064 10013 19073 10047
rect 19073 10013 19107 10047
rect 19107 10013 19116 10047
rect 19064 10004 19116 10013
rect 19248 10047 19300 10056
rect 19248 10013 19257 10047
rect 19257 10013 19291 10047
rect 19291 10013 19300 10047
rect 19248 10004 19300 10013
rect 19800 9936 19852 9988
rect 21180 9979 21232 9988
rect 21180 9945 21189 9979
rect 21189 9945 21223 9979
rect 21223 9945 21232 9979
rect 21180 9936 21232 9945
rect 22284 9936 22336 9988
rect 20260 9911 20312 9920
rect 20260 9877 20269 9911
rect 20269 9877 20303 9911
rect 20303 9877 20312 9911
rect 20260 9868 20312 9877
rect 20536 9868 20588 9920
rect 6148 9766 6200 9818
rect 6212 9766 6264 9818
rect 6276 9766 6328 9818
rect 6340 9766 6392 9818
rect 6404 9766 6456 9818
rect 11346 9766 11398 9818
rect 11410 9766 11462 9818
rect 11474 9766 11526 9818
rect 11538 9766 11590 9818
rect 11602 9766 11654 9818
rect 16544 9766 16596 9818
rect 16608 9766 16660 9818
rect 16672 9766 16724 9818
rect 16736 9766 16788 9818
rect 16800 9766 16852 9818
rect 21742 9766 21794 9818
rect 21806 9766 21858 9818
rect 21870 9766 21922 9818
rect 21934 9766 21986 9818
rect 21998 9766 22050 9818
rect 3056 9664 3108 9716
rect 5080 9664 5132 9716
rect 6644 9664 6696 9716
rect 7564 9664 7616 9716
rect 1492 9639 1544 9648
rect 1492 9605 1501 9639
rect 1501 9605 1535 9639
rect 1535 9605 1544 9639
rect 1492 9596 1544 9605
rect 1952 9596 2004 9648
rect 8484 9664 8536 9716
rect 2228 9571 2280 9580
rect 2228 9537 2237 9571
rect 2237 9537 2271 9571
rect 2271 9537 2280 9571
rect 2228 9528 2280 9537
rect 2504 9528 2556 9580
rect 3516 9528 3568 9580
rect 4712 9528 4764 9580
rect 5264 9571 5316 9580
rect 5264 9537 5273 9571
rect 5273 9537 5307 9571
rect 5307 9537 5316 9571
rect 5264 9528 5316 9537
rect 5448 9528 5500 9580
rect 6552 9528 6604 9580
rect 6920 9528 6972 9580
rect 1584 9460 1636 9512
rect 1860 9460 1912 9512
rect 3976 9460 4028 9512
rect 4436 9460 4488 9512
rect 4620 9460 4672 9512
rect 5540 9503 5592 9512
rect 5540 9469 5549 9503
rect 5549 9469 5583 9503
rect 5583 9469 5592 9503
rect 5540 9460 5592 9469
rect 5724 9460 5776 9512
rect 7656 9571 7708 9580
rect 7656 9537 7663 9571
rect 7663 9537 7697 9571
rect 7697 9537 7708 9571
rect 7656 9528 7708 9537
rect 7748 9528 7800 9580
rect 10508 9664 10560 9716
rect 9128 9528 9180 9580
rect 9956 9571 10008 9580
rect 9956 9537 9965 9571
rect 9965 9537 9999 9571
rect 9999 9537 10008 9571
rect 9956 9528 10008 9537
rect 10600 9528 10652 9580
rect 11704 9528 11756 9580
rect 2504 9392 2556 9444
rect 2872 9392 2924 9444
rect 3056 9435 3108 9444
rect 3056 9401 3065 9435
rect 3065 9401 3099 9435
rect 3099 9401 3108 9435
rect 3056 9392 3108 9401
rect 4068 9392 4120 9444
rect 4252 9324 4304 9376
rect 4804 9392 4856 9444
rect 5080 9392 5132 9444
rect 8300 9324 8352 9376
rect 13268 9664 13320 9716
rect 13820 9596 13872 9648
rect 14280 9596 14332 9648
rect 14832 9639 14884 9648
rect 14832 9605 14841 9639
rect 14841 9605 14875 9639
rect 14875 9605 14884 9639
rect 14832 9596 14884 9605
rect 13268 9571 13320 9580
rect 13268 9537 13277 9571
rect 13277 9537 13311 9571
rect 13311 9537 13320 9571
rect 13268 9528 13320 9537
rect 15016 9596 15068 9648
rect 15292 9596 15344 9648
rect 15568 9664 15620 9716
rect 16028 9664 16080 9716
rect 11888 9460 11940 9512
rect 12348 9460 12400 9512
rect 12072 9392 12124 9444
rect 15200 9571 15252 9580
rect 15200 9537 15209 9571
rect 15209 9537 15243 9571
rect 15243 9537 15252 9571
rect 15200 9528 15252 9537
rect 15752 9596 15804 9648
rect 16212 9596 16264 9648
rect 16120 9528 16172 9580
rect 16304 9528 16356 9580
rect 18604 9664 18656 9716
rect 18052 9571 18104 9580
rect 18052 9537 18086 9571
rect 18086 9537 18104 9571
rect 18052 9528 18104 9537
rect 18604 9528 18656 9580
rect 19156 9528 19208 9580
rect 19524 9664 19576 9716
rect 19616 9596 19668 9648
rect 19984 9596 20036 9648
rect 19800 9571 19852 9580
rect 19800 9537 19807 9571
rect 19807 9537 19841 9571
rect 19841 9537 19852 9571
rect 19800 9528 19852 9537
rect 19892 9528 19944 9580
rect 20168 9528 20220 9580
rect 20260 9528 20312 9580
rect 21088 9571 21140 9580
rect 21088 9537 21097 9571
rect 21097 9537 21131 9571
rect 21131 9537 21140 9571
rect 21088 9528 21140 9537
rect 21272 9528 21324 9580
rect 15292 9460 15344 9512
rect 12716 9435 12768 9444
rect 12716 9401 12725 9435
rect 12725 9401 12759 9435
rect 12759 9401 12768 9435
rect 12716 9392 12768 9401
rect 14556 9392 14608 9444
rect 17776 9503 17828 9512
rect 17776 9469 17785 9503
rect 17785 9469 17819 9503
rect 17819 9469 17828 9503
rect 17776 9460 17828 9469
rect 16212 9392 16264 9444
rect 9680 9324 9732 9376
rect 9864 9324 9916 9376
rect 10324 9324 10376 9376
rect 10692 9367 10744 9376
rect 10692 9333 10701 9367
rect 10701 9333 10735 9367
rect 10735 9333 10744 9367
rect 10692 9324 10744 9333
rect 11336 9324 11388 9376
rect 12256 9324 12308 9376
rect 13452 9324 13504 9376
rect 17224 9324 17276 9376
rect 18788 9324 18840 9376
rect 20352 9392 20404 9444
rect 22284 9324 22336 9376
rect 3549 9222 3601 9274
rect 3613 9222 3665 9274
rect 3677 9222 3729 9274
rect 3741 9222 3793 9274
rect 3805 9222 3857 9274
rect 8747 9222 8799 9274
rect 8811 9222 8863 9274
rect 8875 9222 8927 9274
rect 8939 9222 8991 9274
rect 9003 9222 9055 9274
rect 13945 9222 13997 9274
rect 14009 9222 14061 9274
rect 14073 9222 14125 9274
rect 14137 9222 14189 9274
rect 14201 9222 14253 9274
rect 19143 9222 19195 9274
rect 19207 9222 19259 9274
rect 19271 9222 19323 9274
rect 19335 9222 19387 9274
rect 19399 9222 19451 9274
rect 1768 9163 1820 9172
rect 1768 9129 1777 9163
rect 1777 9129 1811 9163
rect 1811 9129 1820 9163
rect 1768 9120 1820 9129
rect 4068 9120 4120 9172
rect 4528 9120 4580 9172
rect 5632 9120 5684 9172
rect 6644 9120 6696 9172
rect 7840 9120 7892 9172
rect 1400 8984 1452 9036
rect 2136 9027 2188 9036
rect 2136 8993 2145 9027
rect 2145 8993 2179 9027
rect 2179 8993 2188 9027
rect 2136 8984 2188 8993
rect 3792 9027 3844 9036
rect 3792 8993 3801 9027
rect 3801 8993 3835 9027
rect 3835 8993 3844 9027
rect 3792 8984 3844 8993
rect 4528 8984 4580 9036
rect 5448 8984 5500 9036
rect 6920 8984 6972 9036
rect 8484 8984 8536 9036
rect 9496 9120 9548 9172
rect 10048 9163 10100 9172
rect 10048 9129 10057 9163
rect 10057 9129 10091 9163
rect 10091 9129 10100 9163
rect 10048 9120 10100 9129
rect 2504 8916 2556 8968
rect 3424 8916 3476 8968
rect 3608 8916 3660 8968
rect 4068 8959 4120 8968
rect 4068 8925 4075 8959
rect 4075 8925 4109 8959
rect 4109 8925 4120 8959
rect 4068 8916 4120 8925
rect 4160 8916 4212 8968
rect 6828 8916 6880 8968
rect 7656 8916 7708 8968
rect 8392 8916 8444 8968
rect 1492 8891 1544 8900
rect 1492 8857 1501 8891
rect 1501 8857 1535 8891
rect 1535 8857 1544 8891
rect 1492 8848 1544 8857
rect 2688 8848 2740 8900
rect 10324 8848 10376 8900
rect 480 8780 532 8832
rect 5908 8780 5960 8832
rect 6644 8823 6696 8832
rect 6644 8789 6653 8823
rect 6653 8789 6687 8823
rect 6687 8789 6696 8823
rect 6644 8780 6696 8789
rect 6920 8780 6972 8832
rect 7104 8780 7156 8832
rect 9220 8780 9272 8832
rect 9680 8780 9732 8832
rect 10416 8780 10468 8832
rect 10784 8916 10836 8968
rect 11336 8780 11388 8832
rect 12716 9120 12768 9172
rect 12900 9120 12952 9172
rect 11796 8984 11848 9036
rect 15108 9163 15160 9172
rect 15108 9129 15117 9163
rect 15117 9129 15151 9163
rect 15151 9129 15160 9163
rect 15108 9120 15160 9129
rect 15200 9120 15252 9172
rect 14832 9052 14884 9104
rect 12256 8959 12308 8968
rect 12256 8925 12263 8959
rect 12263 8925 12297 8959
rect 12297 8925 12308 8959
rect 12256 8916 12308 8925
rect 12348 8848 12400 8900
rect 13084 8848 13136 8900
rect 15108 8848 15160 8900
rect 15568 8848 15620 8900
rect 15844 8916 15896 8968
rect 16212 8848 16264 8900
rect 12256 8780 12308 8832
rect 13452 8780 13504 8832
rect 17132 9120 17184 9172
rect 17224 9120 17276 9172
rect 17960 9120 18012 9172
rect 18144 9120 18196 9172
rect 19340 9120 19392 9172
rect 21272 9120 21324 9172
rect 21364 9120 21416 9172
rect 21456 9163 21508 9172
rect 21456 9129 21465 9163
rect 21465 9129 21499 9163
rect 21499 9129 21508 9163
rect 21456 9120 21508 9129
rect 17132 8929 17184 8968
rect 17132 8916 17157 8929
rect 17157 8916 17184 8929
rect 17224 8916 17276 8968
rect 17960 8916 18012 8968
rect 20996 9095 21048 9104
rect 20996 9061 21005 9095
rect 21005 9061 21039 9095
rect 21039 9061 21048 9095
rect 20996 9052 21048 9061
rect 18972 8959 19024 8968
rect 18972 8925 18981 8959
rect 18981 8925 19015 8959
rect 19015 8925 19024 8959
rect 18972 8916 19024 8925
rect 19432 8916 19484 8968
rect 19524 8959 19576 8968
rect 19524 8925 19533 8959
rect 19533 8925 19567 8959
rect 19567 8925 19576 8959
rect 19524 8916 19576 8925
rect 16948 8780 17000 8832
rect 17132 8780 17184 8832
rect 19984 8848 20036 8900
rect 20168 8848 20220 8900
rect 18604 8823 18656 8832
rect 18604 8789 18613 8823
rect 18613 8789 18647 8823
rect 18647 8789 18656 8823
rect 18604 8780 18656 8789
rect 19432 8780 19484 8832
rect 21272 8959 21324 8968
rect 21272 8925 21281 8959
rect 21281 8925 21315 8959
rect 21315 8925 21324 8959
rect 21272 8916 21324 8925
rect 20260 8780 20312 8832
rect 20628 8823 20680 8832
rect 20628 8789 20637 8823
rect 20637 8789 20671 8823
rect 20671 8789 20680 8823
rect 20628 8780 20680 8789
rect 6148 8678 6200 8730
rect 6212 8678 6264 8730
rect 6276 8678 6328 8730
rect 6340 8678 6392 8730
rect 6404 8678 6456 8730
rect 11346 8678 11398 8730
rect 11410 8678 11462 8730
rect 11474 8678 11526 8730
rect 11538 8678 11590 8730
rect 11602 8678 11654 8730
rect 16544 8678 16596 8730
rect 16608 8678 16660 8730
rect 16672 8678 16724 8730
rect 16736 8678 16788 8730
rect 16800 8678 16852 8730
rect 21742 8678 21794 8730
rect 21806 8678 21858 8730
rect 21870 8678 21922 8730
rect 21934 8678 21986 8730
rect 21998 8678 22050 8730
rect 2964 8576 3016 8628
rect 3332 8576 3384 8628
rect 4252 8508 4304 8560
rect 4620 8576 4672 8628
rect 7104 8576 7156 8628
rect 7288 8576 7340 8628
rect 4896 8508 4948 8560
rect 1492 8483 1544 8492
rect 1492 8449 1501 8483
rect 1501 8449 1535 8483
rect 1535 8449 1544 8483
rect 1492 8440 1544 8449
rect 2412 8440 2464 8492
rect 2688 8440 2740 8492
rect 3424 8440 3476 8492
rect 3516 8483 3568 8492
rect 3516 8449 3525 8483
rect 3525 8449 3559 8483
rect 3559 8449 3568 8483
rect 3516 8440 3568 8449
rect 4160 8440 4212 8492
rect 5540 8440 5592 8492
rect 2872 8372 2924 8424
rect 3884 8372 3936 8424
rect 2964 8347 3016 8356
rect 2964 8313 2973 8347
rect 2973 8313 3007 8347
rect 3007 8313 3016 8347
rect 2964 8304 3016 8313
rect 4252 8304 4304 8356
rect 7564 8508 7616 8560
rect 8576 8576 8628 8628
rect 9312 8576 9364 8628
rect 9956 8576 10008 8628
rect 10324 8576 10376 8628
rect 6276 8440 6328 8492
rect 8484 8508 8536 8560
rect 11704 8576 11756 8628
rect 12440 8576 12492 8628
rect 13268 8576 13320 8628
rect 15292 8619 15344 8628
rect 15292 8585 15301 8619
rect 15301 8585 15335 8619
rect 15335 8585 15344 8619
rect 15292 8576 15344 8585
rect 9496 8440 9548 8492
rect 10324 8483 10376 8492
rect 10324 8449 10333 8483
rect 10333 8449 10367 8483
rect 10367 8449 10376 8483
rect 10324 8440 10376 8449
rect 11704 8440 11756 8492
rect 11888 8440 11940 8492
rect 12090 8440 12142 8492
rect 13084 8440 13136 8492
rect 13268 8440 13320 8492
rect 14188 8440 14240 8492
rect 14464 8440 14516 8492
rect 17684 8508 17736 8560
rect 18972 8576 19024 8628
rect 20628 8576 20680 8628
rect 21180 8576 21232 8628
rect 17960 8440 18012 8492
rect 19892 8508 19944 8560
rect 20352 8508 20404 8560
rect 19800 8440 19852 8492
rect 9680 8372 9732 8424
rect 10140 8372 10192 8424
rect 10508 8372 10560 8424
rect 10600 8415 10652 8424
rect 10600 8381 10609 8415
rect 10609 8381 10643 8415
rect 10643 8381 10652 8415
rect 10600 8372 10652 8381
rect 12256 8372 12308 8424
rect 12900 8415 12952 8424
rect 12900 8381 12909 8415
rect 12909 8381 12943 8415
rect 12943 8381 12952 8415
rect 12900 8372 12952 8381
rect 15384 8372 15436 8424
rect 16304 8372 16356 8424
rect 16764 8372 16816 8424
rect 18328 8372 18380 8424
rect 18512 8372 18564 8424
rect 19984 8415 20036 8424
rect 19984 8381 19993 8415
rect 19993 8381 20027 8415
rect 20027 8381 20036 8415
rect 19984 8372 20036 8381
rect 4620 8236 4672 8288
rect 5264 8236 5316 8288
rect 6736 8236 6788 8288
rect 6920 8236 6972 8288
rect 7840 8236 7892 8288
rect 8024 8236 8076 8288
rect 8944 8236 8996 8288
rect 9312 8236 9364 8288
rect 9496 8236 9548 8288
rect 11152 8236 11204 8288
rect 11612 8236 11664 8288
rect 11796 8236 11848 8288
rect 14280 8236 14332 8288
rect 14372 8236 14424 8288
rect 15476 8236 15528 8288
rect 16304 8236 16356 8288
rect 16672 8279 16724 8288
rect 16672 8245 16681 8279
rect 16681 8245 16715 8279
rect 16715 8245 16724 8279
rect 16672 8236 16724 8245
rect 16948 8236 17000 8288
rect 19616 8347 19668 8356
rect 19616 8313 19625 8347
rect 19625 8313 19659 8347
rect 19659 8313 19668 8347
rect 19616 8304 19668 8313
rect 21180 8304 21232 8356
rect 20352 8236 20404 8288
rect 3549 8134 3601 8186
rect 3613 8134 3665 8186
rect 3677 8134 3729 8186
rect 3741 8134 3793 8186
rect 3805 8134 3857 8186
rect 8747 8134 8799 8186
rect 8811 8134 8863 8186
rect 8875 8134 8927 8186
rect 8939 8134 8991 8186
rect 9003 8134 9055 8186
rect 13945 8134 13997 8186
rect 14009 8134 14061 8186
rect 14073 8134 14125 8186
rect 14137 8134 14189 8186
rect 14201 8134 14253 8186
rect 19143 8134 19195 8186
rect 19207 8134 19259 8186
rect 19271 8134 19323 8186
rect 19335 8134 19387 8186
rect 19399 8134 19451 8186
rect 3240 8032 3292 8084
rect 4160 8032 4212 8084
rect 4620 8032 4672 8084
rect 4068 7964 4120 8016
rect 4988 8032 5040 8084
rect 5632 8032 5684 8084
rect 6368 8032 6420 8084
rect 6920 8032 6972 8084
rect 7288 8032 7340 8084
rect 7748 8032 7800 8084
rect 8576 8032 8628 8084
rect 8852 8032 8904 8084
rect 5816 7896 5868 7948
rect 6644 7964 6696 8016
rect 7840 7964 7892 8016
rect 8116 7964 8168 8016
rect 8392 8007 8444 8016
rect 8392 7973 8401 8007
rect 8401 7973 8435 8007
rect 8435 7973 8444 8007
rect 8392 7964 8444 7973
rect 10600 8075 10652 8084
rect 10600 8041 10609 8075
rect 10609 8041 10643 8075
rect 10643 8041 10652 8075
rect 10600 8032 10652 8041
rect 15292 8032 15344 8084
rect 11704 7964 11756 8016
rect 11796 8007 11848 8016
rect 11796 7973 11805 8007
rect 11805 7973 11839 8007
rect 11839 7973 11848 8007
rect 11796 7964 11848 7973
rect 12900 7964 12952 8016
rect 13544 7964 13596 8016
rect 15108 7964 15160 8016
rect 2504 7828 2556 7880
rect 2688 7828 2740 7880
rect 3792 7828 3844 7880
rect 4068 7871 4120 7880
rect 4068 7837 4077 7871
rect 4077 7837 4111 7871
rect 4111 7837 4120 7871
rect 4068 7828 4120 7837
rect 4528 7828 4580 7880
rect 6368 7871 6420 7880
rect 6368 7837 6377 7871
rect 6377 7837 6411 7871
rect 6411 7837 6420 7871
rect 6368 7828 6420 7837
rect 7104 7871 7156 7880
rect 7104 7837 7113 7871
rect 7113 7837 7147 7871
rect 7147 7837 7156 7871
rect 7104 7828 7156 7837
rect 7286 7828 7338 7880
rect 7380 7871 7432 7880
rect 7380 7837 7389 7871
rect 7389 7837 7423 7871
rect 7423 7837 7432 7871
rect 7380 7828 7432 7837
rect 8208 7828 8260 7880
rect 8300 7871 8352 7880
rect 8300 7837 8309 7871
rect 8309 7837 8343 7871
rect 8343 7837 8352 7871
rect 8300 7828 8352 7837
rect 8392 7828 8444 7880
rect 12072 7939 12124 7948
rect 12072 7905 12081 7939
rect 12081 7905 12115 7939
rect 12115 7905 12124 7939
rect 12072 7896 12124 7905
rect 12348 7939 12400 7948
rect 12348 7905 12357 7939
rect 12357 7905 12391 7939
rect 12391 7905 12400 7939
rect 12348 7896 12400 7905
rect 17960 8032 18012 8084
rect 18512 8032 18564 8084
rect 17684 7964 17736 8016
rect 17868 7964 17920 8016
rect 18052 7964 18104 8016
rect 21088 8032 21140 8084
rect 22100 7964 22152 8016
rect 2044 7692 2096 7744
rect 2872 7692 2924 7744
rect 3884 7692 3936 7744
rect 5540 7760 5592 7812
rect 4712 7692 4764 7744
rect 8760 7760 8812 7812
rect 10784 7760 10836 7812
rect 11244 7760 11296 7812
rect 8024 7735 8076 7744
rect 8024 7701 8033 7735
rect 8033 7701 8067 7735
rect 8067 7701 8076 7735
rect 8024 7692 8076 7701
rect 8116 7735 8168 7744
rect 8116 7701 8125 7735
rect 8125 7701 8159 7735
rect 8159 7701 8168 7735
rect 8116 7692 8168 7701
rect 8392 7692 8444 7744
rect 10048 7692 10100 7744
rect 10968 7692 11020 7744
rect 12164 7871 12216 7880
rect 12164 7837 12198 7871
rect 12198 7837 12216 7871
rect 12164 7828 12216 7837
rect 13728 7871 13780 7880
rect 13728 7837 13737 7871
rect 13737 7837 13771 7871
rect 13771 7837 13780 7871
rect 13728 7828 13780 7837
rect 14004 7828 14056 7880
rect 14096 7871 14148 7880
rect 14096 7837 14105 7871
rect 14105 7837 14139 7871
rect 14139 7837 14148 7871
rect 14096 7828 14148 7837
rect 16304 7939 16356 7948
rect 16304 7905 16313 7939
rect 16313 7905 16347 7939
rect 16347 7905 16356 7939
rect 16304 7896 16356 7905
rect 19432 7939 19484 7948
rect 19432 7905 19441 7939
rect 19441 7905 19475 7939
rect 19475 7905 19484 7939
rect 19432 7896 19484 7905
rect 11980 7692 12032 7744
rect 12900 7692 12952 7744
rect 12992 7735 13044 7744
rect 12992 7701 13001 7735
rect 13001 7701 13035 7735
rect 13035 7701 13044 7735
rect 12992 7692 13044 7701
rect 13820 7692 13872 7744
rect 15016 7692 15068 7744
rect 16672 7828 16724 7880
rect 17776 7828 17828 7880
rect 15936 7760 15988 7812
rect 16212 7803 16264 7812
rect 16212 7769 16221 7803
rect 16221 7769 16255 7803
rect 16255 7769 16264 7803
rect 16212 7760 16264 7769
rect 16948 7760 17000 7812
rect 16028 7692 16080 7744
rect 17224 7692 17276 7744
rect 17500 7692 17552 7744
rect 18512 7871 18564 7880
rect 18512 7837 18521 7871
rect 18521 7837 18555 7871
rect 18555 7837 18564 7871
rect 18512 7828 18564 7837
rect 20720 7828 20772 7880
rect 19340 7760 19392 7812
rect 19984 7692 20036 7744
rect 20812 7735 20864 7744
rect 20812 7701 20821 7735
rect 20821 7701 20855 7735
rect 20855 7701 20864 7735
rect 20812 7692 20864 7701
rect 6148 7590 6200 7642
rect 6212 7590 6264 7642
rect 6276 7590 6328 7642
rect 6340 7590 6392 7642
rect 6404 7590 6456 7642
rect 11346 7590 11398 7642
rect 11410 7590 11462 7642
rect 11474 7590 11526 7642
rect 11538 7590 11590 7642
rect 11602 7590 11654 7642
rect 16544 7590 16596 7642
rect 16608 7590 16660 7642
rect 16672 7590 16724 7642
rect 16736 7590 16788 7642
rect 16800 7590 16852 7642
rect 21742 7590 21794 7642
rect 21806 7590 21858 7642
rect 21870 7590 21922 7642
rect 21934 7590 21986 7642
rect 21998 7590 22050 7642
rect 1860 7531 1912 7540
rect 1860 7497 1869 7531
rect 1869 7497 1903 7531
rect 1903 7497 1912 7531
rect 1860 7488 1912 7497
rect 4068 7488 4120 7540
rect 4160 7488 4212 7540
rect 4436 7531 4488 7540
rect 4436 7497 4445 7531
rect 4445 7497 4479 7531
rect 4479 7497 4488 7531
rect 4436 7488 4488 7497
rect 5540 7488 5592 7540
rect 7380 7488 7432 7540
rect 8300 7488 8352 7540
rect 1308 7420 1360 7472
rect 1492 7352 1544 7404
rect 3240 7395 3292 7404
rect 3240 7361 3249 7395
rect 3249 7361 3283 7395
rect 3283 7361 3292 7395
rect 3240 7352 3292 7361
rect 3976 7352 4028 7404
rect 5356 7420 5408 7472
rect 1308 7148 1360 7200
rect 1584 7284 1636 7336
rect 2228 7327 2280 7336
rect 2228 7293 2237 7327
rect 2237 7293 2271 7327
rect 2271 7293 2280 7327
rect 2228 7284 2280 7293
rect 2596 7216 2648 7268
rect 2320 7148 2372 7200
rect 3884 7216 3936 7268
rect 4712 7352 4764 7404
rect 4988 7352 5040 7404
rect 4528 7284 4580 7336
rect 5540 7352 5592 7404
rect 8760 7395 8812 7404
rect 8760 7361 8769 7395
rect 8769 7361 8803 7395
rect 8803 7361 8812 7395
rect 8760 7352 8812 7361
rect 10508 7488 10560 7540
rect 11704 7488 11756 7540
rect 11244 7420 11296 7472
rect 12348 7488 12400 7540
rect 12900 7488 12952 7540
rect 15752 7488 15804 7540
rect 16028 7488 16080 7540
rect 16120 7531 16172 7540
rect 16120 7497 16129 7531
rect 16129 7497 16163 7531
rect 16163 7497 16172 7531
rect 16120 7488 16172 7497
rect 17224 7488 17276 7540
rect 17500 7488 17552 7540
rect 17960 7531 18012 7540
rect 17960 7497 17969 7531
rect 17969 7497 18003 7531
rect 18003 7497 18012 7531
rect 17960 7488 18012 7497
rect 18052 7488 18104 7540
rect 18236 7488 18288 7540
rect 18604 7488 18656 7540
rect 19524 7488 19576 7540
rect 21456 7488 21508 7540
rect 4712 7148 4764 7200
rect 6000 7148 6052 7200
rect 7748 7327 7800 7336
rect 7748 7293 7757 7327
rect 7757 7293 7791 7327
rect 7791 7293 7800 7327
rect 7748 7284 7800 7293
rect 8300 7284 8352 7336
rect 10416 7395 10468 7404
rect 10416 7361 10425 7395
rect 10425 7361 10459 7395
rect 10459 7361 10468 7395
rect 10416 7352 10468 7361
rect 10508 7395 10560 7404
rect 10508 7361 10542 7395
rect 10542 7361 10560 7395
rect 10508 7352 10560 7361
rect 11704 7352 11756 7404
rect 12440 7352 12492 7404
rect 13268 7352 13320 7404
rect 14556 7395 14608 7404
rect 14556 7361 14565 7395
rect 14565 7361 14599 7395
rect 14599 7361 14608 7395
rect 14556 7352 14608 7361
rect 15016 7395 15068 7404
rect 15016 7361 15025 7395
rect 15025 7361 15059 7395
rect 15059 7361 15068 7395
rect 15016 7352 15068 7361
rect 7932 7216 7984 7268
rect 8208 7259 8260 7268
rect 8208 7225 8217 7259
rect 8217 7225 8251 7259
rect 8251 7225 8260 7259
rect 8208 7216 8260 7225
rect 9312 7216 9364 7268
rect 9680 7327 9732 7336
rect 9680 7293 9689 7327
rect 9689 7293 9723 7327
rect 9723 7293 9732 7327
rect 9680 7284 9732 7293
rect 10048 7284 10100 7336
rect 10692 7327 10744 7336
rect 10692 7293 10701 7327
rect 10701 7293 10735 7327
rect 10735 7293 10744 7327
rect 10692 7284 10744 7293
rect 15844 7284 15896 7336
rect 10140 7259 10192 7268
rect 10140 7225 10149 7259
rect 10149 7225 10183 7259
rect 10183 7225 10192 7259
rect 10140 7216 10192 7225
rect 6828 7148 6880 7200
rect 7748 7148 7800 7200
rect 11244 7148 11296 7200
rect 12440 7216 12492 7268
rect 13912 7216 13964 7268
rect 14280 7216 14332 7268
rect 15568 7216 15620 7268
rect 16028 7216 16080 7268
rect 11888 7148 11940 7200
rect 15844 7148 15896 7200
rect 16304 7352 16356 7404
rect 17132 7352 17184 7404
rect 18880 7395 18932 7404
rect 18880 7361 18887 7395
rect 18887 7361 18921 7395
rect 18921 7361 18932 7395
rect 18880 7352 18932 7361
rect 19432 7352 19484 7404
rect 19892 7352 19944 7404
rect 20076 7352 20128 7404
rect 18052 7284 18104 7336
rect 19800 7284 19852 7336
rect 16396 7216 16448 7268
rect 18328 7216 18380 7268
rect 17776 7148 17828 7200
rect 19984 7148 20036 7200
rect 21364 7191 21416 7200
rect 21364 7157 21373 7191
rect 21373 7157 21407 7191
rect 21407 7157 21416 7191
rect 21364 7148 21416 7157
rect 3549 7046 3601 7098
rect 3613 7046 3665 7098
rect 3677 7046 3729 7098
rect 3741 7046 3793 7098
rect 3805 7046 3857 7098
rect 8747 7046 8799 7098
rect 8811 7046 8863 7098
rect 8875 7046 8927 7098
rect 8939 7046 8991 7098
rect 9003 7046 9055 7098
rect 13945 7046 13997 7098
rect 14009 7046 14061 7098
rect 14073 7046 14125 7098
rect 14137 7046 14189 7098
rect 14201 7046 14253 7098
rect 19143 7046 19195 7098
rect 19207 7046 19259 7098
rect 19271 7046 19323 7098
rect 19335 7046 19387 7098
rect 19399 7046 19451 7098
rect 3332 6944 3384 6996
rect 6828 6944 6880 6996
rect 6920 6944 6972 6996
rect 8208 6944 8260 6996
rect 8668 6944 8720 6996
rect 4252 6876 4304 6928
rect 1492 6808 1544 6860
rect 1952 6740 2004 6792
rect 4712 6808 4764 6860
rect 4804 6851 4856 6860
rect 4804 6817 4813 6851
rect 4813 6817 4847 6851
rect 4847 6817 4856 6851
rect 4804 6808 4856 6817
rect 6000 6919 6052 6928
rect 6000 6885 6009 6919
rect 6009 6885 6043 6919
rect 6043 6885 6052 6919
rect 6000 6876 6052 6885
rect 5908 6808 5960 6860
rect 8300 6876 8352 6928
rect 10416 6944 10468 6996
rect 10692 6944 10744 6996
rect 11796 6944 11848 6996
rect 12900 6944 12952 6996
rect 14556 6944 14608 6996
rect 11704 6876 11756 6928
rect 15844 6944 15896 6996
rect 16028 6876 16080 6928
rect 18052 6944 18104 6996
rect 18512 6944 18564 6996
rect 19248 6876 19300 6928
rect 3332 6740 3384 6792
rect 3700 6740 3752 6792
rect 4252 6740 4304 6792
rect 4528 6740 4580 6792
rect 5356 6783 5408 6792
rect 5356 6749 5365 6783
rect 5365 6749 5399 6783
rect 5399 6749 5408 6783
rect 5356 6740 5408 6749
rect 6092 6783 6144 6792
rect 6092 6749 6101 6783
rect 6101 6749 6135 6783
rect 6135 6749 6144 6783
rect 6092 6740 6144 6749
rect 6736 6740 6788 6792
rect 2504 6604 2556 6656
rect 3424 6604 3476 6656
rect 7380 6672 7432 6724
rect 8484 6808 8536 6860
rect 9312 6808 9364 6860
rect 10968 6851 11020 6860
rect 10968 6817 10977 6851
rect 10977 6817 11011 6851
rect 11011 6817 11020 6851
rect 10968 6808 11020 6817
rect 9956 6740 10008 6792
rect 10784 6740 10836 6792
rect 12256 6740 12308 6792
rect 13728 6783 13780 6792
rect 13728 6749 13737 6783
rect 13737 6749 13771 6783
rect 13771 6749 13780 6783
rect 13728 6740 13780 6749
rect 14096 6783 14148 6792
rect 14096 6749 14105 6783
rect 14105 6749 14139 6783
rect 14139 6749 14148 6783
rect 14096 6740 14148 6749
rect 4988 6604 5040 6656
rect 7656 6604 7708 6656
rect 13268 6672 13320 6724
rect 10968 6604 11020 6656
rect 11888 6604 11940 6656
rect 14464 6740 14516 6792
rect 15660 6783 15712 6792
rect 15660 6749 15669 6783
rect 15669 6749 15703 6783
rect 15703 6749 15712 6783
rect 15660 6740 15712 6749
rect 16304 6672 16356 6724
rect 18236 6783 18288 6792
rect 18236 6749 18245 6783
rect 18245 6749 18279 6783
rect 18279 6749 18288 6783
rect 18236 6740 18288 6749
rect 18972 6808 19024 6860
rect 20076 6876 20128 6928
rect 19340 6740 19392 6792
rect 14648 6604 14700 6656
rect 16948 6604 17000 6656
rect 18052 6647 18104 6656
rect 18052 6613 18061 6647
rect 18061 6613 18095 6647
rect 18095 6613 18104 6647
rect 18052 6604 18104 6613
rect 18696 6604 18748 6656
rect 19248 6672 19300 6724
rect 19616 6740 19668 6792
rect 21180 6808 21232 6860
rect 21088 6783 21140 6792
rect 21088 6749 21097 6783
rect 21097 6749 21131 6783
rect 21131 6749 21140 6783
rect 21088 6740 21140 6749
rect 19064 6604 19116 6656
rect 19156 6604 19208 6656
rect 20904 6604 20956 6656
rect 21272 6604 21324 6656
rect 6148 6502 6200 6554
rect 6212 6502 6264 6554
rect 6276 6502 6328 6554
rect 6340 6502 6392 6554
rect 6404 6502 6456 6554
rect 11346 6502 11398 6554
rect 11410 6502 11462 6554
rect 11474 6502 11526 6554
rect 11538 6502 11590 6554
rect 11602 6502 11654 6554
rect 16544 6502 16596 6554
rect 16608 6502 16660 6554
rect 16672 6502 16724 6554
rect 16736 6502 16788 6554
rect 16800 6502 16852 6554
rect 21742 6502 21794 6554
rect 21806 6502 21858 6554
rect 21870 6502 21922 6554
rect 21934 6502 21986 6554
rect 21998 6502 22050 6554
rect 1216 6400 1268 6452
rect 3148 6400 3200 6452
rect 3516 6400 3568 6452
rect 4160 6400 4212 6452
rect 5080 6400 5132 6452
rect 5540 6400 5592 6452
rect 10140 6400 10192 6452
rect 11060 6400 11112 6452
rect 11244 6400 11296 6452
rect 13268 6400 13320 6452
rect 13544 6400 13596 6452
rect 13728 6400 13780 6452
rect 14188 6400 14240 6452
rect 1492 6307 1544 6316
rect 1492 6273 1501 6307
rect 1501 6273 1535 6307
rect 1535 6273 1544 6307
rect 1492 6264 1544 6273
rect 1492 6060 1544 6112
rect 7564 6332 7616 6384
rect 7656 6375 7708 6384
rect 7656 6341 7665 6375
rect 7665 6341 7699 6375
rect 7699 6341 7708 6375
rect 7656 6332 7708 6341
rect 8116 6332 8168 6384
rect 3792 6264 3844 6316
rect 3424 6196 3476 6248
rect 4344 6307 4396 6316
rect 4344 6273 4353 6307
rect 4353 6273 4387 6307
rect 4387 6273 4396 6307
rect 4344 6264 4396 6273
rect 5080 6264 5132 6316
rect 6828 6307 6880 6316
rect 6828 6273 6837 6307
rect 6837 6273 6871 6307
rect 6871 6273 6880 6307
rect 6828 6264 6880 6273
rect 6920 6307 6972 6316
rect 6920 6273 6929 6307
rect 6929 6273 6963 6307
rect 6963 6273 6972 6307
rect 6920 6264 6972 6273
rect 7288 6307 7340 6316
rect 7288 6273 7297 6307
rect 7297 6273 7331 6307
rect 7331 6273 7340 6307
rect 7288 6264 7340 6273
rect 7380 6264 7432 6316
rect 6368 6196 6420 6248
rect 3700 6128 3752 6180
rect 4344 6128 4396 6180
rect 9312 6307 9364 6316
rect 9312 6273 9321 6307
rect 9321 6273 9355 6307
rect 9355 6273 9364 6307
rect 9312 6264 9364 6273
rect 9772 6332 9824 6384
rect 12900 6332 12952 6384
rect 14096 6332 14148 6384
rect 14372 6332 14424 6384
rect 15660 6443 15712 6452
rect 15660 6409 15669 6443
rect 15669 6409 15703 6443
rect 15703 6409 15712 6443
rect 15660 6400 15712 6409
rect 16028 6400 16080 6452
rect 17500 6400 17552 6452
rect 18696 6400 18748 6452
rect 19248 6400 19300 6452
rect 20720 6400 20772 6452
rect 20812 6400 20864 6452
rect 20904 6400 20956 6452
rect 21456 6400 21508 6452
rect 12164 6264 12216 6316
rect 14556 6307 14608 6316
rect 14556 6273 14590 6307
rect 14590 6273 14608 6307
rect 14556 6264 14608 6273
rect 10048 6196 10100 6248
rect 14280 6239 14332 6248
rect 14280 6205 14289 6239
rect 14289 6205 14323 6239
rect 14323 6205 14332 6239
rect 14280 6196 14332 6205
rect 20168 6375 20220 6384
rect 15660 6264 15712 6316
rect 15844 6264 15896 6316
rect 17040 6307 17092 6316
rect 17040 6273 17049 6307
rect 17049 6273 17083 6307
rect 17083 6273 17092 6307
rect 17040 6264 17092 6273
rect 17500 6307 17552 6316
rect 17500 6273 17509 6307
rect 17509 6273 17543 6307
rect 17543 6273 17552 6307
rect 17500 6264 17552 6273
rect 18236 6264 18288 6316
rect 18420 6307 18472 6316
rect 18420 6273 18429 6307
rect 18429 6273 18463 6307
rect 18463 6273 18472 6307
rect 18420 6264 18472 6273
rect 18788 6307 18840 6316
rect 18788 6273 18795 6307
rect 18795 6273 18829 6307
rect 18829 6273 18840 6307
rect 18788 6264 18840 6273
rect 20168 6341 20202 6375
rect 20202 6341 20220 6375
rect 20168 6332 20220 6341
rect 11888 6128 11940 6180
rect 14188 6128 14240 6180
rect 2872 6060 2924 6112
rect 3148 6060 3200 6112
rect 4068 6060 4120 6112
rect 6000 6060 6052 6112
rect 6552 6060 6604 6112
rect 9680 6060 9732 6112
rect 10968 6103 11020 6112
rect 10968 6069 10977 6103
rect 10977 6069 11011 6103
rect 11011 6069 11020 6103
rect 10968 6060 11020 6069
rect 11796 6103 11848 6112
rect 11796 6069 11805 6103
rect 11805 6069 11839 6103
rect 11839 6069 11848 6103
rect 11796 6060 11848 6069
rect 14648 6060 14700 6112
rect 15660 6128 15712 6180
rect 17132 6196 17184 6248
rect 18512 6239 18564 6248
rect 18512 6205 18521 6239
rect 18521 6205 18555 6239
rect 18555 6205 18564 6239
rect 18512 6196 18564 6205
rect 19340 6128 19392 6180
rect 15292 6060 15344 6112
rect 19892 6307 19944 6316
rect 19892 6273 19901 6307
rect 19901 6273 19935 6307
rect 19935 6273 19944 6307
rect 19892 6264 19944 6273
rect 20904 6060 20956 6112
rect 3549 5958 3601 6010
rect 3613 5958 3665 6010
rect 3677 5958 3729 6010
rect 3741 5958 3793 6010
rect 3805 5958 3857 6010
rect 8747 5958 8799 6010
rect 8811 5958 8863 6010
rect 8875 5958 8927 6010
rect 8939 5958 8991 6010
rect 9003 5958 9055 6010
rect 13945 5958 13997 6010
rect 14009 5958 14061 6010
rect 14073 5958 14125 6010
rect 14137 5958 14189 6010
rect 14201 5958 14253 6010
rect 19143 5958 19195 6010
rect 19207 5958 19259 6010
rect 19271 5958 19323 6010
rect 19335 5958 19387 6010
rect 19399 5958 19451 6010
rect 1492 5899 1544 5908
rect 1492 5865 1501 5899
rect 1501 5865 1535 5899
rect 1535 5865 1544 5899
rect 1492 5856 1544 5865
rect 1308 5720 1360 5772
rect 1584 5652 1636 5704
rect 4068 5856 4120 5908
rect 5632 5856 5684 5908
rect 5908 5856 5960 5908
rect 6184 5899 6236 5908
rect 6184 5865 6193 5899
rect 6193 5865 6227 5899
rect 6227 5865 6236 5899
rect 6184 5856 6236 5865
rect 6644 5856 6696 5908
rect 6920 5856 6972 5908
rect 9864 5856 9916 5908
rect 11704 5856 11756 5908
rect 15108 5856 15160 5908
rect 15292 5856 15344 5908
rect 15476 5856 15528 5908
rect 15844 5856 15896 5908
rect 17040 5856 17092 5908
rect 17132 5899 17184 5908
rect 17132 5865 17141 5899
rect 17141 5865 17175 5899
rect 17175 5865 17184 5899
rect 17132 5856 17184 5865
rect 18052 5856 18104 5908
rect 2320 5720 2372 5772
rect 2412 5763 2464 5772
rect 2412 5729 2421 5763
rect 2421 5729 2455 5763
rect 2455 5729 2464 5763
rect 2412 5720 2464 5729
rect 4160 5788 4212 5840
rect 4252 5788 4304 5840
rect 4436 5788 4488 5840
rect 3884 5720 3936 5772
rect 4620 5720 4672 5772
rect 2964 5695 3016 5704
rect 2964 5661 2973 5695
rect 2973 5661 3007 5695
rect 3007 5661 3016 5695
rect 2964 5652 3016 5661
rect 3792 5652 3844 5704
rect 4160 5652 4212 5704
rect 7564 5720 7616 5772
rect 5264 5695 5316 5704
rect 5264 5661 5273 5695
rect 5273 5661 5307 5695
rect 5307 5661 5316 5695
rect 5264 5652 5316 5661
rect 6460 5652 6512 5704
rect 6276 5584 6328 5636
rect 1584 5516 1636 5568
rect 3976 5516 4028 5568
rect 4620 5516 4672 5568
rect 4896 5516 4948 5568
rect 8024 5652 8076 5704
rect 8208 5652 8260 5704
rect 9772 5652 9824 5704
rect 12532 5720 12584 5772
rect 14648 5763 14700 5772
rect 14648 5729 14657 5763
rect 14657 5729 14691 5763
rect 14691 5729 14700 5763
rect 14648 5720 14700 5729
rect 18328 5831 18380 5840
rect 18328 5797 18337 5831
rect 18337 5797 18371 5831
rect 18371 5797 18380 5831
rect 18328 5788 18380 5797
rect 19156 5788 19208 5840
rect 6828 5516 6880 5568
rect 12164 5584 12216 5636
rect 14924 5695 14976 5704
rect 14924 5661 14933 5695
rect 14933 5661 14967 5695
rect 14967 5661 14976 5695
rect 14924 5652 14976 5661
rect 15292 5584 15344 5636
rect 7104 5516 7156 5568
rect 10416 5559 10468 5568
rect 10416 5525 10425 5559
rect 10425 5525 10459 5559
rect 10459 5525 10468 5559
rect 10416 5516 10468 5525
rect 10692 5516 10744 5568
rect 12716 5516 12768 5568
rect 13544 5516 13596 5568
rect 14740 5516 14792 5568
rect 15568 5652 15620 5704
rect 15752 5695 15804 5704
rect 15752 5661 15761 5695
rect 15761 5661 15795 5695
rect 15795 5661 15804 5695
rect 15752 5652 15804 5661
rect 16120 5763 16172 5772
rect 16120 5729 16129 5763
rect 16129 5729 16163 5763
rect 16163 5729 16172 5763
rect 16120 5720 16172 5729
rect 17592 5763 17644 5772
rect 17592 5729 17601 5763
rect 17601 5729 17635 5763
rect 17635 5729 17644 5763
rect 17592 5720 17644 5729
rect 15660 5584 15712 5636
rect 17040 5584 17092 5636
rect 16120 5516 16172 5568
rect 16212 5516 16264 5568
rect 17224 5584 17276 5636
rect 18512 5720 18564 5772
rect 18788 5652 18840 5704
rect 18880 5695 18932 5704
rect 18880 5661 18889 5695
rect 18889 5661 18923 5695
rect 18923 5661 18932 5695
rect 18880 5652 18932 5661
rect 18696 5584 18748 5636
rect 19984 5652 20036 5704
rect 21088 5856 21140 5908
rect 20996 5720 21048 5772
rect 21364 5652 21416 5704
rect 19064 5584 19116 5636
rect 20812 5559 20864 5568
rect 20812 5525 20821 5559
rect 20821 5525 20855 5559
rect 20855 5525 20864 5559
rect 20812 5516 20864 5525
rect 6148 5414 6200 5466
rect 6212 5414 6264 5466
rect 6276 5414 6328 5466
rect 6340 5414 6392 5466
rect 6404 5414 6456 5466
rect 11346 5414 11398 5466
rect 11410 5414 11462 5466
rect 11474 5414 11526 5466
rect 11538 5414 11590 5466
rect 11602 5414 11654 5466
rect 16544 5414 16596 5466
rect 16608 5414 16660 5466
rect 16672 5414 16724 5466
rect 16736 5414 16788 5466
rect 16800 5414 16852 5466
rect 21742 5414 21794 5466
rect 21806 5414 21858 5466
rect 21870 5414 21922 5466
rect 21934 5414 21986 5466
rect 21998 5414 22050 5466
rect 1768 5355 1820 5364
rect 1768 5321 1777 5355
rect 1777 5321 1811 5355
rect 1811 5321 1820 5355
rect 1768 5312 1820 5321
rect 2044 5312 2096 5364
rect 2320 5312 2372 5364
rect 2688 5312 2740 5364
rect 3056 5312 3108 5364
rect 5356 5312 5408 5364
rect 1492 5287 1544 5296
rect 1492 5253 1501 5287
rect 1501 5253 1535 5287
rect 1535 5253 1544 5287
rect 1492 5244 1544 5253
rect 3056 5176 3108 5228
rect 2136 5151 2188 5160
rect 2136 5117 2145 5151
rect 2145 5117 2179 5151
rect 2179 5117 2188 5151
rect 2136 5108 2188 5117
rect 1952 4972 2004 5024
rect 2504 4972 2556 5024
rect 3884 5244 3936 5296
rect 4344 5244 4396 5296
rect 8484 5312 8536 5364
rect 12992 5312 13044 5364
rect 14924 5312 14976 5364
rect 15568 5312 15620 5364
rect 15752 5312 15804 5364
rect 15844 5312 15896 5364
rect 16580 5312 16632 5364
rect 17592 5312 17644 5364
rect 17684 5312 17736 5364
rect 17868 5312 17920 5364
rect 18144 5312 18196 5364
rect 18512 5312 18564 5364
rect 18696 5312 18748 5364
rect 10048 5244 10100 5296
rect 12440 5244 12492 5296
rect 4620 5176 4672 5228
rect 5080 5176 5132 5228
rect 4896 5151 4948 5160
rect 4896 5117 4905 5151
rect 4905 5117 4939 5151
rect 4939 5117 4948 5151
rect 4896 5108 4948 5117
rect 5908 5176 5960 5228
rect 6000 5176 6052 5228
rect 6552 5176 6604 5228
rect 6644 5176 6696 5228
rect 6920 5108 6972 5160
rect 11152 5108 11204 5160
rect 12900 5151 12952 5160
rect 12900 5117 12909 5151
rect 12909 5117 12943 5151
rect 12943 5117 12952 5151
rect 12900 5108 12952 5117
rect 10324 4972 10376 5024
rect 14280 5219 14332 5228
rect 14280 5185 14289 5219
rect 14289 5185 14323 5219
rect 14323 5185 14332 5219
rect 14280 5176 14332 5185
rect 15936 5219 15988 5228
rect 15936 5185 15945 5219
rect 15945 5185 15979 5219
rect 15979 5185 15988 5219
rect 15936 5176 15988 5185
rect 16120 5151 16172 5160
rect 16120 5117 16129 5151
rect 16129 5117 16163 5151
rect 16163 5117 16172 5151
rect 16120 5108 16172 5117
rect 14464 4972 14516 5024
rect 14648 4972 14700 5024
rect 15292 4972 15344 5024
rect 15844 4972 15896 5024
rect 16396 5108 16448 5160
rect 18420 5249 18472 5296
rect 16764 5176 16816 5228
rect 18420 5244 18445 5249
rect 18445 5244 18472 5249
rect 20720 5244 20772 5296
rect 20260 5176 20312 5228
rect 20904 5219 20956 5228
rect 20904 5185 20913 5219
rect 20913 5185 20947 5219
rect 20947 5185 20956 5219
rect 20904 5176 20956 5185
rect 21088 5219 21140 5228
rect 21088 5185 21097 5219
rect 21097 5185 21131 5219
rect 21131 5185 21140 5219
rect 21088 5176 21140 5185
rect 21180 5176 21232 5228
rect 16672 5151 16724 5160
rect 16672 5117 16681 5151
rect 16681 5117 16715 5151
rect 16715 5117 16724 5151
rect 16672 5108 16724 5117
rect 19524 5151 19576 5160
rect 19524 5117 19533 5151
rect 19533 5117 19567 5151
rect 19567 5117 19576 5151
rect 19524 5108 19576 5117
rect 17684 4972 17736 5024
rect 18236 4972 18288 5024
rect 19064 4972 19116 5024
rect 3549 4870 3601 4922
rect 3613 4870 3665 4922
rect 3677 4870 3729 4922
rect 3741 4870 3793 4922
rect 3805 4870 3857 4922
rect 8747 4870 8799 4922
rect 8811 4870 8863 4922
rect 8875 4870 8927 4922
rect 8939 4870 8991 4922
rect 9003 4870 9055 4922
rect 13945 4870 13997 4922
rect 14009 4870 14061 4922
rect 14073 4870 14125 4922
rect 14137 4870 14189 4922
rect 14201 4870 14253 4922
rect 19143 4870 19195 4922
rect 19207 4870 19259 4922
rect 19271 4870 19323 4922
rect 19335 4870 19387 4922
rect 19399 4870 19451 4922
rect 3148 4768 3200 4820
rect 4712 4768 4764 4820
rect 4804 4768 4856 4820
rect 3608 4700 3660 4752
rect 12808 4768 12860 4820
rect 15200 4768 15252 4820
rect 16304 4768 16356 4820
rect 16856 4768 16908 4820
rect 17500 4768 17552 4820
rect 2136 4632 2188 4684
rect 1584 4607 1636 4616
rect 1584 4573 1593 4607
rect 1593 4573 1627 4607
rect 1627 4573 1636 4607
rect 1584 4564 1636 4573
rect 1860 4607 1912 4616
rect 1860 4573 1869 4607
rect 1869 4573 1903 4607
rect 1903 4573 1912 4607
rect 1860 4564 1912 4573
rect 3884 4675 3936 4684
rect 3884 4641 3893 4675
rect 3893 4641 3927 4675
rect 3927 4641 3936 4675
rect 3884 4632 3936 4641
rect 2504 4564 2556 4616
rect 5080 4564 5132 4616
rect 3792 4496 3844 4548
rect 4344 4496 4396 4548
rect 6828 4564 6880 4616
rect 14280 4564 14332 4616
rect 14464 4607 14516 4616
rect 14464 4573 14487 4607
rect 14487 4573 14516 4607
rect 14464 4564 14516 4573
rect 16488 4700 16540 4752
rect 17040 4700 17092 4752
rect 18236 4700 18288 4752
rect 16672 4632 16724 4684
rect 15936 4564 15988 4616
rect 16212 4564 16264 4616
rect 16396 4564 16448 4616
rect 5356 4496 5408 4548
rect 7288 4496 7340 4548
rect 16764 4607 16816 4616
rect 16764 4573 16773 4607
rect 16773 4573 16807 4607
rect 16807 4573 16816 4607
rect 16764 4564 16816 4573
rect 16672 4496 16724 4548
rect 3424 4428 3476 4480
rect 5172 4428 5224 4480
rect 5540 4428 5592 4480
rect 10600 4428 10652 4480
rect 14740 4428 14792 4480
rect 16304 4428 16356 4480
rect 17040 4607 17092 4616
rect 17040 4573 17049 4607
rect 17049 4573 17083 4607
rect 17083 4573 17092 4607
rect 17040 4564 17092 4573
rect 17224 4564 17276 4616
rect 19064 4700 19116 4752
rect 19524 4768 19576 4820
rect 21180 4768 21232 4820
rect 19340 4632 19392 4684
rect 17132 4496 17184 4548
rect 16856 4428 16908 4480
rect 17500 4496 17552 4548
rect 17868 4496 17920 4548
rect 17592 4428 17644 4480
rect 18604 4471 18656 4480
rect 18604 4437 18613 4471
rect 18613 4437 18647 4471
rect 18647 4437 18656 4471
rect 18604 4428 18656 4437
rect 19248 4564 19300 4616
rect 19524 4607 19576 4616
rect 19524 4573 19533 4607
rect 19533 4573 19567 4607
rect 19567 4573 19576 4607
rect 19524 4564 19576 4573
rect 19892 4632 19944 4684
rect 19064 4428 19116 4480
rect 19524 4428 19576 4480
rect 19616 4471 19668 4480
rect 19616 4437 19625 4471
rect 19625 4437 19659 4471
rect 19659 4437 19668 4471
rect 19616 4428 19668 4437
rect 21364 4471 21416 4480
rect 21364 4437 21373 4471
rect 21373 4437 21407 4471
rect 21407 4437 21416 4471
rect 21364 4428 21416 4437
rect 6148 4326 6200 4378
rect 6212 4326 6264 4378
rect 6276 4326 6328 4378
rect 6340 4326 6392 4378
rect 6404 4326 6456 4378
rect 11346 4326 11398 4378
rect 11410 4326 11462 4378
rect 11474 4326 11526 4378
rect 11538 4326 11590 4378
rect 11602 4326 11654 4378
rect 16544 4326 16596 4378
rect 16608 4326 16660 4378
rect 16672 4326 16724 4378
rect 16736 4326 16788 4378
rect 16800 4326 16852 4378
rect 21742 4326 21794 4378
rect 21806 4326 21858 4378
rect 21870 4326 21922 4378
rect 21934 4326 21986 4378
rect 21998 4326 22050 4378
rect 2688 4224 2740 4276
rect 1952 4156 2004 4208
rect 3976 4224 4028 4276
rect 4804 4224 4856 4276
rect 11980 4224 12032 4276
rect 14648 4224 14700 4276
rect 14832 4224 14884 4276
rect 15108 4224 15160 4276
rect 16028 4224 16080 4276
rect 2228 4088 2280 4140
rect 3056 4156 3108 4208
rect 4344 4156 4396 4208
rect 5816 4156 5868 4208
rect 6092 4156 6144 4208
rect 6736 4156 6788 4208
rect 3700 4088 3752 4140
rect 3884 4088 3936 4140
rect 4160 4088 4212 4140
rect 1584 4063 1636 4072
rect 1584 4029 1593 4063
rect 1593 4029 1627 4063
rect 1627 4029 1636 4063
rect 1584 4020 1636 4029
rect 3792 4020 3844 4072
rect 3240 3884 3292 3936
rect 4620 3884 4672 3936
rect 5448 4088 5500 4140
rect 5724 4088 5776 4140
rect 6552 4088 6604 4140
rect 13084 4156 13136 4208
rect 17224 4224 17276 4276
rect 17684 4224 17736 4276
rect 18052 4224 18104 4276
rect 17592 4156 17644 4208
rect 5264 4020 5316 4072
rect 5816 4020 5868 4072
rect 7840 4020 7892 4072
rect 5448 3952 5500 4004
rect 13820 4088 13872 4140
rect 14372 4131 14424 4140
rect 14372 4097 14381 4131
rect 14381 4097 14415 4131
rect 14415 4097 14424 4131
rect 14372 4088 14424 4097
rect 14464 4020 14516 4072
rect 14924 4088 14976 4140
rect 15200 4131 15252 4140
rect 15200 4097 15209 4131
rect 15209 4097 15243 4131
rect 15243 4097 15252 4131
rect 15200 4088 15252 4097
rect 15016 4020 15068 4072
rect 15568 4131 15620 4140
rect 15568 4097 15577 4131
rect 15577 4097 15611 4131
rect 15611 4097 15620 4131
rect 15568 4088 15620 4097
rect 16028 4088 16080 4140
rect 16120 4088 16172 4140
rect 16488 4131 16540 4140
rect 16488 4097 16497 4131
rect 16497 4097 16531 4131
rect 16531 4097 16540 4131
rect 16488 4088 16540 4097
rect 16580 4088 16632 4140
rect 17224 4088 17276 4140
rect 17868 4131 17920 4140
rect 17868 4097 17877 4131
rect 17877 4097 17911 4131
rect 17911 4097 17920 4131
rect 17868 4088 17920 4097
rect 16764 4020 16816 4072
rect 16948 3952 17000 4004
rect 18236 4088 18288 4140
rect 18604 4156 18656 4208
rect 19156 4267 19208 4276
rect 19156 4233 19165 4267
rect 19165 4233 19199 4267
rect 19199 4233 19208 4267
rect 19156 4224 19208 4233
rect 19340 4224 19392 4276
rect 18696 4131 18748 4140
rect 18144 3952 18196 4004
rect 18696 4097 18705 4131
rect 18705 4097 18739 4131
rect 18739 4097 18748 4131
rect 18696 4088 18748 4097
rect 19708 4156 19760 4208
rect 19984 4156 20036 4208
rect 18972 4131 19024 4140
rect 18972 4097 18981 4131
rect 18981 4097 19015 4131
rect 19015 4097 19024 4131
rect 18972 4088 19024 4097
rect 21088 4088 21140 4140
rect 21272 4131 21324 4140
rect 21272 4097 21281 4131
rect 21281 4097 21315 4131
rect 21315 4097 21324 4131
rect 21272 4088 21324 4097
rect 18420 3952 18472 4004
rect 5724 3927 5776 3936
rect 5724 3893 5733 3927
rect 5733 3893 5767 3927
rect 5767 3893 5776 3927
rect 5724 3884 5776 3893
rect 6736 3884 6788 3936
rect 9680 3884 9732 3936
rect 12992 3884 13044 3936
rect 15752 3927 15804 3936
rect 15752 3893 15761 3927
rect 15761 3893 15795 3927
rect 15795 3893 15804 3927
rect 15752 3884 15804 3893
rect 16304 3927 16356 3936
rect 16304 3893 16313 3927
rect 16313 3893 16347 3927
rect 16347 3893 16356 3927
rect 16304 3884 16356 3893
rect 18788 3884 18840 3936
rect 19892 3884 19944 3936
rect 20260 3884 20312 3936
rect 20996 3927 21048 3936
rect 20996 3893 21005 3927
rect 21005 3893 21039 3927
rect 21039 3893 21048 3927
rect 20996 3884 21048 3893
rect 21364 3927 21416 3936
rect 21364 3893 21373 3927
rect 21373 3893 21407 3927
rect 21407 3893 21416 3927
rect 21364 3884 21416 3893
rect 3549 3782 3601 3834
rect 3613 3782 3665 3834
rect 3677 3782 3729 3834
rect 3741 3782 3793 3834
rect 3805 3782 3857 3834
rect 8747 3782 8799 3834
rect 8811 3782 8863 3834
rect 8875 3782 8927 3834
rect 8939 3782 8991 3834
rect 9003 3782 9055 3834
rect 13945 3782 13997 3834
rect 14009 3782 14061 3834
rect 14073 3782 14125 3834
rect 14137 3782 14189 3834
rect 14201 3782 14253 3834
rect 19143 3782 19195 3834
rect 19207 3782 19259 3834
rect 19271 3782 19323 3834
rect 19335 3782 19387 3834
rect 19399 3782 19451 3834
rect 2872 3680 2924 3732
rect 3332 3723 3384 3732
rect 3332 3689 3341 3723
rect 3341 3689 3375 3723
rect 3375 3689 3384 3723
rect 3332 3680 3384 3689
rect 2412 3612 2464 3664
rect 5632 3680 5684 3732
rect 1584 3587 1636 3596
rect 1584 3553 1593 3587
rect 1593 3553 1627 3587
rect 1627 3553 1636 3587
rect 1584 3544 1636 3553
rect 3792 3587 3844 3596
rect 3792 3553 3801 3587
rect 3801 3553 3835 3587
rect 3835 3553 3844 3587
rect 3792 3544 3844 3553
rect 5632 3544 5684 3596
rect 11612 3680 11664 3732
rect 11796 3680 11848 3732
rect 15200 3680 15252 3732
rect 480 3476 532 3528
rect 1032 3408 1084 3460
rect 3240 3451 3292 3460
rect 3240 3417 3249 3451
rect 3249 3417 3283 3451
rect 3283 3417 3292 3451
rect 3240 3408 3292 3417
rect 6736 3544 6788 3596
rect 6920 3544 6972 3596
rect 7196 3544 7248 3596
rect 8668 3544 8720 3596
rect 5908 3519 5960 3528
rect 5908 3485 5917 3519
rect 5917 3485 5951 3519
rect 5951 3485 5960 3519
rect 5908 3476 5960 3485
rect 7656 3519 7708 3528
rect 7656 3485 7665 3519
rect 7665 3485 7699 3519
rect 7699 3485 7708 3519
rect 7656 3476 7708 3485
rect 7748 3476 7800 3528
rect 3148 3340 3200 3392
rect 4436 3340 4488 3392
rect 7012 3408 7064 3460
rect 8760 3519 8812 3528
rect 8760 3485 8769 3519
rect 8769 3485 8803 3519
rect 8803 3485 8812 3519
rect 8760 3476 8812 3485
rect 9772 3544 9824 3596
rect 13176 3612 13228 3664
rect 13728 3612 13780 3664
rect 16396 3680 16448 3732
rect 17868 3680 17920 3732
rect 18420 3723 18472 3732
rect 18420 3689 18429 3723
rect 18429 3689 18463 3723
rect 18463 3689 18472 3723
rect 18420 3680 18472 3689
rect 18512 3680 18564 3732
rect 18788 3680 18840 3732
rect 20444 3680 20496 3732
rect 21272 3680 21324 3732
rect 22652 3680 22704 3732
rect 9404 3519 9456 3528
rect 9404 3485 9413 3519
rect 9413 3485 9447 3519
rect 9447 3485 9456 3519
rect 9404 3476 9456 3485
rect 12624 3544 12676 3596
rect 15844 3612 15896 3664
rect 16580 3544 16632 3596
rect 17408 3612 17460 3664
rect 13452 3476 13504 3528
rect 13820 3476 13872 3528
rect 9312 3408 9364 3460
rect 14464 3476 14516 3528
rect 14740 3476 14792 3528
rect 14832 3519 14884 3528
rect 14832 3485 14841 3519
rect 14841 3485 14875 3519
rect 14875 3485 14884 3519
rect 14832 3476 14884 3485
rect 15108 3519 15160 3528
rect 15108 3485 15117 3519
rect 15117 3485 15151 3519
rect 15151 3485 15160 3519
rect 15108 3476 15160 3485
rect 15200 3476 15252 3528
rect 15568 3476 15620 3528
rect 15660 3519 15712 3528
rect 15660 3485 15669 3519
rect 15669 3485 15703 3519
rect 15703 3485 15712 3519
rect 15660 3476 15712 3485
rect 15936 3476 15988 3528
rect 16488 3476 16540 3528
rect 17316 3544 17368 3596
rect 17408 3476 17460 3528
rect 17776 3544 17828 3596
rect 17868 3544 17920 3596
rect 6920 3340 6972 3392
rect 7564 3340 7616 3392
rect 8300 3383 8352 3392
rect 8300 3349 8309 3383
rect 8309 3349 8343 3383
rect 8343 3349 8352 3383
rect 8300 3340 8352 3349
rect 8576 3383 8628 3392
rect 8576 3349 8585 3383
rect 8585 3349 8619 3383
rect 8619 3349 8628 3383
rect 8576 3340 8628 3349
rect 9220 3383 9272 3392
rect 9220 3349 9229 3383
rect 9229 3349 9263 3383
rect 9263 3349 9272 3383
rect 9220 3340 9272 3349
rect 9864 3383 9916 3392
rect 9864 3349 9873 3383
rect 9873 3349 9907 3383
rect 9907 3349 9916 3383
rect 9864 3340 9916 3349
rect 11612 3340 11664 3392
rect 12900 3383 12952 3392
rect 12900 3349 12909 3383
rect 12909 3349 12943 3383
rect 12943 3349 12952 3383
rect 12900 3340 12952 3349
rect 13452 3340 13504 3392
rect 14648 3408 14700 3460
rect 14464 3340 14516 3392
rect 14556 3340 14608 3392
rect 15292 3408 15344 3460
rect 14924 3383 14976 3392
rect 14924 3349 14933 3383
rect 14933 3349 14967 3383
rect 14967 3349 14976 3383
rect 14924 3340 14976 3349
rect 15200 3383 15252 3392
rect 15200 3349 15209 3383
rect 15209 3349 15243 3383
rect 15243 3349 15252 3383
rect 15200 3340 15252 3349
rect 15752 3340 15804 3392
rect 16396 3340 16448 3392
rect 16764 3340 16816 3392
rect 18328 3519 18380 3528
rect 18328 3485 18337 3519
rect 18337 3485 18371 3519
rect 18371 3485 18380 3519
rect 18328 3476 18380 3485
rect 22468 3544 22520 3596
rect 18604 3519 18656 3528
rect 18604 3485 18613 3519
rect 18613 3485 18647 3519
rect 18647 3485 18656 3519
rect 18604 3476 18656 3485
rect 18696 3519 18748 3528
rect 18696 3485 18705 3519
rect 18705 3485 18739 3519
rect 18739 3485 18748 3519
rect 18696 3476 18748 3485
rect 19892 3476 19944 3528
rect 20720 3476 20772 3528
rect 21548 3408 21600 3460
rect 18052 3340 18104 3392
rect 18420 3340 18472 3392
rect 19984 3340 20036 3392
rect 20904 3340 20956 3392
rect 22560 3340 22612 3392
rect 6148 3238 6200 3290
rect 6212 3238 6264 3290
rect 6276 3238 6328 3290
rect 6340 3238 6392 3290
rect 6404 3238 6456 3290
rect 11346 3238 11398 3290
rect 11410 3238 11462 3290
rect 11474 3238 11526 3290
rect 11538 3238 11590 3290
rect 11602 3238 11654 3290
rect 16544 3238 16596 3290
rect 16608 3238 16660 3290
rect 16672 3238 16724 3290
rect 16736 3238 16788 3290
rect 16800 3238 16852 3290
rect 21742 3238 21794 3290
rect 21806 3238 21858 3290
rect 21870 3238 21922 3290
rect 21934 3238 21986 3290
rect 21998 3238 22050 3290
rect 1584 3136 1636 3188
rect 2320 3000 2372 3052
rect 2596 3136 2648 3188
rect 3148 3136 3200 3188
rect 3240 3136 3292 3188
rect 2504 3068 2556 3120
rect 3056 3043 3108 3052
rect 3056 3009 3065 3043
rect 3065 3009 3099 3043
rect 3099 3009 3108 3043
rect 3056 3000 3108 3009
rect 3424 3068 3476 3120
rect 4436 3068 4488 3120
rect 6000 3136 6052 3188
rect 6828 3136 6880 3188
rect 9772 3136 9824 3188
rect 10416 3136 10468 3188
rect 2596 2932 2648 2984
rect 2872 2932 2924 2984
rect 2964 2932 3016 2984
rect 5448 3043 5500 3052
rect 5448 3009 5457 3043
rect 5457 3009 5491 3043
rect 5491 3009 5500 3043
rect 5448 3000 5500 3009
rect 6736 3043 6788 3052
rect 6736 3009 6745 3043
rect 6745 3009 6779 3043
rect 6779 3009 6788 3043
rect 6736 3000 6788 3009
rect 7012 3043 7064 3052
rect 7012 3009 7021 3043
rect 7021 3009 7055 3043
rect 7055 3009 7064 3043
rect 7012 3000 7064 3009
rect 7196 3000 7248 3052
rect 7380 3000 7432 3052
rect 7840 3043 7892 3052
rect 7840 3009 7849 3043
rect 7849 3009 7883 3043
rect 7883 3009 7892 3043
rect 7840 3000 7892 3009
rect 8300 3000 8352 3052
rect 8392 3043 8444 3052
rect 8392 3009 8401 3043
rect 8401 3009 8435 3043
rect 8435 3009 8444 3043
rect 8392 3000 8444 3009
rect 8944 3043 8996 3052
rect 8944 3009 8953 3043
rect 8953 3009 8987 3043
rect 8987 3009 8996 3043
rect 8944 3000 8996 3009
rect 9220 3043 9272 3052
rect 9220 3009 9229 3043
rect 9229 3009 9263 3043
rect 9263 3009 9272 3043
rect 9220 3000 9272 3009
rect 9496 3043 9548 3052
rect 9496 3009 9505 3043
rect 9505 3009 9539 3043
rect 9539 3009 9548 3043
rect 9496 3000 9548 3009
rect 6644 2932 6696 2984
rect 8484 2932 8536 2984
rect 10232 3043 10284 3052
rect 10232 3009 10241 3043
rect 10241 3009 10275 3043
rect 10275 3009 10284 3043
rect 10232 3000 10284 3009
rect 10784 3000 10836 3052
rect 11060 3043 11112 3052
rect 11060 3009 11069 3043
rect 11069 3009 11103 3043
rect 11103 3009 11112 3043
rect 11060 3000 11112 3009
rect 12072 3000 12124 3052
rect 13360 3068 13412 3120
rect 13636 3136 13688 3188
rect 14096 3179 14148 3188
rect 14096 3145 14105 3179
rect 14105 3145 14139 3179
rect 14139 3145 14148 3179
rect 14096 3136 14148 3145
rect 14556 3136 14608 3188
rect 15016 3136 15068 3188
rect 15384 3136 15436 3188
rect 12808 3043 12860 3052
rect 12808 3009 12817 3043
rect 12817 3009 12851 3043
rect 12851 3009 12860 3043
rect 12808 3000 12860 3009
rect 14372 3000 14424 3052
rect 14740 3000 14792 3052
rect 14832 3043 14884 3052
rect 14832 3009 14841 3043
rect 14841 3009 14875 3043
rect 14875 3009 14884 3043
rect 14832 3000 14884 3009
rect 3976 2864 4028 2916
rect 7104 2864 7156 2916
rect 9496 2864 9548 2916
rect 14464 2932 14516 2984
rect 15200 3000 15252 3052
rect 15476 3000 15528 3052
rect 15936 3068 15988 3120
rect 16304 3043 16356 3052
rect 16304 3009 16313 3043
rect 16313 3009 16347 3043
rect 16347 3009 16356 3043
rect 16304 3000 16356 3009
rect 18144 3136 18196 3188
rect 18512 3179 18564 3188
rect 18512 3145 18521 3179
rect 18521 3145 18555 3179
rect 18555 3145 18564 3179
rect 18512 3136 18564 3145
rect 17960 3043 18012 3052
rect 17960 3009 17969 3043
rect 17969 3009 18003 3043
rect 18003 3009 18012 3043
rect 17960 3000 18012 3009
rect 10324 2864 10376 2916
rect 4252 2796 4304 2848
rect 6828 2839 6880 2848
rect 6828 2805 6837 2839
rect 6837 2805 6871 2839
rect 6871 2805 6880 2839
rect 6828 2796 6880 2805
rect 7380 2839 7432 2848
rect 7380 2805 7389 2839
rect 7389 2805 7423 2839
rect 7423 2805 7432 2839
rect 7380 2796 7432 2805
rect 7656 2839 7708 2848
rect 7656 2805 7665 2839
rect 7665 2805 7699 2839
rect 7699 2805 7708 2839
rect 7656 2796 7708 2805
rect 7748 2796 7800 2848
rect 7932 2839 7984 2848
rect 7932 2805 7941 2839
rect 7941 2805 7975 2839
rect 7975 2805 7984 2839
rect 7932 2796 7984 2805
rect 8208 2839 8260 2848
rect 8208 2805 8217 2839
rect 8217 2805 8251 2839
rect 8251 2805 8260 2839
rect 8208 2796 8260 2805
rect 8484 2839 8536 2848
rect 8484 2805 8493 2839
rect 8493 2805 8527 2839
rect 8527 2805 8536 2839
rect 8484 2796 8536 2805
rect 8576 2796 8628 2848
rect 9128 2796 9180 2848
rect 9680 2796 9732 2848
rect 10508 2839 10560 2848
rect 10508 2805 10517 2839
rect 10517 2805 10551 2839
rect 10551 2805 10560 2839
rect 10508 2796 10560 2805
rect 11888 2864 11940 2916
rect 13636 2864 13688 2916
rect 18052 2932 18104 2984
rect 18236 3043 18288 3052
rect 18236 3009 18245 3043
rect 18245 3009 18279 3043
rect 18279 3009 18288 3043
rect 18236 3000 18288 3009
rect 18420 3043 18472 3052
rect 18420 3009 18429 3043
rect 18429 3009 18463 3043
rect 18463 3009 18472 3043
rect 18420 3000 18472 3009
rect 19064 3000 19116 3052
rect 19616 3136 19668 3188
rect 20076 3179 20128 3188
rect 20076 3145 20085 3179
rect 20085 3145 20119 3179
rect 20119 3145 20128 3179
rect 20076 3136 20128 3145
rect 20628 3136 20680 3188
rect 20904 3136 20956 3188
rect 21364 3136 21416 3188
rect 19524 3043 19576 3052
rect 19524 3009 19533 3043
rect 19533 3009 19567 3043
rect 19567 3009 19576 3043
rect 19524 3000 19576 3009
rect 20444 3000 20496 3052
rect 20812 3000 20864 3052
rect 19800 2932 19852 2984
rect 22192 2932 22244 2984
rect 15016 2864 15068 2916
rect 12072 2796 12124 2848
rect 12624 2839 12676 2848
rect 12624 2805 12633 2839
rect 12633 2805 12667 2839
rect 12667 2805 12676 2839
rect 12624 2796 12676 2805
rect 13820 2839 13872 2848
rect 13820 2805 13829 2839
rect 13829 2805 13863 2839
rect 13863 2805 13872 2839
rect 13820 2796 13872 2805
rect 14372 2839 14424 2848
rect 14372 2805 14381 2839
rect 14381 2805 14415 2839
rect 14415 2805 14424 2839
rect 14372 2796 14424 2805
rect 14740 2796 14792 2848
rect 15476 2796 15528 2848
rect 15844 2864 15896 2916
rect 17224 2864 17276 2916
rect 19340 2864 19392 2916
rect 20536 2864 20588 2916
rect 16028 2796 16080 2848
rect 17776 2839 17828 2848
rect 17776 2805 17785 2839
rect 17785 2805 17819 2839
rect 17819 2805 17828 2839
rect 17776 2796 17828 2805
rect 18880 2796 18932 2848
rect 19064 2796 19116 2848
rect 21364 2839 21416 2848
rect 21364 2805 21373 2839
rect 21373 2805 21407 2839
rect 21407 2805 21416 2839
rect 21364 2796 21416 2805
rect 3549 2694 3601 2746
rect 3613 2694 3665 2746
rect 3677 2694 3729 2746
rect 3741 2694 3793 2746
rect 3805 2694 3857 2746
rect 8747 2694 8799 2746
rect 8811 2694 8863 2746
rect 8875 2694 8927 2746
rect 8939 2694 8991 2746
rect 9003 2694 9055 2746
rect 13945 2694 13997 2746
rect 14009 2694 14061 2746
rect 14073 2694 14125 2746
rect 14137 2694 14189 2746
rect 14201 2694 14253 2746
rect 19143 2694 19195 2746
rect 19207 2694 19259 2746
rect 19271 2694 19323 2746
rect 19335 2694 19387 2746
rect 19399 2694 19451 2746
rect 2320 2635 2372 2644
rect 2320 2601 2329 2635
rect 2329 2601 2363 2635
rect 2363 2601 2372 2635
rect 2320 2592 2372 2601
rect 1308 2524 1360 2576
rect 4160 2635 4212 2644
rect 4160 2601 4169 2635
rect 4169 2601 4203 2635
rect 4203 2601 4212 2635
rect 4160 2592 4212 2601
rect 4528 2635 4580 2644
rect 4528 2601 4537 2635
rect 4537 2601 4571 2635
rect 4571 2601 4580 2635
rect 4528 2592 4580 2601
rect 5172 2635 5224 2644
rect 5172 2601 5181 2635
rect 5181 2601 5215 2635
rect 5215 2601 5224 2635
rect 5172 2592 5224 2601
rect 5356 2592 5408 2644
rect 7196 2592 7248 2644
rect 7932 2635 7984 2644
rect 7932 2601 7941 2635
rect 7941 2601 7975 2635
rect 7975 2601 7984 2635
rect 7932 2592 7984 2601
rect 10692 2592 10744 2644
rect 10968 2592 11020 2644
rect 10876 2524 10928 2576
rect 11060 2524 11112 2576
rect 14832 2592 14884 2644
rect 15568 2635 15620 2644
rect 15568 2601 15577 2635
rect 15577 2601 15611 2635
rect 15611 2601 15620 2635
rect 15568 2592 15620 2601
rect 15660 2592 15712 2644
rect 21640 2592 21692 2644
rect 1216 2456 1268 2508
rect 2044 2431 2096 2440
rect 2044 2397 2053 2431
rect 2053 2397 2087 2431
rect 2087 2397 2096 2431
rect 2044 2388 2096 2397
rect 2596 2431 2648 2440
rect 2596 2397 2605 2431
rect 2605 2397 2639 2431
rect 2639 2397 2648 2431
rect 2596 2388 2648 2397
rect 664 2320 716 2372
rect 3884 2431 3936 2440
rect 3884 2397 3893 2431
rect 3893 2397 3927 2431
rect 3927 2397 3936 2431
rect 3884 2388 3936 2397
rect 4160 2388 4212 2440
rect 940 2252 992 2304
rect 3700 2252 3752 2304
rect 4160 2252 4212 2304
rect 4436 2388 4488 2440
rect 4804 2388 4856 2440
rect 10784 2456 10836 2508
rect 4620 2320 4672 2372
rect 5632 2431 5684 2440
rect 5632 2397 5641 2431
rect 5641 2397 5675 2431
rect 5675 2397 5684 2431
rect 5632 2388 5684 2397
rect 5908 2320 5960 2372
rect 6276 2363 6328 2372
rect 6276 2329 6285 2363
rect 6285 2329 6319 2363
rect 6319 2329 6328 2363
rect 6276 2320 6328 2329
rect 6000 2252 6052 2304
rect 6920 2431 6972 2440
rect 6920 2397 6929 2431
rect 6929 2397 6963 2431
rect 6963 2397 6972 2431
rect 6920 2388 6972 2397
rect 7564 2388 7616 2440
rect 7656 2388 7708 2440
rect 8208 2431 8260 2440
rect 8208 2397 8217 2431
rect 8217 2397 8251 2431
rect 8251 2397 8260 2431
rect 8208 2388 8260 2397
rect 8576 2388 8628 2440
rect 9588 2388 9640 2440
rect 10600 2388 10652 2440
rect 9772 2320 9824 2372
rect 6920 2252 6972 2304
rect 7012 2295 7064 2304
rect 7012 2261 7021 2295
rect 7021 2261 7055 2295
rect 7055 2261 7064 2295
rect 7012 2252 7064 2261
rect 7196 2252 7248 2304
rect 10876 2320 10928 2372
rect 11612 2431 11664 2440
rect 11612 2397 11621 2431
rect 11621 2397 11655 2431
rect 11655 2397 11664 2431
rect 11612 2388 11664 2397
rect 16580 2524 16632 2576
rect 18052 2524 18104 2576
rect 15108 2456 15160 2508
rect 15384 2388 15436 2440
rect 16120 2456 16172 2508
rect 17592 2499 17644 2508
rect 17592 2465 17601 2499
rect 17601 2465 17635 2499
rect 17635 2465 17644 2499
rect 17592 2456 17644 2465
rect 17684 2456 17736 2508
rect 9956 2295 10008 2304
rect 9956 2261 9965 2295
rect 9965 2261 9999 2295
rect 9999 2261 10008 2295
rect 9956 2252 10008 2261
rect 10232 2295 10284 2304
rect 10232 2261 10241 2295
rect 10241 2261 10275 2295
rect 10275 2261 10284 2295
rect 10232 2252 10284 2261
rect 10508 2295 10560 2304
rect 10508 2261 10517 2295
rect 10517 2261 10551 2295
rect 10551 2261 10560 2295
rect 10508 2252 10560 2261
rect 11244 2252 11296 2304
rect 11704 2295 11756 2304
rect 11704 2261 11713 2295
rect 11713 2261 11747 2295
rect 11747 2261 11756 2295
rect 11704 2252 11756 2261
rect 11796 2252 11848 2304
rect 11980 2252 12032 2304
rect 12440 2252 12492 2304
rect 13636 2295 13688 2304
rect 13636 2261 13645 2295
rect 13645 2261 13679 2295
rect 13679 2261 13688 2295
rect 13636 2252 13688 2261
rect 15108 2252 15160 2304
rect 17224 2431 17276 2440
rect 17224 2397 17233 2431
rect 17233 2397 17267 2431
rect 17267 2397 17276 2431
rect 17224 2388 17276 2397
rect 17776 2388 17828 2440
rect 18512 2431 18564 2440
rect 18512 2397 18521 2431
rect 18521 2397 18555 2431
rect 18555 2397 18564 2431
rect 18512 2388 18564 2397
rect 18696 2388 18748 2440
rect 20076 2499 20128 2508
rect 20076 2465 20085 2499
rect 20085 2465 20119 2499
rect 20119 2465 20128 2499
rect 20076 2456 20128 2465
rect 21180 2499 21232 2508
rect 21180 2465 21189 2499
rect 21189 2465 21223 2499
rect 21223 2465 21232 2499
rect 21180 2456 21232 2465
rect 16120 2295 16172 2304
rect 16120 2261 16129 2295
rect 16129 2261 16163 2295
rect 16163 2261 16172 2295
rect 16120 2252 16172 2261
rect 20168 2320 20220 2372
rect 18328 2295 18380 2304
rect 18328 2261 18337 2295
rect 18337 2261 18371 2295
rect 18371 2261 18380 2295
rect 18328 2252 18380 2261
rect 6148 2150 6200 2202
rect 6212 2150 6264 2202
rect 6276 2150 6328 2202
rect 6340 2150 6392 2202
rect 6404 2150 6456 2202
rect 11346 2150 11398 2202
rect 11410 2150 11462 2202
rect 11474 2150 11526 2202
rect 11538 2150 11590 2202
rect 11602 2150 11654 2202
rect 16544 2150 16596 2202
rect 16608 2150 16660 2202
rect 16672 2150 16724 2202
rect 16736 2150 16788 2202
rect 16800 2150 16852 2202
rect 21742 2150 21794 2202
rect 21806 2150 21858 2202
rect 21870 2150 21922 2202
rect 21934 2150 21986 2202
rect 21998 2150 22050 2202
rect 1400 2048 1452 2100
rect 2596 2048 2648 2100
rect 2872 2091 2924 2100
rect 2872 2057 2881 2091
rect 2881 2057 2915 2091
rect 2915 2057 2924 2091
rect 2872 2048 2924 2057
rect 1492 2023 1544 2032
rect 1492 1989 1501 2023
rect 1501 1989 1535 2023
rect 1535 1989 1544 2023
rect 1492 1980 1544 1989
rect 1952 1980 2004 2032
rect 3976 2048 4028 2100
rect 4528 2048 4580 2100
rect 4804 2048 4856 2100
rect 5724 2048 5776 2100
rect 7196 2048 7248 2100
rect 7380 1980 7432 2032
rect 8024 2048 8076 2100
rect 9404 2048 9456 2100
rect 9956 2048 10008 2100
rect 7840 2023 7892 2032
rect 7840 1989 7849 2023
rect 7849 1989 7883 2023
rect 7883 1989 7892 2023
rect 7840 1980 7892 1989
rect 8208 2023 8260 2032
rect 8208 1989 8217 2023
rect 8217 1989 8251 2023
rect 8251 1989 8260 2023
rect 8208 1980 8260 1989
rect 2504 1912 2556 1964
rect 3240 1955 3292 1964
rect 3240 1921 3249 1955
rect 3249 1921 3283 1955
rect 3283 1921 3292 1955
rect 3240 1912 3292 1921
rect 3424 1912 3476 1964
rect 3884 1912 3936 1964
rect 4620 1955 4672 1964
rect 4620 1921 4629 1955
rect 4629 1921 4663 1955
rect 4663 1921 4672 1955
rect 4620 1912 4672 1921
rect 4804 1912 4856 1964
rect 4896 1955 4948 1964
rect 4896 1921 4905 1955
rect 4905 1921 4939 1955
rect 4939 1921 4948 1955
rect 4896 1912 4948 1921
rect 6552 1912 6604 1964
rect 6828 1912 6880 1964
rect 9128 1980 9180 2032
rect 9680 1980 9732 2032
rect 10416 2023 10468 2032
rect 10416 1989 10425 2023
rect 10425 1989 10459 2023
rect 10459 1989 10468 2023
rect 10416 1980 10468 1989
rect 12992 2091 13044 2100
rect 12992 2057 13001 2091
rect 13001 2057 13035 2091
rect 13035 2057 13044 2091
rect 12992 2048 13044 2057
rect 11244 1980 11296 2032
rect 13636 1980 13688 2032
rect 15200 1980 15252 2032
rect 572 1844 624 1896
rect 296 1776 348 1828
rect 3148 1776 3200 1828
rect 3700 1776 3752 1828
rect 4988 1776 5040 1828
rect 5264 1887 5316 1896
rect 5264 1853 5273 1887
rect 5273 1853 5307 1887
rect 5307 1853 5316 1887
rect 5264 1844 5316 1853
rect 5448 1844 5500 1896
rect 8024 1844 8076 1896
rect 10140 1844 10192 1896
rect 10508 1844 10560 1896
rect 12716 1912 12768 1964
rect 12900 1912 12952 1964
rect 14924 1955 14976 1964
rect 14924 1921 14933 1955
rect 14933 1921 14967 1955
rect 14967 1921 14976 1955
rect 14924 1912 14976 1921
rect 10048 1776 10100 1828
rect 10600 1776 10652 1828
rect 10784 1776 10836 1828
rect 14464 1844 14516 1896
rect 17132 2048 17184 2100
rect 18880 2048 18932 2100
rect 20996 2048 21048 2100
rect 21364 2048 21416 2100
rect 15476 2023 15528 2032
rect 15476 1989 15485 2023
rect 15485 1989 15519 2023
rect 15519 1989 15528 2023
rect 15476 1980 15528 1989
rect 15752 1980 15804 2032
rect 17040 1980 17092 2032
rect 18788 1980 18840 2032
rect 20352 1980 20404 2032
rect 21456 1980 21508 2032
rect 16856 1912 16908 1964
rect 17132 1912 17184 1964
rect 17868 1912 17920 1964
rect 20720 1912 20772 1964
rect 14372 1776 14424 1828
rect 7196 1751 7248 1760
rect 7196 1717 7205 1751
rect 7205 1717 7239 1751
rect 7239 1717 7248 1751
rect 7196 1708 7248 1717
rect 7656 1708 7708 1760
rect 8760 1708 8812 1760
rect 9588 1751 9640 1760
rect 9588 1717 9597 1751
rect 9597 1717 9631 1751
rect 9631 1717 9640 1751
rect 9588 1708 9640 1717
rect 10140 1751 10192 1760
rect 10140 1717 10149 1751
rect 10149 1717 10183 1751
rect 10183 1717 10192 1751
rect 10140 1708 10192 1717
rect 10232 1708 10284 1760
rect 10508 1751 10560 1760
rect 10508 1717 10517 1751
rect 10517 1717 10551 1751
rect 10551 1717 10560 1751
rect 10508 1708 10560 1717
rect 11060 1751 11112 1760
rect 11060 1717 11069 1751
rect 11069 1717 11103 1751
rect 11103 1717 11112 1751
rect 11060 1708 11112 1717
rect 11244 1708 11296 1760
rect 11980 1708 12032 1760
rect 13084 1708 13136 1760
rect 13452 1708 13504 1760
rect 14096 1708 14148 1760
rect 14648 1776 14700 1828
rect 15752 1708 15804 1760
rect 17040 1887 17092 1896
rect 17040 1853 17049 1887
rect 17049 1853 17083 1887
rect 17083 1853 17092 1887
rect 17040 1844 17092 1853
rect 18328 1844 18380 1896
rect 22836 1844 22888 1896
rect 3549 1606 3601 1658
rect 3613 1606 3665 1658
rect 3677 1606 3729 1658
rect 3741 1606 3793 1658
rect 3805 1606 3857 1658
rect 8747 1606 8799 1658
rect 8811 1606 8863 1658
rect 8875 1606 8927 1658
rect 8939 1606 8991 1658
rect 9003 1606 9055 1658
rect 13945 1606 13997 1658
rect 14009 1606 14061 1658
rect 14073 1606 14125 1658
rect 14137 1606 14189 1658
rect 14201 1606 14253 1658
rect 19143 1606 19195 1658
rect 19207 1606 19259 1658
rect 19271 1606 19323 1658
rect 19335 1606 19387 1658
rect 19399 1606 19451 1658
rect 1584 1547 1636 1556
rect 1584 1513 1593 1547
rect 1593 1513 1627 1547
rect 1627 1513 1636 1547
rect 1584 1504 1636 1513
rect 388 1300 440 1352
rect 5816 1504 5868 1556
rect 6644 1547 6696 1556
rect 6644 1513 6653 1547
rect 6653 1513 6687 1547
rect 6687 1513 6696 1547
rect 6644 1504 6696 1513
rect 7104 1504 7156 1556
rect 7564 1504 7616 1556
rect 8024 1547 8076 1556
rect 8024 1513 8033 1547
rect 8033 1513 8067 1547
rect 8067 1513 8076 1547
rect 8024 1504 8076 1513
rect 9036 1504 9088 1556
rect 9312 1504 9364 1556
rect 3148 1436 3200 1488
rect 10968 1504 11020 1556
rect 12348 1504 12400 1556
rect 13268 1504 13320 1556
rect 1492 1275 1544 1284
rect 1492 1241 1501 1275
rect 1501 1241 1535 1275
rect 1535 1241 1544 1275
rect 1492 1232 1544 1241
rect 2596 1232 2648 1284
rect 2780 1300 2832 1352
rect 3332 1368 3384 1420
rect 4252 1368 4304 1420
rect 10048 1368 10100 1420
rect 10416 1368 10468 1420
rect 3700 1300 3752 1352
rect 4528 1300 4580 1352
rect 3332 1232 3384 1284
rect 2504 1164 2556 1216
rect 3516 1207 3568 1216
rect 3516 1173 3525 1207
rect 3525 1173 3559 1207
rect 3559 1173 3568 1207
rect 3516 1164 3568 1173
rect 4988 1300 5040 1352
rect 5080 1343 5132 1352
rect 5080 1309 5089 1343
rect 5089 1309 5123 1343
rect 5123 1309 5132 1343
rect 5080 1300 5132 1309
rect 5356 1300 5408 1352
rect 5540 1300 5592 1352
rect 5448 1232 5500 1284
rect 6828 1300 6880 1352
rect 7104 1343 7156 1352
rect 7104 1309 7113 1343
rect 7113 1309 7147 1343
rect 7147 1309 7156 1343
rect 7104 1300 7156 1309
rect 7380 1343 7432 1352
rect 7380 1309 7389 1343
rect 7389 1309 7423 1343
rect 7423 1309 7432 1343
rect 7380 1300 7432 1309
rect 8208 1343 8260 1352
rect 8208 1309 8217 1343
rect 8217 1309 8251 1343
rect 8251 1309 8260 1343
rect 8208 1300 8260 1309
rect 8576 1300 8628 1352
rect 9404 1343 9456 1352
rect 9404 1309 9413 1343
rect 9413 1309 9447 1343
rect 9447 1309 9456 1343
rect 9404 1300 9456 1309
rect 9864 1300 9916 1352
rect 10600 1300 10652 1352
rect 4252 1164 4304 1216
rect 4804 1164 4856 1216
rect 6552 1275 6604 1284
rect 6552 1241 6561 1275
rect 6561 1241 6595 1275
rect 6595 1241 6604 1275
rect 6552 1232 6604 1241
rect 7288 1232 7340 1284
rect 7840 1232 7892 1284
rect 8392 1275 8444 1284
rect 8392 1241 8401 1275
rect 8401 1241 8435 1275
rect 8435 1241 8444 1275
rect 8392 1232 8444 1241
rect 8668 1232 8720 1284
rect 9036 1232 9088 1284
rect 7196 1164 7248 1216
rect 10692 1232 10744 1284
rect 11704 1436 11756 1488
rect 11152 1368 11204 1420
rect 11060 1232 11112 1284
rect 12072 1300 12124 1352
rect 13636 1436 13688 1488
rect 15200 1547 15252 1556
rect 15200 1513 15209 1547
rect 15209 1513 15243 1547
rect 15243 1513 15252 1547
rect 15200 1504 15252 1513
rect 16856 1547 16908 1556
rect 16856 1513 16865 1547
rect 16865 1513 16899 1547
rect 16899 1513 16908 1547
rect 16856 1504 16908 1513
rect 22100 1504 22152 1556
rect 14924 1436 14976 1488
rect 16120 1436 16172 1488
rect 12440 1368 12492 1420
rect 12808 1343 12860 1352
rect 12808 1309 12817 1343
rect 12817 1309 12851 1343
rect 12851 1309 12860 1343
rect 12808 1300 12860 1309
rect 13176 1343 13228 1352
rect 13176 1309 13185 1343
rect 13185 1309 13219 1343
rect 13219 1309 13228 1343
rect 13176 1300 13228 1309
rect 13360 1300 13412 1352
rect 14004 1368 14056 1420
rect 15108 1368 15160 1420
rect 9404 1164 9456 1216
rect 9772 1164 9824 1216
rect 9864 1164 9916 1216
rect 12716 1232 12768 1284
rect 13820 1300 13872 1352
rect 14740 1343 14792 1352
rect 14740 1309 14749 1343
rect 14749 1309 14783 1343
rect 14783 1309 14792 1343
rect 14740 1300 14792 1309
rect 15936 1368 15988 1420
rect 16304 1368 16356 1420
rect 17960 1368 18012 1420
rect 18512 1368 18564 1420
rect 15384 1343 15436 1352
rect 15384 1309 15393 1343
rect 15393 1309 15427 1343
rect 15427 1309 15436 1343
rect 15384 1300 15436 1309
rect 11704 1207 11756 1216
rect 11704 1173 11713 1207
rect 11713 1173 11747 1207
rect 11747 1173 11756 1207
rect 11704 1164 11756 1173
rect 12072 1207 12124 1216
rect 12072 1173 12081 1207
rect 12081 1173 12115 1207
rect 12115 1173 12124 1207
rect 12072 1164 12124 1173
rect 12532 1164 12584 1216
rect 13728 1207 13780 1216
rect 13728 1173 13737 1207
rect 13737 1173 13771 1207
rect 13771 1173 13780 1207
rect 13728 1164 13780 1173
rect 16396 1300 16448 1352
rect 18696 1300 18748 1352
rect 17040 1232 17092 1284
rect 17684 1232 17736 1284
rect 22744 1300 22796 1352
rect 22192 1232 22244 1284
rect 17408 1164 17460 1216
rect 18144 1164 18196 1216
rect 18604 1164 18656 1216
rect 6148 1062 6200 1114
rect 6212 1062 6264 1114
rect 6276 1062 6328 1114
rect 6340 1062 6392 1114
rect 6404 1062 6456 1114
rect 11346 1062 11398 1114
rect 11410 1062 11462 1114
rect 11474 1062 11526 1114
rect 11538 1062 11590 1114
rect 11602 1062 11654 1114
rect 16544 1062 16596 1114
rect 16608 1062 16660 1114
rect 16672 1062 16724 1114
rect 16736 1062 16788 1114
rect 16800 1062 16852 1114
rect 21742 1062 21794 1114
rect 21806 1062 21858 1114
rect 21870 1062 21922 1114
rect 21934 1062 21986 1114
rect 21998 1062 22050 1114
rect 2504 960 2556 1012
rect 4344 960 4396 1012
rect 6460 960 6512 1012
rect 6736 960 6788 1012
rect 6920 960 6972 1012
rect 9864 960 9916 1012
rect 14464 960 14516 1012
rect 17500 960 17552 1012
rect 22928 960 22980 1012
rect 848 892 900 944
rect 4712 892 4764 944
rect 8392 892 8444 944
rect 9404 892 9456 944
rect 11796 892 11848 944
rect 11520 756 11572 808
rect 11888 756 11940 808
rect 2780 688 2832 740
rect 3332 688 3384 740
rect 4528 688 4580 740
rect 5724 688 5776 740
rect 5448 620 5500 672
rect 6184 620 6236 672
rect 9956 620 10008 672
rect 10416 620 10468 672
rect 12900 620 12952 672
rect 13728 620 13780 672
<< metal2 >>
rect 2962 44540 3018 45000
rect 3146 44540 3202 45000
rect 3330 44540 3386 45000
rect 3514 44540 3570 45000
rect 3698 44540 3754 45000
rect 3882 44540 3938 45000
rect 4066 44540 4122 45000
rect 4250 44540 4306 45000
rect 4434 44540 4490 45000
rect 4618 44540 4674 45000
rect 4802 44540 4858 45000
rect 4986 44540 5042 45000
rect 5170 44540 5226 45000
rect 5354 44540 5410 45000
rect 5538 44540 5594 45000
rect 5722 44540 5778 45000
rect 5906 44540 5962 45000
rect 6090 44540 6146 45000
rect 6274 44540 6330 45000
rect 6458 44540 6514 45000
rect 6642 44540 6698 45000
rect 6826 44540 6882 45000
rect 7010 44540 7066 45000
rect 7194 44540 7250 45000
rect 7378 44540 7434 45000
rect 7562 44540 7618 45000
rect 7746 44540 7802 45000
rect 7930 44540 7986 45000
rect 8114 44540 8170 45000
rect 8298 44540 8354 45000
rect 8482 44540 8538 45000
rect 8666 44540 8722 45000
rect 8850 44540 8906 45000
rect 9034 44540 9090 45000
rect 9218 44540 9274 45000
rect 9402 44540 9458 45000
rect 9586 44540 9642 45000
rect 9770 44540 9826 45000
rect 9954 44540 10010 45000
rect 10138 44540 10194 45000
rect 10322 44540 10378 45000
rect 10506 44540 10562 45000
rect 10690 44540 10746 45000
rect 10874 44540 10930 45000
rect 11058 44540 11114 45000
rect 11242 44540 11298 45000
rect 11426 44540 11482 45000
rect 11610 44540 11666 45000
rect 11794 44540 11850 45000
rect 11978 44540 12034 45000
rect 12162 44540 12218 45000
rect 12346 44540 12402 45000
rect 12530 44540 12586 45000
rect 12714 44540 12770 45000
rect 12898 44540 12954 45000
rect 13082 44540 13138 45000
rect 13266 44540 13322 45000
rect 13450 44540 13506 45000
rect 13634 44540 13690 45000
rect 13818 44540 13874 45000
rect 14002 44540 14058 45000
rect 14186 44540 14242 45000
rect 14370 44540 14426 45000
rect 14554 44540 14610 45000
rect 14738 44540 14794 45000
rect 14922 44540 14978 45000
rect 15106 44540 15162 45000
rect 15290 44540 15346 45000
rect 15474 44540 15530 45000
rect 15658 44540 15714 45000
rect 15842 44540 15898 45000
rect 16026 44540 16082 45000
rect 16210 44540 16266 45000
rect 16394 44540 16450 45000
rect 16578 44540 16634 45000
rect 16762 44540 16818 45000
rect 16946 44540 17002 45000
rect 17130 44540 17186 45000
rect 17314 44540 17370 45000
rect 17498 44540 17554 45000
rect 17682 44540 17738 45000
rect 17866 44540 17922 45000
rect 18050 44540 18106 45000
rect 18234 44540 18290 45000
rect 18418 44540 18474 45000
rect 18602 44540 18658 45000
rect 18786 44540 18842 45000
rect 18970 44540 19026 45000
rect 19154 44540 19210 45000
rect 19338 44540 19394 45000
rect 19522 44540 19578 45000
rect 19706 44540 19762 45000
rect 19890 44540 19946 45000
rect 2226 43888 2282 43897
rect 2226 43823 2282 43832
rect 1400 43784 1452 43790
rect 1400 43726 1452 43732
rect 1412 42634 1440 43726
rect 2240 43450 2268 43823
rect 2976 43636 3004 44540
rect 2884 43608 3004 43636
rect 2228 43444 2280 43450
rect 2228 43386 2280 43392
rect 2044 43308 2096 43314
rect 2044 43250 2096 43256
rect 2504 43308 2556 43314
rect 2504 43250 2556 43256
rect 1952 42696 2004 42702
rect 1952 42638 2004 42644
rect 388 42628 440 42634
rect 388 42570 440 42576
rect 1400 42628 1452 42634
rect 1400 42570 1452 42576
rect 18 41440 74 41449
rect 18 41375 74 41384
rect 32 29306 60 41375
rect 296 40520 348 40526
rect 296 40462 348 40468
rect 308 35737 336 40462
rect 294 35728 350 35737
rect 294 35663 350 35672
rect 400 34406 428 42570
rect 938 42256 994 42265
rect 938 42191 994 42200
rect 1860 42220 1912 42226
rect 664 42152 716 42158
rect 664 42094 716 42100
rect 846 42120 902 42129
rect 572 36780 624 36786
rect 572 36722 624 36728
rect 478 35592 534 35601
rect 478 35527 534 35536
rect 388 34400 440 34406
rect 388 34342 440 34348
rect 388 32768 440 32774
rect 388 32710 440 32716
rect 294 29608 350 29617
rect 124 29566 294 29594
rect 20 29300 72 29306
rect 20 29242 72 29248
rect 124 25242 152 29566
rect 294 29543 350 29552
rect 294 29064 350 29073
rect 294 28999 350 29008
rect 32 25214 152 25242
rect 32 25090 60 25214
rect 308 25208 336 28999
rect 216 25180 336 25208
rect 20 25084 72 25090
rect 20 25026 72 25032
rect 216 21350 244 25180
rect 296 25084 348 25090
rect 296 25026 348 25032
rect 204 21344 256 21350
rect 204 21286 256 21292
rect 308 1834 336 25026
rect 296 1828 348 1834
rect 296 1770 348 1776
rect 400 1358 428 32710
rect 492 26926 520 35527
rect 480 26920 532 26926
rect 480 26862 532 26868
rect 480 22092 532 22098
rect 480 22034 532 22040
rect 492 17649 520 22034
rect 478 17640 534 17649
rect 478 17575 534 17584
rect 480 16516 532 16522
rect 480 16458 532 16464
rect 492 13682 520 16458
rect 584 13802 612 36722
rect 676 27441 704 42094
rect 846 42055 902 42064
rect 756 41608 808 41614
rect 756 41550 808 41556
rect 768 37913 796 41550
rect 754 37904 810 37913
rect 754 37839 810 37848
rect 756 32496 808 32502
rect 756 32438 808 32444
rect 768 31929 796 32438
rect 754 31920 810 31929
rect 754 31855 810 31864
rect 754 30016 810 30025
rect 754 29951 810 29960
rect 768 29646 796 29951
rect 756 29640 808 29646
rect 756 29582 808 29588
rect 754 28928 810 28937
rect 754 28863 810 28872
rect 768 28558 796 28863
rect 756 28552 808 28558
rect 756 28494 808 28500
rect 756 28076 808 28082
rect 756 28018 808 28024
rect 768 27849 796 28018
rect 754 27840 810 27849
rect 754 27775 810 27784
rect 756 27736 808 27742
rect 756 27678 808 27684
rect 662 27432 718 27441
rect 662 27367 718 27376
rect 768 24698 796 27678
rect 860 26217 888 42055
rect 846 26208 902 26217
rect 846 26143 902 26152
rect 846 24848 902 24857
rect 846 24783 848 24792
rect 900 24783 902 24792
rect 848 24754 900 24760
rect 768 24670 888 24698
rect 756 24200 808 24206
rect 756 24142 808 24148
rect 768 23769 796 24142
rect 754 23760 810 23769
rect 754 23695 810 23704
rect 664 23520 716 23526
rect 664 23462 716 23468
rect 676 22098 704 23462
rect 664 22092 716 22098
rect 664 22034 716 22040
rect 662 21992 718 22001
rect 662 21927 718 21936
rect 756 21956 808 21962
rect 676 20890 704 21927
rect 756 21898 808 21904
rect 768 21593 796 21898
rect 754 21584 810 21593
rect 754 21519 810 21528
rect 754 21040 810 21049
rect 754 20975 756 20984
rect 808 20975 810 20984
rect 756 20946 808 20952
rect 676 20862 796 20890
rect 768 20058 796 20862
rect 756 20052 808 20058
rect 756 19994 808 20000
rect 754 19952 810 19961
rect 754 19887 810 19896
rect 768 19854 796 19887
rect 756 19848 808 19854
rect 756 19790 808 19796
rect 756 19712 808 19718
rect 756 19654 808 19660
rect 664 19576 716 19582
rect 664 19518 716 19524
rect 676 14657 704 19518
rect 662 14648 718 14657
rect 662 14583 718 14592
rect 572 13796 624 13802
rect 572 13738 624 13744
rect 492 13654 704 13682
rect 572 13592 624 13598
rect 572 13534 624 13540
rect 480 8832 532 8838
rect 480 8774 532 8780
rect 492 3534 520 8774
rect 480 3528 532 3534
rect 480 3470 532 3476
rect 584 1902 612 13534
rect 676 2378 704 13654
rect 664 2372 716 2378
rect 664 2314 716 2320
rect 572 1896 624 1902
rect 572 1838 624 1844
rect 768 1465 796 19654
rect 754 1456 810 1465
rect 754 1391 810 1400
rect 388 1352 440 1358
rect 388 1294 440 1300
rect 860 950 888 24670
rect 952 20602 980 42191
rect 1860 42162 1912 42168
rect 1032 42016 1084 42022
rect 1032 41958 1084 41964
rect 1044 27690 1072 41958
rect 1412 41546 1532 41562
rect 1412 41540 1544 41546
rect 1412 41534 1492 41540
rect 1216 41132 1268 41138
rect 1216 41074 1268 41080
rect 1124 39908 1176 39914
rect 1124 39850 1176 39856
rect 1136 38729 1164 39850
rect 1122 38720 1178 38729
rect 1122 38655 1178 38664
rect 1124 38412 1176 38418
rect 1124 38354 1176 38360
rect 1136 36174 1164 38354
rect 1228 36961 1256 41074
rect 1412 39817 1440 41534
rect 1492 41482 1544 41488
rect 1872 41290 1900 42162
rect 1504 41262 1900 41290
rect 1398 39808 1454 39817
rect 1398 39743 1454 39752
rect 1504 39658 1532 41262
rect 1584 41064 1636 41070
rect 1584 41006 1636 41012
rect 1412 39630 1532 39658
rect 1308 39364 1360 39370
rect 1308 39306 1360 39312
rect 1320 39001 1348 39306
rect 1306 38992 1362 39001
rect 1306 38927 1362 38936
rect 1308 38276 1360 38282
rect 1308 38218 1360 38224
rect 1320 37641 1348 38218
rect 1306 37632 1362 37641
rect 1306 37567 1362 37576
rect 1214 36952 1270 36961
rect 1214 36887 1270 36896
rect 1216 36372 1268 36378
rect 1216 36314 1268 36320
rect 1124 36168 1176 36174
rect 1124 36110 1176 36116
rect 1136 34932 1164 36110
rect 1228 35057 1256 36314
rect 1412 36258 1440 39630
rect 1596 39098 1624 41006
rect 1964 40662 1992 42638
rect 2056 42362 2084 43250
rect 2136 42628 2188 42634
rect 2136 42570 2188 42576
rect 2044 42356 2096 42362
rect 2044 42298 2096 42304
rect 2148 41041 2176 42570
rect 2226 41576 2282 41585
rect 2226 41511 2228 41520
rect 2280 41511 2282 41520
rect 2228 41482 2280 41488
rect 2516 41274 2544 43250
rect 2596 43240 2648 43246
rect 2596 43182 2648 43188
rect 2504 41268 2556 41274
rect 2504 41210 2556 41216
rect 2134 41032 2190 41041
rect 2134 40967 2190 40976
rect 1952 40656 2004 40662
rect 1952 40598 2004 40604
rect 1952 40520 2004 40526
rect 1952 40462 2004 40468
rect 2044 40520 2096 40526
rect 2044 40462 2096 40468
rect 1676 40452 1728 40458
rect 1676 40394 1728 40400
rect 1688 40089 1716 40394
rect 1674 40080 1730 40089
rect 1674 40015 1730 40024
rect 1768 40044 1820 40050
rect 1768 39986 1820 39992
rect 1676 39432 1728 39438
rect 1676 39374 1728 39380
rect 1584 39092 1636 39098
rect 1584 39034 1636 39040
rect 1688 38894 1716 39374
rect 1676 38888 1728 38894
rect 1676 38830 1728 38836
rect 1492 38752 1544 38758
rect 1676 38752 1728 38758
rect 1544 38712 1624 38740
rect 1492 38694 1544 38700
rect 1492 37868 1544 37874
rect 1492 37810 1544 37816
rect 1320 36230 1440 36258
rect 1320 35494 1348 36230
rect 1400 36168 1452 36174
rect 1400 36110 1452 36116
rect 1308 35488 1360 35494
rect 1308 35430 1360 35436
rect 1214 35048 1270 35057
rect 1214 34983 1270 34992
rect 1308 34944 1360 34950
rect 1136 34904 1256 34932
rect 1124 32972 1176 32978
rect 1124 32914 1176 32920
rect 1136 30734 1164 32914
rect 1124 30728 1176 30734
rect 1124 30670 1176 30676
rect 1228 30410 1256 34904
rect 1308 34886 1360 34892
rect 1320 32348 1348 34886
rect 1412 33674 1440 36110
rect 1504 35057 1532 37810
rect 1596 36378 1624 38712
rect 1676 38694 1728 38700
rect 1688 36786 1716 38694
rect 1676 36780 1728 36786
rect 1676 36722 1728 36728
rect 1584 36372 1636 36378
rect 1584 36314 1636 36320
rect 1584 36032 1636 36038
rect 1584 35974 1636 35980
rect 1490 35048 1546 35057
rect 1490 34983 1546 34992
rect 1412 33646 1532 33674
rect 1400 33516 1452 33522
rect 1400 33458 1452 33464
rect 1412 32586 1440 33458
rect 1504 33289 1532 33646
rect 1490 33280 1546 33289
rect 1490 33215 1546 33224
rect 1596 32978 1624 35974
rect 1688 35329 1716 36722
rect 1780 36145 1808 39986
rect 1860 39432 1912 39438
rect 1860 39374 1912 39380
rect 1872 39030 1900 39374
rect 1860 39024 1912 39030
rect 1860 38966 1912 38972
rect 1872 38350 1900 38966
rect 1860 38344 1912 38350
rect 1860 38286 1912 38292
rect 1860 37800 1912 37806
rect 1860 37742 1912 37748
rect 1872 37466 1900 37742
rect 1860 37460 1912 37466
rect 1860 37402 1912 37408
rect 1964 37233 1992 40462
rect 2056 38593 2084 40462
rect 2228 40452 2280 40458
rect 2228 40394 2280 40400
rect 2136 40180 2188 40186
rect 2136 40122 2188 40128
rect 2042 38584 2098 38593
rect 2042 38519 2098 38528
rect 2148 38434 2176 40122
rect 2056 38406 2176 38434
rect 1950 37224 2006 37233
rect 1950 37159 2006 37168
rect 1860 37120 1912 37126
rect 1860 37062 1912 37068
rect 1872 36718 1900 37062
rect 1860 36712 1912 36718
rect 1860 36654 1912 36660
rect 1766 36136 1822 36145
rect 1766 36071 1822 36080
rect 1768 35624 1820 35630
rect 1768 35566 1820 35572
rect 1674 35320 1730 35329
rect 1674 35255 1730 35264
rect 1780 35222 1808 35566
rect 1768 35216 1820 35222
rect 1768 35158 1820 35164
rect 1768 35080 1820 35086
rect 1768 35022 1820 35028
rect 1676 35012 1728 35018
rect 1676 34954 1728 34960
rect 1688 33969 1716 34954
rect 1674 33960 1730 33969
rect 1674 33895 1730 33904
rect 1780 32994 1808 35022
rect 1872 34950 1900 36654
rect 1860 34944 1912 34950
rect 2056 34932 2084 38406
rect 2240 36038 2268 40394
rect 2608 40100 2636 43182
rect 2884 42770 2912 43608
rect 3160 43450 3188 44540
rect 3344 43874 3372 44540
rect 3252 43846 3372 43874
rect 3148 43444 3200 43450
rect 3148 43386 3200 43392
rect 3056 43308 3108 43314
rect 3056 43250 3108 43256
rect 2964 43172 3016 43178
rect 2964 43114 3016 43120
rect 2872 42764 2924 42770
rect 2872 42706 2924 42712
rect 2976 42702 3004 43114
rect 2964 42696 3016 42702
rect 2964 42638 3016 42644
rect 2688 42628 2740 42634
rect 2688 42570 2740 42576
rect 2780 42628 2832 42634
rect 2780 42570 2832 42576
rect 2700 41818 2728 42570
rect 2792 42362 2820 42570
rect 3068 42566 3096 43250
rect 3252 42922 3280 43846
rect 3528 43738 3556 44540
rect 3344 43710 3556 43738
rect 3344 43450 3372 43710
rect 3712 43602 3740 44540
rect 3896 43897 3924 44540
rect 3882 43888 3938 43897
rect 3882 43823 3938 43832
rect 3436 43574 3740 43602
rect 3332 43444 3384 43450
rect 3332 43386 3384 43392
rect 3160 42894 3280 42922
rect 3160 42770 3188 42894
rect 3436 42770 3464 43574
rect 3976 43308 4028 43314
rect 3976 43250 4028 43256
rect 3549 43004 3857 43013
rect 3549 43002 3555 43004
rect 3611 43002 3635 43004
rect 3691 43002 3715 43004
rect 3771 43002 3795 43004
rect 3851 43002 3857 43004
rect 3611 42950 3613 43002
rect 3793 42950 3795 43002
rect 3549 42948 3555 42950
rect 3611 42948 3635 42950
rect 3691 42948 3715 42950
rect 3771 42948 3795 42950
rect 3851 42948 3857 42950
rect 3549 42939 3857 42948
rect 3148 42764 3200 42770
rect 3148 42706 3200 42712
rect 3424 42764 3476 42770
rect 3424 42706 3476 42712
rect 3056 42560 3108 42566
rect 3056 42502 3108 42508
rect 2780 42356 2832 42362
rect 2780 42298 2832 42304
rect 3240 42220 3292 42226
rect 3240 42162 3292 42168
rect 3332 42220 3384 42226
rect 3332 42162 3384 42168
rect 3884 42220 3936 42226
rect 3884 42162 3936 42168
rect 2688 41812 2740 41818
rect 2688 41754 2740 41760
rect 2964 41608 3016 41614
rect 2964 41550 3016 41556
rect 2780 41132 2832 41138
rect 2780 41074 2832 41080
rect 2516 40072 2636 40100
rect 2410 39808 2466 39817
rect 2410 39743 2466 39752
rect 2320 38752 2372 38758
rect 2320 38694 2372 38700
rect 2332 37482 2360 38694
rect 2424 37913 2452 39743
rect 2516 39681 2544 40072
rect 2688 40044 2740 40050
rect 2688 39986 2740 39992
rect 2596 39976 2648 39982
rect 2596 39918 2648 39924
rect 2502 39672 2558 39681
rect 2502 39607 2558 39616
rect 2504 39296 2556 39302
rect 2504 39238 2556 39244
rect 2410 37904 2466 37913
rect 2410 37839 2466 37848
rect 2516 37806 2544 39238
rect 2608 39114 2636 39918
rect 2700 39386 2728 39986
rect 2792 39545 2820 41074
rect 2872 40996 2924 41002
rect 2872 40938 2924 40944
rect 2778 39536 2834 39545
rect 2778 39471 2834 39480
rect 2700 39358 2820 39386
rect 2608 39086 2728 39114
rect 2596 38956 2648 38962
rect 2596 38898 2648 38904
rect 2504 37800 2556 37806
rect 2410 37768 2466 37777
rect 2504 37742 2556 37748
rect 2410 37703 2412 37712
rect 2464 37703 2466 37712
rect 2412 37674 2464 37680
rect 2332 37454 2452 37482
rect 2320 37392 2372 37398
rect 2320 37334 2372 37340
rect 2228 36032 2280 36038
rect 2228 35974 2280 35980
rect 2136 35624 2188 35630
rect 2136 35566 2188 35572
rect 2148 35086 2176 35566
rect 2228 35556 2280 35562
rect 2228 35498 2280 35504
rect 2136 35080 2188 35086
rect 2136 35022 2188 35028
rect 2056 34904 2176 34932
rect 1860 34886 1912 34892
rect 2148 34746 2176 34904
rect 2240 34762 2268 35498
rect 2332 34950 2360 37334
rect 2424 36961 2452 37454
rect 2410 36952 2466 36961
rect 2410 36887 2466 36896
rect 2424 36718 2452 36887
rect 2504 36780 2556 36786
rect 2504 36722 2556 36728
rect 2412 36712 2464 36718
rect 2412 36654 2464 36660
rect 2412 36576 2464 36582
rect 2412 36518 2464 36524
rect 2424 35630 2452 36518
rect 2412 35624 2464 35630
rect 2412 35566 2464 35572
rect 2320 34944 2372 34950
rect 2516 34932 2544 36722
rect 2608 36174 2636 38898
rect 2700 38729 2728 39086
rect 2686 38720 2742 38729
rect 2686 38655 2742 38664
rect 2688 38208 2740 38214
rect 2688 38150 2740 38156
rect 2596 36168 2648 36174
rect 2596 36110 2648 36116
rect 2596 36032 2648 36038
rect 2596 35974 2648 35980
rect 2608 35086 2636 35974
rect 2700 35154 2728 38150
rect 2792 37369 2820 39358
rect 2884 38321 2912 40938
rect 2976 39273 3004 41550
rect 3148 40112 3200 40118
rect 3148 40054 3200 40060
rect 3056 39500 3108 39506
rect 3056 39442 3108 39448
rect 2962 39264 3018 39273
rect 2962 39199 3018 39208
rect 2964 39024 3016 39030
rect 2964 38966 3016 38972
rect 2976 38894 3004 38966
rect 2964 38888 3016 38894
rect 2964 38830 3016 38836
rect 2976 38457 3004 38830
rect 2962 38448 3018 38457
rect 2962 38383 3018 38392
rect 2870 38312 2926 38321
rect 2870 38247 2926 38256
rect 3068 38162 3096 39442
rect 3160 39030 3188 40054
rect 3148 39024 3200 39030
rect 3148 38966 3200 38972
rect 3148 38752 3200 38758
rect 3148 38694 3200 38700
rect 2976 38134 3096 38162
rect 2872 37800 2924 37806
rect 2872 37742 2924 37748
rect 2884 37398 2912 37742
rect 2872 37392 2924 37398
rect 2778 37360 2834 37369
rect 2872 37334 2924 37340
rect 2778 37295 2834 37304
rect 2976 37210 3004 38134
rect 3160 37874 3188 38694
rect 3252 38010 3280 42162
rect 3344 41818 3372 42162
rect 3549 41916 3857 41925
rect 3549 41914 3555 41916
rect 3611 41914 3635 41916
rect 3691 41914 3715 41916
rect 3771 41914 3795 41916
rect 3851 41914 3857 41916
rect 3611 41862 3613 41914
rect 3793 41862 3795 41914
rect 3549 41860 3555 41862
rect 3611 41860 3635 41862
rect 3691 41860 3715 41862
rect 3771 41860 3795 41862
rect 3851 41860 3857 41862
rect 3549 41851 3857 41860
rect 3896 41818 3924 42162
rect 3988 41818 4016 43250
rect 4080 42362 4108 44540
rect 4160 43172 4212 43178
rect 4160 43114 4212 43120
rect 4068 42356 4120 42362
rect 4068 42298 4120 42304
rect 4172 42242 4200 43114
rect 4264 42362 4292 44540
rect 4344 43308 4396 43314
rect 4448 43296 4476 44540
rect 4448 43268 4568 43296
rect 4344 43250 4396 43256
rect 4356 42945 4384 43250
rect 4342 42936 4398 42945
rect 4342 42871 4398 42880
rect 4436 42832 4488 42838
rect 4356 42780 4436 42786
rect 4356 42774 4488 42780
rect 4356 42758 4476 42774
rect 4252 42356 4304 42362
rect 4252 42298 4304 42304
rect 4080 42214 4200 42242
rect 3332 41812 3384 41818
rect 3332 41754 3384 41760
rect 3884 41812 3936 41818
rect 3884 41754 3936 41760
rect 3976 41812 4028 41818
rect 3976 41754 4028 41760
rect 4080 41750 4108 42214
rect 4068 41744 4120 41750
rect 4068 41686 4120 41692
rect 4250 41712 4306 41721
rect 4250 41647 4306 41656
rect 4264 41614 4292 41647
rect 3608 41608 3660 41614
rect 3608 41550 3660 41556
rect 3976 41608 4028 41614
rect 3976 41550 4028 41556
rect 4252 41608 4304 41614
rect 4252 41550 4304 41556
rect 3620 41449 3648 41550
rect 3606 41440 3662 41449
rect 3606 41375 3662 41384
rect 3549 40828 3857 40837
rect 3549 40826 3555 40828
rect 3611 40826 3635 40828
rect 3691 40826 3715 40828
rect 3771 40826 3795 40828
rect 3851 40826 3857 40828
rect 3611 40774 3613 40826
rect 3793 40774 3795 40826
rect 3549 40772 3555 40774
rect 3611 40772 3635 40774
rect 3691 40772 3715 40774
rect 3771 40772 3795 40774
rect 3851 40772 3857 40774
rect 3549 40763 3857 40772
rect 3988 40497 4016 41550
rect 4160 41540 4212 41546
rect 4160 41482 4212 41488
rect 4172 41414 4200 41482
rect 4356 41414 4384 42758
rect 4540 42362 4568 43268
rect 4632 42770 4660 44540
rect 4712 43308 4764 43314
rect 4712 43250 4764 43256
rect 4620 42764 4672 42770
rect 4620 42706 4672 42712
rect 4528 42356 4580 42362
rect 4528 42298 4580 42304
rect 4724 41818 4752 43250
rect 4816 42362 4844 44540
rect 5000 42770 5028 44540
rect 5080 43852 5132 43858
rect 5080 43794 5132 43800
rect 5092 43246 5120 43794
rect 5184 43450 5212 44540
rect 5172 43444 5224 43450
rect 5172 43386 5224 43392
rect 5264 43444 5316 43450
rect 5368 43432 5396 44540
rect 5552 43466 5580 44540
rect 5460 43450 5580 43466
rect 5316 43404 5396 43432
rect 5448 43444 5580 43450
rect 5264 43386 5316 43392
rect 5500 43438 5580 43444
rect 5448 43386 5500 43392
rect 5540 43308 5592 43314
rect 5736 43296 5764 44540
rect 5816 43444 5868 43450
rect 5920 43432 5948 44540
rect 6104 43636 6132 44540
rect 6288 43858 6316 44540
rect 6276 43852 6328 43858
rect 6276 43794 6328 43800
rect 5868 43404 5948 43432
rect 6012 43608 6132 43636
rect 6472 43636 6500 44540
rect 6472 43608 6592 43636
rect 5816 43386 5868 43392
rect 5540 43250 5592 43256
rect 5644 43268 5764 43296
rect 5080 43240 5132 43246
rect 5080 43182 5132 43188
rect 4988 42764 5040 42770
rect 4988 42706 5040 42712
rect 4896 42628 4948 42634
rect 4896 42570 4948 42576
rect 5080 42628 5132 42634
rect 5080 42570 5132 42576
rect 4804 42356 4856 42362
rect 4804 42298 4856 42304
rect 4712 41812 4764 41818
rect 4712 41754 4764 41760
rect 4528 41608 4580 41614
rect 4526 41576 4528 41585
rect 4804 41608 4856 41614
rect 4580 41576 4582 41585
rect 4804 41550 4856 41556
rect 4526 41511 4582 41520
rect 4172 41386 4292 41414
rect 4356 41386 4660 41414
rect 4160 41132 4212 41138
rect 4160 41074 4212 41080
rect 4068 41064 4120 41070
rect 4068 41006 4120 41012
rect 3974 40488 4030 40497
rect 3974 40423 4030 40432
rect 3424 39976 3476 39982
rect 3424 39918 3476 39924
rect 3332 39024 3384 39030
rect 3332 38966 3384 38972
rect 3240 38004 3292 38010
rect 3240 37946 3292 37952
rect 3148 37868 3200 37874
rect 3148 37810 3200 37816
rect 3148 37664 3200 37670
rect 3148 37606 3200 37612
rect 3160 37262 3188 37606
rect 2884 37182 3004 37210
rect 3056 37256 3108 37262
rect 3056 37198 3108 37204
rect 3148 37256 3200 37262
rect 3148 37198 3200 37204
rect 2884 36281 2912 37182
rect 2964 37120 3016 37126
rect 2964 37062 3016 37068
rect 2870 36272 2926 36281
rect 2870 36207 2926 36216
rect 2872 35828 2924 35834
rect 2872 35770 2924 35776
rect 2780 35624 2832 35630
rect 2780 35566 2832 35572
rect 2688 35148 2740 35154
rect 2688 35090 2740 35096
rect 2596 35080 2648 35086
rect 2596 35022 2648 35028
rect 2516 34904 2636 34932
rect 2320 34886 2372 34892
rect 2136 34740 2188 34746
rect 2240 34734 2544 34762
rect 2136 34682 2188 34688
rect 2320 34672 2372 34678
rect 2320 34614 2372 34620
rect 2044 34604 2096 34610
rect 2096 34564 2176 34592
rect 2044 34546 2096 34552
rect 1860 33924 1912 33930
rect 1860 33866 1912 33872
rect 1872 33697 1900 33866
rect 1858 33688 1914 33697
rect 1858 33623 1914 33632
rect 1952 33516 2004 33522
rect 1952 33458 2004 33464
rect 1584 32972 1636 32978
rect 1780 32966 1900 32994
rect 1584 32914 1636 32920
rect 1492 32836 1544 32842
rect 1492 32778 1544 32784
rect 1768 32836 1820 32842
rect 1768 32778 1820 32784
rect 1504 32722 1532 32778
rect 1504 32694 1716 32722
rect 1412 32558 1532 32586
rect 1400 32360 1452 32366
rect 1320 32320 1400 32348
rect 1320 31414 1348 32320
rect 1400 32302 1452 32308
rect 1400 31816 1452 31822
rect 1400 31758 1452 31764
rect 1308 31408 1360 31414
rect 1308 31350 1360 31356
rect 1412 30433 1440 31758
rect 1504 31657 1532 32558
rect 1584 32224 1636 32230
rect 1584 32166 1636 32172
rect 1490 31648 1546 31657
rect 1490 31583 1546 31592
rect 1492 31408 1544 31414
rect 1492 31350 1544 31356
rect 1504 31249 1532 31350
rect 1490 31240 1546 31249
rect 1490 31175 1546 31184
rect 1492 31136 1544 31142
rect 1492 31078 1544 31084
rect 1504 30938 1532 31078
rect 1492 30932 1544 30938
rect 1492 30874 1544 30880
rect 1398 30424 1454 30433
rect 1228 30382 1348 30410
rect 1320 29102 1348 30382
rect 1398 30359 1454 30368
rect 1504 30258 1532 30874
rect 1400 30252 1452 30258
rect 1400 30194 1452 30200
rect 1492 30252 1544 30258
rect 1492 30194 1544 30200
rect 1308 29096 1360 29102
rect 1308 29038 1360 29044
rect 1412 28506 1440 30194
rect 1490 29880 1546 29889
rect 1490 29815 1546 29824
rect 1504 29209 1532 29815
rect 1490 29200 1546 29209
rect 1490 29135 1546 29144
rect 1596 28558 1624 32166
rect 1688 30569 1716 32694
rect 1780 32337 1808 32778
rect 1872 32473 1900 32966
rect 1858 32464 1914 32473
rect 1858 32399 1914 32408
rect 1766 32328 1822 32337
rect 1964 32314 1992 33458
rect 2044 33448 2096 33454
rect 2044 33390 2096 33396
rect 1766 32263 1822 32272
rect 1872 32286 1992 32314
rect 1872 32201 1900 32286
rect 1858 32192 1914 32201
rect 1858 32127 1914 32136
rect 1950 31920 2006 31929
rect 1950 31855 2006 31864
rect 1768 31816 1820 31822
rect 1860 31816 1912 31822
rect 1768 31758 1820 31764
rect 1858 31784 1860 31793
rect 1912 31784 1914 31793
rect 1674 30560 1730 30569
rect 1674 30495 1730 30504
rect 1780 30394 1808 31758
rect 1858 31719 1914 31728
rect 1860 31680 1912 31686
rect 1860 31622 1912 31628
rect 1768 30388 1820 30394
rect 1768 30330 1820 30336
rect 1872 29578 1900 31622
rect 1964 30326 1992 31855
rect 2056 31634 2084 33390
rect 2148 32978 2176 34564
rect 2228 33448 2280 33454
rect 2228 33390 2280 33396
rect 2136 32972 2188 32978
rect 2136 32914 2188 32920
rect 2148 31793 2176 32914
rect 2240 32473 2268 33390
rect 2226 32464 2282 32473
rect 2332 32434 2360 34614
rect 2412 33856 2464 33862
rect 2412 33798 2464 33804
rect 2424 33114 2452 33798
rect 2412 33108 2464 33114
rect 2412 33050 2464 33056
rect 2226 32399 2282 32408
rect 2320 32428 2372 32434
rect 2134 31784 2190 31793
rect 2134 31719 2190 31728
rect 2056 31606 2176 31634
rect 2148 31414 2176 31606
rect 2136 31408 2188 31414
rect 2136 31350 2188 31356
rect 2044 31340 2096 31346
rect 2044 31282 2096 31288
rect 1952 30320 2004 30326
rect 1952 30262 2004 30268
rect 1676 29572 1728 29578
rect 1676 29514 1728 29520
rect 1860 29572 1912 29578
rect 1860 29514 1912 29520
rect 1688 29209 1716 29514
rect 1768 29504 1820 29510
rect 1768 29446 1820 29452
rect 1674 29200 1730 29209
rect 1674 29135 1730 29144
rect 1780 28642 1808 29446
rect 1950 29336 2006 29345
rect 1950 29271 2006 29280
rect 1860 28960 1912 28966
rect 1860 28902 1912 28908
rect 1872 28694 1900 28902
rect 1688 28614 1808 28642
rect 1860 28688 1912 28694
rect 1860 28630 1912 28636
rect 1584 28552 1636 28558
rect 1412 28478 1532 28506
rect 1584 28494 1636 28500
rect 1398 28384 1454 28393
rect 1398 28319 1454 28328
rect 1214 27704 1270 27713
rect 1044 27662 1214 27690
rect 1214 27639 1270 27648
rect 1308 27396 1360 27402
rect 1308 27338 1360 27344
rect 1320 27305 1348 27338
rect 1306 27296 1362 27305
rect 1306 27231 1362 27240
rect 1216 27124 1268 27130
rect 1216 27066 1268 27072
rect 1032 26920 1084 26926
rect 1032 26862 1084 26868
rect 940 20596 992 20602
rect 940 20538 992 20544
rect 1044 18970 1072 26862
rect 1228 26761 1256 27066
rect 1308 27056 1360 27062
rect 1306 27024 1308 27033
rect 1360 27024 1362 27033
rect 1412 26994 1440 28319
rect 1504 27577 1532 28478
rect 1584 28416 1636 28422
rect 1584 28358 1636 28364
rect 1490 27568 1546 27577
rect 1490 27503 1546 27512
rect 1596 27470 1624 28358
rect 1688 28082 1716 28614
rect 1768 28552 1820 28558
rect 1768 28494 1820 28500
rect 1676 28076 1728 28082
rect 1676 28018 1728 28024
rect 1674 27976 1730 27985
rect 1674 27911 1676 27920
rect 1728 27911 1730 27920
rect 1676 27882 1728 27888
rect 1676 27668 1728 27674
rect 1676 27610 1728 27616
rect 1584 27464 1636 27470
rect 1584 27406 1636 27412
rect 1306 26959 1362 26968
rect 1400 26988 1452 26994
rect 1400 26930 1452 26936
rect 1492 26988 1544 26994
rect 1492 26930 1544 26936
rect 1398 26888 1454 26897
rect 1398 26823 1454 26832
rect 1214 26752 1270 26761
rect 1214 26687 1270 26696
rect 1412 26450 1440 26823
rect 1400 26444 1452 26450
rect 1400 26386 1452 26392
rect 1412 25378 1440 26386
rect 1320 25350 1440 25378
rect 1320 24290 1348 25350
rect 1400 25288 1452 25294
rect 1400 25230 1452 25236
rect 1412 24449 1440 25230
rect 1504 25129 1532 26930
rect 1596 26314 1624 27406
rect 1584 26308 1636 26314
rect 1584 26250 1636 26256
rect 1584 25900 1636 25906
rect 1584 25842 1636 25848
rect 1490 25120 1546 25129
rect 1490 25055 1546 25064
rect 1490 24984 1546 24993
rect 1490 24919 1546 24928
rect 1398 24440 1454 24449
rect 1398 24375 1454 24384
rect 1400 24336 1452 24342
rect 1320 24284 1400 24290
rect 1320 24278 1452 24284
rect 1320 24262 1440 24278
rect 1412 23730 1440 24262
rect 1504 24206 1532 24919
rect 1492 24200 1544 24206
rect 1492 24142 1544 24148
rect 1596 24041 1624 25842
rect 1688 25362 1716 27610
rect 1780 26489 1808 28494
rect 1872 28490 1900 28630
rect 1860 28484 1912 28490
rect 1860 28426 1912 28432
rect 1964 28370 1992 29271
rect 2056 29238 2084 31282
rect 2136 30728 2188 30734
rect 2136 30670 2188 30676
rect 2044 29232 2096 29238
rect 2044 29174 2096 29180
rect 1872 28342 1992 28370
rect 1872 27470 1900 28342
rect 1952 28076 2004 28082
rect 1952 28018 2004 28024
rect 1860 27464 1912 27470
rect 1860 27406 1912 27412
rect 1872 27169 1900 27406
rect 1858 27160 1914 27169
rect 1858 27095 1914 27104
rect 1858 26616 1914 26625
rect 1858 26551 1914 26560
rect 1766 26480 1822 26489
rect 1766 26415 1822 26424
rect 1766 26344 1822 26353
rect 1766 26279 1822 26288
rect 1676 25356 1728 25362
rect 1676 25298 1728 25304
rect 1780 24410 1808 26279
rect 1872 25922 1900 26551
rect 1964 26217 1992 28018
rect 2056 26926 2084 29174
rect 2044 26920 2096 26926
rect 2044 26862 2096 26868
rect 2148 26738 2176 30670
rect 2240 29345 2268 32399
rect 2320 32370 2372 32376
rect 2412 32020 2464 32026
rect 2332 31980 2412 32008
rect 2332 30682 2360 31980
rect 2412 31962 2464 31968
rect 2516 31906 2544 34734
rect 2608 34610 2636 34904
rect 2596 34604 2648 34610
rect 2596 34546 2648 34552
rect 2792 34134 2820 35566
rect 2884 34950 2912 35770
rect 2976 35698 3004 37062
rect 2964 35692 3016 35698
rect 2964 35634 3016 35640
rect 3068 35193 3096 37198
rect 3240 37188 3292 37194
rect 3240 37130 3292 37136
rect 3148 35624 3200 35630
rect 3148 35566 3200 35572
rect 3054 35184 3110 35193
rect 3054 35119 3110 35128
rect 3054 35048 3110 35057
rect 2976 35006 3054 35034
rect 2872 34944 2924 34950
rect 2872 34886 2924 34892
rect 2976 34542 3004 35006
rect 3054 34983 3110 34992
rect 3056 34944 3108 34950
rect 3056 34886 3108 34892
rect 2964 34536 3016 34542
rect 2964 34478 3016 34484
rect 2872 34400 2924 34406
rect 2872 34342 2924 34348
rect 2780 34128 2832 34134
rect 2780 34070 2832 34076
rect 2688 34060 2740 34066
rect 2688 34002 2740 34008
rect 2596 33856 2648 33862
rect 2596 33798 2648 33804
rect 2608 32366 2636 33798
rect 2596 32360 2648 32366
rect 2596 32302 2648 32308
rect 2594 31920 2650 31929
rect 2412 31884 2464 31890
rect 2516 31878 2594 31906
rect 2594 31855 2650 31864
rect 2412 31826 2464 31832
rect 2424 31482 2452 31826
rect 2700 31804 2728 34002
rect 2780 33584 2832 33590
rect 2780 33526 2832 33532
rect 2792 32570 2820 33526
rect 2884 33454 2912 34342
rect 2964 33992 3016 33998
rect 2964 33934 3016 33940
rect 2872 33448 2924 33454
rect 2872 33390 2924 33396
rect 2976 32745 3004 33934
rect 2962 32736 3018 32745
rect 2962 32671 3018 32680
rect 2780 32564 2832 32570
rect 2780 32506 2832 32512
rect 2962 32328 3018 32337
rect 2792 32286 2962 32314
rect 2792 31890 2820 32286
rect 2962 32263 3018 32272
rect 2964 32224 3016 32230
rect 2964 32166 3016 32172
rect 2780 31884 2832 31890
rect 2780 31826 2832 31832
rect 2976 31822 3004 32166
rect 2516 31776 2728 31804
rect 2964 31816 3016 31822
rect 2412 31476 2464 31482
rect 2412 31418 2464 31424
rect 2516 31346 2544 31776
rect 2964 31758 3016 31764
rect 2780 31476 2832 31482
rect 2780 31418 2832 31424
rect 2596 31408 2648 31414
rect 2596 31350 2648 31356
rect 2504 31340 2556 31346
rect 2504 31282 2556 31288
rect 2608 31249 2636 31350
rect 2792 31346 2820 31418
rect 2688 31340 2740 31346
rect 2688 31282 2740 31288
rect 2780 31340 2832 31346
rect 2780 31282 2832 31288
rect 2410 31240 2466 31249
rect 2410 31175 2466 31184
rect 2594 31240 2650 31249
rect 2594 31175 2650 31184
rect 2424 30938 2452 31175
rect 2700 31113 2728 31282
rect 2872 31272 2924 31278
rect 2872 31214 2924 31220
rect 2686 31104 2742 31113
rect 2686 31039 2742 31048
rect 2412 30932 2464 30938
rect 2412 30874 2464 30880
rect 2884 30818 2912 31214
rect 2700 30790 2912 30818
rect 2964 30864 3016 30870
rect 2964 30806 3016 30812
rect 2594 30696 2650 30705
rect 2332 30654 2452 30682
rect 2320 30592 2372 30598
rect 2320 30534 2372 30540
rect 2332 29714 2360 30534
rect 2424 30326 2452 30654
rect 2594 30631 2650 30640
rect 2412 30320 2464 30326
rect 2412 30262 2464 30268
rect 2502 30152 2558 30161
rect 2502 30087 2558 30096
rect 2320 29708 2372 29714
rect 2320 29650 2372 29656
rect 2516 29578 2544 30087
rect 2504 29572 2556 29578
rect 2504 29514 2556 29520
rect 2608 29458 2636 30631
rect 2700 30598 2728 30790
rect 2780 30728 2832 30734
rect 2872 30728 2924 30734
rect 2780 30670 2832 30676
rect 2870 30696 2872 30705
rect 2924 30696 2926 30705
rect 2688 30592 2740 30598
rect 2688 30534 2740 30540
rect 2688 30048 2740 30054
rect 2688 29990 2740 29996
rect 2700 29646 2728 29990
rect 2792 29753 2820 30670
rect 2870 30631 2926 30640
rect 2872 30592 2924 30598
rect 2872 30534 2924 30540
rect 2884 30190 2912 30534
rect 2872 30184 2924 30190
rect 2872 30126 2924 30132
rect 2778 29744 2834 29753
rect 2778 29679 2834 29688
rect 2688 29640 2740 29646
rect 2688 29582 2740 29588
rect 2332 29430 2636 29458
rect 2226 29336 2282 29345
rect 2226 29271 2282 29280
rect 2332 29034 2360 29430
rect 2596 29300 2648 29306
rect 2596 29242 2648 29248
rect 2412 29232 2464 29238
rect 2412 29174 2464 29180
rect 2320 29028 2372 29034
rect 2320 28970 2372 28976
rect 2332 27962 2360 28970
rect 2424 28966 2452 29174
rect 2412 28960 2464 28966
rect 2412 28902 2464 28908
rect 2504 28552 2556 28558
rect 2424 28512 2504 28540
rect 2424 28393 2452 28512
rect 2504 28494 2556 28500
rect 2504 28416 2556 28422
rect 2410 28384 2466 28393
rect 2504 28358 2556 28364
rect 2410 28319 2466 28328
rect 2516 28150 2544 28358
rect 2608 28257 2636 29242
rect 2884 29238 2912 30126
rect 2976 29646 3004 30806
rect 3068 30054 3096 34886
rect 3160 33833 3188 35566
rect 3252 34921 3280 37130
rect 3344 36786 3372 38966
rect 3436 38894 3464 39918
rect 4080 39846 4108 41006
rect 4068 39840 4120 39846
rect 4068 39782 4120 39788
rect 3549 39740 3857 39749
rect 3549 39738 3555 39740
rect 3611 39738 3635 39740
rect 3691 39738 3715 39740
rect 3771 39738 3795 39740
rect 3851 39738 3857 39740
rect 3611 39686 3613 39738
rect 3793 39686 3795 39738
rect 3549 39684 3555 39686
rect 3611 39684 3635 39686
rect 3691 39684 3715 39686
rect 3771 39684 3795 39686
rect 3851 39684 3857 39686
rect 3549 39675 3857 39684
rect 3700 39500 3752 39506
rect 3700 39442 3752 39448
rect 3712 38962 3740 39442
rect 3976 39364 4028 39370
rect 3976 39306 4028 39312
rect 3700 38956 3752 38962
rect 3700 38898 3752 38904
rect 3424 38888 3476 38894
rect 3424 38830 3476 38836
rect 3884 38752 3936 38758
rect 3884 38694 3936 38700
rect 3549 38652 3857 38661
rect 3549 38650 3555 38652
rect 3611 38650 3635 38652
rect 3691 38650 3715 38652
rect 3771 38650 3795 38652
rect 3851 38650 3857 38652
rect 3611 38598 3613 38650
rect 3793 38598 3795 38650
rect 3549 38596 3555 38598
rect 3611 38596 3635 38598
rect 3691 38596 3715 38598
rect 3771 38596 3795 38598
rect 3851 38596 3857 38598
rect 3549 38587 3857 38596
rect 3896 38418 3924 38694
rect 3988 38654 4016 39306
rect 4172 39302 4200 41074
rect 4160 39296 4212 39302
rect 4160 39238 4212 39244
rect 3988 38626 4108 38654
rect 3884 38412 3936 38418
rect 3884 38354 3936 38360
rect 4080 38350 4108 38626
rect 4264 38593 4292 41386
rect 4344 40656 4396 40662
rect 4344 40598 4396 40604
rect 4250 38584 4306 38593
rect 4250 38519 4306 38528
rect 4068 38344 4120 38350
rect 4068 38286 4120 38292
rect 3424 38276 3476 38282
rect 3424 38218 3476 38224
rect 3436 37913 3464 38218
rect 3422 37904 3478 37913
rect 3422 37839 3478 37848
rect 3884 37868 3936 37874
rect 3884 37810 3936 37816
rect 3549 37564 3857 37573
rect 3549 37562 3555 37564
rect 3611 37562 3635 37564
rect 3691 37562 3715 37564
rect 3771 37562 3795 37564
rect 3851 37562 3857 37564
rect 3611 37510 3613 37562
rect 3793 37510 3795 37562
rect 3549 37508 3555 37510
rect 3611 37508 3635 37510
rect 3691 37508 3715 37510
rect 3771 37508 3795 37510
rect 3851 37508 3857 37510
rect 3549 37499 3857 37508
rect 3896 37448 3924 37810
rect 3974 37768 4030 37777
rect 3974 37703 4030 37712
rect 3804 37420 3924 37448
rect 3804 36922 3832 37420
rect 3988 37262 4016 37703
rect 4080 37330 4108 38286
rect 4160 37800 4212 37806
rect 4160 37742 4212 37748
rect 4068 37324 4120 37330
rect 4068 37266 4120 37272
rect 3976 37256 4028 37262
rect 3976 37198 4028 37204
rect 3884 37120 3936 37126
rect 3884 37062 3936 37068
rect 3792 36916 3844 36922
rect 3792 36858 3844 36864
rect 3332 36780 3384 36786
rect 3332 36722 3384 36728
rect 3424 36712 3476 36718
rect 3424 36654 3476 36660
rect 3332 36032 3384 36038
rect 3332 35974 3384 35980
rect 3238 34912 3294 34921
rect 3238 34847 3294 34856
rect 3344 34082 3372 35974
rect 3436 35329 3464 36654
rect 3549 36476 3857 36485
rect 3549 36474 3555 36476
rect 3611 36474 3635 36476
rect 3691 36474 3715 36476
rect 3771 36474 3795 36476
rect 3851 36474 3857 36476
rect 3611 36422 3613 36474
rect 3793 36422 3795 36474
rect 3549 36420 3555 36422
rect 3611 36420 3635 36422
rect 3691 36420 3715 36422
rect 3771 36420 3795 36422
rect 3851 36420 3857 36422
rect 3549 36411 3857 36420
rect 3516 35760 3568 35766
rect 3516 35702 3568 35708
rect 3528 35601 3556 35702
rect 3514 35592 3570 35601
rect 3514 35527 3570 35536
rect 3549 35388 3857 35397
rect 3549 35386 3555 35388
rect 3611 35386 3635 35388
rect 3691 35386 3715 35388
rect 3771 35386 3795 35388
rect 3851 35386 3857 35388
rect 3611 35334 3613 35386
rect 3793 35334 3795 35386
rect 3549 35332 3555 35334
rect 3611 35332 3635 35334
rect 3691 35332 3715 35334
rect 3771 35332 3795 35334
rect 3851 35332 3857 35334
rect 3422 35320 3478 35329
rect 3549 35323 3857 35332
rect 3422 35255 3478 35264
rect 3516 35284 3568 35290
rect 3896 35272 3924 37062
rect 4068 36712 4120 36718
rect 4172 36700 4200 37742
rect 4252 37460 4304 37466
rect 4252 37402 4304 37408
rect 4120 36672 4200 36700
rect 4068 36654 4120 36660
rect 4068 36100 4120 36106
rect 4068 36042 4120 36048
rect 3976 35488 4028 35494
rect 3976 35430 4028 35436
rect 3516 35226 3568 35232
rect 3804 35244 3924 35272
rect 3528 35193 3556 35226
rect 3514 35184 3570 35193
rect 3514 35119 3570 35128
rect 3514 35048 3570 35057
rect 3514 34983 3570 34992
rect 3608 35012 3660 35018
rect 3528 34950 3556 34983
rect 3608 34954 3660 34960
rect 3516 34944 3568 34950
rect 3516 34886 3568 34892
rect 3620 34762 3648 34954
rect 3252 34054 3372 34082
rect 3436 34734 3648 34762
rect 3146 33824 3202 33833
rect 3146 33759 3202 33768
rect 3252 33674 3280 34054
rect 3332 33992 3384 33998
rect 3332 33934 3384 33940
rect 3160 33646 3280 33674
rect 3160 32774 3188 33646
rect 3240 33516 3292 33522
rect 3240 33458 3292 33464
rect 3252 33114 3280 33458
rect 3240 33108 3292 33114
rect 3240 33050 3292 33056
rect 3344 33017 3372 33934
rect 3330 33008 3386 33017
rect 3330 32943 3386 32952
rect 3238 32872 3294 32881
rect 3238 32807 3294 32816
rect 3148 32768 3200 32774
rect 3148 32710 3200 32716
rect 3148 32564 3200 32570
rect 3148 32506 3200 32512
rect 3160 31634 3188 32506
rect 3252 32502 3280 32807
rect 3240 32496 3292 32502
rect 3240 32438 3292 32444
rect 3332 32360 3384 32366
rect 3332 32302 3384 32308
rect 3344 32026 3372 32302
rect 3332 32020 3384 32026
rect 3332 31962 3384 31968
rect 3160 31606 3372 31634
rect 3056 30048 3108 30054
rect 3056 29990 3108 29996
rect 2964 29640 3016 29646
rect 2964 29582 3016 29588
rect 3160 29306 3188 31606
rect 3238 31512 3294 31521
rect 3344 31482 3372 31606
rect 3238 31447 3294 31456
rect 3332 31476 3384 31482
rect 3252 30802 3280 31447
rect 3332 31418 3384 31424
rect 3436 30870 3464 34734
rect 3804 34649 3832 35244
rect 3884 35012 3936 35018
rect 3884 34954 3936 34960
rect 3790 34640 3846 34649
rect 3790 34575 3846 34584
rect 3549 34300 3857 34309
rect 3549 34298 3555 34300
rect 3611 34298 3635 34300
rect 3691 34298 3715 34300
rect 3771 34298 3795 34300
rect 3851 34298 3857 34300
rect 3611 34246 3613 34298
rect 3793 34246 3795 34298
rect 3549 34244 3555 34246
rect 3611 34244 3635 34246
rect 3691 34244 3715 34246
rect 3771 34244 3795 34246
rect 3851 34244 3857 34246
rect 3549 34235 3857 34244
rect 3896 33697 3924 34954
rect 3988 34066 4016 35430
rect 4080 35193 4108 36042
rect 4172 35290 4200 36672
rect 4264 35873 4292 37402
rect 4356 36938 4384 40598
rect 4528 38752 4580 38758
rect 4448 38712 4528 38740
rect 4448 37398 4476 38712
rect 4528 38694 4580 38700
rect 4528 37664 4580 37670
rect 4528 37606 4580 37612
rect 4540 37398 4568 37606
rect 4436 37392 4488 37398
rect 4436 37334 4488 37340
rect 4528 37392 4580 37398
rect 4528 37334 4580 37340
rect 4356 36910 4476 36938
rect 4344 36780 4396 36786
rect 4344 36722 4396 36728
rect 4250 35864 4306 35873
rect 4250 35799 4306 35808
rect 4356 35698 4384 36722
rect 4252 35692 4304 35698
rect 4252 35634 4304 35640
rect 4344 35692 4396 35698
rect 4344 35634 4396 35640
rect 4160 35284 4212 35290
rect 4160 35226 4212 35232
rect 4066 35184 4122 35193
rect 4066 35119 4122 35128
rect 4068 35012 4120 35018
rect 4068 34954 4120 34960
rect 4080 34105 4108 34954
rect 4264 34649 4292 35634
rect 4344 35216 4396 35222
rect 4344 35158 4396 35164
rect 4250 34640 4306 34649
rect 4250 34575 4306 34584
rect 4252 34400 4304 34406
rect 4252 34342 4304 34348
rect 4264 34202 4292 34342
rect 4252 34196 4304 34202
rect 4252 34138 4304 34144
rect 4066 34096 4122 34105
rect 3976 34060 4028 34066
rect 4356 34082 4384 35158
rect 4066 34031 4122 34040
rect 4264 34054 4384 34082
rect 3976 34002 4028 34008
rect 3882 33688 3938 33697
rect 3882 33623 3938 33632
rect 3884 33584 3936 33590
rect 3884 33526 3936 33532
rect 3549 33212 3857 33221
rect 3549 33210 3555 33212
rect 3611 33210 3635 33212
rect 3691 33210 3715 33212
rect 3771 33210 3795 33212
rect 3851 33210 3857 33212
rect 3611 33158 3613 33210
rect 3793 33158 3795 33210
rect 3549 33156 3555 33158
rect 3611 33156 3635 33158
rect 3691 33156 3715 33158
rect 3771 33156 3795 33158
rect 3851 33156 3857 33158
rect 3549 33147 3857 33156
rect 3790 33008 3846 33017
rect 3790 32943 3846 32952
rect 3804 32842 3832 32943
rect 3792 32836 3844 32842
rect 3792 32778 3844 32784
rect 3896 32502 3924 33526
rect 4264 33454 4292 34054
rect 4344 33924 4396 33930
rect 4344 33866 4396 33872
rect 3976 33448 4028 33454
rect 3976 33390 4028 33396
rect 4252 33448 4304 33454
rect 4252 33390 4304 33396
rect 3884 32496 3936 32502
rect 3884 32438 3936 32444
rect 3549 32124 3857 32133
rect 3549 32122 3555 32124
rect 3611 32122 3635 32124
rect 3691 32122 3715 32124
rect 3771 32122 3795 32124
rect 3851 32122 3857 32124
rect 3611 32070 3613 32122
rect 3793 32070 3795 32122
rect 3549 32068 3555 32070
rect 3611 32068 3635 32070
rect 3691 32068 3715 32070
rect 3771 32068 3795 32070
rect 3851 32068 3857 32070
rect 3549 32059 3857 32068
rect 3896 32008 3924 32438
rect 3712 31980 3924 32008
rect 3712 31521 3740 31980
rect 3792 31816 3844 31822
rect 3792 31758 3844 31764
rect 3698 31512 3754 31521
rect 3698 31447 3754 31456
rect 3804 31385 3832 31758
rect 3790 31376 3846 31385
rect 3790 31311 3846 31320
rect 3884 31136 3936 31142
rect 3884 31078 3936 31084
rect 3549 31036 3857 31045
rect 3549 31034 3555 31036
rect 3611 31034 3635 31036
rect 3691 31034 3715 31036
rect 3771 31034 3795 31036
rect 3851 31034 3857 31036
rect 3611 30982 3613 31034
rect 3793 30982 3795 31034
rect 3549 30980 3555 30982
rect 3611 30980 3635 30982
rect 3691 30980 3715 30982
rect 3771 30980 3795 30982
rect 3851 30980 3857 30982
rect 3549 30971 3857 30980
rect 3896 30870 3924 31078
rect 3424 30864 3476 30870
rect 3424 30806 3476 30812
rect 3884 30864 3936 30870
rect 3884 30806 3936 30812
rect 3240 30796 3292 30802
rect 3240 30738 3292 30744
rect 3424 30728 3476 30734
rect 3424 30670 3476 30676
rect 3792 30728 3844 30734
rect 3988 30716 4016 33390
rect 4068 32768 4120 32774
rect 4068 32710 4120 32716
rect 4080 32473 4108 32710
rect 4160 32564 4212 32570
rect 4160 32506 4212 32512
rect 4066 32464 4122 32473
rect 4066 32399 4122 32408
rect 4068 31816 4120 31822
rect 4066 31784 4068 31793
rect 4120 31784 4122 31793
rect 4066 31719 4122 31728
rect 4172 31686 4200 32506
rect 4252 32292 4304 32298
rect 4252 32234 4304 32240
rect 4264 32065 4292 32234
rect 4250 32056 4306 32065
rect 4250 31991 4306 32000
rect 4160 31680 4212 31686
rect 4160 31622 4212 31628
rect 4252 31680 4304 31686
rect 4252 31622 4304 31628
rect 4068 31136 4120 31142
rect 4068 31078 4120 31084
rect 4080 30841 4108 31078
rect 4066 30832 4122 30841
rect 4172 30802 4200 31622
rect 4264 31521 4292 31622
rect 4250 31512 4306 31521
rect 4250 31447 4306 31456
rect 4066 30767 4122 30776
rect 4160 30796 4212 30802
rect 4160 30738 4212 30744
rect 3844 30688 4016 30716
rect 3792 30670 3844 30676
rect 3240 30252 3292 30258
rect 3240 30194 3292 30200
rect 3252 29889 3280 30194
rect 3332 30048 3384 30054
rect 3332 29990 3384 29996
rect 3238 29880 3294 29889
rect 3238 29815 3294 29824
rect 3240 29504 3292 29510
rect 3344 29492 3372 29990
rect 3292 29464 3372 29492
rect 3240 29446 3292 29452
rect 3148 29300 3200 29306
rect 3148 29242 3200 29248
rect 2872 29232 2924 29238
rect 2872 29174 2924 29180
rect 3054 29200 3110 29209
rect 2964 29164 3016 29170
rect 3054 29135 3110 29144
rect 2964 29106 3016 29112
rect 2688 28960 2740 28966
rect 2688 28902 2740 28908
rect 2594 28248 2650 28257
rect 2594 28183 2650 28192
rect 2504 28144 2556 28150
rect 2504 28086 2556 28092
rect 2700 28014 2728 28902
rect 2872 28552 2924 28558
rect 2792 28512 2872 28540
rect 2056 26710 2176 26738
rect 2240 27934 2360 27962
rect 2688 28008 2740 28014
rect 2688 27950 2740 27956
rect 2056 26489 2084 26710
rect 2042 26480 2098 26489
rect 2042 26415 2098 26424
rect 2044 26376 2096 26382
rect 2044 26318 2096 26324
rect 1950 26208 2006 26217
rect 1950 26143 2006 26152
rect 1872 25894 1992 25922
rect 2056 25906 2084 26318
rect 2134 26072 2190 26081
rect 2134 26007 2190 26016
rect 1860 24880 1912 24886
rect 1860 24822 1912 24828
rect 1872 24721 1900 24822
rect 1858 24712 1914 24721
rect 1858 24647 1914 24656
rect 1768 24404 1820 24410
rect 1768 24346 1820 24352
rect 1582 24032 1638 24041
rect 1582 23967 1638 23976
rect 1400 23724 1452 23730
rect 1400 23666 1452 23672
rect 1768 23724 1820 23730
rect 1964 23712 1992 25894
rect 2044 25900 2096 25906
rect 2044 25842 2096 25848
rect 1820 23684 1992 23712
rect 1768 23666 1820 23672
rect 1412 23610 1440 23666
rect 1412 23582 1532 23610
rect 1398 23488 1454 23497
rect 1398 23423 1454 23432
rect 1124 23316 1176 23322
rect 1124 23258 1176 23264
rect 1136 22681 1164 23258
rect 1412 23118 1440 23423
rect 1504 23186 1532 23582
rect 1492 23180 1544 23186
rect 1492 23122 1544 23128
rect 1400 23112 1452 23118
rect 1400 23054 1452 23060
rect 1582 23080 1638 23089
rect 1308 23044 1360 23050
rect 1582 23015 1638 23024
rect 1308 22986 1360 22992
rect 1320 22953 1348 22986
rect 1596 22982 1624 23015
rect 1584 22976 1636 22982
rect 1306 22944 1362 22953
rect 1584 22918 1636 22924
rect 1306 22879 1362 22888
rect 1674 22808 1730 22817
rect 1674 22743 1676 22752
rect 1728 22743 1730 22752
rect 1676 22714 1728 22720
rect 1122 22672 1178 22681
rect 1122 22607 1178 22616
rect 1122 22536 1178 22545
rect 1122 22471 1178 22480
rect 1032 18964 1084 18970
rect 1032 18906 1084 18912
rect 938 18592 994 18601
rect 938 18527 994 18536
rect 952 18358 980 18527
rect 940 18352 992 18358
rect 940 18294 992 18300
rect 938 14784 994 14793
rect 938 14719 994 14728
rect 952 14006 980 14719
rect 940 14000 992 14006
rect 940 13942 992 13948
rect 938 13832 994 13841
rect 938 13767 994 13776
rect 952 13530 980 13767
rect 940 13524 992 13530
rect 940 13466 992 13472
rect 938 13016 994 13025
rect 938 12951 994 12960
rect 952 11286 980 12951
rect 1030 11520 1086 11529
rect 1030 11455 1086 11464
rect 940 11280 992 11286
rect 940 11222 992 11228
rect 940 11076 992 11082
rect 940 11018 992 11024
rect 952 3641 980 11018
rect 1044 10305 1072 11455
rect 1030 10296 1086 10305
rect 1030 10231 1086 10240
rect 1030 7304 1086 7313
rect 1030 7239 1086 7248
rect 938 3632 994 3641
rect 938 3567 994 3576
rect 1044 3466 1072 7239
rect 1032 3460 1084 3466
rect 1032 3402 1084 3408
rect 1136 2774 1164 22471
rect 1398 22128 1454 22137
rect 1398 22063 1400 22072
rect 1452 22063 1454 22072
rect 1400 22034 1452 22040
rect 1216 22024 1268 22030
rect 1216 21966 1268 21972
rect 1676 22024 1728 22030
rect 1676 21966 1728 21972
rect 1228 21865 1256 21966
rect 1214 21856 1270 21865
rect 1214 21791 1270 21800
rect 1688 21729 1716 21966
rect 1674 21720 1730 21729
rect 1674 21655 1730 21664
rect 1676 21548 1728 21554
rect 1780 21536 1808 23666
rect 1860 23112 1912 23118
rect 1860 23054 1912 23060
rect 1728 21508 1808 21536
rect 1676 21490 1728 21496
rect 1216 21480 1268 21486
rect 1216 21422 1268 21428
rect 1228 19922 1256 21422
rect 1490 21312 1546 21321
rect 1490 21247 1546 21256
rect 1308 20868 1360 20874
rect 1308 20810 1360 20816
rect 1320 20777 1348 20810
rect 1306 20768 1362 20777
rect 1306 20703 1362 20712
rect 1320 20602 1440 20618
rect 1308 20596 1440 20602
rect 1360 20590 1440 20596
rect 1308 20538 1360 20544
rect 1216 19916 1268 19922
rect 1216 19858 1268 19864
rect 1306 17368 1362 17377
rect 1306 17303 1362 17312
rect 1216 16992 1268 16998
rect 1216 16934 1268 16940
rect 1228 14414 1256 16934
rect 1320 16250 1348 17303
rect 1308 16244 1360 16250
rect 1308 16186 1360 16192
rect 1412 15201 1440 20590
rect 1504 20466 1532 21247
rect 1492 20460 1544 20466
rect 1492 20402 1544 20408
rect 1582 20360 1638 20369
rect 1582 20295 1584 20304
rect 1636 20295 1638 20304
rect 1584 20266 1636 20272
rect 1490 20224 1546 20233
rect 1490 20159 1546 20168
rect 1504 18834 1532 20159
rect 1688 19700 1716 21490
rect 1766 21448 1822 21457
rect 1766 21383 1822 21392
rect 1780 20058 1808 21383
rect 1768 20052 1820 20058
rect 1768 19994 1820 20000
rect 1872 19938 1900 23054
rect 1952 22636 2004 22642
rect 1952 22578 2004 22584
rect 1964 22166 1992 22578
rect 1952 22160 2004 22166
rect 1952 22102 2004 22108
rect 2056 21865 2084 25842
rect 2148 25498 2176 26007
rect 2240 25974 2268 27934
rect 2320 27872 2372 27878
rect 2320 27814 2372 27820
rect 2332 27010 2360 27814
rect 2412 27464 2464 27470
rect 2412 27406 2464 27412
rect 2424 27130 2452 27406
rect 2504 27396 2556 27402
rect 2504 27338 2556 27344
rect 2516 27130 2544 27338
rect 2596 27328 2648 27334
rect 2596 27270 2648 27276
rect 2608 27130 2636 27270
rect 2686 27160 2742 27169
rect 2412 27124 2464 27130
rect 2412 27066 2464 27072
rect 2504 27124 2556 27130
rect 2504 27066 2556 27072
rect 2596 27124 2648 27130
rect 2686 27095 2688 27104
rect 2596 27066 2648 27072
rect 2740 27095 2742 27104
rect 2688 27066 2740 27072
rect 2332 26994 2728 27010
rect 2332 26988 2740 26994
rect 2332 26982 2688 26988
rect 2688 26930 2740 26936
rect 2502 26888 2558 26897
rect 2792 26874 2820 28512
rect 2872 28494 2924 28500
rect 2976 28121 3004 29106
rect 2962 28112 3018 28121
rect 2872 28076 2924 28082
rect 2962 28047 3018 28056
rect 2872 28018 2924 28024
rect 2884 27674 2912 28018
rect 2872 27668 2924 27674
rect 2872 27610 2924 27616
rect 2502 26823 2504 26832
rect 2556 26823 2558 26832
rect 2700 26846 2820 26874
rect 2504 26794 2556 26800
rect 2320 26784 2372 26790
rect 2320 26726 2372 26732
rect 2596 26784 2648 26790
rect 2596 26726 2648 26732
rect 2332 25974 2360 26726
rect 2504 26512 2556 26518
rect 2502 26480 2504 26489
rect 2556 26480 2558 26489
rect 2502 26415 2558 26424
rect 2412 26240 2464 26246
rect 2412 26182 2464 26188
rect 2228 25968 2280 25974
rect 2228 25910 2280 25916
rect 2320 25968 2372 25974
rect 2320 25910 2372 25916
rect 2240 25537 2268 25910
rect 2226 25528 2282 25537
rect 2136 25492 2188 25498
rect 2226 25463 2282 25472
rect 2136 25434 2188 25440
rect 2240 25362 2268 25463
rect 2228 25356 2280 25362
rect 2228 25298 2280 25304
rect 2134 25120 2190 25129
rect 2134 25055 2190 25064
rect 2148 24886 2176 25055
rect 2136 24880 2188 24886
rect 2136 24822 2188 24828
rect 2042 21856 2098 21865
rect 2042 21791 2098 21800
rect 1950 21312 2006 21321
rect 1950 21247 2006 21256
rect 1964 20942 1992 21247
rect 2044 21140 2096 21146
rect 2044 21082 2096 21088
rect 1952 20936 2004 20942
rect 1952 20878 2004 20884
rect 1780 19910 1900 19938
rect 1780 19854 1808 19910
rect 1768 19848 1820 19854
rect 1768 19790 1820 19796
rect 1860 19780 1912 19786
rect 1860 19722 1912 19728
rect 1688 19672 1808 19700
rect 1674 18864 1730 18873
rect 1492 18828 1544 18834
rect 1674 18799 1676 18808
rect 1492 18770 1544 18776
rect 1728 18799 1730 18808
rect 1676 18770 1728 18776
rect 1674 18592 1730 18601
rect 1674 18527 1730 18536
rect 1584 18080 1636 18086
rect 1490 18048 1546 18057
rect 1584 18022 1636 18028
rect 1490 17983 1546 17992
rect 1504 17762 1532 17983
rect 1596 17921 1624 18022
rect 1582 17912 1638 17921
rect 1582 17847 1638 17856
rect 1504 17734 1624 17762
rect 1596 17270 1624 17734
rect 1688 17678 1716 18527
rect 1780 18204 1808 19672
rect 1872 18329 1900 19722
rect 1964 19689 1992 20878
rect 2056 19990 2084 21082
rect 2148 20806 2176 24822
rect 2332 24596 2360 25910
rect 2424 24750 2452 26182
rect 2504 25288 2556 25294
rect 2504 25230 2556 25236
rect 2516 24993 2544 25230
rect 2502 24984 2558 24993
rect 2502 24919 2558 24928
rect 2504 24812 2556 24818
rect 2504 24754 2556 24760
rect 2412 24744 2464 24750
rect 2412 24686 2464 24692
rect 2332 24568 2452 24596
rect 2320 23520 2372 23526
rect 2320 23462 2372 23468
rect 2226 22672 2282 22681
rect 2226 22607 2282 22616
rect 2240 21078 2268 22607
rect 2332 22574 2360 23462
rect 2424 22817 2452 24568
rect 2516 24410 2544 24754
rect 2504 24404 2556 24410
rect 2504 24346 2556 24352
rect 2608 24206 2636 26726
rect 2596 24200 2648 24206
rect 2596 24142 2648 24148
rect 2504 22976 2556 22982
rect 2504 22918 2556 22924
rect 2410 22808 2466 22817
rect 2410 22743 2466 22752
rect 2516 22710 2544 22918
rect 2504 22704 2556 22710
rect 2504 22646 2556 22652
rect 2412 22636 2464 22642
rect 2412 22578 2464 22584
rect 2320 22568 2372 22574
rect 2320 22510 2372 22516
rect 2318 22400 2374 22409
rect 2318 22335 2374 22344
rect 2332 22030 2360 22335
rect 2424 22166 2452 22578
rect 2608 22216 2636 24142
rect 2700 23118 2728 26846
rect 2780 26240 2832 26246
rect 2780 26182 2832 26188
rect 2792 25401 2820 26182
rect 2778 25392 2834 25401
rect 2778 25327 2834 25336
rect 2884 24954 2912 27610
rect 2962 27024 3018 27033
rect 2962 26959 2964 26968
rect 3016 26959 3018 26968
rect 2964 26930 3016 26936
rect 2962 26752 3018 26761
rect 2962 26687 3018 26696
rect 2976 26586 3004 26687
rect 2964 26580 3016 26586
rect 2964 26522 3016 26528
rect 3068 26466 3096 29135
rect 3148 29028 3200 29034
rect 3148 28970 3200 28976
rect 3160 28626 3188 28970
rect 3148 28620 3200 28626
rect 3148 28562 3200 28568
rect 3146 28112 3202 28121
rect 3146 28047 3202 28056
rect 3160 27606 3188 28047
rect 3148 27600 3200 27606
rect 3148 27542 3200 27548
rect 3148 27328 3200 27334
rect 3146 27296 3148 27305
rect 3200 27296 3202 27305
rect 3146 27231 3202 27240
rect 3148 26988 3200 26994
rect 3148 26930 3200 26936
rect 3160 26586 3188 26930
rect 3148 26580 3200 26586
rect 3148 26522 3200 26528
rect 3252 26466 3280 29446
rect 3332 28960 3384 28966
rect 3332 28902 3384 28908
rect 3344 28762 3372 28902
rect 3332 28756 3384 28762
rect 3332 28698 3384 28704
rect 3332 28212 3384 28218
rect 3332 28154 3384 28160
rect 3344 27334 3372 28154
rect 3332 27328 3384 27334
rect 3332 27270 3384 27276
rect 3332 27124 3384 27130
rect 3332 27066 3384 27072
rect 3344 26625 3372 27066
rect 3330 26616 3386 26625
rect 3330 26551 3386 26560
rect 3436 26518 3464 30670
rect 4252 30592 4304 30598
rect 4252 30534 4304 30540
rect 3976 30388 4028 30394
rect 3976 30330 4028 30336
rect 3884 30320 3936 30326
rect 3606 30288 3662 30297
rect 3606 30223 3608 30232
rect 3660 30223 3662 30232
rect 3882 30288 3884 30297
rect 3936 30288 3938 30297
rect 3882 30223 3938 30232
rect 3608 30194 3660 30200
rect 3549 29948 3857 29957
rect 3549 29946 3555 29948
rect 3611 29946 3635 29948
rect 3691 29946 3715 29948
rect 3771 29946 3795 29948
rect 3851 29946 3857 29948
rect 3611 29894 3613 29946
rect 3793 29894 3795 29946
rect 3549 29892 3555 29894
rect 3611 29892 3635 29894
rect 3691 29892 3715 29894
rect 3771 29892 3795 29894
rect 3851 29892 3857 29894
rect 3549 29883 3857 29892
rect 3516 29640 3568 29646
rect 3516 29582 3568 29588
rect 3528 29481 3556 29582
rect 3514 29472 3570 29481
rect 3514 29407 3570 29416
rect 3549 28860 3857 28869
rect 3549 28858 3555 28860
rect 3611 28858 3635 28860
rect 3691 28858 3715 28860
rect 3771 28858 3795 28860
rect 3851 28858 3857 28860
rect 3611 28806 3613 28858
rect 3793 28806 3795 28858
rect 3549 28804 3555 28806
rect 3611 28804 3635 28806
rect 3691 28804 3715 28806
rect 3771 28804 3795 28806
rect 3851 28804 3857 28806
rect 3549 28795 3857 28804
rect 3792 28756 3844 28762
rect 3792 28698 3844 28704
rect 3804 28665 3832 28698
rect 3790 28656 3846 28665
rect 3790 28591 3846 28600
rect 3700 28416 3752 28422
rect 3606 28384 3662 28393
rect 3700 28358 3752 28364
rect 3606 28319 3662 28328
rect 3620 28082 3648 28319
rect 3712 28082 3740 28358
rect 3896 28150 3924 30223
rect 3988 28422 4016 30330
rect 4160 30252 4212 30258
rect 4160 30194 4212 30200
rect 4172 29850 4200 30194
rect 4264 30025 4292 30534
rect 4250 30016 4306 30025
rect 4250 29951 4306 29960
rect 4160 29844 4212 29850
rect 4160 29786 4212 29792
rect 4160 29572 4212 29578
rect 4160 29514 4212 29520
rect 4068 29028 4120 29034
rect 4068 28970 4120 28976
rect 3976 28416 4028 28422
rect 3976 28358 4028 28364
rect 3884 28144 3936 28150
rect 3936 28104 4016 28132
rect 3884 28086 3936 28092
rect 3608 28076 3660 28082
rect 3608 28018 3660 28024
rect 3700 28076 3752 28082
rect 3700 28018 3752 28024
rect 3884 27872 3936 27878
rect 3884 27814 3936 27820
rect 3549 27772 3857 27781
rect 3549 27770 3555 27772
rect 3611 27770 3635 27772
rect 3691 27770 3715 27772
rect 3771 27770 3795 27772
rect 3851 27770 3857 27772
rect 3611 27718 3613 27770
rect 3793 27718 3795 27770
rect 3549 27716 3555 27718
rect 3611 27716 3635 27718
rect 3691 27716 3715 27718
rect 3771 27716 3795 27718
rect 3851 27716 3857 27718
rect 3549 27707 3857 27716
rect 3700 27396 3752 27402
rect 3700 27338 3752 27344
rect 3712 27130 3740 27338
rect 3700 27124 3752 27130
rect 3896 27112 3924 27814
rect 3988 27282 4016 28104
rect 4080 28082 4108 28970
rect 4172 28665 4200 29514
rect 4158 28656 4214 28665
rect 4158 28591 4214 28600
rect 4252 28416 4304 28422
rect 4252 28358 4304 28364
rect 4068 28076 4120 28082
rect 4264 28064 4292 28358
rect 4068 28018 4120 28024
rect 4172 28036 4292 28064
rect 4172 27962 4200 28036
rect 4080 27934 4200 27962
rect 4250 27976 4306 27985
rect 4080 27402 4108 27934
rect 4250 27911 4306 27920
rect 4264 27606 4292 27911
rect 4252 27600 4304 27606
rect 4252 27542 4304 27548
rect 4160 27464 4212 27470
rect 4160 27406 4212 27412
rect 4068 27396 4120 27402
rect 4068 27338 4120 27344
rect 4066 27296 4122 27305
rect 3988 27254 4066 27282
rect 4066 27231 4122 27240
rect 4066 27160 4122 27169
rect 3976 27124 4028 27130
rect 3896 27084 3976 27112
rect 3700 27066 3752 27072
rect 4066 27095 4122 27104
rect 3976 27066 4028 27072
rect 3792 27056 3844 27062
rect 3844 27004 3924 27010
rect 3792 26998 3924 27004
rect 3804 26982 3924 26998
rect 3549 26684 3857 26693
rect 3549 26682 3555 26684
rect 3611 26682 3635 26684
rect 3691 26682 3715 26684
rect 3771 26682 3795 26684
rect 3851 26682 3857 26684
rect 3611 26630 3613 26682
rect 3793 26630 3795 26682
rect 3549 26628 3555 26630
rect 3611 26628 3635 26630
rect 3691 26628 3715 26630
rect 3771 26628 3795 26630
rect 3851 26628 3857 26630
rect 3549 26619 3857 26628
rect 3332 26512 3384 26518
rect 2976 26438 3096 26466
rect 3160 26438 3280 26466
rect 3330 26480 3332 26489
rect 3424 26512 3476 26518
rect 3384 26480 3386 26489
rect 2872 24948 2924 24954
rect 2872 24890 2924 24896
rect 2780 23656 2832 23662
rect 2780 23598 2832 23604
rect 2792 23225 2820 23598
rect 2976 23576 3004 26438
rect 3056 26376 3108 26382
rect 3056 26318 3108 26324
rect 3068 25673 3096 26318
rect 3054 25664 3110 25673
rect 3054 25599 3110 25608
rect 2976 23548 3096 23576
rect 2962 23488 3018 23497
rect 2884 23446 2962 23474
rect 2778 23216 2834 23225
rect 2778 23151 2834 23160
rect 2688 23112 2740 23118
rect 2688 23054 2740 23060
rect 2884 22778 2912 23446
rect 2962 23423 3018 23432
rect 3068 22778 3096 23548
rect 2872 22772 2924 22778
rect 2872 22714 2924 22720
rect 3056 22772 3108 22778
rect 3056 22714 3108 22720
rect 2780 22704 2832 22710
rect 3068 22658 3096 22714
rect 2780 22646 2832 22652
rect 2516 22188 2636 22216
rect 2412 22160 2464 22166
rect 2412 22102 2464 22108
rect 2320 22024 2372 22030
rect 2320 21966 2372 21972
rect 2516 21468 2544 22188
rect 2594 22128 2650 22137
rect 2594 22063 2650 22072
rect 2332 21440 2544 21468
rect 2228 21072 2280 21078
rect 2228 21014 2280 21020
rect 2136 20800 2188 20806
rect 2332 20754 2360 21440
rect 2608 21400 2636 22063
rect 2688 21888 2740 21894
rect 2688 21830 2740 21836
rect 2516 21372 2636 21400
rect 2412 21344 2464 21350
rect 2516 21332 2544 21372
rect 2464 21304 2544 21332
rect 2412 21286 2464 21292
rect 2410 21176 2466 21185
rect 2410 21111 2466 21120
rect 2136 20742 2188 20748
rect 2240 20726 2360 20754
rect 2044 19984 2096 19990
rect 2044 19926 2096 19932
rect 1950 19680 2006 19689
rect 1950 19615 2006 19624
rect 1964 19446 1992 19615
rect 1952 19440 2004 19446
rect 1952 19382 2004 19388
rect 2240 18766 2268 20726
rect 2318 20632 2374 20641
rect 2318 20567 2320 20576
rect 2372 20567 2374 20576
rect 2320 20538 2372 20544
rect 2318 19952 2374 19961
rect 2318 19887 2320 19896
rect 2372 19887 2374 19896
rect 2320 19858 2372 19864
rect 2318 19816 2374 19825
rect 2318 19751 2320 19760
rect 2372 19751 2374 19760
rect 2320 19722 2372 19728
rect 2424 19281 2452 21111
rect 2516 20942 2544 21304
rect 2700 21185 2728 21830
rect 2686 21176 2742 21185
rect 2686 21111 2742 21120
rect 2504 20936 2556 20942
rect 2504 20878 2556 20884
rect 2504 20800 2556 20806
rect 2504 20742 2556 20748
rect 2688 20800 2740 20806
rect 2688 20742 2740 20748
rect 2516 20534 2544 20742
rect 2594 20632 2650 20641
rect 2594 20567 2650 20576
rect 2504 20528 2556 20534
rect 2504 20470 2556 20476
rect 2504 20392 2556 20398
rect 2504 20334 2556 20340
rect 2608 20346 2636 20567
rect 2700 20466 2728 20742
rect 2688 20460 2740 20466
rect 2688 20402 2740 20408
rect 2516 19514 2544 20334
rect 2608 20318 2728 20346
rect 2594 19816 2650 19825
rect 2594 19751 2650 19760
rect 2504 19508 2556 19514
rect 2504 19450 2556 19456
rect 2608 19378 2636 19751
rect 2700 19378 2728 20318
rect 2792 20058 2820 22646
rect 2884 22630 3096 22658
rect 2884 21894 2912 22630
rect 2964 22568 3016 22574
rect 2964 22510 3016 22516
rect 2872 21888 2924 21894
rect 2872 21830 2924 21836
rect 2976 20992 3004 22510
rect 3056 21548 3108 21554
rect 3056 21490 3108 21496
rect 3068 21321 3096 21490
rect 3054 21312 3110 21321
rect 3054 21247 3110 21256
rect 3160 21146 3188 26438
rect 3424 26454 3476 26460
rect 3330 26415 3386 26424
rect 3332 26376 3384 26382
rect 3332 26318 3384 26324
rect 3514 26344 3570 26353
rect 3344 26217 3372 26318
rect 3514 26279 3570 26288
rect 3330 26208 3386 26217
rect 3330 26143 3386 26152
rect 3332 25968 3384 25974
rect 3332 25910 3384 25916
rect 3344 25498 3372 25910
rect 3528 25906 3556 26279
rect 3896 26042 3924 26982
rect 3976 26988 4028 26994
rect 3976 26930 4028 26936
rect 3884 26036 3936 26042
rect 3884 25978 3936 25984
rect 3988 25974 4016 26930
rect 4080 26926 4108 27095
rect 4172 27062 4200 27406
rect 4356 27169 4384 33866
rect 4448 31822 4476 36910
rect 4632 35834 4660 41386
rect 4712 41200 4764 41206
rect 4712 41142 4764 41148
rect 4724 39914 4752 41142
rect 4712 39908 4764 39914
rect 4712 39850 4764 39856
rect 4712 37120 4764 37126
rect 4712 37062 4764 37068
rect 4620 35828 4672 35834
rect 4620 35770 4672 35776
rect 4528 35624 4580 35630
rect 4580 35584 4660 35612
rect 4528 35566 4580 35572
rect 4528 35148 4580 35154
rect 4528 35090 4580 35096
rect 4540 34950 4568 35090
rect 4528 34944 4580 34950
rect 4528 34886 4580 34892
rect 4540 34678 4568 34886
rect 4528 34672 4580 34678
rect 4632 34649 4660 35584
rect 4528 34614 4580 34620
rect 4618 34640 4674 34649
rect 4618 34575 4674 34584
rect 4620 34400 4672 34406
rect 4620 34342 4672 34348
rect 4528 34128 4580 34134
rect 4528 34070 4580 34076
rect 4540 33266 4568 34070
rect 4632 33561 4660 34342
rect 4618 33552 4674 33561
rect 4618 33487 4674 33496
rect 4540 33238 4660 33266
rect 4436 31816 4488 31822
rect 4436 31758 4488 31764
rect 4528 31816 4580 31822
rect 4528 31758 4580 31764
rect 4436 31272 4488 31278
rect 4436 31214 4488 31220
rect 4342 27160 4398 27169
rect 4252 27124 4304 27130
rect 4342 27095 4398 27104
rect 4252 27066 4304 27072
rect 4160 27056 4212 27062
rect 4160 26998 4212 27004
rect 4068 26920 4120 26926
rect 4068 26862 4120 26868
rect 4068 26784 4120 26790
rect 4068 26726 4120 26732
rect 3976 25968 4028 25974
rect 3976 25910 4028 25916
rect 3516 25900 3568 25906
rect 3516 25842 3568 25848
rect 3549 25596 3857 25605
rect 3549 25594 3555 25596
rect 3611 25594 3635 25596
rect 3691 25594 3715 25596
rect 3771 25594 3795 25596
rect 3851 25594 3857 25596
rect 3611 25542 3613 25594
rect 3793 25542 3795 25594
rect 3549 25540 3555 25542
rect 3611 25540 3635 25542
rect 3691 25540 3715 25542
rect 3771 25540 3795 25542
rect 3851 25540 3857 25542
rect 3549 25531 3857 25540
rect 3332 25492 3384 25498
rect 3332 25434 3384 25440
rect 3606 25392 3662 25401
rect 3606 25327 3662 25336
rect 3240 25288 3292 25294
rect 3240 25230 3292 25236
rect 3252 24585 3280 25230
rect 3332 24880 3384 24886
rect 3332 24822 3384 24828
rect 3238 24576 3294 24585
rect 3238 24511 3294 24520
rect 3240 24404 3292 24410
rect 3240 24346 3292 24352
rect 3252 23254 3280 24346
rect 3240 23248 3292 23254
rect 3240 23190 3292 23196
rect 3344 22166 3372 24822
rect 3424 24812 3476 24818
rect 3424 24754 3476 24760
rect 3436 23322 3464 24754
rect 3620 24614 3648 25327
rect 4080 25106 4108 26726
rect 3988 25078 4108 25106
rect 3884 24744 3936 24750
rect 3884 24686 3936 24692
rect 3608 24608 3660 24614
rect 3608 24550 3660 24556
rect 3549 24508 3857 24517
rect 3549 24506 3555 24508
rect 3611 24506 3635 24508
rect 3691 24506 3715 24508
rect 3771 24506 3795 24508
rect 3851 24506 3857 24508
rect 3611 24454 3613 24506
rect 3793 24454 3795 24506
rect 3549 24452 3555 24454
rect 3611 24452 3635 24454
rect 3691 24452 3715 24454
rect 3771 24452 3795 24454
rect 3851 24452 3857 24454
rect 3549 24443 3857 24452
rect 3896 23730 3924 24686
rect 3988 23769 4016 25078
rect 4068 24948 4120 24954
rect 4068 24890 4120 24896
rect 3974 23760 4030 23769
rect 3884 23724 3936 23730
rect 3974 23695 4030 23704
rect 3884 23666 3936 23672
rect 3549 23420 3857 23429
rect 3549 23418 3555 23420
rect 3611 23418 3635 23420
rect 3691 23418 3715 23420
rect 3771 23418 3795 23420
rect 3851 23418 3857 23420
rect 3611 23366 3613 23418
rect 3793 23366 3795 23418
rect 3549 23364 3555 23366
rect 3611 23364 3635 23366
rect 3691 23364 3715 23366
rect 3771 23364 3795 23366
rect 3851 23364 3857 23366
rect 3549 23355 3857 23364
rect 3424 23316 3476 23322
rect 3476 23276 3556 23304
rect 3424 23258 3476 23264
rect 3424 23112 3476 23118
rect 3424 23054 3476 23060
rect 3436 22642 3464 23054
rect 3528 22710 3556 23276
rect 3606 23216 3662 23225
rect 3606 23151 3662 23160
rect 3620 22710 3648 23151
rect 3792 23112 3844 23118
rect 3896 23100 3924 23666
rect 3976 23656 4028 23662
rect 3974 23624 3976 23633
rect 4028 23624 4030 23633
rect 3974 23559 4030 23568
rect 3974 23488 4030 23497
rect 3974 23423 4030 23432
rect 3988 23118 4016 23423
rect 3844 23072 3924 23100
rect 3976 23112 4028 23118
rect 3792 23054 3844 23060
rect 3976 23054 4028 23060
rect 4080 22982 4108 24890
rect 4264 24585 4292 27066
rect 4448 26874 4476 31214
rect 4540 28082 4568 31758
rect 4632 29782 4660 33238
rect 4724 33130 4752 37062
rect 4816 36378 4844 41550
rect 4908 41274 4936 42570
rect 4988 41472 5040 41478
rect 4988 41414 5040 41420
rect 4896 41268 4948 41274
rect 4896 41210 4948 41216
rect 4896 38344 4948 38350
rect 4896 38286 4948 38292
rect 5000 38298 5028 41414
rect 5092 41206 5120 42570
rect 5264 42220 5316 42226
rect 5264 42162 5316 42168
rect 5276 41818 5304 42162
rect 5354 42120 5410 42129
rect 5354 42055 5410 42064
rect 5264 41812 5316 41818
rect 5264 41754 5316 41760
rect 5368 41614 5396 42055
rect 5552 41834 5580 43250
rect 5644 42362 5672 43268
rect 6012 42906 6040 43608
rect 6148 43548 6456 43557
rect 6148 43546 6154 43548
rect 6210 43546 6234 43548
rect 6290 43546 6314 43548
rect 6370 43546 6394 43548
rect 6450 43546 6456 43548
rect 6210 43494 6212 43546
rect 6392 43494 6394 43546
rect 6148 43492 6154 43494
rect 6210 43492 6234 43494
rect 6290 43492 6314 43494
rect 6370 43492 6394 43494
rect 6450 43492 6456 43494
rect 6148 43483 6456 43492
rect 6000 42900 6052 42906
rect 6000 42842 6052 42848
rect 6564 42702 6592 43608
rect 6552 42696 6604 42702
rect 6552 42638 6604 42644
rect 5816 42628 5868 42634
rect 5816 42570 5868 42576
rect 5908 42628 5960 42634
rect 5908 42570 5960 42576
rect 5632 42356 5684 42362
rect 5632 42298 5684 42304
rect 5724 42152 5776 42158
rect 5724 42094 5776 42100
rect 5460 41806 5580 41834
rect 5736 41818 5764 42094
rect 5724 41812 5776 41818
rect 5172 41608 5224 41614
rect 5172 41550 5224 41556
rect 5356 41608 5408 41614
rect 5356 41550 5408 41556
rect 5080 41200 5132 41206
rect 5080 41142 5132 41148
rect 5080 39092 5132 39098
rect 5080 39034 5132 39040
rect 5092 38654 5120 39034
rect 5184 38758 5212 41550
rect 5264 41540 5316 41546
rect 5264 41482 5316 41488
rect 5276 41414 5304 41482
rect 5276 41386 5396 41414
rect 5264 41132 5316 41138
rect 5264 41074 5316 41080
rect 5276 40225 5304 41074
rect 5262 40216 5318 40225
rect 5262 40151 5318 40160
rect 5264 38820 5316 38826
rect 5264 38762 5316 38768
rect 5172 38752 5224 38758
rect 5172 38694 5224 38700
rect 5092 38626 5212 38654
rect 4908 37874 4936 38286
rect 5000 38270 5120 38298
rect 4988 38208 5040 38214
rect 4988 38150 5040 38156
rect 4896 37868 4948 37874
rect 4896 37810 4948 37816
rect 4908 37641 4936 37810
rect 4894 37632 4950 37641
rect 4894 37567 4950 37576
rect 5000 37330 5028 38150
rect 4988 37324 5040 37330
rect 4988 37266 5040 37272
rect 4896 37256 4948 37262
rect 4896 37198 4948 37204
rect 4908 36786 4936 37198
rect 4896 36780 4948 36786
rect 4896 36722 4948 36728
rect 4988 36576 5040 36582
rect 4988 36518 5040 36524
rect 4804 36372 4856 36378
rect 4804 36314 4856 36320
rect 4896 35624 4948 35630
rect 4894 35592 4896 35601
rect 4948 35592 4950 35601
rect 4894 35527 4950 35536
rect 4896 35488 4948 35494
rect 4896 35430 4948 35436
rect 4804 35284 4856 35290
rect 4804 35226 4856 35232
rect 4816 34678 4844 35226
rect 4908 34746 4936 35430
rect 4896 34740 4948 34746
rect 4896 34682 4948 34688
rect 4804 34672 4856 34678
rect 4804 34614 4856 34620
rect 4816 33930 4844 34614
rect 4896 34604 4948 34610
rect 4896 34546 4948 34552
rect 4804 33924 4856 33930
rect 4804 33866 4856 33872
rect 4804 33516 4856 33522
rect 4804 33458 4856 33464
rect 4816 33289 4844 33458
rect 4802 33280 4858 33289
rect 4802 33215 4858 33224
rect 4724 33102 4844 33130
rect 4908 33114 4936 34546
rect 5000 34542 5028 36518
rect 5092 34678 5120 38270
rect 5184 35306 5212 38626
rect 5276 38418 5304 38762
rect 5264 38412 5316 38418
rect 5264 38354 5316 38360
rect 5264 38208 5316 38214
rect 5264 38150 5316 38156
rect 5276 36553 5304 38150
rect 5368 37777 5396 41386
rect 5460 40730 5488 41806
rect 5724 41754 5776 41760
rect 5540 41744 5592 41750
rect 5540 41686 5592 41692
rect 5552 41154 5580 41686
rect 5552 41138 5764 41154
rect 5552 41132 5776 41138
rect 5552 41126 5724 41132
rect 5724 41074 5776 41080
rect 5448 40724 5500 40730
rect 5448 40666 5500 40672
rect 5632 40520 5684 40526
rect 5632 40462 5684 40468
rect 5540 39908 5592 39914
rect 5540 39850 5592 39856
rect 5552 38350 5580 39850
rect 5540 38344 5592 38350
rect 5540 38286 5592 38292
rect 5354 37768 5410 37777
rect 5354 37703 5410 37712
rect 5540 37664 5592 37670
rect 5446 37632 5502 37641
rect 5540 37606 5592 37612
rect 5446 37567 5502 37576
rect 5460 37466 5488 37567
rect 5448 37460 5500 37466
rect 5448 37402 5500 37408
rect 5448 37120 5500 37126
rect 5368 37080 5448 37108
rect 5262 36544 5318 36553
rect 5262 36479 5318 36488
rect 5262 35320 5318 35329
rect 5184 35278 5262 35306
rect 5368 35290 5396 37080
rect 5448 37062 5500 37068
rect 5448 36780 5500 36786
rect 5448 36722 5500 36728
rect 5460 36650 5488 36722
rect 5448 36644 5500 36650
rect 5448 36586 5500 36592
rect 5448 36236 5500 36242
rect 5448 36178 5500 36184
rect 5460 36145 5488 36178
rect 5446 36136 5502 36145
rect 5446 36071 5502 36080
rect 5552 35986 5580 37606
rect 5644 36922 5672 40462
rect 5828 39642 5856 42570
rect 5920 41818 5948 42570
rect 6000 42560 6052 42566
rect 6000 42502 6052 42508
rect 6012 42362 6040 42502
rect 6148 42460 6456 42469
rect 6148 42458 6154 42460
rect 6210 42458 6234 42460
rect 6290 42458 6314 42460
rect 6370 42458 6394 42460
rect 6450 42458 6456 42460
rect 6210 42406 6212 42458
rect 6392 42406 6394 42458
rect 6148 42404 6154 42406
rect 6210 42404 6234 42406
rect 6290 42404 6314 42406
rect 6370 42404 6394 42406
rect 6450 42404 6456 42406
rect 6148 42395 6456 42404
rect 6656 42362 6684 44540
rect 6840 42770 6868 44540
rect 7024 42770 7052 44540
rect 6828 42764 6880 42770
rect 6828 42706 6880 42712
rect 7012 42764 7064 42770
rect 7012 42706 7064 42712
rect 6736 42628 6788 42634
rect 6736 42570 6788 42576
rect 6000 42356 6052 42362
rect 6000 42298 6052 42304
rect 6644 42356 6696 42362
rect 6644 42298 6696 42304
rect 6458 42256 6514 42265
rect 6184 42220 6236 42226
rect 6458 42191 6514 42200
rect 6184 42162 6236 42168
rect 6000 42084 6052 42090
rect 6000 42026 6052 42032
rect 5908 41812 5960 41818
rect 5908 41754 5960 41760
rect 5908 41608 5960 41614
rect 5908 41550 5960 41556
rect 5920 41002 5948 41550
rect 6012 41274 6040 42026
rect 6196 41818 6224 42162
rect 6472 41818 6500 42191
rect 6184 41812 6236 41818
rect 6184 41754 6236 41760
rect 6460 41812 6512 41818
rect 6460 41754 6512 41760
rect 6148 41372 6456 41381
rect 6148 41370 6154 41372
rect 6210 41370 6234 41372
rect 6290 41370 6314 41372
rect 6370 41370 6394 41372
rect 6450 41370 6456 41372
rect 6210 41318 6212 41370
rect 6392 41318 6394 41370
rect 6148 41316 6154 41318
rect 6210 41316 6234 41318
rect 6290 41316 6314 41318
rect 6370 41316 6394 41318
rect 6450 41316 6456 41318
rect 6148 41307 6456 41316
rect 6748 41274 6776 42570
rect 7208 42362 7236 44540
rect 7392 43450 7420 44540
rect 7380 43444 7432 43450
rect 7380 43386 7432 43392
rect 7380 43308 7432 43314
rect 7380 43250 7432 43256
rect 7196 42356 7248 42362
rect 7196 42298 7248 42304
rect 7288 42220 7340 42226
rect 7288 42162 7340 42168
rect 7300 41313 7328 42162
rect 7392 41818 7420 43250
rect 7472 43172 7524 43178
rect 7472 43114 7524 43120
rect 7380 41812 7432 41818
rect 7380 41754 7432 41760
rect 7380 41608 7432 41614
rect 7378 41576 7380 41585
rect 7432 41576 7434 41585
rect 7378 41511 7434 41520
rect 7286 41304 7342 41313
rect 6000 41268 6052 41274
rect 6000 41210 6052 41216
rect 6736 41268 6788 41274
rect 7286 41239 7342 41248
rect 6736 41210 6788 41216
rect 7286 41168 7342 41177
rect 6552 41132 6604 41138
rect 7484 41154 7512 43114
rect 7576 42770 7604 44540
rect 7656 43308 7708 43314
rect 7656 43250 7708 43256
rect 7668 42906 7696 43250
rect 7656 42900 7708 42906
rect 7656 42842 7708 42848
rect 7564 42764 7616 42770
rect 7564 42706 7616 42712
rect 7760 42158 7788 44540
rect 7840 42628 7892 42634
rect 7840 42570 7892 42576
rect 7748 42152 7800 42158
rect 7748 42094 7800 42100
rect 7748 42016 7800 42022
rect 7748 41958 7800 41964
rect 7760 41682 7788 41958
rect 7852 41818 7880 42570
rect 7840 41812 7892 41818
rect 7840 41754 7892 41760
rect 7748 41676 7800 41682
rect 7748 41618 7800 41624
rect 7944 41478 7972 44540
rect 8128 43110 8156 44540
rect 8116 43104 8168 43110
rect 8116 43046 8168 43052
rect 8208 43104 8260 43110
rect 8208 43046 8260 43052
rect 8220 42922 8248 43046
rect 8128 42894 8248 42922
rect 8024 42560 8076 42566
rect 8024 42502 8076 42508
rect 7932 41472 7984 41478
rect 7562 41440 7618 41449
rect 7932 41414 7984 41420
rect 8036 41414 8064 42502
rect 8128 42242 8156 42894
rect 8312 42786 8340 44540
rect 8392 43376 8444 43382
rect 8496 43364 8524 44540
rect 8680 43738 8708 44540
rect 8588 43710 8708 43738
rect 8588 43450 8616 43710
rect 8864 43602 8892 44540
rect 8680 43574 8892 43602
rect 8576 43444 8628 43450
rect 8576 43386 8628 43392
rect 8444 43336 8524 43364
rect 8392 43318 8444 43324
rect 8484 43172 8536 43178
rect 8484 43114 8536 43120
rect 8576 43172 8628 43178
rect 8576 43114 8628 43120
rect 8220 42770 8340 42786
rect 8208 42764 8340 42770
rect 8260 42758 8340 42764
rect 8208 42706 8260 42712
rect 8392 42628 8444 42634
rect 8392 42570 8444 42576
rect 8128 42214 8248 42242
rect 8036 41386 8156 41414
rect 7562 41375 7618 41384
rect 7286 41103 7288 41112
rect 6552 41074 6604 41080
rect 7340 41103 7342 41112
rect 7392 41126 7512 41154
rect 7288 41074 7340 41080
rect 5908 40996 5960 41002
rect 5908 40938 5960 40944
rect 6564 40633 6592 41074
rect 7392 41002 7420 41126
rect 7380 40996 7432 41002
rect 7380 40938 7432 40944
rect 7472 40656 7524 40662
rect 6550 40624 6606 40633
rect 7472 40598 7524 40604
rect 6550 40559 6606 40568
rect 7380 40588 7432 40594
rect 7380 40530 7432 40536
rect 7010 40488 7066 40497
rect 6552 40452 6604 40458
rect 7010 40423 7066 40432
rect 6552 40394 6604 40400
rect 6148 40284 6456 40293
rect 6148 40282 6154 40284
rect 6210 40282 6234 40284
rect 6290 40282 6314 40284
rect 6370 40282 6394 40284
rect 6450 40282 6456 40284
rect 6210 40230 6212 40282
rect 6392 40230 6394 40282
rect 6148 40228 6154 40230
rect 6210 40228 6234 40230
rect 6290 40228 6314 40230
rect 6370 40228 6394 40230
rect 6450 40228 6456 40230
rect 6148 40219 6456 40228
rect 5998 39944 6054 39953
rect 5998 39879 6054 39888
rect 5816 39636 5868 39642
rect 5816 39578 5868 39584
rect 5724 39432 5776 39438
rect 5724 39374 5776 39380
rect 5736 37466 5764 39374
rect 6012 39098 6040 39879
rect 6148 39196 6456 39205
rect 6148 39194 6154 39196
rect 6210 39194 6234 39196
rect 6290 39194 6314 39196
rect 6370 39194 6394 39196
rect 6450 39194 6456 39196
rect 6210 39142 6212 39194
rect 6392 39142 6394 39194
rect 6148 39140 6154 39142
rect 6210 39140 6234 39142
rect 6290 39140 6314 39142
rect 6370 39140 6394 39142
rect 6450 39140 6456 39142
rect 6148 39131 6456 39140
rect 6000 39092 6052 39098
rect 6000 39034 6052 39040
rect 6564 38962 6592 40394
rect 6828 39840 6880 39846
rect 6828 39782 6880 39788
rect 6000 38956 6052 38962
rect 6000 38898 6052 38904
rect 6552 38956 6604 38962
rect 6552 38898 6604 38904
rect 6736 38956 6788 38962
rect 6736 38898 6788 38904
rect 5908 38752 5960 38758
rect 5908 38694 5960 38700
rect 5724 37460 5776 37466
rect 5724 37402 5776 37408
rect 5632 36916 5684 36922
rect 5632 36858 5684 36864
rect 5724 36576 5776 36582
rect 5724 36518 5776 36524
rect 5632 36372 5684 36378
rect 5632 36314 5684 36320
rect 5460 35958 5580 35986
rect 5262 35255 5318 35264
rect 5356 35284 5408 35290
rect 5356 35226 5408 35232
rect 5080 34672 5132 34678
rect 5080 34614 5132 34620
rect 4988 34536 5040 34542
rect 4988 34478 5040 34484
rect 5092 33998 5120 34614
rect 5460 33998 5488 35958
rect 5538 34096 5594 34105
rect 5644 34082 5672 36314
rect 5736 36038 5764 36518
rect 5816 36372 5868 36378
rect 5816 36314 5868 36320
rect 5724 36032 5776 36038
rect 5724 35974 5776 35980
rect 5828 35834 5856 36314
rect 5816 35828 5868 35834
rect 5816 35770 5868 35776
rect 5814 35592 5870 35601
rect 5724 35556 5776 35562
rect 5814 35527 5870 35536
rect 5724 35498 5776 35504
rect 5594 34054 5672 34082
rect 5538 34031 5594 34040
rect 5080 33992 5132 33998
rect 5080 33934 5132 33940
rect 5448 33992 5500 33998
rect 5448 33934 5500 33940
rect 4988 33856 5040 33862
rect 4988 33798 5040 33804
rect 4712 32564 4764 32570
rect 4712 32506 4764 32512
rect 4724 32366 4752 32506
rect 4712 32360 4764 32366
rect 4712 32302 4764 32308
rect 4710 32192 4766 32201
rect 4710 32127 4766 32136
rect 4724 31822 4752 32127
rect 4712 31816 4764 31822
rect 4712 31758 4764 31764
rect 4712 31680 4764 31686
rect 4712 31622 4764 31628
rect 4724 30734 4752 31622
rect 4712 30728 4764 30734
rect 4712 30670 4764 30676
rect 4620 29776 4672 29782
rect 4620 29718 4672 29724
rect 4618 29336 4674 29345
rect 4618 29271 4674 29280
rect 4632 29170 4660 29271
rect 4620 29164 4672 29170
rect 4620 29106 4672 29112
rect 4632 28937 4660 29106
rect 4618 28928 4674 28937
rect 4618 28863 4674 28872
rect 4632 28422 4660 28863
rect 4620 28416 4672 28422
rect 4620 28358 4672 28364
rect 4528 28076 4580 28082
rect 4528 28018 4580 28024
rect 4540 27554 4568 28018
rect 4522 27526 4568 27554
rect 4522 27316 4550 27526
rect 4522 27288 4566 27316
rect 4538 27282 4566 27288
rect 4538 27254 4568 27282
rect 4356 26846 4476 26874
rect 4356 24614 4384 26846
rect 4436 26784 4488 26790
rect 4436 26726 4488 26732
rect 4344 24608 4396 24614
rect 4250 24576 4306 24585
rect 4344 24550 4396 24556
rect 4250 24511 4306 24520
rect 4250 24440 4306 24449
rect 4250 24375 4252 24384
rect 4304 24375 4306 24384
rect 4252 24346 4304 24352
rect 4356 24290 4384 24550
rect 4172 24262 4384 24290
rect 4068 22976 4120 22982
rect 3988 22936 4068 22964
rect 3516 22704 3568 22710
rect 3516 22646 3568 22652
rect 3608 22704 3660 22710
rect 3608 22646 3660 22652
rect 3424 22636 3476 22642
rect 3424 22578 3476 22584
rect 3332 22160 3384 22166
rect 3332 22102 3384 22108
rect 3240 21888 3292 21894
rect 3240 21830 3292 21836
rect 3148 21140 3200 21146
rect 3148 21082 3200 21088
rect 2884 20964 3004 20992
rect 2884 20913 2912 20964
rect 2870 20904 2926 20913
rect 2870 20839 2926 20848
rect 2964 20868 3016 20874
rect 2884 20466 2912 20839
rect 2964 20810 3016 20816
rect 2872 20460 2924 20466
rect 2872 20402 2924 20408
rect 2780 20052 2832 20058
rect 2780 19994 2832 20000
rect 2780 19780 2832 19786
rect 2780 19722 2832 19728
rect 2792 19553 2820 19722
rect 2778 19544 2834 19553
rect 2778 19479 2834 19488
rect 2596 19372 2648 19378
rect 2596 19314 2648 19320
rect 2688 19372 2740 19378
rect 2688 19314 2740 19320
rect 2872 19372 2924 19378
rect 2872 19314 2924 19320
rect 2410 19272 2466 19281
rect 2410 19207 2466 19216
rect 2320 18828 2372 18834
rect 2320 18770 2372 18776
rect 2228 18760 2280 18766
rect 2228 18702 2280 18708
rect 1858 18320 1914 18329
rect 1858 18255 1914 18264
rect 1952 18284 2004 18290
rect 1952 18226 2004 18232
rect 1780 18176 1900 18204
rect 1872 17921 1900 18176
rect 1858 17912 1914 17921
rect 1768 17876 1820 17882
rect 1858 17847 1914 17856
rect 1768 17818 1820 17824
rect 1676 17672 1728 17678
rect 1676 17614 1728 17620
rect 1676 17536 1728 17542
rect 1676 17478 1728 17484
rect 1584 17264 1636 17270
rect 1584 17206 1636 17212
rect 1492 16448 1544 16454
rect 1492 16390 1544 16396
rect 1504 16182 1532 16390
rect 1492 16176 1544 16182
rect 1492 16118 1544 16124
rect 1582 15872 1638 15881
rect 1582 15807 1638 15816
rect 1490 15736 1546 15745
rect 1490 15671 1546 15680
rect 1398 15192 1454 15201
rect 1398 15127 1454 15136
rect 1216 14408 1268 14414
rect 1216 14350 1268 14356
rect 1216 14272 1268 14278
rect 1216 14214 1268 14220
rect 1228 10742 1256 14214
rect 1398 13832 1454 13841
rect 1398 13767 1400 13776
rect 1452 13767 1454 13776
rect 1400 13738 1452 13744
rect 1400 13388 1452 13394
rect 1400 13330 1452 13336
rect 1308 13184 1360 13190
rect 1308 13126 1360 13132
rect 1216 10736 1268 10742
rect 1216 10678 1268 10684
rect 1216 10532 1268 10538
rect 1216 10474 1268 10480
rect 1228 6458 1256 10474
rect 1320 7478 1348 13126
rect 1412 12782 1440 13330
rect 1400 12776 1452 12782
rect 1400 12718 1452 12724
rect 1412 11762 1440 12718
rect 1504 12646 1532 15671
rect 1492 12640 1544 12646
rect 1492 12582 1544 12588
rect 1596 12442 1624 15807
rect 1688 15502 1716 17478
rect 1780 17338 1808 17818
rect 1768 17332 1820 17338
rect 1768 17274 1820 17280
rect 1964 17241 1992 18226
rect 2332 18222 2360 18770
rect 2596 18760 2648 18766
rect 2596 18702 2648 18708
rect 2320 18216 2372 18222
rect 2320 18158 2372 18164
rect 2502 18184 2558 18193
rect 2228 18080 2280 18086
rect 2228 18022 2280 18028
rect 2044 17740 2096 17746
rect 2044 17682 2096 17688
rect 1950 17232 2006 17241
rect 1950 17167 2006 17176
rect 1860 17060 1912 17066
rect 1860 17002 1912 17008
rect 1766 16960 1822 16969
rect 1766 16895 1822 16904
rect 1676 15496 1728 15502
rect 1676 15438 1728 15444
rect 1780 14618 1808 16895
rect 1872 14822 1900 17002
rect 1952 16788 2004 16794
rect 1952 16730 2004 16736
rect 1964 15484 1992 16730
rect 2056 16046 2084 17682
rect 2136 17672 2188 17678
rect 2134 17640 2136 17649
rect 2188 17640 2190 17649
rect 2134 17575 2190 17584
rect 2044 16040 2096 16046
rect 2044 15982 2096 15988
rect 2044 15496 2096 15502
rect 1964 15456 2044 15484
rect 2044 15438 2096 15444
rect 1860 14816 1912 14822
rect 1912 14776 1992 14804
rect 1860 14758 1912 14764
rect 1768 14612 1820 14618
rect 1768 14554 1820 14560
rect 1858 14512 1914 14521
rect 1858 14447 1914 14456
rect 1674 14240 1730 14249
rect 1674 14175 1730 14184
rect 1584 12436 1636 12442
rect 1584 12378 1636 12384
rect 1490 12200 1546 12209
rect 1490 12135 1492 12144
rect 1544 12135 1546 12144
rect 1492 12106 1544 12112
rect 1582 11928 1638 11937
rect 1582 11863 1584 11872
rect 1636 11863 1638 11872
rect 1584 11834 1636 11840
rect 1582 11792 1638 11801
rect 1400 11756 1452 11762
rect 1582 11727 1638 11736
rect 1400 11698 1452 11704
rect 1412 10130 1440 11698
rect 1490 11656 1546 11665
rect 1490 11591 1546 11600
rect 1504 10962 1532 11591
rect 1596 11150 1624 11727
rect 1688 11506 1716 14175
rect 1766 13968 1822 13977
rect 1766 13903 1768 13912
rect 1820 13903 1822 13912
rect 1768 13874 1820 13880
rect 1766 13560 1822 13569
rect 1766 13495 1822 13504
rect 1780 12186 1808 13495
rect 1872 12322 1900 14447
rect 1964 13870 1992 14776
rect 1952 13864 2004 13870
rect 1952 13806 2004 13812
rect 1964 13394 1992 13806
rect 1952 13388 2004 13394
rect 1952 13330 2004 13336
rect 2056 12730 2084 15438
rect 2148 15416 2176 17575
rect 2240 16590 2268 18022
rect 2332 17066 2360 18158
rect 2502 18119 2558 18128
rect 2516 17814 2544 18119
rect 2504 17808 2556 17814
rect 2504 17750 2556 17756
rect 2412 17740 2464 17746
rect 2412 17682 2464 17688
rect 2320 17060 2372 17066
rect 2320 17002 2372 17008
rect 2318 16824 2374 16833
rect 2318 16759 2374 16768
rect 2228 16584 2280 16590
rect 2228 16526 2280 16532
rect 2332 16114 2360 16759
rect 2320 16108 2372 16114
rect 2320 16050 2372 16056
rect 2424 15706 2452 17682
rect 2608 17542 2636 18702
rect 2700 18290 2728 19314
rect 2884 19145 2912 19314
rect 2870 19136 2926 19145
rect 2870 19071 2926 19080
rect 2976 18358 3004 20810
rect 3146 20768 3202 20777
rect 3068 20726 3146 20754
rect 3068 19718 3096 20726
rect 3146 20703 3202 20712
rect 3148 20528 3200 20534
rect 3252 20505 3280 21830
rect 3344 20788 3372 22102
rect 3436 21690 3464 22578
rect 3884 22568 3936 22574
rect 3884 22510 3936 22516
rect 3549 22332 3857 22341
rect 3549 22330 3555 22332
rect 3611 22330 3635 22332
rect 3691 22330 3715 22332
rect 3771 22330 3795 22332
rect 3851 22330 3857 22332
rect 3611 22278 3613 22330
rect 3793 22278 3795 22330
rect 3549 22276 3555 22278
rect 3611 22276 3635 22278
rect 3691 22276 3715 22278
rect 3771 22276 3795 22278
rect 3851 22276 3857 22278
rect 3549 22267 3857 22276
rect 3896 21690 3924 22510
rect 3424 21684 3476 21690
rect 3424 21626 3476 21632
rect 3884 21684 3936 21690
rect 3884 21626 3936 21632
rect 3884 21344 3936 21350
rect 3884 21286 3936 21292
rect 3549 21244 3857 21253
rect 3549 21242 3555 21244
rect 3611 21242 3635 21244
rect 3691 21242 3715 21244
rect 3771 21242 3795 21244
rect 3851 21242 3857 21244
rect 3611 21190 3613 21242
rect 3793 21190 3795 21242
rect 3549 21188 3555 21190
rect 3611 21188 3635 21190
rect 3691 21188 3715 21190
rect 3771 21188 3795 21190
rect 3851 21188 3857 21190
rect 3549 21179 3857 21188
rect 3424 20800 3476 20806
rect 3344 20760 3424 20788
rect 3344 20534 3372 20760
rect 3424 20742 3476 20748
rect 3332 20528 3384 20534
rect 3148 20470 3200 20476
rect 3238 20496 3294 20505
rect 3160 19718 3188 20470
rect 3332 20470 3384 20476
rect 3238 20431 3294 20440
rect 3896 20398 3924 21286
rect 3884 20392 3936 20398
rect 3884 20334 3936 20340
rect 3516 20256 3568 20262
rect 3436 20216 3516 20244
rect 3238 19952 3294 19961
rect 3238 19887 3240 19896
rect 3292 19887 3294 19896
rect 3240 19858 3292 19864
rect 3056 19712 3108 19718
rect 3056 19654 3108 19660
rect 3148 19712 3200 19718
rect 3148 19654 3200 19660
rect 3160 19334 3188 19654
rect 3330 19544 3386 19553
rect 3330 19479 3386 19488
rect 3238 19408 3294 19417
rect 3344 19378 3372 19479
rect 3238 19343 3294 19352
rect 3332 19372 3384 19378
rect 3068 19306 3188 19334
rect 2964 18352 3016 18358
rect 2964 18294 3016 18300
rect 2688 18284 2740 18290
rect 2688 18226 2740 18232
rect 2778 18048 2834 18057
rect 2778 17983 2834 17992
rect 2686 17912 2742 17921
rect 2792 17898 2820 17983
rect 2742 17870 2820 17898
rect 2686 17847 2742 17856
rect 2778 17776 2834 17785
rect 2688 17740 2740 17746
rect 2740 17720 2778 17728
rect 3068 17762 3096 19306
rect 3252 18834 3280 19343
rect 3332 19314 3384 19320
rect 3240 18828 3292 18834
rect 3240 18770 3292 18776
rect 3436 18714 3464 20216
rect 3516 20198 3568 20204
rect 3549 20156 3857 20165
rect 3549 20154 3555 20156
rect 3611 20154 3635 20156
rect 3691 20154 3715 20156
rect 3771 20154 3795 20156
rect 3851 20154 3857 20156
rect 3611 20102 3613 20154
rect 3793 20102 3795 20154
rect 3549 20100 3555 20102
rect 3611 20100 3635 20102
rect 3691 20100 3715 20102
rect 3771 20100 3795 20102
rect 3851 20100 3857 20102
rect 3549 20091 3857 20100
rect 3549 19068 3857 19077
rect 3549 19066 3555 19068
rect 3611 19066 3635 19068
rect 3691 19066 3715 19068
rect 3771 19066 3795 19068
rect 3851 19066 3857 19068
rect 3611 19014 3613 19066
rect 3793 19014 3795 19066
rect 3549 19012 3555 19014
rect 3611 19012 3635 19014
rect 3691 19012 3715 19014
rect 3771 19012 3795 19014
rect 3851 19012 3857 19014
rect 3549 19003 3857 19012
rect 3988 18816 4016 22936
rect 4068 22918 4120 22924
rect 4172 22794 4200 24262
rect 4342 24168 4398 24177
rect 4342 24103 4344 24112
rect 4396 24103 4398 24112
rect 4344 24074 4396 24080
rect 4448 23594 4476 26726
rect 4540 26364 4568 27254
rect 4620 26920 4672 26926
rect 4620 26862 4672 26868
rect 4632 26518 4660 26862
rect 4620 26512 4672 26518
rect 4620 26454 4672 26460
rect 4540 26336 4660 26364
rect 4526 25800 4582 25809
rect 4526 25735 4528 25744
rect 4580 25735 4582 25744
rect 4528 25706 4580 25712
rect 4526 25664 4582 25673
rect 4526 25599 4582 25608
rect 4540 25226 4568 25599
rect 4528 25220 4580 25226
rect 4528 25162 4580 25168
rect 4540 24886 4568 25162
rect 4528 24880 4580 24886
rect 4528 24822 4580 24828
rect 4528 24200 4580 24206
rect 4528 24142 4580 24148
rect 4436 23588 4488 23594
rect 4436 23530 4488 23536
rect 4250 23216 4306 23225
rect 4250 23151 4306 23160
rect 4080 22766 4200 22794
rect 4080 21554 4108 22766
rect 4160 22228 4212 22234
rect 4160 22170 4212 22176
rect 4068 21548 4120 21554
rect 4068 21490 4120 21496
rect 4172 20602 4200 22170
rect 4264 22166 4292 23151
rect 4344 22976 4396 22982
rect 4344 22918 4396 22924
rect 4356 22710 4384 22918
rect 4344 22704 4396 22710
rect 4344 22646 4396 22652
rect 4436 22704 4488 22710
rect 4436 22646 4488 22652
rect 4342 22264 4398 22273
rect 4342 22199 4398 22208
rect 4252 22160 4304 22166
rect 4252 22102 4304 22108
rect 4250 21720 4306 21729
rect 4250 21655 4306 21664
rect 4264 21350 4292 21655
rect 4356 21622 4384 22199
rect 4344 21616 4396 21622
rect 4344 21558 4396 21564
rect 4252 21344 4304 21350
rect 4448 21321 4476 22646
rect 4540 21690 4568 24142
rect 4632 23050 4660 26336
rect 4724 23118 4752 30670
rect 4816 28994 4844 33102
rect 4896 33108 4948 33114
rect 4896 33050 4948 33056
rect 4896 32768 4948 32774
rect 4896 32710 4948 32716
rect 4908 32366 4936 32710
rect 4896 32360 4948 32366
rect 4896 32302 4948 32308
rect 4896 31884 4948 31890
rect 4896 31826 4948 31832
rect 4908 31686 4936 31826
rect 4896 31680 4948 31686
rect 4896 31622 4948 31628
rect 5000 30818 5028 33798
rect 5092 33590 5120 33934
rect 5172 33856 5224 33862
rect 5172 33798 5224 33804
rect 5264 33856 5316 33862
rect 5264 33798 5316 33804
rect 5080 33584 5132 33590
rect 5080 33526 5132 33532
rect 5080 33108 5132 33114
rect 5080 33050 5132 33056
rect 5092 33017 5120 33050
rect 5078 33008 5134 33017
rect 5078 32943 5134 32952
rect 4908 30790 5028 30818
rect 4908 30598 4936 30790
rect 4988 30728 5040 30734
rect 4988 30670 5040 30676
rect 4896 30592 4948 30598
rect 4896 30534 4948 30540
rect 5000 30394 5028 30670
rect 4988 30388 5040 30394
rect 4988 30330 5040 30336
rect 4896 30184 4948 30190
rect 4896 30126 4948 30132
rect 4908 29170 4936 30126
rect 4896 29164 4948 29170
rect 4896 29106 4948 29112
rect 4816 28966 5028 28994
rect 4896 28416 4948 28422
rect 4896 28358 4948 28364
rect 4908 28150 4936 28358
rect 4896 28144 4948 28150
rect 4896 28086 4948 28092
rect 4804 28076 4856 28082
rect 4804 28018 4856 28024
rect 4816 27334 4844 28018
rect 4894 27976 4950 27985
rect 4894 27911 4950 27920
rect 4908 27402 4936 27911
rect 4896 27396 4948 27402
rect 4896 27338 4948 27344
rect 4804 27328 4856 27334
rect 4804 27270 4856 27276
rect 4894 27296 4950 27305
rect 4816 24206 4844 27270
rect 4894 27231 4950 27240
rect 4908 24206 4936 27231
rect 5000 24954 5028 28966
rect 5092 27713 5120 32943
rect 5184 32842 5212 33798
rect 5172 32836 5224 32842
rect 5172 32778 5224 32784
rect 5170 32056 5226 32065
rect 5170 31991 5172 32000
rect 5224 31991 5226 32000
rect 5172 31962 5224 31968
rect 5276 31890 5304 33798
rect 5540 33584 5592 33590
rect 5540 33526 5592 33532
rect 5356 33448 5408 33454
rect 5356 33390 5408 33396
rect 5368 33046 5396 33390
rect 5356 33040 5408 33046
rect 5356 32982 5408 32988
rect 5552 32910 5580 33526
rect 5632 33312 5684 33318
rect 5632 33254 5684 33260
rect 5644 32978 5672 33254
rect 5632 32972 5684 32978
rect 5632 32914 5684 32920
rect 5540 32904 5592 32910
rect 5592 32852 5672 32858
rect 5540 32846 5672 32852
rect 5356 32836 5408 32842
rect 5552 32830 5672 32846
rect 5356 32778 5408 32784
rect 5264 31884 5316 31890
rect 5264 31826 5316 31832
rect 5368 31686 5396 32778
rect 5448 32768 5500 32774
rect 5448 32710 5500 32716
rect 5356 31680 5408 31686
rect 5356 31622 5408 31628
rect 5262 31512 5318 31521
rect 5262 31447 5318 31456
rect 5276 31346 5304 31447
rect 5264 31340 5316 31346
rect 5264 31282 5316 31288
rect 5170 31104 5226 31113
rect 5170 31039 5226 31048
rect 5184 30841 5212 31039
rect 5354 30968 5410 30977
rect 5354 30903 5356 30912
rect 5408 30903 5410 30912
rect 5356 30874 5408 30880
rect 5170 30832 5226 30841
rect 5170 30767 5226 30776
rect 5356 30796 5408 30802
rect 5184 30258 5212 30767
rect 5356 30738 5408 30744
rect 5264 30592 5316 30598
rect 5264 30534 5316 30540
rect 5172 30252 5224 30258
rect 5172 30194 5224 30200
rect 5184 30161 5212 30194
rect 5170 30152 5226 30161
rect 5170 30087 5226 30096
rect 5172 29844 5224 29850
rect 5172 29786 5224 29792
rect 5184 29170 5212 29786
rect 5172 29164 5224 29170
rect 5172 29106 5224 29112
rect 5184 29073 5212 29106
rect 5170 29064 5226 29073
rect 5170 28999 5226 29008
rect 5276 28994 5304 30534
rect 5368 30161 5396 30738
rect 5354 30152 5410 30161
rect 5354 30087 5410 30096
rect 5460 29578 5488 32710
rect 5540 32020 5592 32026
rect 5540 31962 5592 31968
rect 5448 29572 5500 29578
rect 5448 29514 5500 29520
rect 5276 28966 5396 28994
rect 5172 28688 5224 28694
rect 5224 28665 5304 28676
rect 5224 28656 5318 28665
rect 5224 28648 5262 28656
rect 5172 28630 5224 28636
rect 5262 28591 5318 28600
rect 5172 28552 5224 28558
rect 5172 28494 5224 28500
rect 5184 28218 5212 28494
rect 5172 28212 5224 28218
rect 5172 28154 5224 28160
rect 5172 28076 5224 28082
rect 5172 28018 5224 28024
rect 5078 27704 5134 27713
rect 5078 27639 5134 27648
rect 5184 27606 5212 28018
rect 5276 27878 5304 28591
rect 5264 27872 5316 27878
rect 5264 27814 5316 27820
rect 5172 27600 5224 27606
rect 5172 27542 5224 27548
rect 5368 27441 5396 28966
rect 5078 27432 5134 27441
rect 5078 27367 5134 27376
rect 5354 27432 5410 27441
rect 5354 27367 5410 27376
rect 5092 26908 5120 27367
rect 5368 27062 5396 27367
rect 5264 27056 5316 27062
rect 5264 26998 5316 27004
rect 5356 27056 5408 27062
rect 5356 26998 5408 27004
rect 5092 26880 5212 26908
rect 5184 26382 5212 26880
rect 5276 26625 5304 26998
rect 5262 26616 5318 26625
rect 5262 26551 5318 26560
rect 5172 26376 5224 26382
rect 5172 26318 5224 26324
rect 5078 25256 5134 25265
rect 5078 25191 5134 25200
rect 4988 24948 5040 24954
rect 4988 24890 5040 24896
rect 4986 24440 5042 24449
rect 4986 24375 5042 24384
rect 5000 24342 5028 24375
rect 4988 24336 5040 24342
rect 4988 24278 5040 24284
rect 4804 24200 4856 24206
rect 4804 24142 4856 24148
rect 4896 24200 4948 24206
rect 4896 24142 4948 24148
rect 5000 24052 5028 24278
rect 4802 24032 4858 24041
rect 4802 23967 4858 23976
rect 4908 24024 5028 24052
rect 4816 23322 4844 23967
rect 4804 23316 4856 23322
rect 4804 23258 4856 23264
rect 4712 23112 4764 23118
rect 4712 23054 4764 23060
rect 4620 23044 4672 23050
rect 4620 22986 4672 22992
rect 4804 22976 4856 22982
rect 4804 22918 4856 22924
rect 4816 22778 4844 22918
rect 4804 22772 4856 22778
rect 4804 22714 4856 22720
rect 4908 22658 4936 24024
rect 5092 23361 5120 25191
rect 5184 24857 5212 26318
rect 5276 25276 5304 26551
rect 5356 26376 5408 26382
rect 5356 26318 5408 26324
rect 5368 26042 5396 26318
rect 5356 26036 5408 26042
rect 5356 25978 5408 25984
rect 5356 25288 5408 25294
rect 5276 25248 5356 25276
rect 5356 25230 5408 25236
rect 5170 24848 5226 24857
rect 5368 24834 5396 25230
rect 5460 24954 5488 29514
rect 5552 28626 5580 31962
rect 5644 29578 5672 32830
rect 5736 31890 5764 35498
rect 5828 35290 5856 35527
rect 5816 35284 5868 35290
rect 5816 35226 5868 35232
rect 5816 34944 5868 34950
rect 5816 34886 5868 34892
rect 5828 34678 5856 34886
rect 5920 34762 5948 38694
rect 6012 38010 6040 38898
rect 6644 38752 6696 38758
rect 6644 38694 6696 38700
rect 6656 38350 6684 38694
rect 6644 38344 6696 38350
rect 6644 38286 6696 38292
rect 6552 38208 6604 38214
rect 6552 38150 6604 38156
rect 6148 38108 6456 38117
rect 6148 38106 6154 38108
rect 6210 38106 6234 38108
rect 6290 38106 6314 38108
rect 6370 38106 6394 38108
rect 6450 38106 6456 38108
rect 6210 38054 6212 38106
rect 6392 38054 6394 38106
rect 6148 38052 6154 38054
rect 6210 38052 6234 38054
rect 6290 38052 6314 38054
rect 6370 38052 6394 38054
rect 6450 38052 6456 38054
rect 6148 38043 6456 38052
rect 6000 38004 6052 38010
rect 6000 37946 6052 37952
rect 6276 37868 6328 37874
rect 6276 37810 6328 37816
rect 6288 37126 6316 37810
rect 6564 37330 6592 38150
rect 6644 37664 6696 37670
rect 6644 37606 6696 37612
rect 6552 37324 6604 37330
rect 6552 37266 6604 37272
rect 6656 37262 6684 37606
rect 6368 37256 6420 37262
rect 6644 37256 6696 37262
rect 6420 37216 6500 37244
rect 6368 37198 6420 37204
rect 6472 37210 6500 37216
rect 6472 37182 6592 37210
rect 6644 37198 6696 37204
rect 6276 37120 6328 37126
rect 6564 37097 6592 37182
rect 6276 37062 6328 37068
rect 6550 37088 6606 37097
rect 6148 37020 6456 37029
rect 6550 37023 6606 37032
rect 6148 37018 6154 37020
rect 6210 37018 6234 37020
rect 6290 37018 6314 37020
rect 6370 37018 6394 37020
rect 6450 37018 6456 37020
rect 6210 36966 6212 37018
rect 6392 36966 6394 37018
rect 6148 36964 6154 36966
rect 6210 36964 6234 36966
rect 6290 36964 6314 36966
rect 6370 36964 6394 36966
rect 6450 36964 6456 36966
rect 5998 36952 6054 36961
rect 6148 36955 6456 36964
rect 6054 36896 6224 36904
rect 5998 36887 6224 36896
rect 6012 36876 6224 36887
rect 6090 36816 6146 36825
rect 6000 36780 6052 36786
rect 6090 36751 6146 36760
rect 6000 36722 6052 36728
rect 6012 35601 6040 36722
rect 6104 36174 6132 36751
rect 6092 36168 6144 36174
rect 6092 36110 6144 36116
rect 6196 36038 6224 36876
rect 6368 36780 6420 36786
rect 6368 36722 6420 36728
rect 6380 36553 6408 36722
rect 6366 36544 6422 36553
rect 6366 36479 6422 36488
rect 6184 36032 6236 36038
rect 6184 35974 6236 35980
rect 6148 35932 6456 35941
rect 6148 35930 6154 35932
rect 6210 35930 6234 35932
rect 6290 35930 6314 35932
rect 6370 35930 6394 35932
rect 6450 35930 6456 35932
rect 6210 35878 6212 35930
rect 6392 35878 6394 35930
rect 6148 35876 6154 35878
rect 6210 35876 6234 35878
rect 6290 35876 6314 35878
rect 6370 35876 6394 35878
rect 6450 35876 6456 35878
rect 6148 35867 6456 35876
rect 5998 35592 6054 35601
rect 5998 35527 6054 35536
rect 6644 35556 6696 35562
rect 6644 35498 6696 35504
rect 6656 35290 6684 35498
rect 6644 35284 6696 35290
rect 6644 35226 6696 35232
rect 6748 35034 6776 38898
rect 6840 38554 6868 39782
rect 6828 38548 6880 38554
rect 6828 38490 6880 38496
rect 6920 38344 6972 38350
rect 6840 38304 6920 38332
rect 6840 36718 6868 38304
rect 6920 38286 6972 38292
rect 6920 37664 6972 37670
rect 6920 37606 6972 37612
rect 6932 37194 6960 37606
rect 6920 37188 6972 37194
rect 6920 37130 6972 37136
rect 6932 36825 6960 37130
rect 6918 36816 6974 36825
rect 6918 36751 6974 36760
rect 6828 36712 6880 36718
rect 6828 36654 6880 36660
rect 6920 36644 6972 36650
rect 6920 36586 6972 36592
rect 6932 36242 6960 36586
rect 6920 36236 6972 36242
rect 6840 36196 6920 36224
rect 6840 35630 6868 36196
rect 6920 36178 6972 36184
rect 6918 36136 6974 36145
rect 6918 36071 6974 36080
rect 6932 36038 6960 36071
rect 6920 36032 6972 36038
rect 6920 35974 6972 35980
rect 6828 35624 6880 35630
rect 6828 35566 6880 35572
rect 7024 35222 7052 40423
rect 7392 38842 7420 40530
rect 7300 38814 7420 38842
rect 7196 38208 7248 38214
rect 7102 38176 7158 38185
rect 7196 38150 7248 38156
rect 7102 38111 7158 38120
rect 7116 37942 7144 38111
rect 7104 37936 7156 37942
rect 7104 37878 7156 37884
rect 7104 37120 7156 37126
rect 7104 37062 7156 37068
rect 7012 35216 7064 35222
rect 7012 35158 7064 35164
rect 6644 35012 6696 35018
rect 6748 35006 6868 35034
rect 6644 34954 6696 34960
rect 6000 34944 6052 34950
rect 5998 34912 6000 34921
rect 6052 34912 6054 34921
rect 5998 34847 6054 34856
rect 6148 34844 6456 34853
rect 6148 34842 6154 34844
rect 6210 34842 6234 34844
rect 6290 34842 6314 34844
rect 6370 34842 6394 34844
rect 6450 34842 6456 34844
rect 6210 34790 6212 34842
rect 6392 34790 6394 34842
rect 6148 34788 6154 34790
rect 6210 34788 6234 34790
rect 6290 34788 6314 34790
rect 6370 34788 6394 34790
rect 6450 34788 6456 34790
rect 6148 34779 6456 34788
rect 5920 34746 6040 34762
rect 5920 34740 6052 34746
rect 5920 34734 6000 34740
rect 6000 34682 6052 34688
rect 6460 34740 6512 34746
rect 6460 34682 6512 34688
rect 5816 34672 5868 34678
rect 5816 34614 5868 34620
rect 6092 34672 6144 34678
rect 6092 34614 6144 34620
rect 6000 34604 6052 34610
rect 6000 34546 6052 34552
rect 5908 34536 5960 34542
rect 5908 34478 5960 34484
rect 5920 33522 5948 34478
rect 6012 33998 6040 34546
rect 6000 33992 6052 33998
rect 6000 33934 6052 33940
rect 5908 33516 5960 33522
rect 5908 33458 5960 33464
rect 5816 33312 5868 33318
rect 5816 33254 5868 33260
rect 5828 32910 5856 33254
rect 5816 32904 5868 32910
rect 5816 32846 5868 32852
rect 5816 32564 5868 32570
rect 5816 32506 5868 32512
rect 5724 31884 5776 31890
rect 5724 31826 5776 31832
rect 5736 31793 5764 31826
rect 5722 31784 5778 31793
rect 5722 31719 5778 31728
rect 5724 31340 5776 31346
rect 5724 31282 5776 31288
rect 5736 30172 5764 31282
rect 5828 30326 5856 32506
rect 5920 32298 5948 33458
rect 6012 32842 6040 33934
rect 6104 33862 6132 34614
rect 6472 34241 6500 34682
rect 6458 34232 6514 34241
rect 6458 34167 6514 34176
rect 6472 33980 6500 34167
rect 6552 33992 6604 33998
rect 6472 33952 6552 33980
rect 6552 33934 6604 33940
rect 6656 33946 6684 34954
rect 6840 34746 6868 35006
rect 7116 34746 7144 37062
rect 7208 36718 7236 38150
rect 7300 37874 7328 38814
rect 7380 38752 7432 38758
rect 7380 38694 7432 38700
rect 7288 37868 7340 37874
rect 7288 37810 7340 37816
rect 7392 37330 7420 38694
rect 7380 37324 7432 37330
rect 7380 37266 7432 37272
rect 7196 36712 7248 36718
rect 7196 36654 7248 36660
rect 7208 36242 7236 36654
rect 7196 36236 7248 36242
rect 7196 36178 7248 36184
rect 7208 35290 7236 36178
rect 7288 36168 7340 36174
rect 7288 36110 7340 36116
rect 7300 35290 7328 36110
rect 7196 35284 7248 35290
rect 7196 35226 7248 35232
rect 7288 35284 7340 35290
rect 7288 35226 7340 35232
rect 6828 34740 6880 34746
rect 6828 34682 6880 34688
rect 7104 34740 7156 34746
rect 7104 34682 7156 34688
rect 6826 34640 6882 34649
rect 7208 34610 7236 35226
rect 7288 35080 7340 35086
rect 7288 35022 7340 35028
rect 6826 34575 6882 34584
rect 7196 34604 7248 34610
rect 6840 34474 6868 34575
rect 7196 34546 7248 34552
rect 6828 34468 6880 34474
rect 6828 34410 6880 34416
rect 6656 33918 6776 33946
rect 6092 33856 6144 33862
rect 6644 33856 6696 33862
rect 6144 33816 6592 33844
rect 6092 33798 6144 33804
rect 6148 33756 6456 33765
rect 6148 33754 6154 33756
rect 6210 33754 6234 33756
rect 6290 33754 6314 33756
rect 6370 33754 6394 33756
rect 6450 33754 6456 33756
rect 6210 33702 6212 33754
rect 6392 33702 6394 33754
rect 6148 33700 6154 33702
rect 6210 33700 6234 33702
rect 6290 33700 6314 33702
rect 6370 33700 6394 33702
rect 6450 33700 6456 33702
rect 6148 33691 6456 33700
rect 6000 32836 6052 32842
rect 6000 32778 6052 32784
rect 6012 32552 6040 32778
rect 6564 32774 6592 33816
rect 6644 33798 6696 33804
rect 6656 33114 6684 33798
rect 6748 33590 6776 33918
rect 6736 33584 6788 33590
rect 6736 33526 6788 33532
rect 6736 33448 6788 33454
rect 6736 33390 6788 33396
rect 6644 33108 6696 33114
rect 6644 33050 6696 33056
rect 6748 32994 6776 33390
rect 6656 32966 6776 32994
rect 6656 32858 6684 32966
rect 6654 32830 6684 32858
rect 6552 32768 6604 32774
rect 6654 32756 6682 32830
rect 6736 32768 6788 32774
rect 6654 32728 6684 32756
rect 6552 32710 6604 32716
rect 6148 32668 6456 32677
rect 6148 32666 6154 32668
rect 6210 32666 6234 32668
rect 6290 32666 6314 32668
rect 6370 32666 6394 32668
rect 6450 32666 6456 32668
rect 6210 32614 6212 32666
rect 6392 32614 6394 32666
rect 6148 32612 6154 32614
rect 6210 32612 6234 32614
rect 6290 32612 6314 32614
rect 6370 32612 6394 32614
rect 6450 32612 6456 32614
rect 6148 32603 6456 32612
rect 6012 32524 6316 32552
rect 6184 32360 6236 32366
rect 5998 32328 6054 32337
rect 5908 32292 5960 32298
rect 6184 32302 6236 32308
rect 5998 32263 6054 32272
rect 5908 32234 5960 32240
rect 5920 31346 5948 32234
rect 6012 32230 6040 32263
rect 6000 32224 6052 32230
rect 6000 32166 6052 32172
rect 6012 31890 6040 32166
rect 6000 31884 6052 31890
rect 6000 31826 6052 31832
rect 6196 31822 6224 32302
rect 6184 31816 6236 31822
rect 6184 31758 6236 31764
rect 6288 31686 6316 32524
rect 6000 31680 6052 31686
rect 6000 31622 6052 31628
rect 6276 31680 6328 31686
rect 6276 31622 6328 31628
rect 5908 31340 5960 31346
rect 5908 31282 5960 31288
rect 5908 31136 5960 31142
rect 5908 31078 5960 31084
rect 5920 30802 5948 31078
rect 5908 30796 5960 30802
rect 5908 30738 5960 30744
rect 5906 30560 5962 30569
rect 5906 30495 5962 30504
rect 5920 30394 5948 30495
rect 5908 30388 5960 30394
rect 5908 30330 5960 30336
rect 5816 30320 5868 30326
rect 5816 30262 5868 30268
rect 5736 30144 5856 30172
rect 5632 29572 5684 29578
rect 5632 29514 5684 29520
rect 5724 29572 5776 29578
rect 5724 29514 5776 29520
rect 5540 28620 5592 28626
rect 5540 28562 5592 28568
rect 5540 28416 5592 28422
rect 5540 28358 5592 28364
rect 5552 28121 5580 28358
rect 5538 28112 5594 28121
rect 5538 28047 5594 28056
rect 5540 27464 5592 27470
rect 5540 27406 5592 27412
rect 5552 27130 5580 27406
rect 5540 27124 5592 27130
rect 5540 27066 5592 27072
rect 5538 27024 5594 27033
rect 5538 26959 5594 26968
rect 5552 25480 5580 26959
rect 5644 26926 5672 29514
rect 5736 29306 5764 29514
rect 5724 29300 5776 29306
rect 5724 29242 5776 29248
rect 5722 27976 5778 27985
rect 5722 27911 5778 27920
rect 5632 26920 5684 26926
rect 5632 26862 5684 26868
rect 5552 25452 5672 25480
rect 5644 25294 5672 25452
rect 5632 25288 5684 25294
rect 5632 25230 5684 25236
rect 5736 25106 5764 27911
rect 5552 25078 5764 25106
rect 5448 24948 5500 24954
rect 5448 24890 5500 24896
rect 5368 24806 5488 24834
rect 5170 24783 5226 24792
rect 5356 23792 5408 23798
rect 5356 23734 5408 23740
rect 5172 23724 5224 23730
rect 5224 23684 5304 23712
rect 5172 23666 5224 23672
rect 5276 23497 5304 23684
rect 5262 23488 5318 23497
rect 5262 23423 5318 23432
rect 5078 23352 5134 23361
rect 5078 23287 5134 23296
rect 5368 23202 5396 23734
rect 5184 23174 5396 23202
rect 4988 23044 5040 23050
rect 4988 22986 5040 22992
rect 4724 22630 4936 22658
rect 4618 22536 4674 22545
rect 4618 22471 4620 22480
rect 4672 22471 4674 22480
rect 4620 22442 4672 22448
rect 4620 22228 4672 22234
rect 4620 22170 4672 22176
rect 4632 22030 4660 22170
rect 4620 22024 4672 22030
rect 4620 21966 4672 21972
rect 4618 21856 4674 21865
rect 4618 21791 4674 21800
rect 4528 21684 4580 21690
rect 4528 21626 4580 21632
rect 4252 21286 4304 21292
rect 4434 21312 4490 21321
rect 4434 21247 4490 21256
rect 4252 20936 4304 20942
rect 4252 20878 4304 20884
rect 4342 20904 4398 20913
rect 4160 20596 4212 20602
rect 4160 20538 4212 20544
rect 4066 20496 4122 20505
rect 4066 20431 4122 20440
rect 4080 20233 4108 20431
rect 4066 20224 4122 20233
rect 4066 20159 4122 20168
rect 4068 18828 4120 18834
rect 3988 18788 4068 18816
rect 4068 18770 4120 18776
rect 3252 18686 3464 18714
rect 3148 18420 3200 18426
rect 3148 18362 3200 18368
rect 2740 17711 2834 17720
rect 2884 17734 3096 17762
rect 2740 17700 2820 17711
rect 2688 17682 2740 17688
rect 2596 17536 2648 17542
rect 2596 17478 2648 17484
rect 2608 17202 2636 17478
rect 2686 17368 2742 17377
rect 2686 17303 2688 17312
rect 2740 17303 2742 17312
rect 2688 17274 2740 17280
rect 2596 17196 2648 17202
rect 2596 17138 2648 17144
rect 2596 16584 2648 16590
rect 2596 16526 2648 16532
rect 2608 16046 2636 16526
rect 2596 16040 2648 16046
rect 2596 15982 2648 15988
rect 2504 15972 2556 15978
rect 2504 15914 2556 15920
rect 2412 15700 2464 15706
rect 2412 15642 2464 15648
rect 2148 15388 2268 15416
rect 2134 15328 2190 15337
rect 2134 15263 2190 15272
rect 2148 13326 2176 15263
rect 2136 13320 2188 13326
rect 2136 13262 2188 13268
rect 2240 12850 2268 15388
rect 2410 15192 2466 15201
rect 2410 15127 2466 15136
rect 2424 14278 2452 15127
rect 2412 14272 2464 14278
rect 2412 14214 2464 14220
rect 2516 13954 2544 15914
rect 2608 15065 2636 15982
rect 2594 15056 2650 15065
rect 2594 14991 2650 15000
rect 2700 14346 2728 17274
rect 2780 17196 2832 17202
rect 2780 17138 2832 17144
rect 2792 16590 2820 17138
rect 2780 16584 2832 16590
rect 2780 16526 2832 16532
rect 2780 16244 2832 16250
rect 2780 16186 2832 16192
rect 2688 14340 2740 14346
rect 2688 14282 2740 14288
rect 2516 13926 2728 13954
rect 2412 13728 2464 13734
rect 2412 13670 2464 13676
rect 2228 12844 2280 12850
rect 2228 12786 2280 12792
rect 2320 12776 2372 12782
rect 2056 12702 2268 12730
rect 2320 12718 2372 12724
rect 2240 12374 2268 12702
rect 2136 12368 2188 12374
rect 1872 12294 1992 12322
rect 2136 12310 2188 12316
rect 2228 12368 2280 12374
rect 2228 12310 2280 12316
rect 1780 12158 1900 12186
rect 1768 11824 1820 11830
rect 1766 11792 1768 11801
rect 1820 11792 1822 11801
rect 1766 11727 1822 11736
rect 1688 11478 1808 11506
rect 1674 11384 1730 11393
rect 1674 11319 1730 11328
rect 1584 11144 1636 11150
rect 1584 11086 1636 11092
rect 1504 10934 1624 10962
rect 1492 10260 1544 10266
rect 1492 10202 1544 10208
rect 1400 10124 1452 10130
rect 1400 10066 1452 10072
rect 1412 9042 1440 10066
rect 1504 9654 1532 10202
rect 1492 9648 1544 9654
rect 1492 9590 1544 9596
rect 1596 9518 1624 10934
rect 1688 10266 1716 11319
rect 1780 10470 1808 11478
rect 1768 10464 1820 10470
rect 1768 10406 1820 10412
rect 1676 10260 1728 10266
rect 1676 10202 1728 10208
rect 1674 9888 1730 9897
rect 1674 9823 1730 9832
rect 1584 9512 1636 9518
rect 1490 9480 1546 9489
rect 1584 9454 1636 9460
rect 1490 9415 1546 9424
rect 1400 9036 1452 9042
rect 1400 8978 1452 8984
rect 1504 8906 1532 9415
rect 1582 9344 1638 9353
rect 1582 9279 1638 9288
rect 1492 8900 1544 8906
rect 1492 8842 1544 8848
rect 1398 8800 1454 8809
rect 1398 8735 1454 8744
rect 1412 8401 1440 8735
rect 1492 8492 1544 8498
rect 1492 8434 1544 8440
rect 1398 8392 1454 8401
rect 1398 8327 1454 8336
rect 1504 7993 1532 8434
rect 1490 7984 1546 7993
rect 1490 7919 1546 7928
rect 1596 7834 1624 9279
rect 1412 7806 1624 7834
rect 1308 7472 1360 7478
rect 1308 7414 1360 7420
rect 1308 7200 1360 7206
rect 1308 7142 1360 7148
rect 1216 6452 1268 6458
rect 1216 6394 1268 6400
rect 1214 6352 1270 6361
rect 1214 6287 1270 6296
rect 952 2746 1164 2774
rect 952 2310 980 2746
rect 1228 2514 1256 6287
rect 1320 5778 1348 7142
rect 1308 5772 1360 5778
rect 1308 5714 1360 5720
rect 1306 4720 1362 4729
rect 1306 4655 1362 4664
rect 1320 2582 1348 4655
rect 1308 2576 1360 2582
rect 1308 2518 1360 2524
rect 1216 2508 1268 2514
rect 1216 2450 1268 2456
rect 940 2304 992 2310
rect 940 2246 992 2252
rect 1412 2106 1440 7806
rect 1490 7576 1546 7585
rect 1490 7511 1546 7520
rect 1504 7410 1532 7511
rect 1492 7404 1544 7410
rect 1492 7346 1544 7352
rect 1584 7336 1636 7342
rect 1584 7278 1636 7284
rect 1492 6860 1544 6866
rect 1492 6802 1544 6808
rect 1504 6322 1532 6802
rect 1492 6316 1544 6322
rect 1492 6258 1544 6264
rect 1492 6112 1544 6118
rect 1492 6054 1544 6060
rect 1504 5914 1532 6054
rect 1492 5908 1544 5914
rect 1492 5850 1544 5856
rect 1596 5710 1624 7278
rect 1584 5704 1636 5710
rect 1584 5646 1636 5652
rect 1584 5568 1636 5574
rect 1584 5510 1636 5516
rect 1490 5400 1546 5409
rect 1490 5335 1546 5344
rect 1504 5302 1532 5335
rect 1492 5296 1544 5302
rect 1492 5238 1544 5244
rect 1596 4622 1624 5510
rect 1688 5352 1716 9823
rect 1872 9602 1900 12158
rect 1964 9654 1992 12294
rect 2044 12096 2096 12102
rect 2044 12038 2096 12044
rect 1780 9574 1900 9602
rect 1952 9648 2004 9654
rect 1952 9590 2004 9596
rect 1780 9178 1808 9574
rect 1860 9512 1912 9518
rect 2056 9466 2084 12038
rect 2148 10062 2176 12310
rect 2240 11354 2268 12310
rect 2332 11762 2360 12718
rect 2320 11756 2372 11762
rect 2320 11698 2372 11704
rect 2332 11665 2360 11698
rect 2318 11656 2374 11665
rect 2318 11591 2374 11600
rect 2228 11348 2280 11354
rect 2228 11290 2280 11296
rect 2226 11112 2282 11121
rect 2424 11082 2452 13670
rect 2594 13560 2650 13569
rect 2594 13495 2650 13504
rect 2608 13326 2636 13495
rect 2596 13320 2648 13326
rect 2596 13262 2648 13268
rect 2504 12844 2556 12850
rect 2504 12786 2556 12792
rect 2516 11132 2544 12786
rect 2594 12744 2650 12753
rect 2594 12679 2650 12688
rect 2608 11393 2636 12679
rect 2700 11898 2728 13926
rect 2792 13716 2820 16186
rect 2884 16028 2912 17734
rect 2964 17672 3016 17678
rect 2964 17614 3016 17620
rect 2976 16794 3004 17614
rect 3056 17536 3108 17542
rect 3056 17478 3108 17484
rect 2964 16788 3016 16794
rect 2964 16730 3016 16736
rect 2964 16040 3016 16046
rect 2884 16000 2964 16028
rect 2884 13870 2912 16000
rect 3068 16017 3096 17478
rect 2964 15982 3016 15988
rect 3054 16008 3110 16017
rect 3054 15943 3110 15952
rect 3160 15638 3188 18362
rect 3252 16522 3280 18686
rect 3332 18624 3384 18630
rect 3332 18566 3384 18572
rect 3344 17134 3372 18566
rect 4066 18320 4122 18329
rect 4066 18255 4122 18264
rect 4080 18222 4108 18255
rect 4172 18222 4200 20538
rect 4264 19378 4292 20878
rect 4448 20874 4476 21247
rect 4540 21146 4568 21626
rect 4632 21185 4660 21791
rect 4618 21176 4674 21185
rect 4528 21140 4580 21146
rect 4618 21111 4674 21120
rect 4528 21082 4580 21088
rect 4342 20839 4398 20848
rect 4436 20868 4488 20874
rect 4356 20602 4384 20839
rect 4436 20810 4488 20816
rect 4528 20800 4580 20806
rect 4528 20742 4580 20748
rect 4540 20602 4568 20742
rect 4344 20596 4396 20602
rect 4344 20538 4396 20544
rect 4528 20596 4580 20602
rect 4528 20538 4580 20544
rect 4436 20460 4488 20466
rect 4436 20402 4488 20408
rect 4528 20460 4580 20466
rect 4528 20402 4580 20408
rect 4448 20058 4476 20402
rect 4436 20052 4488 20058
rect 4436 19994 4488 20000
rect 4540 19922 4568 20402
rect 4528 19916 4580 19922
rect 4528 19858 4580 19864
rect 4436 19848 4488 19854
rect 4632 19802 4660 21111
rect 4488 19796 4660 19802
rect 4436 19790 4660 19796
rect 4448 19774 4660 19790
rect 4632 19553 4660 19774
rect 4618 19544 4674 19553
rect 4618 19479 4674 19488
rect 4436 19440 4488 19446
rect 4436 19382 4488 19388
rect 4252 19372 4304 19378
rect 4252 19314 4304 19320
rect 4344 19236 4396 19242
rect 4344 19178 4396 19184
rect 3424 18216 3476 18222
rect 3424 18158 3476 18164
rect 4068 18216 4120 18222
rect 4068 18158 4120 18164
rect 4160 18216 4212 18222
rect 4160 18158 4212 18164
rect 3436 17626 3464 18158
rect 3884 18148 3936 18154
rect 3884 18090 3936 18096
rect 3549 17980 3857 17989
rect 3549 17978 3555 17980
rect 3611 17978 3635 17980
rect 3691 17978 3715 17980
rect 3771 17978 3795 17980
rect 3851 17978 3857 17980
rect 3611 17926 3613 17978
rect 3793 17926 3795 17978
rect 3549 17924 3555 17926
rect 3611 17924 3635 17926
rect 3691 17924 3715 17926
rect 3771 17924 3795 17926
rect 3851 17924 3857 17926
rect 3549 17915 3857 17924
rect 3700 17672 3752 17678
rect 3514 17640 3570 17649
rect 3436 17598 3514 17626
rect 3700 17614 3752 17620
rect 3514 17575 3570 17584
rect 3712 17270 3740 17614
rect 3896 17338 3924 18090
rect 3976 18080 4028 18086
rect 4080 18068 4108 18158
rect 4080 18040 4200 18068
rect 3976 18022 4028 18028
rect 3988 17338 4016 18022
rect 4066 17912 4122 17921
rect 4066 17847 4122 17856
rect 4080 17746 4108 17847
rect 4068 17740 4120 17746
rect 4068 17682 4120 17688
rect 4172 17377 4200 18040
rect 4356 17785 4384 19178
rect 4342 17776 4398 17785
rect 4342 17711 4398 17720
rect 4252 17672 4304 17678
rect 4252 17614 4304 17620
rect 4158 17368 4214 17377
rect 3884 17332 3936 17338
rect 3884 17274 3936 17280
rect 3976 17332 4028 17338
rect 4158 17303 4214 17312
rect 3976 17274 4028 17280
rect 3700 17264 3752 17270
rect 3700 17206 3752 17212
rect 3804 17156 4108 17184
rect 3332 17128 3384 17134
rect 3332 17070 3384 17076
rect 3804 17066 3832 17156
rect 4080 17105 4108 17156
rect 3882 17096 3938 17105
rect 3792 17060 3844 17066
rect 3882 17031 3938 17040
rect 4066 17096 4122 17105
rect 4066 17031 4122 17040
rect 3792 17002 3844 17008
rect 3424 16992 3476 16998
rect 3424 16934 3476 16940
rect 3436 16833 3464 16934
rect 3549 16892 3857 16901
rect 3549 16890 3555 16892
rect 3611 16890 3635 16892
rect 3691 16890 3715 16892
rect 3771 16890 3795 16892
rect 3851 16890 3857 16892
rect 3611 16838 3613 16890
rect 3793 16838 3795 16890
rect 3549 16836 3555 16838
rect 3611 16836 3635 16838
rect 3691 16836 3715 16838
rect 3771 16836 3795 16838
rect 3851 16836 3857 16838
rect 3422 16824 3478 16833
rect 3549 16827 3857 16836
rect 3422 16759 3478 16768
rect 3608 16788 3660 16794
rect 3896 16776 3924 17031
rect 3976 16992 4028 16998
rect 3976 16934 4028 16940
rect 4068 16992 4120 16998
rect 4068 16934 4120 16940
rect 3608 16730 3660 16736
rect 3804 16748 3924 16776
rect 3620 16697 3648 16730
rect 3606 16688 3662 16697
rect 3606 16623 3662 16632
rect 3240 16516 3292 16522
rect 3240 16458 3292 16464
rect 3332 16516 3384 16522
rect 3332 16458 3384 16464
rect 3344 15688 3372 16458
rect 3424 16108 3476 16114
rect 3424 16050 3476 16056
rect 3252 15660 3372 15688
rect 3148 15632 3200 15638
rect 3148 15574 3200 15580
rect 3056 15360 3108 15366
rect 3056 15302 3108 15308
rect 2964 14952 3016 14958
rect 2964 14894 3016 14900
rect 2872 13864 2924 13870
rect 2872 13806 2924 13812
rect 2872 13728 2924 13734
rect 2792 13696 2872 13716
rect 2924 13696 2926 13705
rect 2792 13688 2870 13696
rect 2870 13631 2926 13640
rect 2976 13326 3004 14894
rect 3068 14113 3096 15302
rect 3148 15156 3200 15162
rect 3148 15098 3200 15104
rect 3054 14104 3110 14113
rect 3054 14039 3110 14048
rect 3056 13864 3108 13870
rect 3056 13806 3108 13812
rect 3068 13512 3096 13806
rect 3160 13580 3188 15098
rect 3252 14385 3280 15660
rect 3436 14482 3464 16050
rect 3804 15910 3832 16748
rect 3988 16658 4016 16934
rect 3976 16652 4028 16658
rect 3976 16594 4028 16600
rect 3976 16448 4028 16454
rect 3974 16416 3976 16425
rect 4028 16416 4030 16425
rect 3974 16351 4030 16360
rect 4080 16232 4108 16934
rect 4264 16232 4292 17614
rect 4356 17066 4384 17711
rect 4344 17060 4396 17066
rect 4344 17002 4396 17008
rect 4344 16584 4396 16590
rect 4344 16526 4396 16532
rect 3988 16204 4108 16232
rect 4172 16204 4292 16232
rect 3792 15904 3844 15910
rect 3792 15846 3844 15852
rect 3884 15904 3936 15910
rect 3884 15846 3936 15852
rect 3549 15804 3857 15813
rect 3549 15802 3555 15804
rect 3611 15802 3635 15804
rect 3691 15802 3715 15804
rect 3771 15802 3795 15804
rect 3851 15802 3857 15804
rect 3611 15750 3613 15802
rect 3793 15750 3795 15802
rect 3549 15748 3555 15750
rect 3611 15748 3635 15750
rect 3691 15748 3715 15750
rect 3771 15748 3795 15750
rect 3851 15748 3857 15750
rect 3549 15739 3857 15748
rect 3549 14716 3857 14725
rect 3549 14714 3555 14716
rect 3611 14714 3635 14716
rect 3691 14714 3715 14716
rect 3771 14714 3795 14716
rect 3851 14714 3857 14716
rect 3611 14662 3613 14714
rect 3793 14662 3795 14714
rect 3549 14660 3555 14662
rect 3611 14660 3635 14662
rect 3691 14660 3715 14662
rect 3771 14660 3795 14662
rect 3851 14660 3857 14662
rect 3549 14651 3857 14660
rect 3896 14521 3924 15846
rect 3988 15638 4016 16204
rect 3976 15632 4028 15638
rect 3976 15574 4028 15580
rect 4172 15570 4200 16204
rect 4252 16108 4304 16114
rect 4252 16050 4304 16056
rect 4264 15706 4292 16050
rect 4356 15706 4384 16526
rect 4252 15700 4304 15706
rect 4252 15642 4304 15648
rect 4344 15700 4396 15706
rect 4344 15642 4396 15648
rect 4160 15564 4212 15570
rect 4160 15506 4212 15512
rect 4344 15564 4396 15570
rect 4344 15506 4396 15512
rect 4172 15450 4200 15506
rect 3988 15422 4200 15450
rect 4252 15496 4304 15502
rect 4252 15438 4304 15444
rect 3988 15026 4016 15422
rect 4068 15360 4120 15366
rect 4068 15302 4120 15308
rect 3976 15020 4028 15026
rect 3976 14962 4028 14968
rect 3976 14816 4028 14822
rect 3976 14758 4028 14764
rect 3882 14512 3938 14521
rect 3424 14476 3476 14482
rect 3424 14418 3476 14424
rect 3608 14476 3660 14482
rect 3882 14447 3938 14456
rect 3608 14418 3660 14424
rect 3238 14376 3294 14385
rect 3238 14311 3294 14320
rect 3240 14272 3292 14278
rect 3620 14226 3648 14418
rect 3240 14214 3292 14220
rect 3252 13938 3280 14214
rect 3528 14198 3648 14226
rect 3882 14240 3938 14249
rect 3240 13932 3292 13938
rect 3424 13932 3476 13938
rect 3240 13874 3292 13880
rect 3344 13892 3424 13920
rect 3240 13728 3292 13734
rect 3344 13716 3372 13892
rect 3424 13874 3476 13880
rect 3528 13716 3556 14198
rect 3882 14175 3938 14184
rect 3292 13688 3372 13716
rect 3436 13688 3556 13716
rect 3240 13670 3292 13676
rect 3160 13552 3372 13580
rect 3068 13484 3280 13512
rect 2964 13320 3016 13326
rect 2964 13262 3016 13268
rect 2870 13152 2926 13161
rect 2870 13087 2926 13096
rect 2778 12880 2834 12889
rect 2778 12815 2834 12824
rect 2688 11892 2740 11898
rect 2688 11834 2740 11840
rect 2686 11656 2742 11665
rect 2686 11591 2742 11600
rect 2594 11384 2650 11393
rect 2594 11319 2650 11328
rect 2516 11104 2602 11132
rect 2700 11121 2728 11591
rect 2226 11047 2282 11056
rect 2412 11076 2464 11082
rect 2136 10056 2188 10062
rect 2136 9998 2188 10004
rect 2240 10010 2268 11047
rect 2412 11018 2464 11024
rect 2574 10996 2602 11104
rect 2686 11112 2742 11121
rect 2686 11047 2742 11056
rect 2516 10968 2602 10996
rect 2412 10600 2464 10606
rect 2412 10542 2464 10548
rect 2240 9982 2360 10010
rect 2136 9920 2188 9926
rect 2136 9862 2188 9868
rect 1860 9454 1912 9460
rect 1768 9172 1820 9178
rect 1768 9114 1820 9120
rect 1766 8664 1822 8673
rect 1766 8599 1822 8608
rect 1780 7426 1808 8599
rect 1872 7546 1900 9454
rect 1964 9438 2084 9466
rect 1860 7540 1912 7546
rect 1860 7482 1912 7488
rect 1780 7398 1900 7426
rect 1766 7032 1822 7041
rect 1766 6967 1822 6976
rect 1780 5522 1808 6967
rect 1872 6610 1900 7398
rect 1964 6798 1992 9438
rect 2148 9042 2176 9862
rect 2226 9752 2282 9761
rect 2226 9687 2282 9696
rect 2240 9586 2268 9687
rect 2228 9580 2280 9586
rect 2228 9522 2280 9528
rect 2332 9466 2360 9982
rect 2240 9438 2360 9466
rect 2136 9036 2188 9042
rect 2136 8978 2188 8984
rect 2134 7848 2190 7857
rect 2134 7783 2190 7792
rect 2044 7744 2096 7750
rect 2044 7686 2096 7692
rect 1952 6792 2004 6798
rect 1952 6734 2004 6740
rect 1872 6582 1992 6610
rect 1780 5494 1900 5522
rect 1768 5364 1820 5370
rect 1688 5324 1768 5352
rect 1768 5306 1820 5312
rect 1872 5250 1900 5494
rect 1780 5222 1900 5250
rect 1584 4616 1636 4622
rect 1584 4558 1636 4564
rect 1584 4072 1636 4078
rect 1584 4014 1636 4020
rect 1596 3602 1624 4014
rect 1584 3596 1636 3602
rect 1584 3538 1636 3544
rect 1490 3360 1546 3369
rect 1490 3295 1546 3304
rect 1400 2100 1452 2106
rect 1400 2042 1452 2048
rect 1504 2038 1532 3295
rect 1596 3194 1624 3538
rect 1584 3188 1636 3194
rect 1584 3130 1636 3136
rect 1780 2774 1808 5222
rect 1858 5128 1914 5137
rect 1858 5063 1914 5072
rect 1872 4622 1900 5063
rect 1964 5030 1992 6582
rect 2056 5370 2084 7686
rect 2044 5364 2096 5370
rect 2044 5306 2096 5312
rect 2148 5250 2176 7783
rect 2240 7342 2268 9438
rect 2424 8498 2452 10542
rect 2516 9586 2544 10968
rect 2686 10840 2742 10849
rect 2686 10775 2742 10784
rect 2700 10606 2728 10775
rect 2688 10600 2740 10606
rect 2688 10542 2740 10548
rect 2504 9580 2556 9586
rect 2504 9522 2556 9528
rect 2504 9444 2556 9450
rect 2504 9386 2556 9392
rect 2516 9353 2544 9386
rect 2502 9344 2558 9353
rect 2502 9279 2558 9288
rect 2504 8968 2556 8974
rect 2504 8910 2556 8916
rect 2412 8492 2464 8498
rect 2412 8434 2464 8440
rect 2410 8120 2466 8129
rect 2410 8055 2466 8064
rect 2228 7336 2280 7342
rect 2228 7278 2280 7284
rect 2320 7200 2372 7206
rect 2226 7168 2282 7177
rect 2320 7142 2372 7148
rect 2226 7103 2282 7112
rect 2056 5222 2176 5250
rect 1952 5024 2004 5030
rect 1952 4966 2004 4972
rect 1860 4616 1912 4622
rect 1860 4558 1912 4564
rect 1952 4208 2004 4214
rect 1952 4150 2004 4156
rect 1596 2746 1808 2774
rect 1492 2032 1544 2038
rect 1492 1974 1544 1980
rect 1596 1562 1624 2746
rect 1964 2038 1992 4150
rect 2056 4128 2084 5222
rect 2136 5160 2188 5166
rect 2136 5102 2188 5108
rect 2148 4690 2176 5102
rect 2136 4684 2188 4690
rect 2136 4626 2188 4632
rect 2240 4146 2268 7103
rect 2332 5778 2360 7142
rect 2424 6225 2452 8055
rect 2516 7886 2544 8910
rect 2700 8906 2728 10542
rect 2792 10266 2820 12815
rect 2884 12356 2912 13087
rect 3054 12880 3110 12889
rect 3252 12850 3280 13484
rect 3344 12968 3372 13552
rect 3436 13530 3464 13688
rect 3549 13628 3857 13637
rect 3549 13626 3555 13628
rect 3611 13626 3635 13628
rect 3691 13626 3715 13628
rect 3771 13626 3795 13628
rect 3851 13626 3857 13628
rect 3611 13574 3613 13626
rect 3793 13574 3795 13626
rect 3549 13572 3555 13574
rect 3611 13572 3635 13574
rect 3691 13572 3715 13574
rect 3771 13572 3795 13574
rect 3851 13572 3857 13574
rect 3549 13563 3857 13572
rect 3424 13524 3476 13530
rect 3896 13512 3924 14175
rect 3424 13466 3476 13472
rect 3712 13484 3924 13512
rect 3344 12940 3648 12968
rect 3054 12815 3110 12824
rect 3240 12844 3292 12850
rect 2964 12708 3016 12714
rect 2964 12650 3016 12656
rect 2976 12424 3004 12650
rect 3068 12617 3096 12815
rect 3516 12844 3568 12850
rect 3240 12786 3292 12792
rect 3344 12804 3516 12832
rect 3054 12608 3110 12617
rect 3054 12543 3110 12552
rect 2976 12396 3096 12424
rect 2884 12328 3004 12356
rect 2872 11756 2924 11762
rect 2872 11698 2924 11704
rect 2884 11014 2912 11698
rect 2872 11008 2924 11014
rect 2872 10950 2924 10956
rect 2872 10600 2924 10606
rect 2872 10542 2924 10548
rect 2780 10260 2832 10266
rect 2780 10202 2832 10208
rect 2778 10160 2834 10169
rect 2778 10095 2834 10104
rect 2688 8900 2740 8906
rect 2688 8842 2740 8848
rect 2700 8498 2728 8842
rect 2688 8492 2740 8498
rect 2688 8434 2740 8440
rect 2504 7880 2556 7886
rect 2504 7822 2556 7828
rect 2688 7880 2740 7886
rect 2688 7822 2740 7828
rect 2596 7268 2648 7274
rect 2596 7210 2648 7216
rect 2608 6848 2636 7210
rect 2700 7018 2728 7822
rect 2792 7154 2820 10095
rect 2884 9926 2912 10542
rect 2872 9920 2924 9926
rect 2872 9862 2924 9868
rect 2884 9450 2912 9862
rect 2872 9444 2924 9450
rect 2872 9386 2924 9392
rect 2884 8430 2912 9386
rect 2976 8634 3004 12328
rect 3068 11694 3096 12396
rect 3252 12102 3280 12786
rect 3240 12096 3292 12102
rect 3240 12038 3292 12044
rect 3056 11688 3108 11694
rect 3056 11630 3108 11636
rect 3240 11688 3292 11694
rect 3240 11630 3292 11636
rect 3056 11552 3108 11558
rect 3056 11494 3108 11500
rect 3068 11082 3096 11494
rect 3056 11076 3108 11082
rect 3056 11018 3108 11024
rect 3056 10532 3108 10538
rect 3108 10492 3188 10520
rect 3056 10474 3108 10480
rect 3054 10296 3110 10305
rect 3054 10231 3110 10240
rect 3068 10198 3096 10231
rect 3056 10192 3108 10198
rect 3056 10134 3108 10140
rect 3056 10056 3108 10062
rect 3056 9998 3108 10004
rect 3068 9722 3096 9998
rect 3056 9716 3108 9722
rect 3056 9658 3108 9664
rect 3056 9444 3108 9450
rect 3056 9386 3108 9392
rect 2964 8628 3016 8634
rect 2964 8570 3016 8576
rect 2872 8424 2924 8430
rect 2872 8366 2924 8372
rect 2964 8356 3016 8362
rect 2964 8298 3016 8304
rect 2872 7744 2924 7750
rect 2872 7686 2924 7692
rect 2884 7313 2912 7686
rect 2870 7304 2926 7313
rect 2870 7239 2926 7248
rect 2792 7126 2912 7154
rect 2700 6990 2820 7018
rect 2606 6820 2636 6848
rect 2502 6760 2558 6769
rect 2502 6695 2558 6704
rect 2606 6712 2634 6820
rect 2516 6662 2544 6695
rect 2606 6684 2636 6712
rect 2504 6656 2556 6662
rect 2504 6598 2556 6604
rect 2502 6352 2558 6361
rect 2502 6287 2558 6296
rect 2410 6216 2466 6225
rect 2410 6151 2466 6160
rect 2320 5772 2372 5778
rect 2320 5714 2372 5720
rect 2412 5772 2464 5778
rect 2412 5714 2464 5720
rect 2320 5364 2372 5370
rect 2320 5306 2372 5312
rect 2228 4140 2280 4146
rect 2056 4100 2176 4128
rect 2042 3224 2098 3233
rect 2042 3159 2098 3168
rect 2056 2446 2084 3159
rect 2148 2774 2176 4100
rect 2228 4082 2280 4088
rect 2332 3058 2360 5306
rect 2424 3670 2452 5714
rect 2516 5681 2544 6287
rect 2502 5672 2558 5681
rect 2502 5607 2558 5616
rect 2504 5024 2556 5030
rect 2504 4966 2556 4972
rect 2516 4622 2544 4966
rect 2504 4616 2556 4622
rect 2504 4558 2556 4564
rect 2412 3664 2464 3670
rect 2412 3606 2464 3612
rect 2608 3194 2636 6684
rect 2792 6610 2820 6990
rect 2700 6582 2820 6610
rect 2700 5370 2728 6582
rect 2778 6216 2834 6225
rect 2778 6151 2834 6160
rect 2688 5364 2740 5370
rect 2688 5306 2740 5312
rect 2686 4584 2742 4593
rect 2686 4519 2742 4528
rect 2700 4282 2728 4519
rect 2688 4276 2740 4282
rect 2688 4218 2740 4224
rect 2596 3188 2648 3194
rect 2596 3130 2648 3136
rect 2504 3120 2556 3126
rect 2504 3062 2556 3068
rect 2320 3052 2372 3058
rect 2320 2994 2372 3000
rect 2148 2746 2360 2774
rect 2332 2650 2360 2746
rect 2320 2644 2372 2650
rect 2320 2586 2372 2592
rect 2044 2440 2096 2446
rect 2044 2382 2096 2388
rect 1952 2032 2004 2038
rect 1952 1974 2004 1980
rect 2516 1970 2544 3062
rect 2596 2984 2648 2990
rect 2596 2926 2648 2932
rect 2608 2446 2636 2926
rect 2792 2802 2820 6151
rect 2884 6118 2912 7126
rect 2872 6112 2924 6118
rect 2872 6054 2924 6060
rect 2976 5794 3004 8298
rect 2884 5766 3004 5794
rect 2884 3738 2912 5766
rect 2964 5704 3016 5710
rect 2964 5646 3016 5652
rect 2872 3732 2924 3738
rect 2872 3674 2924 3680
rect 2870 3360 2926 3369
rect 2870 3295 2926 3304
rect 2884 2990 2912 3295
rect 2976 2990 3004 5646
rect 3068 5370 3096 9386
rect 3160 6458 3188 10492
rect 3252 8090 3280 11630
rect 3344 10266 3372 12804
rect 3516 12786 3568 12792
rect 3620 12628 3648 12940
rect 3712 12782 3740 13484
rect 3884 13388 3936 13394
rect 3884 13330 3936 13336
rect 3792 13320 3844 13326
rect 3790 13288 3792 13297
rect 3844 13288 3846 13297
rect 3790 13223 3846 13232
rect 3700 12776 3752 12782
rect 3700 12718 3752 12724
rect 3436 12600 3648 12628
rect 3436 12186 3464 12600
rect 3549 12540 3857 12549
rect 3549 12538 3555 12540
rect 3611 12538 3635 12540
rect 3691 12538 3715 12540
rect 3771 12538 3795 12540
rect 3851 12538 3857 12540
rect 3611 12486 3613 12538
rect 3793 12486 3795 12538
rect 3549 12484 3555 12486
rect 3611 12484 3635 12486
rect 3691 12484 3715 12486
rect 3771 12484 3795 12486
rect 3851 12484 3857 12486
rect 3549 12475 3857 12484
rect 3896 12442 3924 13330
rect 3988 13326 4016 14758
rect 3976 13320 4028 13326
rect 3976 13262 4028 13268
rect 3988 12617 4016 13262
rect 3974 12608 4030 12617
rect 3974 12543 4030 12552
rect 3884 12436 3936 12442
rect 3884 12378 3936 12384
rect 3976 12436 4028 12442
rect 3976 12378 4028 12384
rect 3988 12345 4016 12378
rect 4080 12374 4108 15302
rect 4160 15020 4212 15026
rect 4160 14962 4212 14968
rect 4172 14074 4200 14962
rect 4264 14822 4292 15438
rect 4252 14816 4304 14822
rect 4252 14758 4304 14764
rect 4250 14648 4306 14657
rect 4356 14618 4384 15506
rect 4448 15314 4476 19382
rect 4620 19168 4672 19174
rect 4620 19110 4672 19116
rect 4528 18964 4580 18970
rect 4528 18906 4580 18912
rect 4540 16833 4568 18906
rect 4632 18698 4660 19110
rect 4620 18692 4672 18698
rect 4620 18634 4672 18640
rect 4724 17678 4752 22630
rect 5000 22420 5028 22986
rect 5078 22944 5134 22953
rect 5078 22879 5134 22888
rect 5092 22574 5120 22879
rect 5080 22568 5132 22574
rect 5080 22510 5132 22516
rect 5000 22392 5120 22420
rect 4804 22160 4856 22166
rect 4804 22102 4856 22108
rect 4816 19242 4844 22102
rect 4896 22092 4948 22098
rect 4896 22034 4948 22040
rect 4908 21554 4936 22034
rect 4988 22024 5040 22030
rect 4988 21966 5040 21972
rect 5000 21894 5028 21966
rect 4988 21888 5040 21894
rect 4988 21830 5040 21836
rect 4896 21548 4948 21554
rect 4896 21490 4948 21496
rect 4896 20800 4948 20806
rect 4896 20742 4948 20748
rect 4804 19236 4856 19242
rect 4804 19178 4856 19184
rect 4804 18692 4856 18698
rect 4804 18634 4856 18640
rect 4816 18442 4844 18634
rect 4908 18630 4936 20742
rect 5000 19718 5028 21830
rect 4988 19712 5040 19718
rect 4988 19654 5040 19660
rect 4896 18624 4948 18630
rect 4896 18566 4948 18572
rect 4816 18414 5028 18442
rect 5000 18290 5028 18414
rect 4988 18284 5040 18290
rect 4988 18226 5040 18232
rect 4804 18216 4856 18222
rect 4856 18176 4936 18204
rect 4804 18158 4856 18164
rect 4804 18080 4856 18086
rect 4804 18022 4856 18028
rect 4712 17672 4764 17678
rect 4712 17614 4764 17620
rect 4620 17536 4672 17542
rect 4620 17478 4672 17484
rect 4526 16824 4582 16833
rect 4526 16759 4582 16768
rect 4528 16516 4580 16522
rect 4528 16458 4580 16464
rect 4540 15638 4568 16458
rect 4528 15632 4580 15638
rect 4526 15600 4528 15609
rect 4580 15600 4582 15609
rect 4526 15535 4582 15544
rect 4632 15337 4660 17478
rect 4712 17128 4764 17134
rect 4712 17070 4764 17076
rect 4724 16522 4752 17070
rect 4712 16516 4764 16522
rect 4712 16458 4764 16464
rect 4710 16144 4766 16153
rect 4710 16079 4766 16088
rect 4618 15328 4674 15337
rect 4448 15286 4568 15314
rect 4434 14784 4490 14793
rect 4434 14719 4490 14728
rect 4250 14583 4306 14592
rect 4344 14612 4396 14618
rect 4264 14550 4292 14583
rect 4344 14554 4396 14560
rect 4252 14544 4304 14550
rect 4252 14486 4304 14492
rect 4344 14340 4396 14346
rect 4344 14282 4396 14288
rect 4160 14068 4212 14074
rect 4160 14010 4212 14016
rect 4356 13870 4384 14282
rect 4448 14074 4476 14719
rect 4436 14068 4488 14074
rect 4436 14010 4488 14016
rect 4436 13932 4488 13938
rect 4436 13874 4488 13880
rect 4344 13864 4396 13870
rect 4344 13806 4396 13812
rect 4252 13796 4304 13802
rect 4252 13738 4304 13744
rect 4160 13524 4212 13530
rect 4160 13466 4212 13472
rect 4068 12368 4120 12374
rect 3974 12336 4030 12345
rect 4068 12310 4120 12316
rect 3974 12271 4030 12280
rect 4172 12186 4200 13466
rect 4264 12374 4292 13738
rect 4252 12368 4304 12374
rect 4252 12310 4304 12316
rect 3436 12158 3556 12186
rect 3424 12096 3476 12102
rect 3424 12038 3476 12044
rect 3436 11354 3464 12038
rect 3528 11762 3556 12158
rect 3884 12164 3936 12170
rect 4172 12158 4292 12186
rect 3884 12106 3936 12112
rect 3516 11756 3568 11762
rect 3516 11698 3568 11704
rect 3549 11452 3857 11461
rect 3549 11450 3555 11452
rect 3611 11450 3635 11452
rect 3691 11450 3715 11452
rect 3771 11450 3795 11452
rect 3851 11450 3857 11452
rect 3611 11398 3613 11450
rect 3793 11398 3795 11450
rect 3549 11396 3555 11398
rect 3611 11396 3635 11398
rect 3691 11396 3715 11398
rect 3771 11396 3795 11398
rect 3851 11396 3857 11398
rect 3549 11387 3857 11396
rect 3424 11348 3476 11354
rect 3424 11290 3476 11296
rect 3608 11348 3660 11354
rect 3608 11290 3660 11296
rect 3516 10668 3568 10674
rect 3516 10610 3568 10616
rect 3528 10520 3556 10610
rect 3436 10492 3556 10520
rect 3332 10260 3384 10266
rect 3332 10202 3384 10208
rect 3330 9616 3386 9625
rect 3330 9551 3386 9560
rect 3344 8650 3372 9551
rect 3436 8974 3464 10492
rect 3620 10470 3648 11290
rect 3896 11257 3924 12106
rect 4066 12064 4122 12073
rect 4066 11999 4122 12008
rect 3976 11756 4028 11762
rect 3976 11698 4028 11704
rect 3988 11354 4016 11698
rect 4080 11354 4108 11999
rect 4158 11928 4214 11937
rect 4158 11863 4214 11872
rect 3976 11348 4028 11354
rect 3976 11290 4028 11296
rect 4068 11348 4120 11354
rect 4068 11290 4120 11296
rect 3882 11248 3938 11257
rect 4172 11200 4200 11863
rect 4264 11218 4292 12158
rect 3882 11183 3938 11192
rect 3988 11172 4200 11200
rect 4252 11212 4304 11218
rect 3792 11076 3844 11082
rect 3792 11018 3844 11024
rect 3804 10810 3832 11018
rect 3792 10804 3844 10810
rect 3988 10792 4016 11172
rect 4252 11154 4304 11160
rect 4160 11076 4212 11082
rect 4160 11018 4212 11024
rect 4252 11076 4304 11082
rect 4252 11018 4304 11024
rect 4066 10976 4122 10985
rect 4066 10911 4122 10920
rect 3792 10746 3844 10752
rect 3896 10764 4016 10792
rect 3896 10606 3924 10764
rect 3974 10704 4030 10713
rect 3974 10639 4030 10648
rect 3884 10600 3936 10606
rect 3884 10542 3936 10548
rect 3608 10464 3660 10470
rect 3608 10406 3660 10412
rect 3549 10364 3857 10373
rect 3549 10362 3555 10364
rect 3611 10362 3635 10364
rect 3691 10362 3715 10364
rect 3771 10362 3795 10364
rect 3851 10362 3857 10364
rect 3611 10310 3613 10362
rect 3793 10310 3795 10362
rect 3549 10308 3555 10310
rect 3611 10308 3635 10310
rect 3691 10308 3715 10310
rect 3771 10308 3795 10310
rect 3851 10308 3857 10310
rect 3549 10299 3857 10308
rect 3896 10248 3924 10542
rect 3988 10266 4016 10639
rect 3712 10220 3924 10248
rect 3976 10260 4028 10266
rect 3712 9602 3740 10220
rect 3976 10202 4028 10208
rect 3974 10160 4030 10169
rect 4080 10130 4108 10911
rect 4172 10713 4200 11018
rect 4158 10704 4214 10713
rect 4158 10639 4214 10648
rect 4160 10464 4212 10470
rect 4160 10406 4212 10412
rect 3974 10095 4030 10104
rect 4068 10124 4120 10130
rect 3988 10010 4016 10095
rect 4068 10066 4120 10072
rect 3884 9988 3936 9994
rect 3988 9982 4108 10010
rect 3884 9930 3936 9936
rect 3896 9761 3924 9930
rect 3882 9752 3938 9761
rect 3882 9687 3938 9696
rect 3516 9580 3568 9586
rect 3712 9574 3924 9602
rect 3712 9568 3740 9574
rect 3568 9540 3740 9568
rect 3516 9522 3568 9528
rect 3549 9276 3857 9285
rect 3549 9274 3555 9276
rect 3611 9274 3635 9276
rect 3691 9274 3715 9276
rect 3771 9274 3795 9276
rect 3851 9274 3857 9276
rect 3611 9222 3613 9274
rect 3793 9222 3795 9274
rect 3549 9220 3555 9222
rect 3611 9220 3635 9222
rect 3691 9220 3715 9222
rect 3771 9220 3795 9222
rect 3851 9220 3857 9222
rect 3549 9211 3857 9220
rect 3896 9160 3924 9574
rect 3976 9512 4028 9518
rect 3976 9454 4028 9460
rect 3988 9217 4016 9454
rect 4080 9450 4108 9982
rect 4068 9444 4120 9450
rect 4068 9386 4120 9392
rect 3528 9132 3924 9160
rect 3974 9208 4030 9217
rect 3974 9143 4030 9152
rect 4068 9172 4120 9178
rect 3424 8968 3476 8974
rect 3424 8910 3476 8916
rect 3528 8820 3556 9132
rect 4068 9114 4120 9120
rect 3792 9036 3844 9042
rect 3792 8978 3844 8984
rect 3608 8968 3660 8974
rect 3608 8910 3660 8916
rect 3326 8634 3372 8650
rect 3436 8792 3556 8820
rect 3326 8628 3384 8634
rect 3326 8588 3332 8628
rect 3332 8570 3384 8576
rect 3436 8498 3464 8792
rect 3424 8492 3476 8498
rect 3424 8434 3476 8440
rect 3516 8492 3568 8498
rect 3516 8434 3568 8440
rect 3528 8344 3556 8434
rect 3344 8316 3556 8344
rect 3344 8265 3372 8316
rect 3620 8276 3648 8910
rect 3804 8412 3832 8978
rect 4080 8974 4108 9114
rect 4172 8974 4200 10406
rect 4264 9382 4292 11018
rect 4356 10985 4384 13806
rect 4448 13512 4476 13874
rect 4540 13705 4568 15286
rect 4618 15263 4674 15272
rect 4620 14884 4672 14890
rect 4620 14826 4672 14832
rect 4632 14414 4660 14826
rect 4620 14408 4672 14414
rect 4620 14350 4672 14356
rect 4632 13802 4660 14350
rect 4724 14346 4752 16079
rect 4712 14340 4764 14346
rect 4712 14282 4764 14288
rect 4620 13796 4672 13802
rect 4620 13738 4672 13744
rect 4526 13696 4582 13705
rect 4526 13631 4582 13640
rect 4448 13484 4568 13512
rect 4434 13424 4490 13433
rect 4434 13359 4490 13368
rect 4448 11150 4476 13359
rect 4540 11898 4568 13484
rect 4712 13388 4764 13394
rect 4816 13376 4844 18022
rect 4908 17921 4936 18176
rect 4894 17912 4950 17921
rect 4894 17847 4950 17856
rect 4908 16658 4936 17847
rect 4988 17536 5040 17542
rect 4986 17504 4988 17513
rect 5040 17504 5042 17513
rect 4986 17439 5042 17448
rect 4988 17332 5040 17338
rect 4988 17274 5040 17280
rect 5000 17202 5028 17274
rect 4988 17196 5040 17202
rect 4988 17138 5040 17144
rect 4896 16652 4948 16658
rect 4896 16594 4948 16600
rect 4894 16416 4950 16425
rect 4894 16351 4950 16360
rect 4908 16182 4936 16351
rect 4896 16176 4948 16182
rect 4896 16118 4948 16124
rect 4988 16176 5040 16182
rect 4988 16118 5040 16124
rect 5000 16028 5028 16118
rect 4908 16000 5028 16028
rect 4908 15881 4936 16000
rect 4988 15904 5040 15910
rect 4894 15872 4950 15881
rect 4988 15846 5040 15852
rect 4894 15807 4950 15816
rect 4894 15736 4950 15745
rect 4894 15671 4950 15680
rect 4908 14822 4936 15671
rect 4896 14816 4948 14822
rect 4896 14758 4948 14764
rect 5000 13784 5028 15846
rect 5092 15570 5120 22392
rect 5184 20806 5212 23174
rect 5264 23112 5316 23118
rect 5264 23054 5316 23060
rect 5356 23112 5408 23118
rect 5356 23054 5408 23060
rect 5172 20800 5224 20806
rect 5172 20742 5224 20748
rect 5276 20346 5304 23054
rect 5368 22030 5396 23054
rect 5460 22982 5488 24806
rect 5448 22976 5500 22982
rect 5448 22918 5500 22924
rect 5446 22808 5502 22817
rect 5446 22743 5502 22752
rect 5460 22574 5488 22743
rect 5448 22568 5500 22574
rect 5448 22510 5500 22516
rect 5356 22024 5408 22030
rect 5408 21984 5488 22012
rect 5356 21966 5408 21972
rect 5356 21888 5408 21894
rect 5356 21830 5408 21836
rect 5368 20398 5396 21830
rect 5460 21010 5488 21984
rect 5552 21457 5580 25078
rect 5724 24676 5776 24682
rect 5724 24618 5776 24624
rect 5632 24608 5684 24614
rect 5632 24550 5684 24556
rect 5644 24410 5672 24550
rect 5736 24410 5764 24618
rect 5828 24449 5856 30144
rect 5908 30048 5960 30054
rect 5908 29990 5960 29996
rect 5920 29714 5948 29990
rect 5908 29708 5960 29714
rect 5908 29650 5960 29656
rect 6012 29578 6040 31622
rect 6148 31580 6456 31589
rect 6148 31578 6154 31580
rect 6210 31578 6234 31580
rect 6290 31578 6314 31580
rect 6370 31578 6394 31580
rect 6450 31578 6456 31580
rect 6210 31526 6212 31578
rect 6392 31526 6394 31578
rect 6148 31524 6154 31526
rect 6210 31524 6234 31526
rect 6290 31524 6314 31526
rect 6370 31524 6394 31526
rect 6450 31524 6456 31526
rect 6148 31515 6456 31524
rect 6460 31476 6512 31482
rect 6460 31418 6512 31424
rect 6472 31346 6500 31418
rect 6460 31340 6512 31346
rect 6460 31282 6512 31288
rect 6366 31240 6422 31249
rect 6366 31175 6422 31184
rect 6092 31136 6144 31142
rect 6092 31078 6144 31084
rect 6104 30841 6132 31078
rect 6090 30832 6146 30841
rect 6090 30767 6146 30776
rect 6380 30666 6408 31175
rect 6368 30660 6420 30666
rect 6368 30602 6420 30608
rect 6564 30546 6592 32710
rect 6656 32348 6684 32728
rect 6736 32710 6788 32716
rect 6748 32502 6776 32710
rect 6736 32496 6788 32502
rect 6736 32438 6788 32444
rect 6840 32450 6868 34410
rect 7012 33992 7064 33998
rect 7012 33934 7064 33940
rect 7104 33992 7156 33998
rect 7104 33934 7156 33940
rect 6920 33856 6972 33862
rect 6920 33798 6972 33804
rect 6932 33318 6960 33798
rect 7024 33386 7052 33934
rect 7012 33380 7064 33386
rect 7012 33322 7064 33328
rect 6920 33312 6972 33318
rect 6920 33254 6972 33260
rect 6920 32904 6972 32910
rect 6920 32846 6972 32852
rect 6932 32570 6960 32846
rect 6920 32564 6972 32570
rect 6920 32506 6972 32512
rect 6840 32422 6960 32450
rect 6656 32320 6776 32348
rect 6644 32224 6696 32230
rect 6644 32166 6696 32172
rect 6656 30734 6684 32166
rect 6748 31414 6776 32320
rect 6826 32328 6882 32337
rect 6826 32263 6882 32272
rect 6736 31408 6788 31414
rect 6736 31350 6788 31356
rect 6840 31278 6868 32263
rect 6828 31272 6880 31278
rect 6828 31214 6880 31220
rect 6644 30728 6696 30734
rect 6644 30670 6696 30676
rect 6546 30518 6592 30546
rect 6148 30492 6456 30501
rect 6148 30490 6154 30492
rect 6210 30490 6234 30492
rect 6290 30490 6314 30492
rect 6370 30490 6394 30492
rect 6450 30490 6456 30492
rect 6210 30438 6212 30490
rect 6392 30438 6394 30490
rect 6148 30436 6154 30438
rect 6210 30436 6234 30438
rect 6290 30436 6314 30438
rect 6370 30436 6394 30438
rect 6450 30436 6456 30438
rect 6148 30427 6456 30436
rect 6092 30388 6144 30394
rect 6546 30376 6574 30518
rect 6092 30330 6144 30336
rect 6472 30348 6574 30376
rect 6104 30297 6132 30330
rect 6090 30288 6146 30297
rect 6090 30223 6146 30232
rect 6368 30184 6420 30190
rect 6368 30126 6420 30132
rect 6380 29889 6408 30126
rect 6366 29880 6422 29889
rect 6366 29815 6422 29824
rect 6000 29572 6052 29578
rect 6000 29514 6052 29520
rect 6472 29510 6500 30348
rect 6552 29572 6604 29578
rect 6552 29514 6604 29520
rect 5908 29504 5960 29510
rect 6460 29504 6512 29510
rect 5908 29446 5960 29452
rect 5998 29472 6054 29481
rect 5920 26217 5948 29446
rect 6460 29446 6512 29452
rect 5998 29407 6054 29416
rect 6012 29073 6040 29407
rect 6148 29404 6456 29413
rect 6148 29402 6154 29404
rect 6210 29402 6234 29404
rect 6290 29402 6314 29404
rect 6370 29402 6394 29404
rect 6450 29402 6456 29404
rect 6210 29350 6212 29402
rect 6392 29350 6394 29402
rect 6148 29348 6154 29350
rect 6210 29348 6234 29350
rect 6290 29348 6314 29350
rect 6370 29348 6394 29350
rect 6450 29348 6456 29350
rect 6148 29339 6456 29348
rect 5998 29064 6054 29073
rect 5998 28999 6054 29008
rect 6148 28316 6456 28325
rect 6148 28314 6154 28316
rect 6210 28314 6234 28316
rect 6290 28314 6314 28316
rect 6370 28314 6394 28316
rect 6450 28314 6456 28316
rect 6210 28262 6212 28314
rect 6392 28262 6394 28314
rect 6148 28260 6154 28262
rect 6210 28260 6234 28262
rect 6290 28260 6314 28262
rect 6370 28260 6394 28262
rect 6450 28260 6456 28262
rect 6148 28251 6456 28260
rect 6000 27872 6052 27878
rect 6000 27814 6052 27820
rect 6012 27470 6040 27814
rect 6000 27464 6052 27470
rect 6000 27406 6052 27412
rect 6000 27328 6052 27334
rect 6000 27270 6052 27276
rect 6012 27062 6040 27270
rect 6148 27228 6456 27237
rect 6148 27226 6154 27228
rect 6210 27226 6234 27228
rect 6290 27226 6314 27228
rect 6370 27226 6394 27228
rect 6450 27226 6456 27228
rect 6210 27174 6212 27226
rect 6392 27174 6394 27226
rect 6148 27172 6154 27174
rect 6210 27172 6234 27174
rect 6290 27172 6314 27174
rect 6370 27172 6394 27174
rect 6450 27172 6456 27174
rect 6148 27163 6456 27172
rect 6000 27056 6052 27062
rect 6000 26998 6052 27004
rect 6564 26926 6592 29514
rect 6656 29510 6684 30670
rect 6828 30660 6880 30666
rect 6828 30602 6880 30608
rect 6734 30152 6790 30161
rect 6840 30138 6868 30602
rect 6790 30110 6868 30138
rect 6734 30087 6790 30096
rect 6736 29776 6788 29782
rect 6736 29718 6788 29724
rect 6644 29504 6696 29510
rect 6644 29446 6696 29452
rect 6656 28801 6684 29446
rect 6642 28792 6698 28801
rect 6642 28727 6698 28736
rect 6552 26920 6604 26926
rect 6552 26862 6604 26868
rect 6000 26784 6052 26790
rect 6000 26726 6052 26732
rect 6012 26450 6040 26726
rect 6000 26444 6052 26450
rect 6000 26386 6052 26392
rect 5906 26208 5962 26217
rect 5906 26143 5962 26152
rect 6012 25430 6040 26386
rect 6276 26376 6328 26382
rect 6366 26344 6422 26353
rect 6328 26324 6366 26330
rect 6276 26318 6366 26324
rect 6288 26302 6366 26318
rect 6366 26279 6422 26288
rect 6148 26140 6456 26149
rect 6148 26138 6154 26140
rect 6210 26138 6234 26140
rect 6290 26138 6314 26140
rect 6370 26138 6394 26140
rect 6450 26138 6456 26140
rect 6210 26086 6212 26138
rect 6392 26086 6394 26138
rect 6148 26084 6154 26086
rect 6210 26084 6234 26086
rect 6290 26084 6314 26086
rect 6370 26084 6394 26086
rect 6450 26084 6456 26086
rect 6148 26075 6456 26084
rect 6000 25424 6052 25430
rect 6000 25366 6052 25372
rect 5908 25356 5960 25362
rect 5908 25298 5960 25304
rect 6092 25356 6144 25362
rect 6564 25344 6592 26862
rect 6644 26240 6696 26246
rect 6644 26182 6696 26188
rect 6656 25838 6684 26182
rect 6644 25832 6696 25838
rect 6644 25774 6696 25780
rect 6656 25537 6684 25774
rect 6748 25673 6776 29718
rect 6828 29572 6880 29578
rect 6828 29514 6880 29520
rect 6840 26761 6868 29514
rect 6932 28529 6960 32422
rect 7024 32366 7052 33322
rect 7116 33318 7144 33934
rect 7104 33312 7156 33318
rect 7104 33254 7156 33260
rect 7116 32910 7144 33254
rect 7104 32904 7156 32910
rect 7104 32846 7156 32852
rect 7104 32768 7156 32774
rect 7104 32710 7156 32716
rect 7012 32360 7064 32366
rect 7012 32302 7064 32308
rect 7116 31793 7144 32710
rect 7196 32428 7248 32434
rect 7196 32370 7248 32376
rect 7208 32026 7236 32370
rect 7196 32020 7248 32026
rect 7196 31962 7248 31968
rect 7102 31784 7158 31793
rect 7102 31719 7158 31728
rect 7300 31754 7328 35022
rect 7380 34060 7432 34066
rect 7380 34002 7432 34008
rect 7392 33114 7420 34002
rect 7380 33108 7432 33114
rect 7380 33050 7432 33056
rect 7380 32904 7432 32910
rect 7380 32846 7432 32852
rect 7392 32570 7420 32846
rect 7380 32564 7432 32570
rect 7380 32506 7432 32512
rect 7380 32438 7432 32444
rect 7380 32380 7432 32386
rect 7392 31890 7420 32380
rect 7380 31884 7432 31890
rect 7380 31826 7432 31832
rect 7300 31726 7420 31754
rect 7288 31680 7340 31686
rect 7288 31622 7340 31628
rect 7012 31340 7064 31346
rect 7012 31282 7064 31288
rect 7196 31340 7248 31346
rect 7196 31282 7248 31288
rect 7024 29889 7052 31282
rect 7102 30968 7158 30977
rect 7102 30903 7158 30912
rect 7116 30258 7144 30903
rect 7208 30598 7236 31282
rect 7196 30592 7248 30598
rect 7196 30534 7248 30540
rect 7208 30394 7236 30534
rect 7196 30388 7248 30394
rect 7196 30330 7248 30336
rect 7194 30288 7250 30297
rect 7104 30252 7156 30258
rect 7194 30223 7250 30232
rect 7104 30194 7156 30200
rect 7010 29880 7066 29889
rect 7010 29815 7066 29824
rect 6918 28520 6974 28529
rect 6918 28455 6974 28464
rect 6826 26752 6882 26761
rect 6826 26687 6882 26696
rect 7024 26625 7052 29815
rect 7116 29714 7144 30194
rect 7104 29708 7156 29714
rect 7104 29650 7156 29656
rect 7116 28558 7144 29650
rect 7208 29578 7236 30223
rect 7196 29572 7248 29578
rect 7196 29514 7248 29520
rect 7300 28558 7328 31622
rect 7392 31482 7420 31726
rect 7380 31476 7432 31482
rect 7380 31418 7432 31424
rect 7380 30728 7432 30734
rect 7380 30670 7432 30676
rect 7392 30394 7420 30670
rect 7380 30388 7432 30394
rect 7380 30330 7432 30336
rect 7484 29782 7512 40598
rect 7576 38758 7604 41375
rect 7656 41200 7708 41206
rect 7654 41168 7656 41177
rect 7708 41168 7710 41177
rect 7654 41103 7710 41112
rect 7748 41064 7800 41070
rect 7748 41006 7800 41012
rect 7760 40934 7788 41006
rect 7748 40928 7800 40934
rect 7748 40870 7800 40876
rect 7760 40662 7788 40870
rect 7748 40656 7800 40662
rect 7748 40598 7800 40604
rect 8128 40202 8156 41386
rect 8220 40594 8248 42214
rect 8404 41721 8432 42570
rect 8390 41712 8446 41721
rect 8390 41647 8446 41656
rect 8496 41546 8524 43114
rect 8588 42838 8616 43114
rect 8576 42832 8628 42838
rect 8576 42774 8628 42780
rect 8680 42770 8708 43574
rect 9048 43450 9076 44540
rect 9036 43444 9088 43450
rect 9036 43386 9088 43392
rect 8944 43308 8996 43314
rect 8944 43250 8996 43256
rect 8956 43217 8984 43250
rect 8942 43208 8998 43217
rect 8942 43143 8998 43152
rect 8747 43004 9055 43013
rect 8747 43002 8753 43004
rect 8809 43002 8833 43004
rect 8889 43002 8913 43004
rect 8969 43002 8993 43004
rect 9049 43002 9055 43004
rect 8809 42950 8811 43002
rect 8991 42950 8993 43002
rect 8747 42948 8753 42950
rect 8809 42948 8833 42950
rect 8889 42948 8913 42950
rect 8969 42948 8993 42950
rect 9049 42948 9055 42950
rect 8747 42939 9055 42948
rect 9232 42770 9260 44540
rect 9416 43450 9444 44540
rect 9404 43444 9456 43450
rect 9404 43386 9456 43392
rect 8668 42764 8720 42770
rect 8668 42706 8720 42712
rect 8760 42764 8812 42770
rect 8760 42706 8812 42712
rect 9220 42764 9272 42770
rect 9220 42706 9272 42712
rect 8574 42664 8630 42673
rect 8772 42634 8800 42706
rect 9600 42702 9628 44540
rect 9784 43874 9812 44540
rect 9692 43846 9812 43874
rect 9692 43314 9720 43846
rect 9772 43376 9824 43382
rect 9968 43364 9996 44540
rect 10048 43444 10100 43450
rect 10048 43386 10100 43392
rect 9824 43336 9996 43364
rect 9772 43318 9824 43324
rect 9680 43308 9732 43314
rect 9680 43250 9732 43256
rect 9680 42900 9732 42906
rect 9680 42842 9732 42848
rect 9128 42696 9180 42702
rect 9588 42696 9640 42702
rect 9128 42638 9180 42644
rect 9402 42664 9458 42673
rect 8574 42599 8630 42608
rect 8760 42628 8812 42634
rect 8588 42022 8616 42599
rect 8760 42570 8812 42576
rect 8668 42560 8720 42566
rect 8668 42502 8720 42508
rect 8576 42016 8628 42022
rect 8576 41958 8628 41964
rect 8484 41540 8536 41546
rect 8484 41482 8536 41488
rect 8390 41304 8446 41313
rect 8390 41239 8392 41248
rect 8444 41239 8446 41248
rect 8588 41256 8616 41958
rect 8680 41614 8708 42502
rect 9140 42401 9168 42638
rect 9312 42628 9364 42634
rect 9588 42638 9640 42644
rect 9402 42599 9458 42608
rect 9496 42628 9548 42634
rect 9312 42570 9364 42576
rect 9220 42560 9272 42566
rect 9220 42502 9272 42508
rect 9126 42392 9182 42401
rect 9126 42327 9182 42336
rect 8942 42120 8998 42129
rect 8942 42055 8944 42064
rect 8996 42055 8998 42064
rect 9036 42084 9088 42090
rect 8944 42026 8996 42032
rect 9088 42044 9168 42072
rect 9036 42026 9088 42032
rect 8747 41916 9055 41925
rect 8747 41914 8753 41916
rect 8809 41914 8833 41916
rect 8889 41914 8913 41916
rect 8969 41914 8993 41916
rect 9049 41914 9055 41916
rect 8809 41862 8811 41914
rect 8991 41862 8993 41914
rect 8747 41860 8753 41862
rect 8809 41860 8833 41862
rect 8889 41860 8913 41862
rect 8969 41860 8993 41862
rect 9049 41860 9055 41862
rect 8747 41851 9055 41860
rect 9140 41750 9168 42044
rect 9128 41744 9180 41750
rect 9128 41686 9180 41692
rect 8668 41608 8720 41614
rect 8668 41550 8720 41556
rect 8588 41228 8708 41256
rect 8392 41210 8444 41216
rect 8576 41132 8628 41138
rect 8576 41074 8628 41080
rect 8588 40730 8616 41074
rect 8576 40724 8628 40730
rect 8576 40666 8628 40672
rect 8208 40588 8260 40594
rect 8208 40530 8260 40536
rect 8208 40384 8260 40390
rect 8208 40326 8260 40332
rect 7668 40174 8156 40202
rect 7564 38752 7616 38758
rect 7564 38694 7616 38700
rect 7562 38584 7618 38593
rect 7562 38519 7618 38528
rect 7576 38418 7604 38519
rect 7564 38412 7616 38418
rect 7564 38354 7616 38360
rect 7562 37904 7618 37913
rect 7668 37874 7696 40174
rect 8022 40080 8078 40089
rect 8022 40015 8078 40024
rect 7840 38276 7892 38282
rect 7840 38218 7892 38224
rect 7748 38208 7800 38214
rect 7852 38185 7880 38218
rect 7748 38150 7800 38156
rect 7838 38176 7894 38185
rect 7562 37839 7618 37848
rect 7656 37868 7708 37874
rect 7576 36938 7604 37839
rect 7656 37810 7708 37816
rect 7760 37806 7788 38150
rect 7838 38111 7894 38120
rect 7840 37868 7892 37874
rect 7840 37810 7892 37816
rect 7748 37800 7800 37806
rect 7748 37742 7800 37748
rect 7852 37369 7880 37810
rect 7838 37360 7894 37369
rect 7838 37295 7894 37304
rect 7748 37120 7800 37126
rect 7746 37088 7748 37097
rect 7800 37088 7802 37097
rect 7746 37023 7802 37032
rect 7576 36910 7788 36938
rect 7562 36816 7618 36825
rect 7562 36751 7564 36760
rect 7616 36751 7618 36760
rect 7656 36780 7708 36786
rect 7564 36722 7616 36728
rect 7656 36722 7708 36728
rect 7668 36174 7696 36722
rect 7760 36174 7788 36910
rect 7656 36168 7708 36174
rect 7656 36110 7708 36116
rect 7748 36168 7800 36174
rect 7748 36110 7800 36116
rect 7760 36009 7788 36110
rect 8036 36106 8064 40015
rect 8116 39568 8168 39574
rect 8116 39510 8168 39516
rect 8024 36100 8076 36106
rect 8024 36042 8076 36048
rect 7840 36032 7892 36038
rect 7746 36000 7802 36009
rect 7840 35974 7892 35980
rect 7746 35935 7802 35944
rect 7564 35760 7616 35766
rect 7564 35702 7616 35708
rect 7576 34134 7604 35702
rect 7748 35692 7800 35698
rect 7748 35634 7800 35640
rect 7654 35184 7710 35193
rect 7654 35119 7710 35128
rect 7564 34128 7616 34134
rect 7564 34070 7616 34076
rect 7668 32960 7696 35119
rect 7576 32932 7696 32960
rect 7576 32842 7604 32932
rect 7654 32872 7710 32881
rect 7564 32836 7616 32842
rect 7654 32807 7710 32816
rect 7564 32778 7616 32784
rect 7564 32428 7616 32434
rect 7564 32370 7616 32376
rect 7576 31210 7604 32370
rect 7668 32065 7696 32807
rect 7654 32056 7710 32065
rect 7654 31991 7710 32000
rect 7656 31748 7708 31754
rect 7656 31690 7708 31696
rect 7564 31204 7616 31210
rect 7564 31146 7616 31152
rect 7562 31104 7618 31113
rect 7562 31039 7618 31048
rect 7576 30274 7604 31039
rect 7668 30394 7696 31690
rect 7656 30388 7708 30394
rect 7656 30330 7708 30336
rect 7576 30246 7696 30274
rect 7562 30016 7618 30025
rect 7562 29951 7618 29960
rect 7472 29776 7524 29782
rect 7472 29718 7524 29724
rect 7380 29640 7432 29646
rect 7432 29588 7512 29594
rect 7380 29582 7512 29588
rect 7392 29566 7512 29582
rect 7576 29578 7604 29951
rect 7380 29504 7432 29510
rect 7380 29446 7432 29452
rect 7392 29170 7420 29446
rect 7380 29164 7432 29170
rect 7380 29106 7432 29112
rect 7378 29064 7434 29073
rect 7378 28999 7434 29008
rect 7104 28552 7156 28558
rect 7104 28494 7156 28500
rect 7288 28552 7340 28558
rect 7288 28494 7340 28500
rect 7116 27996 7144 28494
rect 7288 28008 7340 28014
rect 7116 27968 7288 27996
rect 7288 27950 7340 27956
rect 7102 27840 7158 27849
rect 7158 27798 7236 27826
rect 7102 27775 7158 27784
rect 7104 27328 7156 27334
rect 7104 27270 7156 27276
rect 7116 26926 7144 27270
rect 7104 26920 7156 26926
rect 7104 26862 7156 26868
rect 7010 26616 7066 26625
rect 7010 26551 7066 26560
rect 6920 26444 6972 26450
rect 6920 26386 6972 26392
rect 6826 26344 6882 26353
rect 6826 26279 6882 26288
rect 6734 25664 6790 25673
rect 6734 25599 6790 25608
rect 6642 25528 6698 25537
rect 6642 25463 6698 25472
rect 6736 25492 6788 25498
rect 6736 25434 6788 25440
rect 6564 25316 6684 25344
rect 6092 25298 6144 25304
rect 5920 24886 5948 25298
rect 6104 25140 6132 25298
rect 6550 25256 6606 25265
rect 6550 25191 6606 25200
rect 6012 25129 6132 25140
rect 5998 25120 6132 25129
rect 6054 25112 6132 25120
rect 5998 25055 6054 25064
rect 6148 25052 6456 25061
rect 6148 25050 6154 25052
rect 6210 25050 6234 25052
rect 6290 25050 6314 25052
rect 6370 25050 6394 25052
rect 6450 25050 6456 25052
rect 6210 24998 6212 25050
rect 6392 24998 6394 25050
rect 6148 24996 6154 24998
rect 6210 24996 6234 24998
rect 6290 24996 6314 24998
rect 6370 24996 6394 24998
rect 6450 24996 6456 24998
rect 6148 24987 6456 24996
rect 6000 24948 6052 24954
rect 6000 24890 6052 24896
rect 5908 24880 5960 24886
rect 5908 24822 5960 24828
rect 5814 24440 5870 24449
rect 5632 24404 5684 24410
rect 5632 24346 5684 24352
rect 5724 24404 5776 24410
rect 5814 24375 5870 24384
rect 5724 24346 5776 24352
rect 5644 23254 5672 24346
rect 5814 24304 5870 24313
rect 5814 24239 5870 24248
rect 5828 23322 5856 24239
rect 5908 24200 5960 24206
rect 5908 24142 5960 24148
rect 5920 23526 5948 24142
rect 5908 23520 5960 23526
rect 5908 23462 5960 23468
rect 5724 23316 5776 23322
rect 5724 23258 5776 23264
rect 5816 23316 5868 23322
rect 5816 23258 5868 23264
rect 5632 23248 5684 23254
rect 5632 23190 5684 23196
rect 5736 22545 5764 23258
rect 5722 22536 5778 22545
rect 5722 22471 5778 22480
rect 5632 21888 5684 21894
rect 5632 21830 5684 21836
rect 5644 21690 5672 21830
rect 5736 21690 5764 22471
rect 5632 21684 5684 21690
rect 5632 21626 5684 21632
rect 5724 21684 5776 21690
rect 5724 21626 5776 21632
rect 5538 21448 5594 21457
rect 5538 21383 5594 21392
rect 5632 21344 5684 21350
rect 5632 21286 5684 21292
rect 5448 21004 5500 21010
rect 5448 20946 5500 20952
rect 5448 20460 5500 20466
rect 5448 20402 5500 20408
rect 5184 20318 5304 20346
rect 5356 20392 5408 20398
rect 5356 20334 5408 20340
rect 5080 15564 5132 15570
rect 5080 15506 5132 15512
rect 5078 15192 5134 15201
rect 5078 15127 5134 15136
rect 5092 15094 5120 15127
rect 5080 15088 5132 15094
rect 5080 15030 5132 15036
rect 5184 14822 5212 20318
rect 5264 20256 5316 20262
rect 5264 20198 5316 20204
rect 5276 19553 5304 20198
rect 5368 20058 5396 20334
rect 5356 20052 5408 20058
rect 5356 19994 5408 20000
rect 5354 19952 5410 19961
rect 5354 19887 5410 19896
rect 5262 19544 5318 19553
rect 5262 19479 5318 19488
rect 5368 19446 5396 19887
rect 5356 19440 5408 19446
rect 5356 19382 5408 19388
rect 5356 19168 5408 19174
rect 5356 19110 5408 19116
rect 5262 18728 5318 18737
rect 5368 18714 5396 19110
rect 5460 18970 5488 20402
rect 5538 19680 5594 19689
rect 5538 19615 5594 19624
rect 5552 19378 5580 19615
rect 5540 19372 5592 19378
rect 5540 19314 5592 19320
rect 5448 18964 5500 18970
rect 5448 18906 5500 18912
rect 5552 18834 5580 19314
rect 5540 18828 5592 18834
rect 5540 18770 5592 18776
rect 5368 18686 5580 18714
rect 5262 18663 5264 18672
rect 5316 18663 5318 18672
rect 5264 18634 5316 18640
rect 5276 16250 5304 18634
rect 5356 18624 5408 18630
rect 5356 18566 5408 18572
rect 5448 18624 5500 18630
rect 5448 18566 5500 18572
rect 5368 18222 5396 18566
rect 5356 18216 5408 18222
rect 5460 18193 5488 18566
rect 5552 18222 5580 18686
rect 5540 18216 5592 18222
rect 5356 18158 5408 18164
rect 5446 18184 5502 18193
rect 5540 18158 5592 18164
rect 5446 18119 5502 18128
rect 5552 18068 5580 18158
rect 5368 18040 5580 18068
rect 5264 16244 5316 16250
rect 5264 16186 5316 16192
rect 5368 15910 5396 18040
rect 5446 17912 5502 17921
rect 5502 17870 5580 17898
rect 5446 17847 5502 17856
rect 5552 17134 5580 17870
rect 5540 17128 5592 17134
rect 5540 17070 5592 17076
rect 5448 17060 5500 17066
rect 5448 17002 5500 17008
rect 5460 16454 5488 17002
rect 5644 16810 5672 21286
rect 5736 20942 5764 21626
rect 5724 20936 5776 20942
rect 5724 20878 5776 20884
rect 5736 20330 5764 20878
rect 5724 20324 5776 20330
rect 5724 20266 5776 20272
rect 5724 20052 5776 20058
rect 5724 19994 5776 20000
rect 5736 18970 5764 19994
rect 5724 18964 5776 18970
rect 5724 18906 5776 18912
rect 5722 18184 5778 18193
rect 5722 18119 5778 18128
rect 5736 17746 5764 18119
rect 5724 17740 5776 17746
rect 5724 17682 5776 17688
rect 5828 17320 5856 23258
rect 5908 22772 5960 22778
rect 5908 22714 5960 22720
rect 5920 21350 5948 22714
rect 5908 21344 5960 21350
rect 5908 21286 5960 21292
rect 5908 20936 5960 20942
rect 5908 20878 5960 20884
rect 5920 19514 5948 20878
rect 5908 19508 5960 19514
rect 5908 19450 5960 19456
rect 5908 17672 5960 17678
rect 5908 17614 5960 17620
rect 5920 17542 5948 17614
rect 5908 17536 5960 17542
rect 5908 17478 5960 17484
rect 5552 16782 5672 16810
rect 5736 17292 5856 17320
rect 5552 16454 5580 16782
rect 5632 16652 5684 16658
rect 5632 16594 5684 16600
rect 5448 16448 5500 16454
rect 5540 16448 5592 16454
rect 5448 16390 5500 16396
rect 5538 16416 5540 16425
rect 5592 16416 5594 16425
rect 5538 16351 5594 16360
rect 5356 15904 5408 15910
rect 5356 15846 5408 15852
rect 5448 15564 5500 15570
rect 5448 15506 5500 15512
rect 5264 15496 5316 15502
rect 5264 15438 5316 15444
rect 5172 14816 5224 14822
rect 5172 14758 5224 14764
rect 5078 14104 5134 14113
rect 5078 14039 5134 14048
rect 5092 13938 5120 14039
rect 5080 13932 5132 13938
rect 5184 13920 5212 14758
rect 5276 14618 5304 15438
rect 5264 14612 5316 14618
rect 5264 14554 5316 14560
rect 5356 14340 5408 14346
rect 5356 14282 5408 14288
rect 5262 14240 5318 14249
rect 5262 14175 5318 14184
rect 5276 14074 5304 14175
rect 5368 14074 5396 14282
rect 5264 14068 5316 14074
rect 5264 14010 5316 14016
rect 5356 14068 5408 14074
rect 5356 14010 5408 14016
rect 5184 13892 5396 13920
rect 5080 13874 5132 13880
rect 5000 13756 5212 13784
rect 4894 13560 4950 13569
rect 4894 13495 4950 13504
rect 4908 13394 4936 13495
rect 4764 13348 4844 13376
rect 4896 13388 4948 13394
rect 4712 13330 4764 13336
rect 4896 13330 4948 13336
rect 4618 13288 4674 13297
rect 4618 13223 4674 13232
rect 4632 12850 4660 13223
rect 4620 12844 4672 12850
rect 4620 12786 4672 12792
rect 4632 12306 4660 12786
rect 4724 12442 4752 13330
rect 4986 13288 5042 13297
rect 4986 13223 5042 13232
rect 4804 12640 4856 12646
rect 5000 12594 5028 13223
rect 5184 12594 5212 13756
rect 5368 13410 5396 13892
rect 4804 12582 4856 12588
rect 4712 12436 4764 12442
rect 4712 12378 4764 12384
rect 4620 12300 4672 12306
rect 4620 12242 4672 12248
rect 4712 12300 4764 12306
rect 4816 12288 4844 12582
rect 4764 12260 4844 12288
rect 4908 12566 5028 12594
rect 5090 12566 5212 12594
rect 5276 13382 5396 13410
rect 4712 12242 4764 12248
rect 4528 11892 4580 11898
rect 4528 11834 4580 11840
rect 4712 11892 4764 11898
rect 4712 11834 4764 11840
rect 4724 11762 4752 11834
rect 4712 11756 4764 11762
rect 4712 11698 4764 11704
rect 4436 11144 4488 11150
rect 4436 11086 4488 11092
rect 4804 11076 4856 11082
rect 4804 11018 4856 11024
rect 4342 10976 4398 10985
rect 4342 10911 4398 10920
rect 4618 10976 4674 10985
rect 4816 10962 4844 11018
rect 4618 10911 4674 10920
rect 4724 10934 4844 10962
rect 4342 10840 4398 10849
rect 4342 10775 4398 10784
rect 4252 9376 4304 9382
rect 4252 9318 4304 9324
rect 4068 8968 4120 8974
rect 4068 8910 4120 8916
rect 4160 8968 4212 8974
rect 4160 8910 4212 8916
rect 4080 8809 4108 8910
rect 4066 8800 4122 8809
rect 4066 8735 4122 8744
rect 4252 8560 4304 8566
rect 4252 8502 4304 8508
rect 4160 8492 4212 8498
rect 4160 8434 4212 8440
rect 3884 8424 3936 8430
rect 3804 8384 3884 8412
rect 3884 8366 3936 8372
rect 3330 8256 3386 8265
rect 3330 8191 3386 8200
rect 3436 8248 3648 8276
rect 3896 8294 3924 8366
rect 3896 8266 4108 8294
rect 3240 8084 3292 8090
rect 3240 8026 3292 8032
rect 3238 7848 3294 7857
rect 3294 7806 3372 7834
rect 3238 7783 3294 7792
rect 3240 7404 3292 7410
rect 3240 7346 3292 7352
rect 3148 6452 3200 6458
rect 3148 6394 3200 6400
rect 3148 6112 3200 6118
rect 3148 6054 3200 6060
rect 3056 5364 3108 5370
rect 3056 5306 3108 5312
rect 3056 5228 3108 5234
rect 3056 5170 3108 5176
rect 3068 5137 3096 5170
rect 3054 5128 3110 5137
rect 3054 5063 3110 5072
rect 3160 4826 3188 6054
rect 3148 4820 3200 4826
rect 3148 4762 3200 4768
rect 3056 4208 3108 4214
rect 3056 4150 3108 4156
rect 3068 3058 3096 4150
rect 3252 3942 3280 7346
rect 3344 7002 3372 7806
rect 3332 6996 3384 7002
rect 3332 6938 3384 6944
rect 3332 6792 3384 6798
rect 3330 6760 3332 6769
rect 3384 6760 3386 6769
rect 3330 6695 3386 6704
rect 3436 6662 3464 8248
rect 3549 8188 3857 8197
rect 3549 8186 3555 8188
rect 3611 8186 3635 8188
rect 3691 8186 3715 8188
rect 3771 8186 3795 8188
rect 3851 8186 3857 8188
rect 3611 8134 3613 8186
rect 3793 8134 3795 8186
rect 3549 8132 3555 8134
rect 3611 8132 3635 8134
rect 3691 8132 3715 8134
rect 3771 8132 3795 8134
rect 3851 8132 3857 8134
rect 3549 8123 3857 8132
rect 4080 8022 4108 8266
rect 4172 8090 4200 8434
rect 4264 8362 4292 8502
rect 4252 8356 4304 8362
rect 4252 8298 4304 8304
rect 4160 8084 4212 8090
rect 4160 8026 4212 8032
rect 4068 8016 4120 8022
rect 4120 7964 4292 7970
rect 4068 7958 4292 7964
rect 4080 7942 4292 7958
rect 3792 7880 3844 7886
rect 3790 7848 3792 7857
rect 4068 7880 4120 7886
rect 3844 7848 3846 7857
rect 4068 7822 4120 7828
rect 3790 7783 3846 7792
rect 3884 7744 3936 7750
rect 3884 7686 3936 7692
rect 3896 7274 3924 7686
rect 4080 7546 4108 7822
rect 4158 7712 4214 7721
rect 4158 7647 4214 7656
rect 4172 7546 4200 7647
rect 4068 7540 4120 7546
rect 4068 7482 4120 7488
rect 4160 7540 4212 7546
rect 4160 7482 4212 7488
rect 4264 7460 4292 7942
rect 4356 7528 4384 10775
rect 4436 10736 4488 10742
rect 4436 10678 4488 10684
rect 4448 9518 4476 10678
rect 4528 10056 4580 10062
rect 4528 9998 4580 10004
rect 4436 9512 4488 9518
rect 4436 9454 4488 9460
rect 4448 7732 4476 9454
rect 4540 9178 4568 9998
rect 4632 9926 4660 10911
rect 4724 10674 4752 10934
rect 4712 10668 4764 10674
rect 4712 10610 4764 10616
rect 4620 9920 4672 9926
rect 4620 9862 4672 9868
rect 4724 9738 4752 10610
rect 4802 10568 4858 10577
rect 4802 10503 4858 10512
rect 4816 10033 4844 10503
rect 4802 10024 4858 10033
rect 4802 9959 4858 9968
rect 4632 9710 4752 9738
rect 4632 9518 4660 9710
rect 4712 9580 4764 9586
rect 4712 9522 4764 9528
rect 4620 9512 4672 9518
rect 4620 9454 4672 9460
rect 4528 9172 4580 9178
rect 4528 9114 4580 9120
rect 4528 9036 4580 9042
rect 4528 8978 4580 8984
rect 4540 8401 4568 8978
rect 4632 8634 4660 9454
rect 4724 9353 4752 9522
rect 4804 9444 4856 9450
rect 4804 9386 4856 9392
rect 4710 9344 4766 9353
rect 4710 9279 4766 9288
rect 4710 9072 4766 9081
rect 4710 9007 4766 9016
rect 4620 8628 4672 8634
rect 4620 8570 4672 8576
rect 4526 8392 4582 8401
rect 4526 8327 4582 8336
rect 4620 8288 4672 8294
rect 4620 8230 4672 8236
rect 4526 8120 4582 8129
rect 4632 8090 4660 8230
rect 4526 8055 4582 8064
rect 4620 8084 4672 8090
rect 4540 7886 4568 8055
rect 4620 8026 4672 8032
rect 4528 7880 4580 7886
rect 4528 7822 4580 7828
rect 4724 7750 4752 9007
rect 4712 7744 4764 7750
rect 4448 7704 4660 7732
rect 4436 7540 4488 7546
rect 4356 7500 4436 7528
rect 4436 7482 4488 7488
rect 4158 7440 4214 7449
rect 3976 7404 4028 7410
rect 4264 7432 4384 7460
rect 4158 7375 4214 7384
rect 3976 7346 4028 7352
rect 3884 7268 3936 7274
rect 3884 7210 3936 7216
rect 3549 7100 3857 7109
rect 3549 7098 3555 7100
rect 3611 7098 3635 7100
rect 3691 7098 3715 7100
rect 3771 7098 3795 7100
rect 3851 7098 3857 7100
rect 3611 7046 3613 7098
rect 3793 7046 3795 7098
rect 3549 7044 3555 7046
rect 3611 7044 3635 7046
rect 3691 7044 3715 7046
rect 3771 7044 3795 7046
rect 3851 7044 3857 7046
rect 3549 7035 3857 7044
rect 3700 6792 3752 6798
rect 3700 6734 3752 6740
rect 3790 6760 3846 6769
rect 3424 6656 3476 6662
rect 3424 6598 3476 6604
rect 3516 6452 3568 6458
rect 3516 6394 3568 6400
rect 3424 6248 3476 6254
rect 3528 6225 3556 6394
rect 3424 6190 3476 6196
rect 3514 6216 3570 6225
rect 3330 5672 3386 5681
rect 3330 5607 3386 5616
rect 3240 3936 3292 3942
rect 3240 3878 3292 3884
rect 3344 3738 3372 5607
rect 3436 4486 3464 6190
rect 3712 6186 3740 6734
rect 3790 6695 3846 6704
rect 3804 6322 3832 6695
rect 3882 6488 3938 6497
rect 3882 6423 3938 6432
rect 3792 6316 3844 6322
rect 3792 6258 3844 6264
rect 3514 6151 3570 6160
rect 3700 6180 3752 6186
rect 3700 6122 3752 6128
rect 3549 6012 3857 6021
rect 3549 6010 3555 6012
rect 3611 6010 3635 6012
rect 3691 6010 3715 6012
rect 3771 6010 3795 6012
rect 3851 6010 3857 6012
rect 3611 5958 3613 6010
rect 3793 5958 3795 6010
rect 3549 5956 3555 5958
rect 3611 5956 3635 5958
rect 3691 5956 3715 5958
rect 3771 5956 3795 5958
rect 3851 5956 3857 5958
rect 3549 5947 3857 5956
rect 3896 5896 3924 6423
rect 3804 5868 3924 5896
rect 3804 5710 3832 5868
rect 3884 5772 3936 5778
rect 3988 5760 4016 7346
rect 4066 6896 4122 6905
rect 4066 6831 4122 6840
rect 4080 6118 4108 6831
rect 4172 6458 4200 7375
rect 4252 6928 4304 6934
rect 4250 6896 4252 6905
rect 4304 6896 4306 6905
rect 4250 6831 4306 6840
rect 4252 6792 4304 6798
rect 4250 6760 4252 6769
rect 4304 6760 4306 6769
rect 4250 6695 4306 6704
rect 4160 6452 4212 6458
rect 4160 6394 4212 6400
rect 4158 6352 4214 6361
rect 4158 6287 4214 6296
rect 4068 6112 4120 6118
rect 4068 6054 4120 6060
rect 4068 5908 4120 5914
rect 4068 5850 4120 5856
rect 4080 5817 4108 5850
rect 4172 5846 4200 6287
rect 4264 5846 4292 6695
rect 4356 6322 4384 7432
rect 4434 7440 4490 7449
rect 4434 7375 4490 7384
rect 4344 6316 4396 6322
rect 4344 6258 4396 6264
rect 4448 6225 4476 7375
rect 4528 7336 4580 7342
rect 4528 7278 4580 7284
rect 4540 7177 4568 7278
rect 4526 7168 4582 7177
rect 4526 7103 4582 7112
rect 4528 6792 4580 6798
rect 4632 6769 4660 7704
rect 4712 7686 4764 7692
rect 4710 7440 4766 7449
rect 4710 7375 4712 7384
rect 4764 7375 4766 7384
rect 4712 7346 4764 7352
rect 4816 7290 4844 9386
rect 4908 8566 4936 12566
rect 5090 12458 5118 12566
rect 5000 12430 5118 12458
rect 5172 12436 5224 12442
rect 5000 11898 5028 12430
rect 5172 12378 5224 12384
rect 5078 12336 5134 12345
rect 5078 12271 5134 12280
rect 5092 12238 5120 12271
rect 5080 12232 5132 12238
rect 5080 12174 5132 12180
rect 4988 11892 5040 11898
rect 4988 11834 5040 11840
rect 4988 11756 5040 11762
rect 4988 11698 5040 11704
rect 5000 11529 5028 11698
rect 4986 11520 5042 11529
rect 4986 11455 5042 11464
rect 4988 11280 5040 11286
rect 4988 11222 5040 11228
rect 5000 10849 5028 11222
rect 4986 10840 5042 10849
rect 4986 10775 5042 10784
rect 4988 10532 5040 10538
rect 4988 10474 5040 10480
rect 4896 8560 4948 8566
rect 4896 8502 4948 8508
rect 4724 7262 4844 7290
rect 4724 7206 4752 7262
rect 4712 7200 4764 7206
rect 4712 7142 4764 7148
rect 4724 6866 4752 7142
rect 4712 6860 4764 6866
rect 4712 6802 4764 6808
rect 4804 6860 4856 6866
rect 4804 6802 4856 6808
rect 4528 6734 4580 6740
rect 4618 6760 4674 6769
rect 4540 6610 4568 6734
rect 4618 6695 4674 6704
rect 4618 6624 4674 6633
rect 4540 6582 4618 6610
rect 4618 6559 4674 6568
rect 4434 6216 4490 6225
rect 4344 6180 4396 6186
rect 4434 6151 4490 6160
rect 4344 6122 4396 6128
rect 4160 5840 4212 5846
rect 3936 5732 4016 5760
rect 4066 5808 4122 5817
rect 4160 5782 4212 5788
rect 4252 5840 4304 5846
rect 4252 5782 4304 5788
rect 4066 5743 4122 5752
rect 3884 5714 3936 5720
rect 3792 5704 3844 5710
rect 4160 5704 4212 5710
rect 3792 5646 3844 5652
rect 4158 5672 4160 5681
rect 4212 5672 4214 5681
rect 4158 5607 4214 5616
rect 3976 5568 4028 5574
rect 3976 5510 4028 5516
rect 4066 5536 4122 5545
rect 3884 5296 3936 5302
rect 3884 5238 3936 5244
rect 3549 4924 3857 4933
rect 3549 4922 3555 4924
rect 3611 4922 3635 4924
rect 3691 4922 3715 4924
rect 3771 4922 3795 4924
rect 3851 4922 3857 4924
rect 3611 4870 3613 4922
rect 3793 4870 3795 4922
rect 3549 4868 3555 4870
rect 3611 4868 3635 4870
rect 3691 4868 3715 4870
rect 3771 4868 3795 4870
rect 3851 4868 3857 4870
rect 3549 4859 3857 4868
rect 3608 4752 3660 4758
rect 3608 4694 3660 4700
rect 3620 4593 3648 4694
rect 3896 4690 3924 5238
rect 3884 4684 3936 4690
rect 3884 4626 3936 4632
rect 3606 4584 3662 4593
rect 3606 4519 3662 4528
rect 3792 4548 3844 4554
rect 3792 4490 3844 4496
rect 3424 4480 3476 4486
rect 3424 4422 3476 4428
rect 3698 4448 3754 4457
rect 3698 4383 3754 4392
rect 3712 4146 3740 4383
rect 3700 4140 3752 4146
rect 3700 4082 3752 4088
rect 3804 4078 3832 4490
rect 3896 4146 3924 4626
rect 3988 4282 4016 5510
rect 4122 5494 4292 5522
rect 4066 5471 4122 5480
rect 4066 5264 4122 5273
rect 4066 5199 4122 5208
rect 3976 4276 4028 4282
rect 3976 4218 4028 4224
rect 3884 4140 3936 4146
rect 3884 4082 3936 4088
rect 3792 4072 3844 4078
rect 3792 4014 3844 4020
rect 3549 3836 3857 3845
rect 3549 3834 3555 3836
rect 3611 3834 3635 3836
rect 3691 3834 3715 3836
rect 3771 3834 3795 3836
rect 3851 3834 3857 3836
rect 3611 3782 3613 3834
rect 3793 3782 3795 3834
rect 3549 3780 3555 3782
rect 3611 3780 3635 3782
rect 3691 3780 3715 3782
rect 3771 3780 3795 3782
rect 3851 3780 3857 3782
rect 3549 3771 3857 3780
rect 3332 3732 3384 3738
rect 3332 3674 3384 3680
rect 3792 3596 3844 3602
rect 3896 3584 3924 4082
rect 3844 3556 3924 3584
rect 3792 3538 3844 3544
rect 4080 3482 4108 5199
rect 4160 4140 4212 4146
rect 4160 4082 4212 4088
rect 4172 3641 4200 4082
rect 4158 3632 4214 3641
rect 4158 3567 4214 3576
rect 3240 3460 3292 3466
rect 4080 3454 4200 3482
rect 3240 3402 3292 3408
rect 3148 3392 3200 3398
rect 3148 3334 3200 3340
rect 3160 3194 3188 3334
rect 3252 3194 3280 3402
rect 3148 3188 3200 3194
rect 3148 3130 3200 3136
rect 3240 3188 3292 3194
rect 3240 3130 3292 3136
rect 3424 3120 3476 3126
rect 3424 3062 3476 3068
rect 3056 3052 3108 3058
rect 3056 2994 3108 3000
rect 2872 2984 2924 2990
rect 2872 2926 2924 2932
rect 2964 2984 3016 2990
rect 2964 2926 3016 2932
rect 2700 2774 2820 2802
rect 3436 2774 3464 3062
rect 4066 2952 4122 2961
rect 3976 2916 4028 2922
rect 4066 2887 4122 2896
rect 3976 2858 4028 2864
rect 3988 2774 4016 2858
rect 2596 2440 2648 2446
rect 2596 2382 2648 2388
rect 2700 2292 2728 2774
rect 3344 2746 3464 2774
rect 3549 2748 3857 2757
rect 3549 2746 3555 2748
rect 3611 2746 3635 2748
rect 3691 2746 3715 2748
rect 3771 2746 3795 2748
rect 3851 2746 3857 2748
rect 2870 2544 2926 2553
rect 2870 2479 2926 2488
rect 2608 2264 2728 2292
rect 2608 2106 2636 2264
rect 2884 2106 2912 2479
rect 2596 2100 2648 2106
rect 2596 2042 2648 2048
rect 2872 2100 2924 2106
rect 2872 2042 2924 2048
rect 2504 1964 2556 1970
rect 2504 1906 2556 1912
rect 3240 1964 3292 1970
rect 3240 1906 3292 1912
rect 3148 1828 3200 1834
rect 3148 1770 3200 1776
rect 1584 1556 1636 1562
rect 1584 1498 1636 1504
rect 3160 1494 3188 1770
rect 3148 1488 3200 1494
rect 3148 1430 3200 1436
rect 2780 1352 2832 1358
rect 2780 1294 2832 1300
rect 1492 1284 1544 1290
rect 1492 1226 1544 1232
rect 2596 1284 2648 1290
rect 2596 1226 2648 1232
rect 848 944 900 950
rect 848 886 900 892
rect 1504 785 1532 1226
rect 2504 1216 2556 1222
rect 2504 1158 2556 1164
rect 2516 1018 2544 1158
rect 2504 1012 2556 1018
rect 2504 954 2556 960
rect 1490 776 1546 785
rect 1490 711 1546 720
rect 2608 82 2636 1226
rect 2792 746 2820 1294
rect 2780 740 2832 746
rect 2780 682 2832 688
rect 2962 82 3018 160
rect 2608 54 3018 82
rect 2962 -300 3018 54
rect 3146 82 3202 160
rect 3252 82 3280 1906
rect 3344 1426 3372 2746
rect 3611 2694 3613 2746
rect 3793 2694 3795 2746
rect 3549 2692 3555 2694
rect 3611 2692 3635 2694
rect 3691 2692 3715 2694
rect 3771 2692 3795 2694
rect 3851 2692 3857 2694
rect 3549 2683 3857 2692
rect 3896 2746 4016 2774
rect 3896 2446 3924 2746
rect 4080 2666 4108 2887
rect 3988 2638 4108 2666
rect 4172 2650 4200 3454
rect 4264 2854 4292 5494
rect 4356 5302 4384 6122
rect 4724 5896 4752 6802
rect 4632 5868 4752 5896
rect 4436 5840 4488 5846
rect 4436 5782 4488 5788
rect 4448 5658 4476 5782
rect 4632 5778 4660 5868
rect 4620 5772 4672 5778
rect 4620 5714 4672 5720
rect 4448 5630 4752 5658
rect 4620 5568 4672 5574
rect 4620 5510 4672 5516
rect 4344 5296 4396 5302
rect 4344 5238 4396 5244
rect 4632 5234 4660 5510
rect 4620 5228 4672 5234
rect 4620 5170 4672 5176
rect 4724 4826 4752 5630
rect 4816 4826 4844 6802
rect 4908 5574 4936 8502
rect 5000 8090 5028 10474
rect 5092 10033 5120 12174
rect 5184 10112 5212 12378
rect 5276 11830 5304 13382
rect 5354 13288 5410 13297
rect 5354 13223 5410 13232
rect 5366 13212 5396 13223
rect 5368 12850 5396 13212
rect 5356 12844 5408 12850
rect 5356 12786 5408 12792
rect 5354 12064 5410 12073
rect 5354 11999 5410 12008
rect 5264 11824 5316 11830
rect 5264 11766 5316 11772
rect 5276 10656 5304 11766
rect 5368 11529 5396 11999
rect 5354 11520 5410 11529
rect 5354 11455 5410 11464
rect 5460 11218 5488 15506
rect 5540 15360 5592 15366
rect 5540 15302 5592 15308
rect 5552 13530 5580 15302
rect 5644 14074 5672 16594
rect 5736 15026 5764 17292
rect 6012 17218 6040 24890
rect 6564 24886 6592 25191
rect 6552 24880 6604 24886
rect 6552 24822 6604 24828
rect 6090 24576 6146 24585
rect 6090 24511 6146 24520
rect 6104 24274 6132 24511
rect 6092 24268 6144 24274
rect 6092 24210 6144 24216
rect 6552 24064 6604 24070
rect 6552 24006 6604 24012
rect 6148 23964 6456 23973
rect 6148 23962 6154 23964
rect 6210 23962 6234 23964
rect 6290 23962 6314 23964
rect 6370 23962 6394 23964
rect 6450 23962 6456 23964
rect 6210 23910 6212 23962
rect 6392 23910 6394 23962
rect 6148 23908 6154 23910
rect 6210 23908 6234 23910
rect 6290 23908 6314 23910
rect 6370 23908 6394 23910
rect 6450 23908 6456 23910
rect 6148 23899 6456 23908
rect 6564 23730 6592 24006
rect 6552 23724 6604 23730
rect 6552 23666 6604 23672
rect 6460 23520 6512 23526
rect 6460 23462 6512 23468
rect 6552 23520 6604 23526
rect 6552 23462 6604 23468
rect 6276 23316 6328 23322
rect 6276 23258 6328 23264
rect 6288 23186 6316 23258
rect 6472 23186 6500 23462
rect 6564 23225 6592 23462
rect 6550 23216 6606 23225
rect 6276 23180 6328 23186
rect 6276 23122 6328 23128
rect 6460 23180 6512 23186
rect 6550 23151 6606 23160
rect 6460 23122 6512 23128
rect 6552 22976 6604 22982
rect 6552 22918 6604 22924
rect 6148 22876 6456 22885
rect 6148 22874 6154 22876
rect 6210 22874 6234 22876
rect 6290 22874 6314 22876
rect 6370 22874 6394 22876
rect 6450 22874 6456 22876
rect 6210 22822 6212 22874
rect 6392 22822 6394 22874
rect 6148 22820 6154 22822
rect 6210 22820 6234 22822
rect 6290 22820 6314 22822
rect 6370 22820 6394 22822
rect 6450 22820 6456 22822
rect 6148 22811 6456 22820
rect 6564 22760 6592 22918
rect 6472 22732 6592 22760
rect 6472 22273 6500 22732
rect 6552 22568 6604 22574
rect 6552 22510 6604 22516
rect 6458 22264 6514 22273
rect 6458 22199 6514 22208
rect 6368 22160 6420 22166
rect 6288 22120 6368 22148
rect 6288 22001 6316 22120
rect 6368 22102 6420 22108
rect 6472 22098 6500 22199
rect 6460 22092 6512 22098
rect 6460 22034 6512 22040
rect 6274 21992 6330 22001
rect 6274 21927 6330 21936
rect 6148 21788 6456 21797
rect 6148 21786 6154 21788
rect 6210 21786 6234 21788
rect 6290 21786 6314 21788
rect 6370 21786 6394 21788
rect 6450 21786 6456 21788
rect 6210 21734 6212 21786
rect 6392 21734 6394 21786
rect 6148 21732 6154 21734
rect 6210 21732 6234 21734
rect 6290 21732 6314 21734
rect 6370 21732 6394 21734
rect 6450 21732 6456 21734
rect 6148 21723 6456 21732
rect 6184 21344 6236 21350
rect 6184 21286 6236 21292
rect 6196 21146 6224 21286
rect 6184 21140 6236 21146
rect 6184 21082 6236 21088
rect 6182 20904 6238 20913
rect 6182 20839 6238 20848
rect 6196 20806 6224 20839
rect 6184 20800 6236 20806
rect 6184 20742 6236 20748
rect 6148 20700 6456 20709
rect 6148 20698 6154 20700
rect 6210 20698 6234 20700
rect 6290 20698 6314 20700
rect 6370 20698 6394 20700
rect 6450 20698 6456 20700
rect 6210 20646 6212 20698
rect 6392 20646 6394 20698
rect 6148 20644 6154 20646
rect 6210 20644 6234 20646
rect 6290 20644 6314 20646
rect 6370 20644 6394 20646
rect 6450 20644 6456 20646
rect 6148 20635 6456 20644
rect 6564 20534 6592 22510
rect 6460 20528 6512 20534
rect 6458 20496 6460 20505
rect 6552 20528 6604 20534
rect 6512 20496 6514 20505
rect 6552 20470 6604 20476
rect 6458 20431 6514 20440
rect 6656 20346 6684 25316
rect 6748 21962 6776 25434
rect 6840 24818 6868 26279
rect 6932 25294 6960 26386
rect 7208 26330 7236 27798
rect 7300 27713 7328 27950
rect 7286 27704 7342 27713
rect 7286 27639 7342 27648
rect 7288 27464 7340 27470
rect 7288 27406 7340 27412
rect 7116 26302 7236 26330
rect 7116 25786 7144 26302
rect 7196 26240 7248 26246
rect 7196 26182 7248 26188
rect 7208 26042 7236 26182
rect 7300 26042 7328 27406
rect 7392 27112 7420 28999
rect 7484 27470 7512 29566
rect 7564 29572 7616 29578
rect 7564 29514 7616 29520
rect 7576 29073 7604 29514
rect 7562 29064 7618 29073
rect 7562 28999 7618 29008
rect 7668 28150 7696 30246
rect 7656 28144 7708 28150
rect 7656 28086 7708 28092
rect 7668 27713 7696 28086
rect 7760 27985 7788 35634
rect 7852 30682 7880 35974
rect 8024 35488 8076 35494
rect 8024 35430 8076 35436
rect 7930 35184 7986 35193
rect 8036 35154 8064 35430
rect 7930 35119 7986 35128
rect 8024 35148 8076 35154
rect 7944 34610 7972 35119
rect 8024 35090 8076 35096
rect 8024 34944 8076 34950
rect 8024 34886 8076 34892
rect 7932 34604 7984 34610
rect 7932 34546 7984 34552
rect 7944 32774 7972 34546
rect 8036 34048 8064 34886
rect 8128 34202 8156 39510
rect 8220 38214 8248 40326
rect 8392 39296 8444 39302
rect 8392 39238 8444 39244
rect 8300 39024 8352 39030
rect 8300 38966 8352 38972
rect 8312 38457 8340 38966
rect 8298 38448 8354 38457
rect 8298 38383 8354 38392
rect 8208 38208 8260 38214
rect 8208 38150 8260 38156
rect 8300 37868 8352 37874
rect 8300 37810 8352 37816
rect 8312 36922 8340 37810
rect 8300 36916 8352 36922
rect 8300 36858 8352 36864
rect 8300 36100 8352 36106
rect 8300 36042 8352 36048
rect 8312 35737 8340 36042
rect 8298 35728 8354 35737
rect 8298 35663 8354 35672
rect 8300 35216 8352 35222
rect 8300 35158 8352 35164
rect 8206 34776 8262 34785
rect 8206 34711 8262 34720
rect 8116 34196 8168 34202
rect 8116 34138 8168 34144
rect 8116 34060 8168 34066
rect 8036 34020 8116 34048
rect 8116 34002 8168 34008
rect 8220 33969 8248 34711
rect 8022 33960 8078 33969
rect 8022 33895 8024 33904
rect 8076 33895 8078 33904
rect 8206 33960 8262 33969
rect 8206 33895 8262 33904
rect 8024 33866 8076 33872
rect 8036 33522 8064 33866
rect 8024 33516 8076 33522
rect 8024 33458 8076 33464
rect 7932 32768 7984 32774
rect 7932 32710 7984 32716
rect 8024 32224 8076 32230
rect 7930 32192 7986 32201
rect 8024 32166 8076 32172
rect 7930 32127 7986 32136
rect 7944 31754 7972 32127
rect 7932 31748 7984 31754
rect 7932 31690 7984 31696
rect 7932 31272 7984 31278
rect 8036 31260 8064 32166
rect 8114 31784 8170 31793
rect 8114 31719 8170 31728
rect 7984 31232 8064 31260
rect 7932 31214 7984 31220
rect 8024 31136 8076 31142
rect 8024 31078 8076 31084
rect 8036 30802 8064 31078
rect 8024 30796 8076 30802
rect 8024 30738 8076 30744
rect 7852 30654 8064 30682
rect 7932 30592 7984 30598
rect 7932 30534 7984 30540
rect 7840 30048 7892 30054
rect 7840 29990 7892 29996
rect 7852 29850 7880 29990
rect 7840 29844 7892 29850
rect 7840 29786 7892 29792
rect 7840 29640 7892 29646
rect 7840 29582 7892 29588
rect 7852 29034 7880 29582
rect 7840 29028 7892 29034
rect 7840 28970 7892 28976
rect 7840 28688 7892 28694
rect 7838 28656 7840 28665
rect 7892 28656 7894 28665
rect 7838 28591 7894 28600
rect 7840 28552 7892 28558
rect 7840 28494 7892 28500
rect 7746 27976 7802 27985
rect 7746 27911 7802 27920
rect 7748 27872 7800 27878
rect 7748 27814 7800 27820
rect 7654 27704 7710 27713
rect 7654 27639 7710 27648
rect 7472 27464 7524 27470
rect 7472 27406 7524 27412
rect 7760 27402 7788 27814
rect 7564 27396 7616 27402
rect 7564 27338 7616 27344
rect 7656 27396 7708 27402
rect 7656 27338 7708 27344
rect 7748 27396 7800 27402
rect 7748 27338 7800 27344
rect 7392 27084 7512 27112
rect 7378 27024 7434 27033
rect 7378 26959 7380 26968
rect 7432 26959 7434 26968
rect 7380 26930 7432 26936
rect 7392 26330 7420 26930
rect 7484 26432 7512 27084
rect 7576 26994 7604 27338
rect 7564 26988 7616 26994
rect 7564 26930 7616 26936
rect 7484 26404 7604 26432
rect 7392 26302 7512 26330
rect 7196 26036 7248 26042
rect 7196 25978 7248 25984
rect 7288 26036 7340 26042
rect 7288 25978 7340 25984
rect 7116 25758 7236 25786
rect 7104 25696 7156 25702
rect 7104 25638 7156 25644
rect 7010 25528 7066 25537
rect 7116 25498 7144 25638
rect 7010 25463 7066 25472
rect 7104 25492 7156 25498
rect 6920 25288 6972 25294
rect 6920 25230 6972 25236
rect 6932 25158 6960 25230
rect 6920 25152 6972 25158
rect 6920 25094 6972 25100
rect 6828 24812 6880 24818
rect 6828 24754 6880 24760
rect 6828 24200 6880 24206
rect 6828 24142 6880 24148
rect 6840 23186 6868 24142
rect 6828 23180 6880 23186
rect 6828 23122 6880 23128
rect 6840 22642 6868 23122
rect 6828 22636 6880 22642
rect 6828 22578 6880 22584
rect 7024 22522 7052 25463
rect 7104 25434 7156 25440
rect 7104 24676 7156 24682
rect 7104 24618 7156 24624
rect 6840 22494 7052 22522
rect 6736 21956 6788 21962
rect 6736 21898 6788 21904
rect 6736 21344 6788 21350
rect 6736 21286 6788 21292
rect 6748 20942 6776 21286
rect 6736 20936 6788 20942
rect 6736 20878 6788 20884
rect 6840 20874 6868 22494
rect 7116 22386 7144 24618
rect 7208 24177 7236 25758
rect 7300 24818 7328 25978
rect 7288 24812 7340 24818
rect 7288 24754 7340 24760
rect 7380 24744 7432 24750
rect 7380 24686 7432 24692
rect 7194 24168 7250 24177
rect 7194 24103 7250 24112
rect 7392 24052 7420 24686
rect 7114 22358 7144 22386
rect 7208 24024 7420 24052
rect 7114 22250 7142 22358
rect 7114 22222 7144 22250
rect 6920 21480 6972 21486
rect 6920 21422 6972 21428
rect 6828 20868 6880 20874
rect 6828 20810 6880 20816
rect 6932 20777 6960 21422
rect 7116 20924 7144 22222
rect 7208 21298 7236 24024
rect 7484 23730 7512 26302
rect 7576 24206 7604 26404
rect 7668 24426 7696 27338
rect 7852 27282 7880 28494
rect 7760 27254 7880 27282
rect 7760 25906 7788 27254
rect 7840 26376 7892 26382
rect 7838 26344 7840 26353
rect 7892 26344 7894 26353
rect 7838 26279 7894 26288
rect 7840 26240 7892 26246
rect 7840 26182 7892 26188
rect 7852 25906 7880 26182
rect 7748 25900 7800 25906
rect 7748 25842 7800 25848
rect 7840 25900 7892 25906
rect 7840 25842 7892 25848
rect 7760 25673 7788 25842
rect 7746 25664 7802 25673
rect 7746 25599 7802 25608
rect 7852 24750 7880 25842
rect 7840 24744 7892 24750
rect 7840 24686 7892 24692
rect 7668 24398 7880 24426
rect 7564 24200 7616 24206
rect 7564 24142 7616 24148
rect 7748 24064 7800 24070
rect 7748 24006 7800 24012
rect 7472 23724 7524 23730
rect 7392 23684 7472 23712
rect 7286 23216 7342 23225
rect 7286 23151 7342 23160
rect 7300 22166 7328 23151
rect 7392 22778 7420 23684
rect 7472 23666 7524 23672
rect 7564 23724 7616 23730
rect 7564 23666 7616 23672
rect 7472 23520 7524 23526
rect 7472 23462 7524 23468
rect 7380 22772 7432 22778
rect 7380 22714 7432 22720
rect 7484 22642 7512 23462
rect 7472 22636 7524 22642
rect 7472 22578 7524 22584
rect 7576 22522 7604 23666
rect 7656 23520 7708 23526
rect 7656 23462 7708 23468
rect 7484 22494 7604 22522
rect 7380 22228 7432 22234
rect 7380 22170 7432 22176
rect 7288 22160 7340 22166
rect 7288 22102 7340 22108
rect 7392 21554 7420 22170
rect 7380 21548 7432 21554
rect 7380 21490 7432 21496
rect 7286 21312 7342 21321
rect 7208 21270 7286 21298
rect 7286 21247 7342 21256
rect 7116 20896 7236 20924
rect 7104 20800 7156 20806
rect 6918 20768 6974 20777
rect 7104 20742 7156 20748
rect 6918 20703 6974 20712
rect 7116 20618 7144 20742
rect 6840 20602 7144 20618
rect 6828 20596 7144 20602
rect 6880 20590 7144 20596
rect 6828 20538 6880 20544
rect 6736 20528 6788 20534
rect 6736 20470 6788 20476
rect 6564 20330 6684 20346
rect 6460 20324 6512 20330
rect 6460 20266 6512 20272
rect 6552 20324 6684 20330
rect 6604 20318 6684 20324
rect 6552 20266 6604 20272
rect 6092 20052 6144 20058
rect 6092 19994 6144 20000
rect 6104 19768 6132 19994
rect 6184 19780 6236 19786
rect 6104 19740 6184 19768
rect 6472 19768 6500 20266
rect 6644 20256 6696 20262
rect 6644 20198 6696 20204
rect 6656 19854 6684 20198
rect 6644 19848 6696 19854
rect 6644 19790 6696 19796
rect 6472 19740 6592 19768
rect 6184 19722 6236 19728
rect 6564 19700 6592 19740
rect 6564 19672 6684 19700
rect 6148 19612 6456 19621
rect 6148 19610 6154 19612
rect 6210 19610 6234 19612
rect 6290 19610 6314 19612
rect 6370 19610 6394 19612
rect 6450 19610 6456 19612
rect 6210 19558 6212 19610
rect 6392 19558 6394 19610
rect 6148 19556 6154 19558
rect 6210 19556 6234 19558
rect 6290 19556 6314 19558
rect 6370 19556 6394 19558
rect 6450 19556 6456 19558
rect 6148 19547 6456 19556
rect 6552 19508 6604 19514
rect 6552 19450 6604 19456
rect 6148 18524 6456 18533
rect 6148 18522 6154 18524
rect 6210 18522 6234 18524
rect 6290 18522 6314 18524
rect 6370 18522 6394 18524
rect 6450 18522 6456 18524
rect 6210 18470 6212 18522
rect 6392 18470 6394 18522
rect 6148 18468 6154 18470
rect 6210 18468 6234 18470
rect 6290 18468 6314 18470
rect 6370 18468 6394 18470
rect 6450 18468 6456 18470
rect 6148 18459 6456 18468
rect 6564 17954 6592 19450
rect 6656 18601 6684 19672
rect 6642 18592 6698 18601
rect 6642 18527 6698 18536
rect 6748 18426 6776 20470
rect 6736 18420 6788 18426
rect 6736 18362 6788 18368
rect 6472 17926 6592 17954
rect 6182 17912 6238 17921
rect 6092 17876 6144 17882
rect 6182 17847 6184 17856
rect 6092 17818 6144 17824
rect 6236 17847 6238 17856
rect 6184 17818 6236 17824
rect 6104 17542 6132 17818
rect 6472 17796 6500 17926
rect 6736 17808 6788 17814
rect 6472 17768 6592 17796
rect 6092 17536 6144 17542
rect 6092 17478 6144 17484
rect 6148 17436 6456 17445
rect 6148 17434 6154 17436
rect 6210 17434 6234 17436
rect 6290 17434 6314 17436
rect 6370 17434 6394 17436
rect 6450 17434 6456 17436
rect 6210 17382 6212 17434
rect 6392 17382 6394 17434
rect 6148 17380 6154 17382
rect 6210 17380 6234 17382
rect 6290 17380 6314 17382
rect 6370 17380 6394 17382
rect 6450 17380 6456 17382
rect 6148 17371 6456 17380
rect 5828 17190 6040 17218
rect 6564 17218 6592 17768
rect 6736 17750 6788 17756
rect 6564 17190 6684 17218
rect 5724 15020 5776 15026
rect 5724 14962 5776 14968
rect 5722 14920 5778 14929
rect 5722 14855 5778 14864
rect 5632 14068 5684 14074
rect 5632 14010 5684 14016
rect 5540 13524 5592 13530
rect 5540 13466 5592 13472
rect 5736 13410 5764 14855
rect 5552 13382 5764 13410
rect 5828 13410 5856 17190
rect 6000 17128 6052 17134
rect 6000 17070 6052 17076
rect 6552 17128 6604 17134
rect 6552 17070 6604 17076
rect 5906 16688 5962 16697
rect 5906 16623 5908 16632
rect 5960 16623 5962 16632
rect 5908 16594 5960 16600
rect 6012 16182 6040 17070
rect 6092 16584 6144 16590
rect 6092 16526 6144 16532
rect 6104 16454 6132 16526
rect 6092 16448 6144 16454
rect 6092 16390 6144 16396
rect 6148 16348 6456 16357
rect 6148 16346 6154 16348
rect 6210 16346 6234 16348
rect 6290 16346 6314 16348
rect 6370 16346 6394 16348
rect 6450 16346 6456 16348
rect 6210 16294 6212 16346
rect 6392 16294 6394 16346
rect 6148 16292 6154 16294
rect 6210 16292 6234 16294
rect 6290 16292 6314 16294
rect 6370 16292 6394 16294
rect 6450 16292 6456 16294
rect 6148 16283 6456 16292
rect 6000 16176 6052 16182
rect 6000 16118 6052 16124
rect 5908 15496 5960 15502
rect 5908 15438 5960 15444
rect 5920 15162 5948 15438
rect 6000 15360 6052 15366
rect 5998 15328 6000 15337
rect 6052 15328 6054 15337
rect 5998 15263 6054 15272
rect 6148 15260 6456 15269
rect 6148 15258 6154 15260
rect 6210 15258 6234 15260
rect 6290 15258 6314 15260
rect 6370 15258 6394 15260
rect 6450 15258 6456 15260
rect 6210 15206 6212 15258
rect 6392 15206 6394 15258
rect 6148 15204 6154 15206
rect 6210 15204 6234 15206
rect 6290 15204 6314 15206
rect 6370 15204 6394 15206
rect 6450 15204 6456 15206
rect 6148 15195 6456 15204
rect 5908 15156 5960 15162
rect 5908 15098 5960 15104
rect 6092 14952 6144 14958
rect 6092 14894 6144 14900
rect 6368 14952 6420 14958
rect 6368 14894 6420 14900
rect 5908 14408 5960 14414
rect 5908 14350 5960 14356
rect 5920 13734 5948 14350
rect 6104 14260 6132 14894
rect 6380 14550 6408 14894
rect 6564 14822 6592 17070
rect 6552 14816 6604 14822
rect 6458 14784 6514 14793
rect 6552 14758 6604 14764
rect 6458 14719 6514 14728
rect 6472 14618 6500 14719
rect 6460 14612 6512 14618
rect 6460 14554 6512 14560
rect 6368 14544 6420 14550
rect 6368 14486 6420 14492
rect 6552 14476 6604 14482
rect 6552 14418 6604 14424
rect 6058 14232 6132 14260
rect 6058 13988 6086 14232
rect 6148 14172 6456 14181
rect 6148 14170 6154 14172
rect 6210 14170 6234 14172
rect 6290 14170 6314 14172
rect 6370 14170 6394 14172
rect 6450 14170 6456 14172
rect 6210 14118 6212 14170
rect 6392 14118 6394 14170
rect 6148 14116 6154 14118
rect 6210 14116 6234 14118
rect 6290 14116 6314 14118
rect 6370 14116 6394 14118
rect 6450 14116 6456 14118
rect 6148 14107 6456 14116
rect 6564 14006 6592 14418
rect 6012 13960 6086 13988
rect 6276 14000 6328 14006
rect 5908 13728 5960 13734
rect 5908 13670 5960 13676
rect 5906 13560 5962 13569
rect 6012 13546 6040 13960
rect 6552 14000 6604 14006
rect 6276 13942 6328 13948
rect 6472 13960 6552 13988
rect 5962 13518 6040 13546
rect 5906 13495 5962 13504
rect 6288 13433 6316 13942
rect 6274 13424 6330 13433
rect 5828 13382 5948 13410
rect 5552 12356 5580 13382
rect 5724 13320 5776 13326
rect 5722 13288 5724 13297
rect 5816 13320 5868 13326
rect 5776 13288 5778 13297
rect 5816 13262 5868 13268
rect 5722 13223 5778 13232
rect 5632 13184 5684 13190
rect 5632 13126 5684 13132
rect 5724 13184 5776 13190
rect 5724 13126 5776 13132
rect 5644 12646 5672 13126
rect 5736 12850 5764 13126
rect 5828 12918 5856 13262
rect 5816 12912 5868 12918
rect 5816 12854 5868 12860
rect 5724 12844 5776 12850
rect 5724 12786 5776 12792
rect 5920 12764 5948 13382
rect 6274 13359 6330 13368
rect 6288 13326 6316 13359
rect 6276 13320 6328 13326
rect 6276 13262 6328 13268
rect 6472 13190 6500 13960
rect 6552 13942 6604 13948
rect 6552 13864 6604 13870
rect 6552 13806 6604 13812
rect 6460 13184 6512 13190
rect 6460 13126 6512 13132
rect 6148 13084 6456 13093
rect 6148 13082 6154 13084
rect 6210 13082 6234 13084
rect 6290 13082 6314 13084
rect 6370 13082 6394 13084
rect 6450 13082 6456 13084
rect 6210 13030 6212 13082
rect 6392 13030 6394 13082
rect 6148 13028 6154 13030
rect 6210 13028 6234 13030
rect 6290 13028 6314 13030
rect 6370 13028 6394 13030
rect 6450 13028 6456 13030
rect 6148 13019 6456 13028
rect 6564 12900 6592 13806
rect 6472 12872 6592 12900
rect 6276 12844 6328 12850
rect 6276 12786 6328 12792
rect 5828 12736 5948 12764
rect 5724 12708 5776 12714
rect 5724 12650 5776 12656
rect 5632 12640 5684 12646
rect 5632 12582 5684 12588
rect 5736 12481 5764 12650
rect 5722 12472 5778 12481
rect 5722 12407 5778 12416
rect 5552 12328 5764 12356
rect 5632 12232 5684 12238
rect 5632 12174 5684 12180
rect 5644 11898 5672 12174
rect 5632 11892 5684 11898
rect 5632 11834 5684 11840
rect 5644 11801 5672 11834
rect 5630 11792 5686 11801
rect 5630 11727 5686 11736
rect 5736 11558 5764 12328
rect 5724 11552 5776 11558
rect 5724 11494 5776 11500
rect 5828 11506 5856 12736
rect 6288 12345 6316 12786
rect 6368 12640 6420 12646
rect 6368 12582 6420 12588
rect 6274 12336 6330 12345
rect 6274 12271 6330 12280
rect 6380 12102 6408 12582
rect 6472 12442 6500 12872
rect 6552 12776 6604 12782
rect 6552 12718 6604 12724
rect 6460 12436 6512 12442
rect 6460 12378 6512 12384
rect 6368 12096 6420 12102
rect 5998 12064 6054 12073
rect 6368 12038 6420 12044
rect 5998 11999 6054 12008
rect 6012 11830 6040 11999
rect 6148 11996 6456 12005
rect 6148 11994 6154 11996
rect 6210 11994 6234 11996
rect 6290 11994 6314 11996
rect 6370 11994 6394 11996
rect 6450 11994 6456 11996
rect 6210 11942 6212 11994
rect 6392 11942 6394 11994
rect 6148 11940 6154 11942
rect 6210 11940 6234 11942
rect 6290 11940 6314 11942
rect 6370 11940 6394 11942
rect 6450 11940 6456 11942
rect 6148 11931 6456 11940
rect 6564 11898 6592 12718
rect 6552 11892 6604 11898
rect 6552 11834 6604 11840
rect 5908 11824 5960 11830
rect 5908 11766 5960 11772
rect 6000 11824 6052 11830
rect 6000 11766 6052 11772
rect 6656 11778 6684 17190
rect 6748 16794 6776 17750
rect 6840 17728 6868 20538
rect 6920 20392 6972 20398
rect 6920 20334 6972 20340
rect 7012 20392 7064 20398
rect 7012 20334 7064 20340
rect 7104 20392 7156 20398
rect 7104 20334 7156 20340
rect 6932 19854 6960 20334
rect 6920 19848 6972 19854
rect 6920 19790 6972 19796
rect 7024 19514 7052 20334
rect 7012 19508 7064 19514
rect 7012 19450 7064 19456
rect 6920 19168 6972 19174
rect 6920 19110 6972 19116
rect 6932 18426 6960 19110
rect 7116 18970 7144 20334
rect 7104 18964 7156 18970
rect 7104 18906 7156 18912
rect 7104 18692 7156 18698
rect 7104 18634 7156 18640
rect 7116 18465 7144 18634
rect 7102 18456 7158 18465
rect 6920 18420 6972 18426
rect 7102 18391 7158 18400
rect 6920 18362 6972 18368
rect 7208 18329 7236 20896
rect 7286 20632 7342 20641
rect 7286 20567 7342 20576
rect 7300 18902 7328 20567
rect 7392 19825 7420 21490
rect 7378 19816 7434 19825
rect 7378 19751 7434 19760
rect 7288 18896 7340 18902
rect 7288 18838 7340 18844
rect 7194 18320 7250 18329
rect 7104 18284 7156 18290
rect 7194 18255 7250 18264
rect 7104 18226 7156 18232
rect 7116 18193 7144 18226
rect 7102 18184 7158 18193
rect 7102 18119 7158 18128
rect 7010 17912 7066 17921
rect 7010 17847 7066 17856
rect 7024 17746 7052 17847
rect 7012 17740 7064 17746
rect 6840 17700 6960 17728
rect 6828 17604 6880 17610
rect 6828 17546 6880 17552
rect 6840 16794 6868 17546
rect 6736 16788 6788 16794
rect 6736 16730 6788 16736
rect 6828 16788 6880 16794
rect 6828 16730 6880 16736
rect 6932 16674 6960 17700
rect 7012 17682 7064 17688
rect 7010 17640 7066 17649
rect 7010 17575 7012 17584
rect 7064 17575 7066 17584
rect 7012 17546 7064 17552
rect 7024 17270 7052 17546
rect 7012 17264 7064 17270
rect 7012 17206 7064 17212
rect 7024 16726 7052 17206
rect 6840 16646 6960 16674
rect 7012 16720 7064 16726
rect 7012 16662 7064 16668
rect 6736 16516 6788 16522
rect 6736 16458 6788 16464
rect 6748 15434 6776 16458
rect 6736 15428 6788 15434
rect 6736 15370 6788 15376
rect 6748 14482 6776 15370
rect 6736 14476 6788 14482
rect 6736 14418 6788 14424
rect 6734 14376 6790 14385
rect 6734 14311 6790 14320
rect 6748 11898 6776 14311
rect 6840 12374 6868 16646
rect 7012 16584 7064 16590
rect 7012 16526 7064 16532
rect 6920 16516 6972 16522
rect 6920 16458 6972 16464
rect 6932 16114 6960 16458
rect 7024 16114 7052 16526
rect 6920 16108 6972 16114
rect 6920 16050 6972 16056
rect 7012 16108 7064 16114
rect 7012 16050 7064 16056
rect 7012 15360 7064 15366
rect 7012 15302 7064 15308
rect 6920 14884 6972 14890
rect 6920 14826 6972 14832
rect 6932 12481 6960 14826
rect 7024 14550 7052 15302
rect 7012 14544 7064 14550
rect 7012 14486 7064 14492
rect 7024 14006 7052 14486
rect 7116 14346 7144 18119
rect 7288 18080 7340 18086
rect 7288 18022 7340 18028
rect 7196 17740 7248 17746
rect 7196 17682 7248 17688
rect 7208 16250 7236 17682
rect 7300 16250 7328 18022
rect 7392 17513 7420 19751
rect 7484 18290 7512 22494
rect 7562 22264 7618 22273
rect 7562 22199 7618 22208
rect 7576 21486 7604 22199
rect 7564 21480 7616 21486
rect 7564 21422 7616 21428
rect 7668 20534 7696 23462
rect 7760 23322 7788 24006
rect 7748 23316 7800 23322
rect 7748 23258 7800 23264
rect 7748 23112 7800 23118
rect 7748 23054 7800 23060
rect 7760 22438 7788 23054
rect 7748 22432 7800 22438
rect 7748 22374 7800 22380
rect 7748 22024 7800 22030
rect 7748 21966 7800 21972
rect 7760 21690 7788 21966
rect 7748 21684 7800 21690
rect 7748 21626 7800 21632
rect 7748 21004 7800 21010
rect 7748 20946 7800 20952
rect 7656 20528 7708 20534
rect 7656 20470 7708 20476
rect 7564 19168 7616 19174
rect 7564 19110 7616 19116
rect 7576 18698 7604 19110
rect 7564 18692 7616 18698
rect 7564 18634 7616 18640
rect 7564 18420 7616 18426
rect 7564 18362 7616 18368
rect 7472 18284 7524 18290
rect 7472 18226 7524 18232
rect 7484 17678 7512 18226
rect 7576 17678 7604 18362
rect 7472 17672 7524 17678
rect 7472 17614 7524 17620
rect 7564 17672 7616 17678
rect 7564 17614 7616 17620
rect 7378 17504 7434 17513
rect 7378 17439 7434 17448
rect 7472 17332 7524 17338
rect 7392 17292 7472 17320
rect 7196 16244 7248 16250
rect 7196 16186 7248 16192
rect 7288 16244 7340 16250
rect 7288 16186 7340 16192
rect 7288 16108 7340 16114
rect 7288 16050 7340 16056
rect 7194 15600 7250 15609
rect 7194 15535 7250 15544
rect 7104 14340 7156 14346
rect 7104 14282 7156 14288
rect 7012 14000 7064 14006
rect 7012 13942 7064 13948
rect 7024 13002 7052 13942
rect 7104 13932 7156 13938
rect 7104 13874 7156 13880
rect 7116 13530 7144 13874
rect 7104 13524 7156 13530
rect 7104 13466 7156 13472
rect 7024 12974 7144 13002
rect 7116 12918 7144 12974
rect 7104 12912 7156 12918
rect 7104 12854 7156 12860
rect 7012 12844 7064 12850
rect 7012 12786 7064 12792
rect 6918 12472 6974 12481
rect 7024 12442 7052 12786
rect 6918 12407 6974 12416
rect 7012 12436 7064 12442
rect 7012 12378 7064 12384
rect 6828 12368 6880 12374
rect 7208 12322 7236 15535
rect 7300 14793 7328 16050
rect 7392 15434 7420 17292
rect 7472 17274 7524 17280
rect 7564 17264 7616 17270
rect 7564 17206 7616 17212
rect 7472 17196 7524 17202
rect 7472 17138 7524 17144
rect 7484 15434 7512 17138
rect 7576 16794 7604 17206
rect 7564 16788 7616 16794
rect 7564 16730 7616 16736
rect 7564 16448 7616 16454
rect 7564 16390 7616 16396
rect 7380 15428 7432 15434
rect 7380 15370 7432 15376
rect 7472 15428 7524 15434
rect 7472 15370 7524 15376
rect 7392 15162 7420 15370
rect 7576 15366 7604 16390
rect 7564 15360 7616 15366
rect 7564 15302 7616 15308
rect 7380 15156 7432 15162
rect 7380 15098 7432 15104
rect 7286 14784 7342 14793
rect 7286 14719 7342 14728
rect 7288 14272 7340 14278
rect 7288 14214 7340 14220
rect 7300 13462 7328 14214
rect 7392 13938 7420 15098
rect 7472 14952 7524 14958
rect 7472 14894 7524 14900
rect 7564 14952 7616 14958
rect 7564 14894 7616 14900
rect 7484 14822 7512 14894
rect 7472 14816 7524 14822
rect 7472 14758 7524 14764
rect 7576 14634 7604 14894
rect 7484 14618 7604 14634
rect 7472 14612 7604 14618
rect 7524 14606 7604 14612
rect 7472 14554 7524 14560
rect 7380 13932 7432 13938
rect 7380 13874 7432 13880
rect 7564 13932 7616 13938
rect 7564 13874 7616 13880
rect 7288 13456 7340 13462
rect 7288 13398 7340 13404
rect 7286 13016 7342 13025
rect 7286 12951 7342 12960
rect 7300 12850 7328 12951
rect 7392 12918 7420 13874
rect 7472 13388 7524 13394
rect 7472 13330 7524 13336
rect 7380 12912 7432 12918
rect 7378 12880 7380 12889
rect 7432 12880 7434 12889
rect 7288 12844 7340 12850
rect 7378 12815 7434 12824
rect 7288 12786 7340 12792
rect 7484 12594 7512 13330
rect 7576 12918 7604 13874
rect 7564 12912 7616 12918
rect 7564 12854 7616 12860
rect 6828 12310 6880 12316
rect 6932 12294 7236 12322
rect 7300 12566 7512 12594
rect 7300 12306 7328 12566
rect 7472 12436 7524 12442
rect 7472 12378 7524 12384
rect 7378 12336 7434 12345
rect 7288 12300 7340 12306
rect 6828 12096 6880 12102
rect 6828 12038 6880 12044
rect 6736 11892 6788 11898
rect 6736 11834 6788 11840
rect 5920 11608 5948 11766
rect 6276 11756 6328 11762
rect 6656 11750 6776 11778
rect 6328 11716 6592 11744
rect 6276 11698 6328 11704
rect 5920 11580 6040 11608
rect 5828 11478 5930 11506
rect 5448 11212 5500 11218
rect 5448 11154 5500 11160
rect 5540 11212 5592 11218
rect 5592 11172 5672 11200
rect 5540 11154 5592 11160
rect 5460 11098 5488 11154
rect 5460 11070 5580 11098
rect 5552 10996 5580 11070
rect 5460 10968 5580 10996
rect 5356 10668 5408 10674
rect 5276 10628 5356 10656
rect 5356 10610 5408 10616
rect 5184 10084 5304 10112
rect 5078 10024 5134 10033
rect 5078 9959 5134 9968
rect 5078 9888 5134 9897
rect 5078 9823 5134 9832
rect 5092 9722 5120 9823
rect 5080 9716 5132 9722
rect 5080 9658 5132 9664
rect 5276 9586 5304 10084
rect 5460 9586 5488 10968
rect 5644 10792 5672 11172
rect 5902 10996 5930 11478
rect 6012 11218 6040 11580
rect 6564 11540 6592 11716
rect 6644 11552 6696 11558
rect 6366 11520 6422 11529
rect 6564 11512 6644 11540
rect 6422 11478 6500 11506
rect 6644 11494 6696 11500
rect 6366 11455 6422 11464
rect 6472 11218 6500 11478
rect 6000 11212 6052 11218
rect 6000 11154 6052 11160
rect 6460 11212 6512 11218
rect 6460 11154 6512 11160
rect 6092 11144 6144 11150
rect 6092 11086 6144 11092
rect 6104 10996 6132 11086
rect 5828 10968 5930 10996
rect 6012 10968 6132 10996
rect 6644 11008 6696 11014
rect 5644 10764 5764 10792
rect 5630 10704 5686 10713
rect 5540 10668 5592 10674
rect 5630 10639 5686 10648
rect 5540 10610 5592 10616
rect 5552 9602 5580 10610
rect 5644 9761 5672 10639
rect 5736 10470 5764 10764
rect 5724 10464 5776 10470
rect 5724 10406 5776 10412
rect 5630 9752 5686 9761
rect 5630 9687 5686 9696
rect 5722 9616 5778 9625
rect 5264 9580 5316 9586
rect 5264 9522 5316 9528
rect 5448 9580 5500 9586
rect 5552 9574 5672 9602
rect 5448 9522 5500 9528
rect 5540 9512 5592 9518
rect 5540 9454 5592 9460
rect 5080 9444 5132 9450
rect 5080 9386 5132 9392
rect 4988 8084 5040 8090
rect 4988 8026 5040 8032
rect 4988 7404 5040 7410
rect 4988 7346 5040 7352
rect 5000 7041 5028 7346
rect 4986 7032 5042 7041
rect 4986 6967 5042 6976
rect 4988 6656 5040 6662
rect 4988 6598 5040 6604
rect 5000 6474 5028 6598
rect 4966 6446 5028 6474
rect 5092 6458 5120 9386
rect 5448 9036 5500 9042
rect 5448 8978 5500 8984
rect 5354 8664 5410 8673
rect 5354 8599 5410 8608
rect 5264 8288 5316 8294
rect 5184 8236 5264 8242
rect 5184 8230 5316 8236
rect 5184 8214 5304 8230
rect 5080 6452 5132 6458
rect 4966 6338 4994 6446
rect 5080 6394 5132 6400
rect 4966 6310 5028 6338
rect 4896 5568 4948 5574
rect 4896 5510 4948 5516
rect 4896 5160 4948 5166
rect 4896 5102 4948 5108
rect 4908 5001 4936 5102
rect 4894 4992 4950 5001
rect 4894 4927 4950 4936
rect 4712 4820 4764 4826
rect 4712 4762 4764 4768
rect 4804 4820 4856 4826
rect 4804 4762 4856 4768
rect 5000 4706 5028 6310
rect 5080 6316 5132 6322
rect 5080 6258 5132 6264
rect 5092 5234 5120 6258
rect 5080 5228 5132 5234
rect 5080 5170 5132 5176
rect 4540 4678 5028 4706
rect 4342 4584 4398 4593
rect 4342 4519 4344 4528
rect 4396 4519 4398 4528
rect 4344 4490 4396 4496
rect 4344 4208 4396 4214
rect 4344 4150 4396 4156
rect 4252 2848 4304 2854
rect 4252 2790 4304 2796
rect 4356 2666 4384 4150
rect 4436 3392 4488 3398
rect 4436 3334 4488 3340
rect 4448 3126 4476 3334
rect 4436 3120 4488 3126
rect 4436 3062 4488 3068
rect 4160 2644 4212 2650
rect 3884 2440 3936 2446
rect 3884 2382 3936 2388
rect 3700 2304 3752 2310
rect 3700 2246 3752 2252
rect 3424 1964 3476 1970
rect 3424 1906 3476 1912
rect 3332 1420 3384 1426
rect 3332 1362 3384 1368
rect 3332 1284 3384 1290
rect 3332 1226 3384 1232
rect 3344 1193 3372 1226
rect 3330 1184 3386 1193
rect 3330 1119 3386 1128
rect 3332 740 3384 746
rect 3332 682 3384 688
rect 3344 160 3372 682
rect 3146 54 3280 82
rect 3146 -300 3202 54
rect 3330 -300 3386 160
rect 3436 82 3464 1906
rect 3712 1834 3740 2246
rect 3988 2106 4016 2638
rect 4160 2586 4212 2592
rect 4264 2638 4384 2666
rect 4540 2650 4568 4678
rect 5092 4622 5120 5170
rect 5080 4616 5132 4622
rect 4986 4584 5042 4593
rect 5080 4558 5132 4564
rect 4986 4519 5042 4528
rect 4804 4276 4856 4282
rect 4804 4218 4856 4224
rect 4620 3936 4672 3942
rect 4620 3878 4672 3884
rect 4528 2644 4580 2650
rect 4158 2544 4214 2553
rect 4158 2479 4214 2488
rect 4172 2446 4200 2479
rect 4160 2440 4212 2446
rect 4160 2382 4212 2388
rect 4160 2304 4212 2310
rect 4160 2246 4212 2252
rect 3976 2100 4028 2106
rect 3976 2042 4028 2048
rect 3884 1964 3936 1970
rect 3884 1906 3936 1912
rect 3700 1828 3752 1834
rect 3700 1770 3752 1776
rect 3549 1660 3857 1669
rect 3549 1658 3555 1660
rect 3611 1658 3635 1660
rect 3691 1658 3715 1660
rect 3771 1658 3795 1660
rect 3851 1658 3857 1660
rect 3611 1606 3613 1658
rect 3793 1606 3795 1658
rect 3549 1604 3555 1606
rect 3611 1604 3635 1606
rect 3691 1604 3715 1606
rect 3771 1604 3795 1606
rect 3851 1604 3857 1606
rect 3549 1595 3857 1604
rect 3700 1352 3752 1358
rect 3514 1320 3570 1329
rect 3700 1294 3752 1300
rect 3514 1255 3570 1264
rect 3528 1222 3556 1255
rect 3516 1216 3568 1222
rect 3516 1158 3568 1164
rect 3712 160 3740 1294
rect 3896 160 3924 1906
rect 4172 1204 4200 2246
rect 4264 1426 4292 2638
rect 4528 2586 4580 2592
rect 4632 2530 4660 3878
rect 4540 2502 4660 2530
rect 4436 2440 4488 2446
rect 4356 2400 4436 2428
rect 4252 1420 4304 1426
rect 4252 1362 4304 1368
rect 4080 1176 4200 1204
rect 4252 1216 4304 1222
rect 4080 160 4108 1176
rect 4252 1158 4304 1164
rect 4264 160 4292 1158
rect 4356 1018 4384 2400
rect 4436 2382 4488 2388
rect 4540 2106 4568 2502
rect 4816 2446 4844 4218
rect 4804 2440 4856 2446
rect 4804 2382 4856 2388
rect 4620 2372 4672 2378
rect 4620 2314 4672 2320
rect 4528 2100 4580 2106
rect 4632 2088 4660 2314
rect 4802 2272 4858 2281
rect 4802 2207 4858 2216
rect 4816 2106 4844 2207
rect 4804 2100 4856 2106
rect 4632 2060 4752 2088
rect 4528 2042 4580 2048
rect 4620 1964 4672 1970
rect 4448 1924 4620 1952
rect 4344 1012 4396 1018
rect 4344 954 4396 960
rect 4448 160 4476 1924
rect 4620 1906 4672 1912
rect 4724 1408 4752 2060
rect 4804 2042 4856 2048
rect 4804 1964 4856 1970
rect 4804 1906 4856 1912
rect 4896 1964 4948 1970
rect 4896 1906 4948 1912
rect 4632 1380 4752 1408
rect 4528 1352 4580 1358
rect 4528 1294 4580 1300
rect 4540 746 4568 1294
rect 4528 740 4580 746
rect 4528 682 4580 688
rect 4632 160 4660 1380
rect 4816 1340 4844 1906
rect 4724 1312 4844 1340
rect 4724 950 4752 1312
rect 4804 1216 4856 1222
rect 4804 1158 4856 1164
rect 4712 944 4764 950
rect 4712 886 4764 892
rect 4816 785 4844 1158
rect 4802 776 4858 785
rect 4802 711 4858 720
rect 3514 82 3570 160
rect 3436 54 3570 82
rect 3514 -300 3570 54
rect 3698 -300 3754 160
rect 3882 -300 3938 160
rect 4066 -300 4122 160
rect 4250 -300 4306 160
rect 4434 -300 4490 160
rect 4618 -300 4674 160
rect 4802 82 4858 160
rect 4908 82 4936 1906
rect 5000 1834 5028 4519
rect 5184 4486 5212 8214
rect 5262 8120 5318 8129
rect 5262 8055 5318 8064
rect 5276 6361 5304 8055
rect 5368 7478 5396 8599
rect 5356 7472 5408 7478
rect 5356 7414 5408 7420
rect 5460 7177 5488 8978
rect 5552 8498 5580 9454
rect 5644 9178 5672 9574
rect 5722 9551 5778 9560
rect 5736 9518 5764 9551
rect 5724 9512 5776 9518
rect 5724 9454 5776 9460
rect 5722 9344 5778 9353
rect 5722 9279 5778 9288
rect 5632 9172 5684 9178
rect 5632 9114 5684 9120
rect 5540 8492 5592 8498
rect 5540 8434 5592 8440
rect 5632 8084 5684 8090
rect 5632 8026 5684 8032
rect 5540 7812 5592 7818
rect 5540 7754 5592 7760
rect 5552 7546 5580 7754
rect 5540 7540 5592 7546
rect 5540 7482 5592 7488
rect 5540 7404 5592 7410
rect 5540 7346 5592 7352
rect 5446 7168 5502 7177
rect 5446 7103 5502 7112
rect 5446 6896 5502 6905
rect 5446 6831 5502 6840
rect 5356 6792 5408 6798
rect 5356 6734 5408 6740
rect 5262 6352 5318 6361
rect 5262 6287 5318 6296
rect 5264 5704 5316 5710
rect 5264 5646 5316 5652
rect 5172 4480 5224 4486
rect 5172 4422 5224 4428
rect 5276 4078 5304 5646
rect 5368 5370 5396 6734
rect 5460 6633 5488 6831
rect 5446 6624 5502 6633
rect 5446 6559 5502 6568
rect 5552 6458 5580 7346
rect 5540 6452 5592 6458
rect 5540 6394 5592 6400
rect 5644 6338 5672 8026
rect 5552 6310 5672 6338
rect 5552 5658 5580 6310
rect 5632 5908 5684 5914
rect 5632 5850 5684 5856
rect 5460 5630 5580 5658
rect 5356 5364 5408 5370
rect 5356 5306 5408 5312
rect 5356 4548 5408 4554
rect 5356 4490 5408 4496
rect 5264 4072 5316 4078
rect 5170 4040 5226 4049
rect 5264 4014 5316 4020
rect 5170 3975 5226 3984
rect 5184 2650 5212 3975
rect 5262 3632 5318 3641
rect 5262 3567 5318 3576
rect 5172 2644 5224 2650
rect 5172 2586 5224 2592
rect 5276 1986 5304 3567
rect 5368 2650 5396 4490
rect 5460 4146 5488 5630
rect 5540 4480 5592 4486
rect 5540 4422 5592 4428
rect 5448 4140 5500 4146
rect 5448 4082 5500 4088
rect 5448 4004 5500 4010
rect 5448 3946 5500 3952
rect 5460 3233 5488 3946
rect 5446 3224 5502 3233
rect 5446 3159 5502 3168
rect 5446 3088 5502 3097
rect 5446 3023 5448 3032
rect 5500 3023 5502 3032
rect 5448 2994 5500 3000
rect 5356 2644 5408 2650
rect 5356 2586 5408 2592
rect 5446 2272 5502 2281
rect 5446 2207 5502 2216
rect 5184 1958 5304 1986
rect 4988 1828 5040 1834
rect 4988 1770 5040 1776
rect 4988 1352 5040 1358
rect 4988 1294 5040 1300
rect 5080 1352 5132 1358
rect 5184 1340 5212 1958
rect 5460 1902 5488 2207
rect 5264 1896 5316 1902
rect 5264 1838 5316 1844
rect 5448 1896 5500 1902
rect 5448 1838 5500 1844
rect 5132 1312 5212 1340
rect 5080 1294 5132 1300
rect 5000 160 5028 1294
rect 5276 1000 5304 1838
rect 5552 1358 5580 4422
rect 5644 3738 5672 5850
rect 5736 4146 5764 9279
rect 5828 7954 5856 10968
rect 5908 10464 5960 10470
rect 5908 10406 5960 10412
rect 5920 8838 5948 10406
rect 6012 10266 6040 10968
rect 6644 10950 6696 10956
rect 6148 10908 6456 10917
rect 6148 10906 6154 10908
rect 6210 10906 6234 10908
rect 6290 10906 6314 10908
rect 6370 10906 6394 10908
rect 6450 10906 6456 10908
rect 6210 10854 6212 10906
rect 6392 10854 6394 10906
rect 6148 10852 6154 10854
rect 6210 10852 6234 10854
rect 6290 10852 6314 10854
rect 6370 10852 6394 10854
rect 6450 10852 6456 10854
rect 6148 10843 6456 10852
rect 6368 10804 6420 10810
rect 6368 10746 6420 10752
rect 6090 10704 6146 10713
rect 6090 10639 6146 10648
rect 6000 10260 6052 10266
rect 6000 10202 6052 10208
rect 6104 10010 6132 10639
rect 6380 10062 6408 10746
rect 6460 10464 6512 10470
rect 6460 10406 6512 10412
rect 6472 10062 6500 10406
rect 6550 10296 6606 10305
rect 6550 10231 6606 10240
rect 6012 9982 6132 10010
rect 6368 10056 6420 10062
rect 6368 9998 6420 10004
rect 6460 10056 6512 10062
rect 6460 9998 6512 10004
rect 5908 8832 5960 8838
rect 5908 8774 5960 8780
rect 5816 7948 5868 7954
rect 5816 7890 5868 7896
rect 6012 7324 6040 9982
rect 6148 9820 6456 9829
rect 6148 9818 6154 9820
rect 6210 9818 6234 9820
rect 6290 9818 6314 9820
rect 6370 9818 6394 9820
rect 6450 9818 6456 9820
rect 6210 9766 6212 9818
rect 6392 9766 6394 9818
rect 6148 9764 6154 9766
rect 6210 9764 6234 9766
rect 6290 9764 6314 9766
rect 6370 9764 6394 9766
rect 6450 9764 6456 9766
rect 6148 9755 6456 9764
rect 6564 9674 6592 10231
rect 6656 10130 6684 10950
rect 6644 10124 6696 10130
rect 6644 10066 6696 10072
rect 6472 9646 6592 9674
rect 6644 9716 6696 9722
rect 6644 9658 6696 9664
rect 6472 9081 6500 9646
rect 6552 9580 6604 9586
rect 6552 9522 6604 9528
rect 6458 9072 6514 9081
rect 6458 9007 6514 9016
rect 6148 8732 6456 8741
rect 6148 8730 6154 8732
rect 6210 8730 6234 8732
rect 6290 8730 6314 8732
rect 6370 8730 6394 8732
rect 6450 8730 6456 8732
rect 6210 8678 6212 8730
rect 6392 8678 6394 8730
rect 6148 8676 6154 8678
rect 6210 8676 6234 8678
rect 6290 8676 6314 8678
rect 6370 8676 6394 8678
rect 6450 8676 6456 8678
rect 6148 8667 6456 8676
rect 6274 8528 6330 8537
rect 6274 8463 6276 8472
rect 6328 8463 6330 8472
rect 6276 8434 6328 8440
rect 6368 8084 6420 8090
rect 6368 8026 6420 8032
rect 6380 7886 6408 8026
rect 6368 7880 6420 7886
rect 6368 7822 6420 7828
rect 6148 7644 6456 7653
rect 6148 7642 6154 7644
rect 6210 7642 6234 7644
rect 6290 7642 6314 7644
rect 6370 7642 6394 7644
rect 6450 7642 6456 7644
rect 6210 7590 6212 7642
rect 6392 7590 6394 7642
rect 6148 7588 6154 7590
rect 6210 7588 6234 7590
rect 6290 7588 6314 7590
rect 6370 7588 6394 7590
rect 6450 7588 6456 7590
rect 6148 7579 6456 7588
rect 5828 7296 6040 7324
rect 5828 4214 5856 7296
rect 6000 7200 6052 7206
rect 6000 7142 6052 7148
rect 6090 7168 6146 7177
rect 6012 6934 6040 7142
rect 6146 7126 6224 7154
rect 6090 7103 6146 7112
rect 6000 6928 6052 6934
rect 5906 6896 5962 6905
rect 6000 6870 6052 6876
rect 5906 6831 5908 6840
rect 5960 6831 5962 6840
rect 5908 6802 5960 6808
rect 5920 5914 5948 6802
rect 6092 6792 6144 6798
rect 6196 6780 6224 7126
rect 6144 6752 6224 6780
rect 6092 6734 6144 6740
rect 6148 6556 6456 6565
rect 6148 6554 6154 6556
rect 6210 6554 6234 6556
rect 6290 6554 6314 6556
rect 6370 6554 6394 6556
rect 6450 6554 6456 6556
rect 6210 6502 6212 6554
rect 6392 6502 6394 6554
rect 6148 6500 6154 6502
rect 6210 6500 6234 6502
rect 6290 6500 6314 6502
rect 6370 6500 6394 6502
rect 6450 6500 6456 6502
rect 6148 6491 6456 6500
rect 6368 6248 6420 6254
rect 6182 6216 6238 6225
rect 6368 6190 6420 6196
rect 6182 6151 6238 6160
rect 6000 6112 6052 6118
rect 5998 6080 6000 6089
rect 6052 6080 6054 6089
rect 5998 6015 6054 6024
rect 6196 5914 6224 6151
rect 6274 6080 6330 6089
rect 6274 6015 6330 6024
rect 5908 5908 5960 5914
rect 5908 5850 5960 5856
rect 6184 5908 6236 5914
rect 6184 5850 6236 5856
rect 6288 5642 6316 6015
rect 6276 5636 6328 5642
rect 6276 5578 6328 5584
rect 6380 5556 6408 6190
rect 6564 6118 6592 9522
rect 6656 9178 6684 9658
rect 6644 9172 6696 9178
rect 6644 9114 6696 9120
rect 6644 8832 6696 8838
rect 6644 8774 6696 8780
rect 6656 8022 6684 8774
rect 6748 8294 6776 11750
rect 6840 11150 6868 12038
rect 6828 11144 6880 11150
rect 6828 11086 6880 11092
rect 6826 10704 6882 10713
rect 6826 10639 6828 10648
rect 6880 10639 6882 10648
rect 6828 10610 6880 10616
rect 6932 10554 6960 12294
rect 7378 12271 7434 12280
rect 7288 12242 7340 12248
rect 7196 12232 7248 12238
rect 7196 12174 7248 12180
rect 7208 12073 7236 12174
rect 7288 12096 7340 12102
rect 7194 12064 7250 12073
rect 7288 12038 7340 12044
rect 7194 11999 7250 12008
rect 7104 11756 7156 11762
rect 7300 11744 7328 12038
rect 7392 11762 7420 12271
rect 7104 11698 7156 11704
rect 7208 11716 7328 11744
rect 7380 11756 7432 11762
rect 7012 11688 7064 11694
rect 7012 11630 7064 11636
rect 7024 11234 7052 11630
rect 7116 11354 7144 11698
rect 7104 11348 7156 11354
rect 7104 11290 7156 11296
rect 7024 11206 7144 11234
rect 7012 11008 7064 11014
rect 7012 10950 7064 10956
rect 6840 10526 6960 10554
rect 6840 8974 6868 10526
rect 6920 10464 6972 10470
rect 6918 10432 6920 10441
rect 6972 10432 6974 10441
rect 6918 10367 6974 10376
rect 7024 10130 7052 10950
rect 7012 10124 7064 10130
rect 7012 10066 7064 10072
rect 7010 9752 7066 9761
rect 7010 9687 7066 9696
rect 6920 9580 6972 9586
rect 6920 9522 6972 9528
rect 6932 9489 6960 9522
rect 6918 9480 6974 9489
rect 6918 9415 6974 9424
rect 6932 9042 6960 9415
rect 6920 9036 6972 9042
rect 6920 8978 6972 8984
rect 6828 8968 6880 8974
rect 6828 8910 6880 8916
rect 6736 8288 6788 8294
rect 6736 8230 6788 8236
rect 6644 8016 6696 8022
rect 6644 7958 6696 7964
rect 6840 7857 6868 8910
rect 6920 8832 6972 8838
rect 6920 8774 6972 8780
rect 6932 8412 6960 8774
rect 7024 8673 7052 9687
rect 7116 8838 7144 11206
rect 7104 8832 7156 8838
rect 7104 8774 7156 8780
rect 7010 8664 7066 8673
rect 7010 8599 7066 8608
rect 7104 8628 7156 8634
rect 7104 8570 7156 8576
rect 6932 8384 7052 8412
rect 6920 8288 6972 8294
rect 6920 8230 6972 8236
rect 6932 8090 6960 8230
rect 6920 8084 6972 8090
rect 6920 8026 6972 8032
rect 6826 7848 6882 7857
rect 6826 7783 6882 7792
rect 6734 7712 6790 7721
rect 7024 7698 7052 8384
rect 7116 7886 7144 8570
rect 7104 7880 7156 7886
rect 7102 7848 7104 7857
rect 7156 7848 7158 7857
rect 7102 7783 7158 7792
rect 7024 7670 7144 7698
rect 6734 7647 6790 7656
rect 6748 6798 6776 7647
rect 6828 7200 6880 7206
rect 6828 7142 6880 7148
rect 6918 7168 6974 7177
rect 6840 7002 6868 7142
rect 6918 7103 6974 7112
rect 6932 7002 6960 7103
rect 6828 6996 6880 7002
rect 6828 6938 6880 6944
rect 6920 6996 6972 7002
rect 6920 6938 6972 6944
rect 6736 6792 6788 6798
rect 7116 6746 7144 7670
rect 6736 6734 6788 6740
rect 7024 6718 7144 6746
rect 6828 6316 6880 6322
rect 6828 6258 6880 6264
rect 6920 6316 6972 6322
rect 6920 6258 6972 6264
rect 6642 6216 6698 6225
rect 6642 6151 6698 6160
rect 6552 6112 6604 6118
rect 6552 6054 6604 6060
rect 6656 5914 6684 6151
rect 6644 5908 6696 5914
rect 6644 5850 6696 5856
rect 6460 5704 6512 5710
rect 6512 5664 6684 5692
rect 6460 5646 6512 5652
rect 6380 5528 6592 5556
rect 6148 5468 6456 5477
rect 6148 5466 6154 5468
rect 6210 5466 6234 5468
rect 6290 5466 6314 5468
rect 6370 5466 6394 5468
rect 6450 5466 6456 5468
rect 6210 5414 6212 5466
rect 6392 5414 6394 5466
rect 6148 5412 6154 5414
rect 6210 5412 6234 5414
rect 6290 5412 6314 5414
rect 6370 5412 6394 5414
rect 6450 5412 6456 5414
rect 6148 5403 6456 5412
rect 5998 5264 6054 5273
rect 5908 5228 5960 5234
rect 6564 5234 6592 5528
rect 6656 5352 6684 5664
rect 6840 5658 6868 6258
rect 6932 5914 6960 6258
rect 6920 5908 6972 5914
rect 6920 5850 6972 5856
rect 6840 5630 6960 5658
rect 6828 5568 6880 5574
rect 6828 5510 6880 5516
rect 6656 5324 6742 5352
rect 6714 5284 6742 5324
rect 6714 5256 6776 5284
rect 5998 5199 6000 5208
rect 5908 5170 5960 5176
rect 6052 5199 6054 5208
rect 6552 5228 6604 5234
rect 6000 5170 6052 5176
rect 6552 5170 6604 5176
rect 6644 5228 6696 5234
rect 6644 5170 6696 5176
rect 5816 4208 5868 4214
rect 5816 4150 5868 4156
rect 5724 4140 5776 4146
rect 5724 4082 5776 4088
rect 5816 4072 5868 4078
rect 5816 4014 5868 4020
rect 5724 3936 5776 3942
rect 5724 3878 5776 3884
rect 5632 3732 5684 3738
rect 5632 3674 5684 3680
rect 5632 3596 5684 3602
rect 5632 3538 5684 3544
rect 5644 2553 5672 3538
rect 5736 3369 5764 3878
rect 5722 3360 5778 3369
rect 5722 3295 5778 3304
rect 5630 2544 5686 2553
rect 5630 2479 5686 2488
rect 5632 2440 5684 2446
rect 5632 2382 5684 2388
rect 5356 1352 5408 1358
rect 5356 1294 5408 1300
rect 5540 1352 5592 1358
rect 5540 1294 5592 1300
rect 5184 972 5304 1000
rect 5184 160 5212 972
rect 5368 160 5396 1294
rect 5448 1284 5500 1290
rect 5448 1226 5500 1232
rect 5460 678 5488 1226
rect 5448 672 5500 678
rect 5448 614 5500 620
rect 4802 54 4936 82
rect 4802 -300 4858 54
rect 4986 -300 5042 160
rect 5170 -300 5226 160
rect 5354 -300 5410 160
rect 5538 82 5594 160
rect 5644 82 5672 2382
rect 5722 2136 5778 2145
rect 5722 2071 5724 2080
rect 5776 2071 5778 2080
rect 5724 2042 5776 2048
rect 5828 1562 5856 4014
rect 5920 3534 5948 5170
rect 6148 4380 6456 4389
rect 6148 4378 6154 4380
rect 6210 4378 6234 4380
rect 6290 4378 6314 4380
rect 6370 4378 6394 4380
rect 6450 4378 6456 4380
rect 6210 4326 6212 4378
rect 6392 4326 6394 4378
rect 6148 4324 6154 4326
rect 6210 4324 6234 4326
rect 6290 4324 6314 4326
rect 6370 4324 6394 4326
rect 6450 4324 6456 4326
rect 6148 4315 6456 4324
rect 6092 4208 6144 4214
rect 6092 4150 6144 4156
rect 5908 3528 5960 3534
rect 5908 3470 5960 3476
rect 6104 3380 6132 4150
rect 6552 4140 6604 4146
rect 6552 4082 6604 4088
rect 6012 3352 6132 3380
rect 6012 3194 6040 3352
rect 6148 3292 6456 3301
rect 6148 3290 6154 3292
rect 6210 3290 6234 3292
rect 6290 3290 6314 3292
rect 6370 3290 6394 3292
rect 6450 3290 6456 3292
rect 6210 3238 6212 3290
rect 6392 3238 6394 3290
rect 6148 3236 6154 3238
rect 6210 3236 6234 3238
rect 6290 3236 6314 3238
rect 6370 3236 6394 3238
rect 6450 3236 6456 3238
rect 6148 3227 6456 3236
rect 6000 3188 6052 3194
rect 6000 3130 6052 3136
rect 6564 2836 6592 4082
rect 6656 2990 6684 5170
rect 6748 4214 6776 5256
rect 6840 4622 6868 5510
rect 6932 5166 6960 5630
rect 6920 5160 6972 5166
rect 6920 5102 6972 5108
rect 6828 4616 6880 4622
rect 6828 4558 6880 4564
rect 6736 4208 6788 4214
rect 6736 4150 6788 4156
rect 6736 3936 6788 3942
rect 6736 3878 6788 3884
rect 6748 3602 6776 3878
rect 6736 3596 6788 3602
rect 6736 3538 6788 3544
rect 6920 3596 6972 3602
rect 6920 3538 6972 3544
rect 6932 3482 6960 3538
rect 6840 3454 6960 3482
rect 7024 3466 7052 6718
rect 7104 5568 7156 5574
rect 7104 5510 7156 5516
rect 7012 3460 7064 3466
rect 6840 3194 6868 3454
rect 7012 3402 7064 3408
rect 6920 3392 6972 3398
rect 6920 3334 6972 3340
rect 6828 3188 6880 3194
rect 6828 3130 6880 3136
rect 6736 3052 6788 3058
rect 6736 2994 6788 3000
rect 6644 2984 6696 2990
rect 6644 2926 6696 2932
rect 6564 2808 6684 2836
rect 6550 2544 6606 2553
rect 6550 2479 6606 2488
rect 6274 2408 6330 2417
rect 5908 2372 5960 2378
rect 6274 2343 6276 2352
rect 5908 2314 5960 2320
rect 6328 2343 6330 2352
rect 6276 2314 6328 2320
rect 5816 1556 5868 1562
rect 5816 1498 5868 1504
rect 5724 740 5776 746
rect 5724 682 5776 688
rect 5736 160 5764 682
rect 5920 160 5948 2314
rect 6000 2304 6052 2310
rect 6000 2246 6052 2252
rect 6012 1000 6040 2246
rect 6148 2204 6456 2213
rect 6148 2202 6154 2204
rect 6210 2202 6234 2204
rect 6290 2202 6314 2204
rect 6370 2202 6394 2204
rect 6450 2202 6456 2204
rect 6210 2150 6212 2202
rect 6392 2150 6394 2202
rect 6148 2148 6154 2150
rect 6210 2148 6234 2150
rect 6290 2148 6314 2150
rect 6370 2148 6394 2150
rect 6450 2148 6456 2150
rect 6148 2139 6456 2148
rect 6564 1970 6592 2479
rect 6552 1964 6604 1970
rect 6552 1906 6604 1912
rect 6656 1562 6684 2808
rect 6644 1556 6696 1562
rect 6644 1498 6696 1504
rect 6552 1284 6604 1290
rect 6604 1244 6684 1272
rect 6552 1226 6604 1232
rect 6148 1116 6456 1125
rect 6148 1114 6154 1116
rect 6210 1114 6234 1116
rect 6290 1114 6314 1116
rect 6370 1114 6394 1116
rect 6450 1114 6456 1116
rect 6210 1062 6212 1114
rect 6392 1062 6394 1114
rect 6148 1060 6154 1062
rect 6210 1060 6234 1062
rect 6290 1060 6314 1062
rect 6370 1060 6394 1062
rect 6450 1060 6456 1062
rect 6148 1051 6456 1060
rect 6460 1012 6512 1018
rect 6012 972 6132 1000
rect 6104 160 6132 972
rect 6460 954 6512 960
rect 6184 672 6236 678
rect 6184 614 6236 620
rect 5538 54 5672 82
rect 5538 -300 5594 54
rect 5722 -300 5778 160
rect 5906 -300 5962 160
rect 6090 -300 6146 160
rect 6196 82 6224 614
rect 6472 160 6500 954
rect 6656 160 6684 1244
rect 6748 1018 6776 2994
rect 6828 2848 6880 2854
rect 6828 2790 6880 2796
rect 6840 1970 6868 2790
rect 6932 2446 6960 3334
rect 7012 3052 7064 3058
rect 7012 2994 7064 3000
rect 7024 2774 7052 2994
rect 7116 2922 7144 5510
rect 7208 3602 7236 11716
rect 7380 11698 7432 11704
rect 7288 11552 7340 11558
rect 7288 11494 7340 11500
rect 7300 11218 7328 11494
rect 7288 11212 7340 11218
rect 7288 11154 7340 11160
rect 7300 10606 7328 11154
rect 7378 10976 7434 10985
rect 7378 10911 7434 10920
rect 7288 10600 7340 10606
rect 7288 10542 7340 10548
rect 7288 10124 7340 10130
rect 7288 10066 7340 10072
rect 7300 8634 7328 10066
rect 7288 8628 7340 8634
rect 7288 8570 7340 8576
rect 7392 8129 7420 10911
rect 7378 8120 7434 8129
rect 7288 8084 7340 8090
rect 7378 8055 7434 8064
rect 7288 8026 7340 8032
rect 7300 7886 7328 8026
rect 7286 7880 7338 7886
rect 7286 7822 7338 7828
rect 7380 7880 7432 7886
rect 7380 7822 7432 7828
rect 7392 7546 7420 7822
rect 7380 7540 7432 7546
rect 7380 7482 7432 7488
rect 7380 6724 7432 6730
rect 7380 6666 7432 6672
rect 7392 6322 7420 6666
rect 7288 6316 7340 6322
rect 7288 6258 7340 6264
rect 7380 6316 7432 6322
rect 7380 6258 7432 6264
rect 7300 4554 7328 6258
rect 7378 6216 7434 6225
rect 7378 6151 7434 6160
rect 7392 5001 7420 6151
rect 7378 4992 7434 5001
rect 7378 4927 7434 4936
rect 7288 4548 7340 4554
rect 7288 4490 7340 4496
rect 7484 4049 7512 12378
rect 7576 11694 7604 12854
rect 7668 12764 7696 20470
rect 7760 13297 7788 20946
rect 7852 20534 7880 24398
rect 7944 24313 7972 30534
rect 8036 28801 8064 30654
rect 8128 29594 8156 31719
rect 8220 31686 8248 33895
rect 8208 31680 8260 31686
rect 8208 31622 8260 31628
rect 8208 31272 8260 31278
rect 8208 31214 8260 31220
rect 8220 30938 8248 31214
rect 8208 30932 8260 30938
rect 8208 30874 8260 30880
rect 8312 29646 8340 35158
rect 8404 33114 8432 39238
rect 8574 38312 8630 38321
rect 8574 38247 8630 38256
rect 8484 37664 8536 37670
rect 8482 37632 8484 37641
rect 8536 37632 8538 37641
rect 8482 37567 8538 37576
rect 8588 37126 8616 38247
rect 8576 37120 8628 37126
rect 8576 37062 8628 37068
rect 8680 36145 8708 41228
rect 8747 40828 9055 40837
rect 8747 40826 8753 40828
rect 8809 40826 8833 40828
rect 8889 40826 8913 40828
rect 8969 40826 8993 40828
rect 9049 40826 9055 40828
rect 8809 40774 8811 40826
rect 8991 40774 8993 40826
rect 8747 40772 8753 40774
rect 8809 40772 8833 40774
rect 8889 40772 8913 40774
rect 8969 40772 8993 40774
rect 9049 40772 9055 40774
rect 8747 40763 9055 40772
rect 9232 40186 9260 42502
rect 9324 41682 9352 42570
rect 9416 42226 9444 42599
rect 9496 42570 9548 42576
rect 9404 42220 9456 42226
rect 9404 42162 9456 42168
rect 9402 42120 9458 42129
rect 9402 42055 9458 42064
rect 9312 41676 9364 41682
rect 9312 41618 9364 41624
rect 9416 41614 9444 42055
rect 9404 41608 9456 41614
rect 9404 41550 9456 41556
rect 9220 40180 9272 40186
rect 9220 40122 9272 40128
rect 8747 39740 9055 39749
rect 8747 39738 8753 39740
rect 8809 39738 8833 39740
rect 8889 39738 8913 39740
rect 8969 39738 8993 39740
rect 9049 39738 9055 39740
rect 8809 39686 8811 39738
rect 8991 39686 8993 39738
rect 8747 39684 8753 39686
rect 8809 39684 8833 39686
rect 8889 39684 8913 39686
rect 8969 39684 8993 39686
rect 9049 39684 9055 39686
rect 8747 39675 9055 39684
rect 8747 38652 9055 38661
rect 9508 38654 9536 42570
rect 9588 42016 9640 42022
rect 9588 41958 9640 41964
rect 9600 41857 9628 41958
rect 9586 41848 9642 41857
rect 9586 41783 9642 41792
rect 9692 41698 9720 42842
rect 10060 42650 10088 43386
rect 10152 43364 10180 44540
rect 10336 43636 10364 44540
rect 10336 43608 10456 43636
rect 10324 43376 10376 43382
rect 10152 43336 10324 43364
rect 10324 43318 10376 43324
rect 10232 43172 10284 43178
rect 10232 43114 10284 43120
rect 9600 41682 9720 41698
rect 9588 41676 9720 41682
rect 9640 41670 9720 41676
rect 9784 42622 10088 42650
rect 9588 41618 9640 41624
rect 9680 41608 9732 41614
rect 9680 41550 9732 41556
rect 9692 41414 9720 41550
rect 9784 41449 9812 42622
rect 9864 42560 9916 42566
rect 9864 42502 9916 42508
rect 10048 42560 10100 42566
rect 10048 42502 10100 42508
rect 9876 42294 9904 42502
rect 9864 42288 9916 42294
rect 9864 42230 9916 42236
rect 9864 42016 9916 42022
rect 9864 41958 9916 41964
rect 9956 42016 10008 42022
rect 10060 41993 10088 42502
rect 10140 42152 10192 42158
rect 10140 42094 10192 42100
rect 9956 41958 10008 41964
rect 10046 41984 10102 41993
rect 9876 41478 9904 41958
rect 9864 41472 9916 41478
rect 8747 38650 8753 38652
rect 8809 38650 8833 38652
rect 8889 38650 8913 38652
rect 8969 38650 8993 38652
rect 9049 38650 9055 38652
rect 8809 38598 8811 38650
rect 8991 38598 8993 38650
rect 8747 38596 8753 38598
rect 8809 38596 8833 38598
rect 8889 38596 8913 38598
rect 8969 38596 8993 38598
rect 9049 38596 9055 38598
rect 8747 38587 9055 38596
rect 9324 38626 9536 38654
rect 9600 41386 9720 41414
rect 9770 41440 9826 41449
rect 9128 38344 9180 38350
rect 9128 38286 9180 38292
rect 8747 37564 9055 37573
rect 8747 37562 8753 37564
rect 8809 37562 8833 37564
rect 8889 37562 8913 37564
rect 8969 37562 8993 37564
rect 9049 37562 9055 37564
rect 8809 37510 8811 37562
rect 8991 37510 8993 37562
rect 8747 37508 8753 37510
rect 8809 37508 8833 37510
rect 8889 37508 8913 37510
rect 8969 37508 8993 37510
rect 9049 37508 9055 37510
rect 8747 37499 9055 37508
rect 8852 37120 8904 37126
rect 8852 37062 8904 37068
rect 8864 36786 8892 37062
rect 9140 36854 9168 38286
rect 9220 37664 9272 37670
rect 9220 37606 9272 37612
rect 9128 36848 9180 36854
rect 9128 36790 9180 36796
rect 8852 36780 8904 36786
rect 8852 36722 8904 36728
rect 8747 36476 9055 36485
rect 8747 36474 8753 36476
rect 8809 36474 8833 36476
rect 8889 36474 8913 36476
rect 8969 36474 8993 36476
rect 9049 36474 9055 36476
rect 8809 36422 8811 36474
rect 8991 36422 8993 36474
rect 8747 36420 8753 36422
rect 8809 36420 8833 36422
rect 8889 36420 8913 36422
rect 8969 36420 8993 36422
rect 9049 36420 9055 36422
rect 8747 36411 9055 36420
rect 8666 36136 8722 36145
rect 8666 36071 8722 36080
rect 8760 36032 8812 36038
rect 8760 35974 8812 35980
rect 9128 36032 9180 36038
rect 9128 35974 9180 35980
rect 8666 35864 8722 35873
rect 8666 35799 8722 35808
rect 8576 35760 8628 35766
rect 8574 35728 8576 35737
rect 8628 35728 8630 35737
rect 8574 35663 8630 35672
rect 8576 35624 8628 35630
rect 8576 35566 8628 35572
rect 8482 35456 8538 35465
rect 8482 35391 8538 35400
rect 8496 34660 8524 35391
rect 8588 34785 8616 35566
rect 8680 35086 8708 35799
rect 8772 35630 8800 35974
rect 8760 35624 8812 35630
rect 8760 35566 8812 35572
rect 8747 35388 9055 35397
rect 8747 35386 8753 35388
rect 8809 35386 8833 35388
rect 8889 35386 8913 35388
rect 8969 35386 8993 35388
rect 9049 35386 9055 35388
rect 8809 35334 8811 35386
rect 8991 35334 8993 35386
rect 8747 35332 8753 35334
rect 8809 35332 8833 35334
rect 8889 35332 8913 35334
rect 8969 35332 8993 35334
rect 9049 35332 9055 35334
rect 8747 35323 9055 35332
rect 8668 35080 8720 35086
rect 8668 35022 8720 35028
rect 8574 34776 8630 34785
rect 8574 34711 8630 34720
rect 8496 34632 8616 34660
rect 8484 34400 8536 34406
rect 8484 34342 8536 34348
rect 8496 33454 8524 34342
rect 8484 33448 8536 33454
rect 8484 33390 8536 33396
rect 8392 33108 8444 33114
rect 8392 33050 8444 33056
rect 8496 32978 8524 33390
rect 8484 32972 8536 32978
rect 8484 32914 8536 32920
rect 8392 32904 8444 32910
rect 8392 32846 8444 32852
rect 8300 29640 8352 29646
rect 8128 29566 8248 29594
rect 8300 29582 8352 29588
rect 8116 29504 8168 29510
rect 8116 29446 8168 29452
rect 8128 29102 8156 29446
rect 8116 29096 8168 29102
rect 8116 29038 8168 29044
rect 8022 28792 8078 28801
rect 8022 28727 8078 28736
rect 8116 28688 8168 28694
rect 8116 28630 8168 28636
rect 8022 28112 8078 28121
rect 8022 28047 8078 28056
rect 8036 27470 8064 28047
rect 8128 27538 8156 28630
rect 8116 27532 8168 27538
rect 8116 27474 8168 27480
rect 8024 27464 8076 27470
rect 8024 27406 8076 27412
rect 8116 27056 8168 27062
rect 8036 27016 8116 27044
rect 7930 24304 7986 24313
rect 7930 24239 7986 24248
rect 7932 24200 7984 24206
rect 7932 24142 7984 24148
rect 7944 23322 7972 24142
rect 8036 23662 8064 27016
rect 8116 26998 8168 27004
rect 8116 26920 8168 26926
rect 8116 26862 8168 26868
rect 8128 26625 8156 26862
rect 8114 26616 8170 26625
rect 8114 26551 8170 26560
rect 8116 26376 8168 26382
rect 8220 26353 8248 29566
rect 8404 29186 8432 32846
rect 8484 32768 8536 32774
rect 8484 32710 8536 32716
rect 8496 32366 8524 32710
rect 8484 32360 8536 32366
rect 8588 32337 8616 34632
rect 8747 34300 9055 34309
rect 8747 34298 8753 34300
rect 8809 34298 8833 34300
rect 8889 34298 8913 34300
rect 8969 34298 8993 34300
rect 9049 34298 9055 34300
rect 8809 34246 8811 34298
rect 8991 34246 8993 34298
rect 8747 34244 8753 34246
rect 8809 34244 8833 34246
rect 8889 34244 8913 34246
rect 8969 34244 8993 34246
rect 9049 34244 9055 34246
rect 8747 34235 9055 34244
rect 8760 34128 8812 34134
rect 8760 34070 8812 34076
rect 8772 33844 8800 34070
rect 9036 34060 9088 34066
rect 9036 34002 9088 34008
rect 8680 33816 8800 33844
rect 8484 32302 8536 32308
rect 8574 32328 8630 32337
rect 8574 32263 8630 32272
rect 8576 32224 8628 32230
rect 8576 32166 8628 32172
rect 8482 32056 8538 32065
rect 8482 31991 8538 32000
rect 8496 31822 8524 31991
rect 8484 31816 8536 31822
rect 8482 31784 8484 31793
rect 8536 31784 8538 31793
rect 8482 31719 8538 31728
rect 8588 31686 8616 32166
rect 8484 31680 8536 31686
rect 8484 31622 8536 31628
rect 8576 31680 8628 31686
rect 8576 31622 8628 31628
rect 8496 31346 8524 31622
rect 8484 31340 8536 31346
rect 8484 31282 8536 31288
rect 8482 31240 8538 31249
rect 8482 31175 8538 31184
rect 8496 31142 8524 31175
rect 8484 31136 8536 31142
rect 8484 31078 8536 31084
rect 8576 30048 8628 30054
rect 8576 29990 8628 29996
rect 8312 29158 8432 29186
rect 8588 29170 8616 29990
rect 8484 29164 8536 29170
rect 8312 28994 8340 29158
rect 8484 29106 8536 29112
rect 8576 29164 8628 29170
rect 8576 29106 8628 29112
rect 8312 28966 8432 28994
rect 8496 28966 8524 29106
rect 8298 28112 8354 28121
rect 8298 28047 8354 28056
rect 8116 26318 8168 26324
rect 8206 26344 8262 26353
rect 8128 25498 8156 26318
rect 8206 26279 8262 26288
rect 8208 26036 8260 26042
rect 8208 25978 8260 25984
rect 8116 25492 8168 25498
rect 8116 25434 8168 25440
rect 8220 25362 8248 25978
rect 8312 25401 8340 28047
rect 8404 27418 8432 28966
rect 8484 28960 8536 28966
rect 8484 28902 8536 28908
rect 8574 28928 8630 28937
rect 8496 28529 8524 28902
rect 8574 28863 8630 28872
rect 8482 28520 8538 28529
rect 8482 28455 8538 28464
rect 8484 28416 8536 28422
rect 8484 28358 8536 28364
rect 8496 27946 8524 28358
rect 8588 28150 8616 28863
rect 8680 28422 8708 33816
rect 9048 33454 9076 34002
rect 9036 33448 9088 33454
rect 9036 33390 9088 33396
rect 8747 33212 9055 33221
rect 8747 33210 8753 33212
rect 8809 33210 8833 33212
rect 8889 33210 8913 33212
rect 8969 33210 8993 33212
rect 9049 33210 9055 33212
rect 8809 33158 8811 33210
rect 8991 33158 8993 33210
rect 8747 33156 8753 33158
rect 8809 33156 8833 33158
rect 8889 33156 8913 33158
rect 8969 33156 8993 33158
rect 9049 33156 9055 33158
rect 8747 33147 9055 33156
rect 8852 32972 8904 32978
rect 8852 32914 8904 32920
rect 8864 32298 8892 32914
rect 8942 32736 8998 32745
rect 8942 32671 8998 32680
rect 8956 32570 8984 32671
rect 8944 32564 8996 32570
rect 8944 32506 8996 32512
rect 9036 32496 9088 32502
rect 9140 32484 9168 35974
rect 9232 35714 9260 37606
rect 9324 36038 9352 38626
rect 9600 38321 9628 41386
rect 9864 41414 9916 41420
rect 9770 41375 9826 41384
rect 9968 41177 9996 41958
rect 10046 41919 10102 41928
rect 9954 41168 10010 41177
rect 9954 41103 10010 41112
rect 10152 39642 10180 42094
rect 10244 41562 10272 43114
rect 10428 42702 10456 43608
rect 10520 43330 10548 44540
rect 10704 43874 10732 44540
rect 10704 43846 10824 43874
rect 10796 43364 10824 43846
rect 10888 43636 10916 44540
rect 10888 43608 11008 43636
rect 10876 43376 10928 43382
rect 10796 43336 10876 43364
rect 10520 43302 10732 43330
rect 10876 43318 10928 43324
rect 10600 43240 10652 43246
rect 10600 43182 10652 43188
rect 10416 42696 10468 42702
rect 10416 42638 10468 42644
rect 10508 42560 10560 42566
rect 10506 42528 10508 42537
rect 10560 42528 10562 42537
rect 10506 42463 10562 42472
rect 10612 42362 10640 43182
rect 10704 42702 10732 43302
rect 10784 43104 10836 43110
rect 10784 43046 10836 43052
rect 10796 42786 10824 43046
rect 10796 42758 10916 42786
rect 10692 42696 10744 42702
rect 10692 42638 10744 42644
rect 10888 42616 10916 42758
rect 10980 42702 11008 43608
rect 11072 42922 11100 44540
rect 11256 43738 11284 44540
rect 11164 43710 11284 43738
rect 11164 43330 11192 43710
rect 11440 43636 11468 44540
rect 11624 43874 11652 44540
rect 11624 43846 11744 43874
rect 11256 43608 11468 43636
rect 11256 43432 11284 43608
rect 11346 43548 11654 43557
rect 11346 43546 11352 43548
rect 11408 43546 11432 43548
rect 11488 43546 11512 43548
rect 11568 43546 11592 43548
rect 11648 43546 11654 43548
rect 11408 43494 11410 43546
rect 11590 43494 11592 43546
rect 11346 43492 11352 43494
rect 11408 43492 11432 43494
rect 11488 43492 11512 43494
rect 11568 43492 11592 43494
rect 11648 43492 11654 43494
rect 11346 43483 11654 43492
rect 11256 43404 11468 43432
rect 11164 43302 11376 43330
rect 11152 43104 11204 43110
rect 11150 43072 11152 43081
rect 11204 43072 11206 43081
rect 11150 43007 11206 43016
rect 11072 42894 11192 42922
rect 11164 42702 11192 42894
rect 11348 42838 11376 43302
rect 11336 42832 11388 42838
rect 11336 42774 11388 42780
rect 11440 42702 11468 43404
rect 11612 43308 11664 43314
rect 11716 43296 11744 43846
rect 11664 43268 11744 43296
rect 11612 43250 11664 43256
rect 11704 43104 11756 43110
rect 11704 43046 11756 43052
rect 10968 42696 11020 42702
rect 10968 42638 11020 42644
rect 11152 42696 11204 42702
rect 11152 42638 11204 42644
rect 11428 42696 11480 42702
rect 11428 42638 11480 42644
rect 10796 42588 10916 42616
rect 10692 42560 10744 42566
rect 10692 42502 10744 42508
rect 10704 42401 10732 42502
rect 10690 42392 10746 42401
rect 10600 42356 10652 42362
rect 10690 42327 10746 42336
rect 10600 42298 10652 42304
rect 10692 42288 10744 42294
rect 10520 42236 10692 42242
rect 10520 42230 10744 42236
rect 10520 42214 10732 42230
rect 10244 41534 10364 41562
rect 10230 41440 10286 41449
rect 10230 41375 10286 41384
rect 10140 39636 10192 39642
rect 10140 39578 10192 39584
rect 9680 38548 9732 38554
rect 9680 38490 9732 38496
rect 9586 38312 9642 38321
rect 9586 38247 9642 38256
rect 9404 36780 9456 36786
rect 9404 36722 9456 36728
rect 9312 36032 9364 36038
rect 9416 36009 9444 36722
rect 9588 36576 9640 36582
rect 9588 36518 9640 36524
rect 9312 35974 9364 35980
rect 9402 36000 9458 36009
rect 9402 35935 9458 35944
rect 9402 35864 9458 35873
rect 9402 35799 9458 35808
rect 9600 35816 9628 36518
rect 9692 36122 9720 38490
rect 10048 38004 10100 38010
rect 10048 37946 10100 37952
rect 9954 37360 10010 37369
rect 9954 37295 9956 37304
rect 10008 37295 10010 37304
rect 9956 37266 10008 37272
rect 9772 37120 9824 37126
rect 9772 37062 9824 37068
rect 9784 36378 9812 37062
rect 9956 36916 10008 36922
rect 9956 36858 10008 36864
rect 9864 36576 9916 36582
rect 9862 36544 9864 36553
rect 9916 36544 9918 36553
rect 9862 36479 9918 36488
rect 9772 36372 9824 36378
rect 9772 36314 9824 36320
rect 9968 36156 9996 36858
rect 10060 36786 10088 37946
rect 10244 37210 10272 41375
rect 10152 37182 10272 37210
rect 10048 36780 10100 36786
rect 10048 36722 10100 36728
rect 10060 36310 10088 36722
rect 10048 36304 10100 36310
rect 10048 36246 10100 36252
rect 9968 36128 10088 36156
rect 9692 36094 9904 36122
rect 9772 36032 9824 36038
rect 9772 35974 9824 35980
rect 9416 35714 9444 35799
rect 9600 35788 9720 35816
rect 9198 35686 9260 35714
rect 9324 35698 9444 35714
rect 9312 35692 9444 35698
rect 9198 35612 9226 35686
rect 9364 35686 9444 35692
rect 9312 35634 9364 35640
rect 9429 35624 9481 35630
rect 9198 35584 9260 35612
rect 9232 34950 9260 35584
rect 9416 35572 9429 35578
rect 9416 35566 9481 35572
rect 9588 35624 9640 35630
rect 9692 35612 9720 35788
rect 9640 35584 9720 35612
rect 9588 35566 9640 35572
rect 9416 35550 9469 35566
rect 9416 35544 9444 35550
rect 9324 35516 9444 35544
rect 9220 34944 9272 34950
rect 9220 34886 9272 34892
rect 9218 34096 9274 34105
rect 9218 34031 9274 34040
rect 9088 32456 9168 32484
rect 9036 32438 9088 32444
rect 8852 32292 8904 32298
rect 8852 32234 8904 32240
rect 8747 32124 9055 32133
rect 8747 32122 8753 32124
rect 8809 32122 8833 32124
rect 8889 32122 8913 32124
rect 8969 32122 8993 32124
rect 9049 32122 9055 32124
rect 8809 32070 8811 32122
rect 8991 32070 8993 32122
rect 8747 32068 8753 32070
rect 8809 32068 8833 32070
rect 8889 32068 8913 32070
rect 8969 32068 8993 32070
rect 9049 32068 9055 32070
rect 8747 32059 9055 32068
rect 9232 31906 9260 34031
rect 9324 33862 9352 35516
rect 9402 35456 9458 35465
rect 9402 35391 9458 35400
rect 9416 34678 9444 35391
rect 9784 35329 9812 35974
rect 9494 35320 9550 35329
rect 9494 35255 9550 35264
rect 9770 35320 9826 35329
rect 9770 35255 9826 35264
rect 9508 35086 9536 35255
rect 9876 35136 9904 36094
rect 9954 35864 10010 35873
rect 9954 35799 10010 35808
rect 9784 35108 9904 35136
rect 9496 35080 9548 35086
rect 9496 35022 9548 35028
rect 9496 34944 9548 34950
rect 9496 34886 9548 34892
rect 9404 34672 9456 34678
rect 9404 34614 9456 34620
rect 9312 33856 9364 33862
rect 9312 33798 9364 33804
rect 9312 32836 9364 32842
rect 9312 32778 9364 32784
rect 9324 32570 9352 32778
rect 9508 32756 9536 34886
rect 9680 34672 9732 34678
rect 9678 34640 9680 34649
rect 9732 34640 9734 34649
rect 9588 34604 9640 34610
rect 9678 34575 9734 34584
rect 9588 34546 9640 34552
rect 9600 34202 9628 34546
rect 9588 34196 9640 34202
rect 9588 34138 9640 34144
rect 9588 33856 9640 33862
rect 9588 33798 9640 33804
rect 9416 32728 9536 32756
rect 9312 32564 9364 32570
rect 9312 32506 9364 32512
rect 9140 31878 9260 31906
rect 8747 31036 9055 31045
rect 8747 31034 8753 31036
rect 8809 31034 8833 31036
rect 8889 31034 8913 31036
rect 8969 31034 8993 31036
rect 9049 31034 9055 31036
rect 8809 30982 8811 31034
rect 8991 30982 8993 31034
rect 8747 30980 8753 30982
rect 8809 30980 8833 30982
rect 8889 30980 8913 30982
rect 8969 30980 8993 30982
rect 9049 30980 9055 30982
rect 8747 30971 9055 30980
rect 9034 30560 9090 30569
rect 9034 30495 9090 30504
rect 9048 30326 9076 30495
rect 9036 30320 9088 30326
rect 9036 30262 9088 30268
rect 8747 29948 9055 29957
rect 8747 29946 8753 29948
rect 8809 29946 8833 29948
rect 8889 29946 8913 29948
rect 8969 29946 8993 29948
rect 9049 29946 9055 29948
rect 8809 29894 8811 29946
rect 8991 29894 8993 29946
rect 8747 29892 8753 29894
rect 8809 29892 8833 29894
rect 8889 29892 8913 29894
rect 8969 29892 8993 29894
rect 9049 29892 9055 29894
rect 8747 29883 9055 29892
rect 9036 29708 9088 29714
rect 9036 29650 9088 29656
rect 9048 29034 9076 29650
rect 9036 29028 9088 29034
rect 9036 28970 9088 28976
rect 8747 28860 9055 28869
rect 8747 28858 8753 28860
rect 8809 28858 8833 28860
rect 8889 28858 8913 28860
rect 8969 28858 8993 28860
rect 9049 28858 9055 28860
rect 8809 28806 8811 28858
rect 8991 28806 8993 28858
rect 8747 28804 8753 28806
rect 8809 28804 8833 28806
rect 8889 28804 8913 28806
rect 8969 28804 8993 28806
rect 9049 28804 9055 28806
rect 8747 28795 9055 28804
rect 9036 28620 9088 28626
rect 9036 28562 9088 28568
rect 8852 28552 8904 28558
rect 8852 28494 8904 28500
rect 8668 28416 8720 28422
rect 8668 28358 8720 28364
rect 8864 28257 8892 28494
rect 8850 28248 8906 28257
rect 9048 28218 9076 28562
rect 8850 28183 8906 28192
rect 8944 28212 8996 28218
rect 8576 28144 8628 28150
rect 8576 28086 8628 28092
rect 8864 28082 8892 28183
rect 8944 28154 8996 28160
rect 9036 28212 9088 28218
rect 9036 28154 9088 28160
rect 8852 28076 8904 28082
rect 8852 28018 8904 28024
rect 8668 28008 8720 28014
rect 8956 27985 8984 28154
rect 8668 27950 8720 27956
rect 8942 27976 8998 27985
rect 8484 27940 8536 27946
rect 8484 27882 8536 27888
rect 8680 27614 8708 27950
rect 8942 27911 8998 27920
rect 8747 27772 9055 27781
rect 8747 27770 8753 27772
rect 8809 27770 8833 27772
rect 8889 27770 8913 27772
rect 8969 27770 8993 27772
rect 9049 27770 9055 27772
rect 8809 27718 8811 27770
rect 8991 27718 8993 27770
rect 8747 27716 8753 27718
rect 8809 27716 8833 27718
rect 8889 27716 8913 27718
rect 8969 27716 8993 27718
rect 9049 27716 9055 27718
rect 8747 27707 9055 27716
rect 9140 27674 9168 31878
rect 9312 31748 9364 31754
rect 9312 31690 9364 31696
rect 9220 30252 9272 30258
rect 9220 30194 9272 30200
rect 9232 29850 9260 30194
rect 9220 29844 9272 29850
rect 9220 29786 9272 29792
rect 9220 29640 9272 29646
rect 9220 29582 9272 29588
rect 9232 29238 9260 29582
rect 9220 29232 9272 29238
rect 9220 29174 9272 29180
rect 9220 29028 9272 29034
rect 9220 28970 9272 28976
rect 9128 27668 9180 27674
rect 8680 27586 8800 27614
rect 9128 27610 9180 27616
rect 9232 27614 9260 28970
rect 9324 28948 9352 31690
rect 9416 31124 9444 32728
rect 9600 32450 9628 33798
rect 9680 33584 9732 33590
rect 9680 33526 9732 33532
rect 9566 32422 9628 32450
rect 9692 32434 9720 33526
rect 9784 33454 9812 35108
rect 9864 35012 9916 35018
rect 9864 34954 9916 34960
rect 9772 33448 9824 33454
rect 9772 33390 9824 33396
rect 9772 33312 9824 33318
rect 9772 33254 9824 33260
rect 9784 32502 9812 33254
rect 9772 32496 9824 32502
rect 9772 32438 9824 32444
rect 9680 32428 9732 32434
rect 9566 32348 9594 32422
rect 9680 32370 9732 32376
rect 9566 32320 9628 32348
rect 9600 31890 9628 32320
rect 9770 32328 9826 32337
rect 9770 32263 9826 32272
rect 9588 31884 9640 31890
rect 9588 31826 9640 31832
rect 9680 31680 9732 31686
rect 9680 31622 9732 31628
rect 9692 31278 9720 31622
rect 9680 31272 9732 31278
rect 9784 31249 9812 32263
rect 9680 31214 9732 31220
rect 9770 31240 9826 31249
rect 9416 31096 9536 31124
rect 9404 30796 9456 30802
rect 9404 30738 9456 30744
rect 9416 30122 9444 30738
rect 9404 30116 9456 30122
rect 9404 30058 9456 30064
rect 9416 29238 9444 30058
rect 9508 29714 9536 31096
rect 9586 31104 9642 31113
rect 9586 31039 9642 31048
rect 9496 29708 9548 29714
rect 9496 29650 9548 29656
rect 9416 29232 9481 29238
rect 9416 29192 9429 29232
rect 9429 29174 9481 29180
rect 9404 29096 9456 29102
rect 9456 29056 9536 29084
rect 9404 29038 9456 29044
rect 9324 28920 9444 28948
rect 9310 28792 9366 28801
rect 9310 28727 9366 28736
rect 9324 28490 9352 28727
rect 9312 28484 9364 28490
rect 9312 28426 9364 28432
rect 9232 27586 9352 27614
rect 8404 27390 8708 27418
rect 8392 27328 8444 27334
rect 8392 27270 8444 27276
rect 8484 27328 8536 27334
rect 8484 27270 8536 27276
rect 8404 25974 8432 27270
rect 8496 26586 8524 27270
rect 8574 27160 8630 27169
rect 8574 27095 8630 27104
rect 8484 26580 8536 26586
rect 8484 26522 8536 26528
rect 8484 26240 8536 26246
rect 8484 26182 8536 26188
rect 8392 25968 8444 25974
rect 8392 25910 8444 25916
rect 8298 25392 8354 25401
rect 8208 25356 8260 25362
rect 8298 25327 8354 25336
rect 8208 25298 8260 25304
rect 8404 25226 8432 25910
rect 8496 25498 8524 26182
rect 8484 25492 8536 25498
rect 8484 25434 8536 25440
rect 8392 25220 8444 25226
rect 8392 25162 8444 25168
rect 8116 24948 8168 24954
rect 8116 24890 8168 24896
rect 8128 23730 8156 24890
rect 8300 24676 8352 24682
rect 8300 24618 8352 24624
rect 8206 24440 8262 24449
rect 8312 24410 8340 24618
rect 8392 24608 8444 24614
rect 8392 24550 8444 24556
rect 8206 24375 8262 24384
rect 8300 24404 8352 24410
rect 8116 23724 8168 23730
rect 8116 23666 8168 23672
rect 8024 23656 8076 23662
rect 8024 23598 8076 23604
rect 7932 23316 7984 23322
rect 7932 23258 7984 23264
rect 7944 22778 7972 23258
rect 8220 22982 8248 24375
rect 8300 24346 8352 24352
rect 8312 23662 8340 24346
rect 8300 23656 8352 23662
rect 8300 23598 8352 23604
rect 8404 23508 8432 24550
rect 8312 23480 8432 23508
rect 8024 22976 8076 22982
rect 8024 22918 8076 22924
rect 8208 22976 8260 22982
rect 8208 22918 8260 22924
rect 7932 22772 7984 22778
rect 7932 22714 7984 22720
rect 7932 22500 7984 22506
rect 7932 22442 7984 22448
rect 7944 22030 7972 22442
rect 7932 22024 7984 22030
rect 7932 21966 7984 21972
rect 8036 21962 8064 22918
rect 8220 22234 8248 22918
rect 8208 22228 8260 22234
rect 8208 22170 8260 22176
rect 8114 22128 8170 22137
rect 8114 22063 8170 22072
rect 8024 21956 8076 21962
rect 8024 21898 8076 21904
rect 7932 21344 7984 21350
rect 7932 21286 7984 21292
rect 8022 21312 8078 21321
rect 7944 20942 7972 21286
rect 8022 21247 8078 21256
rect 7932 20936 7984 20942
rect 7932 20878 7984 20884
rect 7944 20602 7972 20878
rect 8036 20602 8064 21247
rect 8128 21146 8156 22063
rect 8312 22030 8340 23480
rect 8588 23338 8616 27095
rect 8680 27033 8708 27390
rect 8666 27024 8722 27033
rect 8666 26959 8668 26968
rect 8720 26959 8722 26968
rect 8668 26930 8720 26936
rect 8666 26888 8722 26897
rect 8666 26823 8722 26832
rect 8680 25974 8708 26823
rect 8772 26790 8800 27586
rect 9126 27568 9182 27577
rect 9126 27503 9182 27512
rect 8760 26784 8812 26790
rect 8760 26726 8812 26732
rect 8747 26684 9055 26693
rect 8747 26682 8753 26684
rect 8809 26682 8833 26684
rect 8889 26682 8913 26684
rect 8969 26682 8993 26684
rect 9049 26682 9055 26684
rect 8809 26630 8811 26682
rect 8991 26630 8993 26682
rect 8747 26628 8753 26630
rect 8809 26628 8833 26630
rect 8889 26628 8913 26630
rect 8969 26628 8993 26630
rect 9049 26628 9055 26630
rect 8747 26619 9055 26628
rect 9140 26586 9168 27503
rect 9220 27396 9272 27402
rect 9220 27338 9272 27344
rect 9128 26580 9180 26586
rect 9128 26522 9180 26528
rect 9232 26432 9260 27338
rect 9324 27062 9352 27586
rect 9416 27334 9444 28920
rect 9508 28234 9536 29056
rect 9600 28393 9628 31039
rect 9586 28384 9642 28393
rect 9586 28319 9642 28328
rect 9508 28218 9628 28234
rect 9508 28212 9640 28218
rect 9508 28206 9588 28212
rect 9588 28154 9640 28160
rect 9496 28144 9548 28150
rect 9496 28086 9548 28092
rect 9508 27985 9536 28086
rect 9494 27976 9550 27985
rect 9494 27911 9550 27920
rect 9496 27668 9548 27674
rect 9496 27610 9548 27616
rect 9404 27328 9456 27334
rect 9404 27270 9456 27276
rect 9312 27056 9364 27062
rect 9312 26998 9364 27004
rect 9404 26920 9456 26926
rect 9404 26862 9456 26868
rect 9312 26784 9364 26790
rect 9312 26726 9364 26732
rect 9324 26450 9352 26726
rect 9140 26404 9260 26432
rect 9312 26444 9364 26450
rect 8668 25968 8720 25974
rect 8668 25910 8720 25916
rect 8680 25362 8708 25910
rect 8747 25596 9055 25605
rect 8747 25594 8753 25596
rect 8809 25594 8833 25596
rect 8889 25594 8913 25596
rect 8969 25594 8993 25596
rect 9049 25594 9055 25596
rect 8809 25542 8811 25594
rect 8991 25542 8993 25594
rect 8747 25540 8753 25542
rect 8809 25540 8833 25542
rect 8889 25540 8913 25542
rect 8969 25540 8993 25542
rect 9049 25540 9055 25542
rect 8747 25531 9055 25540
rect 9140 25498 9168 26404
rect 9312 26386 9364 26392
rect 9220 26308 9272 26314
rect 9220 26250 9272 26256
rect 9128 25492 9180 25498
rect 8956 25452 9128 25480
rect 8668 25356 8720 25362
rect 8668 25298 8720 25304
rect 8668 25220 8720 25226
rect 8668 25162 8720 25168
rect 8680 23644 8708 25162
rect 8956 24834 8984 25452
rect 9128 25434 9180 25440
rect 8772 24818 8984 24834
rect 8760 24812 8984 24818
rect 8812 24806 8984 24812
rect 8760 24754 8812 24760
rect 9232 24750 9260 26250
rect 9312 26240 9364 26246
rect 9312 26182 9364 26188
rect 9036 24744 9088 24750
rect 9220 24744 9272 24750
rect 9088 24704 9168 24732
rect 9036 24686 9088 24692
rect 8747 24508 9055 24517
rect 8747 24506 8753 24508
rect 8809 24506 8833 24508
rect 8889 24506 8913 24508
rect 8969 24506 8993 24508
rect 9049 24506 9055 24508
rect 8809 24454 8811 24506
rect 8991 24454 8993 24506
rect 8747 24452 8753 24454
rect 8809 24452 8833 24454
rect 8889 24452 8913 24454
rect 8969 24452 8993 24454
rect 9049 24452 9055 24454
rect 8747 24443 9055 24452
rect 9140 23662 9168 24704
rect 9220 24686 9272 24692
rect 9324 24256 9352 26182
rect 9416 25158 9444 26862
rect 9404 25152 9456 25158
rect 9404 25094 9456 25100
rect 9508 24886 9536 27610
rect 9588 27396 9640 27402
rect 9588 27338 9640 27344
rect 9600 25786 9628 27338
rect 9692 26364 9720 31214
rect 9770 31175 9826 31184
rect 9876 30297 9904 34954
rect 9968 34950 9996 35799
rect 9956 34944 10008 34950
rect 9956 34886 10008 34892
rect 9954 34640 10010 34649
rect 10060 34610 10088 36128
rect 10152 35714 10180 37182
rect 10232 37120 10284 37126
rect 10232 37062 10284 37068
rect 10244 36922 10272 37062
rect 10232 36916 10284 36922
rect 10232 36858 10284 36864
rect 10232 36780 10284 36786
rect 10232 36722 10284 36728
rect 10244 36689 10272 36722
rect 10230 36680 10286 36689
rect 10230 36615 10286 36624
rect 10336 35873 10364 41534
rect 10416 37188 10468 37194
rect 10416 37130 10468 37136
rect 10428 36922 10456 37130
rect 10416 36916 10468 36922
rect 10416 36858 10468 36864
rect 10322 35864 10378 35873
rect 10322 35799 10378 35808
rect 10520 35714 10548 42214
rect 10692 42084 10744 42090
rect 10692 42026 10744 42032
rect 10704 41414 10732 42026
rect 10612 41386 10732 41414
rect 10612 36553 10640 41386
rect 10692 37664 10744 37670
rect 10692 37606 10744 37612
rect 10704 37330 10732 37606
rect 10692 37324 10744 37330
rect 10692 37266 10744 37272
rect 10598 36544 10654 36553
rect 10598 36479 10654 36488
rect 10612 36174 10640 36479
rect 10600 36168 10652 36174
rect 10600 36110 10652 36116
rect 10152 35686 10456 35714
rect 10520 35686 10640 35714
rect 10230 35592 10286 35601
rect 10230 35527 10286 35536
rect 10244 35018 10272 35527
rect 10322 35184 10378 35193
rect 10322 35119 10378 35128
rect 10232 35012 10284 35018
rect 10232 34954 10284 34960
rect 9954 34575 9956 34584
rect 10008 34575 10010 34584
rect 10048 34604 10100 34610
rect 9956 34546 10008 34552
rect 10048 34546 10100 34552
rect 10336 33980 10364 35119
rect 10428 34746 10456 35686
rect 10612 35086 10640 35686
rect 10600 35080 10652 35086
rect 10600 35022 10652 35028
rect 10508 34944 10560 34950
rect 10508 34886 10560 34892
rect 10416 34740 10468 34746
rect 10416 34682 10468 34688
rect 10416 33992 10468 33998
rect 10336 33952 10416 33980
rect 10416 33934 10468 33940
rect 10416 33516 10468 33522
rect 10416 33458 10468 33464
rect 9956 33448 10008 33454
rect 9956 33390 10008 33396
rect 9968 31906 9996 33390
rect 10048 32768 10100 32774
rect 10428 32722 10456 33458
rect 10048 32710 10100 32716
rect 10060 32026 10088 32710
rect 10152 32694 10456 32722
rect 10048 32020 10100 32026
rect 10048 31962 10100 31968
rect 9968 31878 10088 31906
rect 9956 31816 10008 31822
rect 9954 31784 9956 31793
rect 10008 31784 10010 31793
rect 9954 31719 10010 31728
rect 10060 31346 10088 31878
rect 10048 31340 10100 31346
rect 10048 31282 10100 31288
rect 10060 30938 10088 31282
rect 10048 30932 10100 30938
rect 10048 30874 10100 30880
rect 10048 30388 10100 30394
rect 10048 30330 10100 30336
rect 9862 30288 9918 30297
rect 9862 30223 9918 30232
rect 10060 29832 10088 30330
rect 10042 29804 10088 29832
rect 10042 29764 10070 29804
rect 9968 29736 10070 29764
rect 9968 29696 9996 29736
rect 9784 29668 9996 29696
rect 9784 28014 9812 29668
rect 10152 29646 10180 32694
rect 10428 32502 10456 32694
rect 10232 32496 10284 32502
rect 10232 32438 10284 32444
rect 10416 32496 10468 32502
rect 10416 32438 10468 32444
rect 10244 31686 10272 32438
rect 10416 32292 10468 32298
rect 10416 32234 10468 32240
rect 10324 32224 10376 32230
rect 10428 32201 10456 32234
rect 10324 32166 10376 32172
rect 10414 32192 10470 32201
rect 10336 31890 10364 32166
rect 10414 32127 10470 32136
rect 10324 31884 10376 31890
rect 10324 31826 10376 31832
rect 10232 31680 10284 31686
rect 10232 31622 10284 31628
rect 10428 31498 10456 32127
rect 10336 31470 10456 31498
rect 10140 29640 10192 29646
rect 9876 29600 10140 29628
rect 9772 28008 9824 28014
rect 9772 27950 9824 27956
rect 9784 27538 9812 27950
rect 9772 27532 9824 27538
rect 9772 27474 9824 27480
rect 9784 26994 9812 27474
rect 9772 26988 9824 26994
rect 9772 26930 9824 26936
rect 9772 26784 9824 26790
rect 9772 26726 9824 26732
rect 9784 26586 9812 26726
rect 9772 26580 9824 26586
rect 9772 26522 9824 26528
rect 9772 26376 9824 26382
rect 9692 26336 9772 26364
rect 9772 26318 9824 26324
rect 9876 26024 9904 29600
rect 10140 29582 10192 29588
rect 10048 29504 10100 29510
rect 10048 29446 10100 29452
rect 10060 29288 10088 29446
rect 10060 29260 10272 29288
rect 9954 28928 10010 28937
rect 9954 28863 10010 28872
rect 9968 27402 9996 28863
rect 10060 27614 10088 29260
rect 10244 29170 10272 29260
rect 10140 29164 10192 29170
rect 10140 29106 10192 29112
rect 10232 29164 10284 29170
rect 10232 29106 10284 29112
rect 10152 28744 10180 29106
rect 10336 28948 10364 31470
rect 10416 31408 10468 31414
rect 10416 31350 10468 31356
rect 10428 30977 10456 31350
rect 10414 30968 10470 30977
rect 10414 30903 10470 30912
rect 10336 28937 10456 28948
rect 10336 28928 10470 28937
rect 10336 28920 10414 28928
rect 10414 28863 10470 28872
rect 10416 28756 10468 28762
rect 10152 28716 10416 28744
rect 10416 28698 10468 28704
rect 10140 28484 10192 28490
rect 10140 28426 10192 28432
rect 10152 28082 10180 28426
rect 10416 28416 10468 28422
rect 10416 28358 10468 28364
rect 10324 28212 10376 28218
rect 10324 28154 10376 28160
rect 10140 28076 10192 28082
rect 10140 28018 10192 28024
rect 10060 27586 10272 27614
rect 10046 27432 10102 27441
rect 9956 27396 10008 27402
rect 10046 27367 10102 27376
rect 9956 27338 10008 27344
rect 9956 26376 10008 26382
rect 10060 26364 10088 27367
rect 10138 27160 10194 27169
rect 10138 27095 10194 27104
rect 10152 27062 10180 27095
rect 10140 27056 10192 27062
rect 10140 26998 10192 27004
rect 10008 26336 10088 26364
rect 9956 26318 10008 26324
rect 9784 25996 9904 26024
rect 9600 25758 9720 25786
rect 9588 25696 9640 25702
rect 9588 25638 9640 25644
rect 9496 24880 9548 24886
rect 9496 24822 9548 24828
rect 9404 24676 9456 24682
rect 9404 24618 9456 24624
rect 9232 24228 9352 24256
rect 8760 23656 8812 23662
rect 8680 23616 8760 23644
rect 8760 23598 8812 23604
rect 9128 23656 9180 23662
rect 9128 23598 9180 23604
rect 8772 23526 8800 23598
rect 8760 23520 8812 23526
rect 8760 23462 8812 23468
rect 8747 23420 9055 23429
rect 8747 23418 8753 23420
rect 8809 23418 8833 23420
rect 8889 23418 8913 23420
rect 8969 23418 8993 23420
rect 9049 23418 9055 23420
rect 8809 23366 8811 23418
rect 8991 23366 8993 23418
rect 8747 23364 8753 23366
rect 8809 23364 8833 23366
rect 8889 23364 8913 23366
rect 8969 23364 8993 23366
rect 9049 23364 9055 23366
rect 8747 23355 9055 23364
rect 8404 23310 8616 23338
rect 9140 23322 9168 23598
rect 9128 23316 9180 23322
rect 8404 22137 8432 23310
rect 9128 23258 9180 23264
rect 8668 22636 8720 22642
rect 8668 22578 8720 22584
rect 8484 22500 8536 22506
rect 8484 22442 8536 22448
rect 8390 22128 8446 22137
rect 8390 22063 8446 22072
rect 8300 22024 8352 22030
rect 8206 21992 8262 22001
rect 8300 21966 8352 21972
rect 8392 22024 8444 22030
rect 8392 21966 8444 21972
rect 8206 21927 8262 21936
rect 8116 21140 8168 21146
rect 8116 21082 8168 21088
rect 7932 20596 7984 20602
rect 7932 20538 7984 20544
rect 8024 20596 8076 20602
rect 8024 20538 8076 20544
rect 7840 20528 7892 20534
rect 7840 20470 7892 20476
rect 7852 19122 7880 20470
rect 7932 20460 7984 20466
rect 7932 20402 7984 20408
rect 7944 19514 7972 20402
rect 8220 20058 8248 21927
rect 8298 21176 8354 21185
rect 8404 21162 8432 21966
rect 8354 21134 8432 21162
rect 8298 21111 8354 21120
rect 8300 20528 8352 20534
rect 8300 20470 8352 20476
rect 8312 20233 8340 20470
rect 8298 20224 8354 20233
rect 8298 20159 8354 20168
rect 8208 20052 8260 20058
rect 8208 19994 8260 20000
rect 7932 19508 7984 19514
rect 7932 19450 7984 19456
rect 8208 19372 8260 19378
rect 8208 19314 8260 19320
rect 7852 19094 7972 19122
rect 7838 19000 7894 19009
rect 7838 18935 7894 18944
rect 7852 18698 7880 18935
rect 7840 18692 7892 18698
rect 7840 18634 7892 18640
rect 7852 18465 7880 18634
rect 7838 18456 7894 18465
rect 7944 18426 7972 19094
rect 8220 18630 8248 19314
rect 8300 19236 8352 19242
rect 8300 19178 8352 19184
rect 8312 18698 8340 19178
rect 8300 18692 8352 18698
rect 8300 18634 8352 18640
rect 8208 18624 8260 18630
rect 8208 18566 8260 18572
rect 8392 18624 8444 18630
rect 8392 18566 8444 18572
rect 7838 18391 7894 18400
rect 7932 18420 7984 18426
rect 7932 18362 7984 18368
rect 8116 18352 8168 18358
rect 8116 18294 8168 18300
rect 7932 18284 7984 18290
rect 7932 18226 7984 18232
rect 7840 18080 7892 18086
rect 7840 18022 7892 18028
rect 7852 17678 7880 18022
rect 7840 17672 7892 17678
rect 7840 17614 7892 17620
rect 7840 17332 7892 17338
rect 7944 17320 7972 18226
rect 8128 17678 8156 18294
rect 8116 17672 8168 17678
rect 8116 17614 8168 17620
rect 8116 17536 8168 17542
rect 8116 17478 8168 17484
rect 7892 17292 7972 17320
rect 7840 17274 7892 17280
rect 8128 17270 8156 17478
rect 8116 17264 8168 17270
rect 8036 17224 8116 17252
rect 8036 16266 8064 17224
rect 8116 17206 8168 17212
rect 7944 16238 8064 16266
rect 7840 15428 7892 15434
rect 7944 15416 7972 16238
rect 8114 16144 8170 16153
rect 8114 16079 8170 16088
rect 8024 15496 8076 15502
rect 8024 15438 8076 15444
rect 7892 15388 7972 15416
rect 7840 15370 7892 15376
rect 7852 13938 7880 15370
rect 7932 14952 7984 14958
rect 7932 14894 7984 14900
rect 7944 14278 7972 14894
rect 8036 14618 8064 15438
rect 8024 14612 8076 14618
rect 8024 14554 8076 14560
rect 7932 14272 7984 14278
rect 7932 14214 7984 14220
rect 7840 13932 7892 13938
rect 7840 13874 7892 13880
rect 7838 13696 7894 13705
rect 7838 13631 7894 13640
rect 7852 13326 7880 13631
rect 7840 13320 7892 13326
rect 7746 13288 7802 13297
rect 7840 13262 7892 13268
rect 7746 13223 7802 13232
rect 7944 13161 7972 14214
rect 7930 13152 7986 13161
rect 7930 13087 7986 13096
rect 7748 12776 7800 12782
rect 7668 12736 7748 12764
rect 7800 12736 7880 12764
rect 7748 12718 7800 12724
rect 7654 12608 7710 12617
rect 7710 12566 7788 12594
rect 7654 12543 7710 12552
rect 7654 12472 7710 12481
rect 7760 12442 7788 12566
rect 7654 12407 7710 12416
rect 7748 12436 7800 12442
rect 7668 12238 7696 12407
rect 7748 12378 7800 12384
rect 7656 12232 7708 12238
rect 7656 12174 7708 12180
rect 7654 12064 7710 12073
rect 7654 11999 7710 12008
rect 7564 11688 7616 11694
rect 7564 11630 7616 11636
rect 7668 10810 7696 11999
rect 7760 11150 7788 12378
rect 7748 11144 7800 11150
rect 7748 11086 7800 11092
rect 7656 10804 7708 10810
rect 7656 10746 7708 10752
rect 7564 10464 7616 10470
rect 7564 10406 7616 10412
rect 7576 9722 7604 10406
rect 7852 10146 7880 12736
rect 8128 12628 8156 16079
rect 8220 15026 8248 18566
rect 8300 18420 8352 18426
rect 8300 18362 8352 18368
rect 8312 17678 8340 18362
rect 8404 18222 8432 18566
rect 8392 18216 8444 18222
rect 8392 18158 8444 18164
rect 8390 17776 8446 17785
rect 8390 17711 8446 17720
rect 8300 17672 8352 17678
rect 8300 17614 8352 17620
rect 8300 16108 8352 16114
rect 8300 16050 8352 16056
rect 8312 15162 8340 16050
rect 8404 15201 8432 17711
rect 8390 15192 8446 15201
rect 8300 15156 8352 15162
rect 8390 15127 8446 15136
rect 8300 15098 8352 15104
rect 8208 15020 8260 15026
rect 8208 14962 8260 14968
rect 8208 14816 8260 14822
rect 8208 14758 8260 14764
rect 8392 14816 8444 14822
rect 8392 14758 8444 14764
rect 8220 14657 8248 14758
rect 8206 14648 8262 14657
rect 8206 14583 8262 14592
rect 8298 14512 8354 14521
rect 8298 14447 8354 14456
rect 8206 13832 8262 13841
rect 8206 13767 8262 13776
rect 8036 12600 8156 12628
rect 7930 11928 7986 11937
rect 7930 11863 7986 11872
rect 7944 11558 7972 11863
rect 7932 11552 7984 11558
rect 7932 11494 7984 11500
rect 7656 10124 7708 10130
rect 7760 10118 7880 10146
rect 7760 10112 7788 10118
rect 8036 10112 8064 12600
rect 8220 12288 8248 13767
rect 8312 13394 8340 14447
rect 8300 13388 8352 13394
rect 8300 13330 8352 13336
rect 8128 12260 8248 12288
rect 8128 12102 8156 12260
rect 8208 12164 8260 12170
rect 8208 12106 8260 12112
rect 8116 12096 8168 12102
rect 8116 12038 8168 12044
rect 8220 11898 8248 12106
rect 8208 11892 8260 11898
rect 8208 11834 8260 11840
rect 8300 11688 8352 11694
rect 8298 11656 8300 11665
rect 8352 11656 8354 11665
rect 8298 11591 8354 11600
rect 8116 11552 8168 11558
rect 8116 11494 8168 11500
rect 7708 10084 7788 10112
rect 7944 10084 8064 10112
rect 7656 10066 7708 10072
rect 7840 10056 7892 10062
rect 7840 9998 7892 10004
rect 7564 9716 7616 9722
rect 7564 9658 7616 9664
rect 7654 9616 7710 9625
rect 7654 9551 7656 9560
rect 7708 9551 7710 9560
rect 7748 9580 7800 9586
rect 7656 9522 7708 9528
rect 7748 9522 7800 9528
rect 7562 9480 7618 9489
rect 7562 9415 7618 9424
rect 7576 8566 7604 9415
rect 7656 8968 7708 8974
rect 7654 8936 7656 8945
rect 7708 8936 7710 8945
rect 7654 8871 7710 8880
rect 7564 8560 7616 8566
rect 7564 8502 7616 8508
rect 7760 8090 7788 9522
rect 7852 9178 7880 9998
rect 7840 9172 7892 9178
rect 7840 9114 7892 9120
rect 7944 9058 7972 10084
rect 8128 10010 8156 11494
rect 8208 11348 8260 11354
rect 8208 11290 8260 11296
rect 7852 9030 7972 9058
rect 8036 9982 8156 10010
rect 7852 8294 7880 9030
rect 8036 8401 8064 9982
rect 8220 9874 8248 11290
rect 8300 10192 8352 10198
rect 8300 10134 8352 10140
rect 8128 9846 8248 9874
rect 8022 8392 8078 8401
rect 8022 8327 8078 8336
rect 7840 8288 7892 8294
rect 7840 8230 7892 8236
rect 8024 8288 8076 8294
rect 8024 8230 8076 8236
rect 7748 8084 7800 8090
rect 7748 8026 7800 8032
rect 7760 7342 7788 8026
rect 7840 8016 7892 8022
rect 8036 7970 8064 8230
rect 8128 8022 8156 9846
rect 8312 9738 8340 10134
rect 8220 9710 8340 9738
rect 7840 7958 7892 7964
rect 7852 7449 7880 7958
rect 7944 7942 8064 7970
rect 8116 8016 8168 8022
rect 8116 7958 8168 7964
rect 7838 7440 7894 7449
rect 7838 7375 7894 7384
rect 7748 7336 7800 7342
rect 7748 7278 7800 7284
rect 7944 7274 7972 7942
rect 8220 7886 8248 9710
rect 8300 9376 8352 9382
rect 8300 9318 8352 9324
rect 8312 8106 8340 9318
rect 8404 8974 8432 14758
rect 8496 14498 8524 22442
rect 8576 22160 8628 22166
rect 8576 22102 8628 22108
rect 8588 20602 8616 22102
rect 8680 22098 8708 22578
rect 9128 22432 9180 22438
rect 9128 22374 9180 22380
rect 8747 22332 9055 22341
rect 8747 22330 8753 22332
rect 8809 22330 8833 22332
rect 8889 22330 8913 22332
rect 8969 22330 8993 22332
rect 9049 22330 9055 22332
rect 8809 22278 8811 22330
rect 8991 22278 8993 22330
rect 8747 22276 8753 22278
rect 8809 22276 8833 22278
rect 8889 22276 8913 22278
rect 8969 22276 8993 22278
rect 9049 22276 9055 22278
rect 8747 22267 9055 22276
rect 8668 22092 8720 22098
rect 8668 22034 8720 22040
rect 8668 21956 8720 21962
rect 9140 21944 9168 22374
rect 8668 21898 8720 21904
rect 9048 21916 9168 21944
rect 8576 20596 8628 20602
rect 8576 20538 8628 20544
rect 8680 20482 8708 21898
rect 9048 21622 9076 21916
rect 9232 21842 9260 24228
rect 9310 24168 9366 24177
rect 9310 24103 9366 24112
rect 9140 21814 9260 21842
rect 9324 21842 9352 24103
rect 9416 22001 9444 24618
rect 9496 24608 9548 24614
rect 9496 24550 9548 24556
rect 9508 24410 9536 24550
rect 9496 24404 9548 24410
rect 9496 24346 9548 24352
rect 9600 23594 9628 25638
rect 9588 23588 9640 23594
rect 9588 23530 9640 23536
rect 9692 23474 9720 25758
rect 9508 23446 9720 23474
rect 9508 22642 9536 23446
rect 9586 23352 9642 23361
rect 9586 23287 9642 23296
rect 9600 22953 9628 23287
rect 9680 23112 9732 23118
rect 9680 23054 9732 23060
rect 9586 22944 9642 22953
rect 9586 22879 9642 22888
rect 9496 22636 9548 22642
rect 9496 22578 9548 22584
rect 9692 22012 9720 23054
rect 9784 23050 9812 25996
rect 9862 25936 9918 25945
rect 9862 25871 9864 25880
rect 9916 25871 9918 25880
rect 9864 25842 9916 25848
rect 9864 25288 9916 25294
rect 9864 25230 9916 25236
rect 10140 25288 10192 25294
rect 10140 25230 10192 25236
rect 9876 24954 9904 25230
rect 10152 24954 10180 25230
rect 9864 24948 9916 24954
rect 9864 24890 9916 24896
rect 10140 24948 10192 24954
rect 10140 24890 10192 24896
rect 10244 24562 10272 27586
rect 9968 24534 10272 24562
rect 9864 24064 9916 24070
rect 9864 24006 9916 24012
rect 9876 23866 9904 24006
rect 9864 23860 9916 23866
rect 9864 23802 9916 23808
rect 9772 23044 9824 23050
rect 9772 22986 9824 22992
rect 9864 22976 9916 22982
rect 9862 22944 9864 22953
rect 9916 22944 9918 22953
rect 9862 22879 9918 22888
rect 9864 22432 9916 22438
rect 9864 22374 9916 22380
rect 9876 22166 9904 22374
rect 9864 22160 9916 22166
rect 9864 22102 9916 22108
rect 9772 22024 9824 22030
rect 9402 21992 9458 22001
rect 9692 21984 9772 22012
rect 9772 21966 9824 21972
rect 9402 21927 9458 21936
rect 9324 21814 9720 21842
rect 9140 21622 9168 21814
rect 9496 21684 9548 21690
rect 9496 21626 9548 21632
rect 9036 21616 9088 21622
rect 9036 21558 9088 21564
rect 9128 21616 9180 21622
rect 9128 21558 9180 21564
rect 9140 21298 9168 21558
rect 9404 21548 9456 21554
rect 9404 21490 9456 21496
rect 9416 21321 9444 21490
rect 9402 21312 9458 21321
rect 9140 21270 9260 21298
rect 8747 21244 9055 21253
rect 8747 21242 8753 21244
rect 8809 21242 8833 21244
rect 8889 21242 8913 21244
rect 8969 21242 8993 21244
rect 9049 21242 9055 21244
rect 8809 21190 8811 21242
rect 8991 21190 8993 21242
rect 8747 21188 8753 21190
rect 8809 21188 8833 21190
rect 8889 21188 8913 21190
rect 8969 21188 8993 21190
rect 9049 21188 9055 21190
rect 8747 21179 9055 21188
rect 9232 21146 9260 21270
rect 9402 21247 9458 21256
rect 9036 21140 9088 21146
rect 9220 21140 9272 21146
rect 9088 21100 9168 21128
rect 9036 21082 9088 21088
rect 9140 21049 9168 21100
rect 9220 21082 9272 21088
rect 9126 21040 9182 21049
rect 9126 20975 9182 20984
rect 9140 20942 9168 20975
rect 9128 20936 9180 20942
rect 9128 20878 9180 20884
rect 9508 20806 9536 21626
rect 9588 20936 9640 20942
rect 9588 20878 9640 20884
rect 9496 20800 9548 20806
rect 9496 20742 9548 20748
rect 9404 20596 9456 20602
rect 9404 20538 9456 20544
rect 8588 20454 8708 20482
rect 9220 20528 9272 20534
rect 9220 20470 9272 20476
rect 8588 18057 8616 20454
rect 9128 20256 9180 20262
rect 9128 20198 9180 20204
rect 8747 20156 9055 20165
rect 8747 20154 8753 20156
rect 8809 20154 8833 20156
rect 8889 20154 8913 20156
rect 8969 20154 8993 20156
rect 9049 20154 9055 20156
rect 8809 20102 8811 20154
rect 8991 20102 8993 20154
rect 8747 20100 8753 20102
rect 8809 20100 8833 20102
rect 8889 20100 8913 20102
rect 8969 20100 8993 20102
rect 9049 20100 9055 20102
rect 8747 20091 9055 20100
rect 8668 20052 8720 20058
rect 8668 19994 8720 20000
rect 8680 19174 8708 19994
rect 8668 19168 8720 19174
rect 8668 19110 8720 19116
rect 8574 18048 8630 18057
rect 8574 17983 8630 17992
rect 8588 17882 8616 17983
rect 8576 17876 8628 17882
rect 8680 17864 8708 19110
rect 8747 19068 9055 19077
rect 8747 19066 8753 19068
rect 8809 19066 8833 19068
rect 8889 19066 8913 19068
rect 8969 19066 8993 19068
rect 9049 19066 9055 19068
rect 8809 19014 8811 19066
rect 8991 19014 8993 19066
rect 8747 19012 8753 19014
rect 8809 19012 8833 19014
rect 8889 19012 8913 19014
rect 8969 19012 8993 19014
rect 9049 19012 9055 19014
rect 8747 19003 9055 19012
rect 9140 18850 9168 20198
rect 9048 18822 9168 18850
rect 8852 18760 8904 18766
rect 8852 18702 8904 18708
rect 8864 18358 8892 18702
rect 8852 18352 8904 18358
rect 8852 18294 8904 18300
rect 9048 18068 9076 18822
rect 9232 18426 9260 20470
rect 9416 19961 9444 20538
rect 9402 19952 9458 19961
rect 9402 19887 9458 19896
rect 9310 19816 9366 19825
rect 9310 19751 9366 19760
rect 9220 18420 9272 18426
rect 9220 18362 9272 18368
rect 9048 18040 9168 18068
rect 8747 17980 9055 17989
rect 8747 17978 8753 17980
rect 8809 17978 8833 17980
rect 8889 17978 8913 17980
rect 8969 17978 8993 17980
rect 9049 17978 9055 17980
rect 8809 17926 8811 17978
rect 8991 17926 8993 17978
rect 8747 17924 8753 17926
rect 8809 17924 8833 17926
rect 8889 17924 8913 17926
rect 8969 17924 8993 17926
rect 9049 17924 9055 17926
rect 8747 17915 9055 17924
rect 8680 17836 8984 17864
rect 8576 17818 8628 17824
rect 8588 17728 8616 17818
rect 8588 17700 8708 17728
rect 8574 17640 8630 17649
rect 8574 17575 8630 17584
rect 8588 17270 8616 17575
rect 8576 17264 8628 17270
rect 8576 17206 8628 17212
rect 8680 16658 8708 17700
rect 8956 17678 8984 17836
rect 8944 17672 8996 17678
rect 8944 17614 8996 17620
rect 8760 17536 8812 17542
rect 8758 17504 8760 17513
rect 8812 17504 8814 17513
rect 8758 17439 8814 17448
rect 8956 16998 8984 17614
rect 8944 16992 8996 16998
rect 8944 16934 8996 16940
rect 8747 16892 9055 16901
rect 8747 16890 8753 16892
rect 8809 16890 8833 16892
rect 8889 16890 8913 16892
rect 8969 16890 8993 16892
rect 9049 16890 9055 16892
rect 8809 16838 8811 16890
rect 8991 16838 8993 16890
rect 8747 16836 8753 16838
rect 8809 16836 8833 16838
rect 8889 16836 8913 16838
rect 8969 16836 8993 16838
rect 9049 16836 9055 16838
rect 8747 16827 9055 16836
rect 8668 16652 8720 16658
rect 8668 16594 8720 16600
rect 9140 16153 9168 18040
rect 9218 17912 9274 17921
rect 9218 17847 9274 17856
rect 9232 17678 9260 17847
rect 9220 17672 9272 17678
rect 9220 17614 9272 17620
rect 9324 16590 9352 19751
rect 9416 18834 9444 19887
rect 9494 19680 9550 19689
rect 9494 19615 9550 19624
rect 9404 18828 9456 18834
rect 9404 18770 9456 18776
rect 9508 17218 9536 19615
rect 9600 19174 9628 20878
rect 9692 19718 9720 21814
rect 9772 21616 9824 21622
rect 9772 21558 9824 21564
rect 9784 21146 9812 21558
rect 9772 21140 9824 21146
rect 9772 21082 9824 21088
rect 9876 20346 9904 22102
rect 9968 21729 9996 24534
rect 10048 24404 10100 24410
rect 10336 24392 10364 28154
rect 10048 24346 10100 24352
rect 10244 24364 10364 24392
rect 10060 24206 10088 24346
rect 10048 24200 10100 24206
rect 10048 24142 10100 24148
rect 10140 24064 10192 24070
rect 10046 24032 10102 24041
rect 10140 24006 10192 24012
rect 10046 23967 10102 23976
rect 10060 23118 10088 23967
rect 10048 23112 10100 23118
rect 10048 23054 10100 23060
rect 10046 22944 10102 22953
rect 10046 22879 10102 22888
rect 10060 22710 10088 22879
rect 10048 22704 10100 22710
rect 10048 22646 10100 22652
rect 10048 22568 10100 22574
rect 10048 22510 10100 22516
rect 10060 22234 10088 22510
rect 10048 22228 10100 22234
rect 10048 22170 10100 22176
rect 9954 21720 10010 21729
rect 9954 21655 9956 21664
rect 10008 21655 10010 21664
rect 9956 21626 10008 21632
rect 10048 21004 10100 21010
rect 10048 20946 10100 20952
rect 9876 20318 9996 20346
rect 9864 20256 9916 20262
rect 9864 20198 9916 20204
rect 9680 19712 9732 19718
rect 9680 19654 9732 19660
rect 9770 19544 9826 19553
rect 9680 19508 9732 19514
rect 9770 19479 9826 19488
rect 9680 19450 9732 19456
rect 9588 19168 9640 19174
rect 9588 19110 9640 19116
rect 9692 17898 9720 19450
rect 9784 19446 9812 19479
rect 9772 19440 9824 19446
rect 9772 19382 9824 19388
rect 9876 19378 9904 20198
rect 9864 19372 9916 19378
rect 9864 19314 9916 19320
rect 9772 19236 9824 19242
rect 9772 19178 9824 19184
rect 9784 19145 9812 19178
rect 9770 19136 9826 19145
rect 9770 19071 9826 19080
rect 9772 18964 9824 18970
rect 9772 18906 9824 18912
rect 9600 17870 9720 17898
rect 9600 17785 9628 17870
rect 9586 17776 9642 17785
rect 9586 17711 9642 17720
rect 9416 17190 9536 17218
rect 9312 16584 9364 16590
rect 9312 16526 9364 16532
rect 9220 16176 9272 16182
rect 9126 16144 9182 16153
rect 9220 16118 9272 16124
rect 9126 16079 9182 16088
rect 9128 15904 9180 15910
rect 9128 15846 9180 15852
rect 8747 15804 9055 15813
rect 8747 15802 8753 15804
rect 8809 15802 8833 15804
rect 8889 15802 8913 15804
rect 8969 15802 8993 15804
rect 9049 15802 9055 15804
rect 8809 15750 8811 15802
rect 8991 15750 8993 15802
rect 8747 15748 8753 15750
rect 8809 15748 8833 15750
rect 8889 15748 8913 15750
rect 8969 15748 8993 15750
rect 9049 15748 9055 15750
rect 8747 15739 9055 15748
rect 9140 15706 9168 15846
rect 9232 15706 9260 16118
rect 9128 15700 9180 15706
rect 9128 15642 9180 15648
rect 9220 15700 9272 15706
rect 9220 15642 9272 15648
rect 8668 15496 8720 15502
rect 8668 15438 8720 15444
rect 9220 15496 9272 15502
rect 9220 15438 9272 15444
rect 8680 14958 8708 15438
rect 9232 15094 9260 15438
rect 9324 15434 9352 16526
rect 9312 15428 9364 15434
rect 9312 15370 9364 15376
rect 9220 15088 9272 15094
rect 9126 15056 9182 15065
rect 9220 15030 9272 15036
rect 9126 14991 9182 15000
rect 8668 14952 8720 14958
rect 8668 14894 8720 14900
rect 8747 14716 9055 14725
rect 8747 14714 8753 14716
rect 8809 14714 8833 14716
rect 8889 14714 8913 14716
rect 8969 14714 8993 14716
rect 9049 14714 9055 14716
rect 8809 14662 8811 14714
rect 8991 14662 8993 14714
rect 8747 14660 8753 14662
rect 8809 14660 8833 14662
rect 8889 14660 8913 14662
rect 8969 14660 8993 14662
rect 9049 14660 9055 14662
rect 8747 14651 9055 14660
rect 8496 14470 8708 14498
rect 8576 13252 8628 13258
rect 8576 13194 8628 13200
rect 8588 11880 8616 13194
rect 8496 11852 8616 11880
rect 8496 10010 8524 11852
rect 8576 11756 8628 11762
rect 8576 11698 8628 11704
rect 8588 10810 8616 11698
rect 8576 10804 8628 10810
rect 8576 10746 8628 10752
rect 8496 9982 8616 10010
rect 8484 9920 8536 9926
rect 8484 9862 8536 9868
rect 8496 9722 8524 9862
rect 8484 9716 8536 9722
rect 8484 9658 8536 9664
rect 8484 9036 8536 9042
rect 8484 8978 8536 8984
rect 8392 8968 8444 8974
rect 8392 8910 8444 8916
rect 8496 8566 8524 8978
rect 8588 8673 8616 9982
rect 8574 8664 8630 8673
rect 8574 8599 8576 8608
rect 8628 8599 8630 8608
rect 8576 8570 8628 8576
rect 8484 8560 8536 8566
rect 8484 8502 8536 8508
rect 8496 8242 8524 8502
rect 8496 8214 8616 8242
rect 8312 8078 8524 8106
rect 8588 8090 8616 8214
rect 8392 8016 8444 8022
rect 8390 7984 8392 7993
rect 8444 7984 8446 7993
rect 8390 7919 8446 7928
rect 8208 7880 8260 7886
rect 8208 7822 8260 7828
rect 8300 7880 8352 7886
rect 8300 7822 8352 7828
rect 8392 7880 8444 7886
rect 8496 7868 8524 8078
rect 8576 8084 8628 8090
rect 8576 8026 8628 8032
rect 8444 7840 8524 7868
rect 8392 7822 8444 7828
rect 8024 7744 8076 7750
rect 8024 7686 8076 7692
rect 8116 7744 8168 7750
rect 8116 7686 8168 7692
rect 7932 7268 7984 7274
rect 7932 7210 7984 7216
rect 7748 7200 7800 7206
rect 7748 7142 7800 7148
rect 7760 7041 7788 7142
rect 7746 7032 7802 7041
rect 7746 6967 7802 6976
rect 7656 6656 7708 6662
rect 7656 6598 7708 6604
rect 7838 6624 7894 6633
rect 7668 6390 7696 6598
rect 7838 6559 7894 6568
rect 7564 6384 7616 6390
rect 7564 6326 7616 6332
rect 7656 6384 7708 6390
rect 7656 6326 7708 6332
rect 7576 5778 7604 6326
rect 7564 5772 7616 5778
rect 7564 5714 7616 5720
rect 7852 4078 7880 6559
rect 8036 5710 8064 7686
rect 8128 6390 8156 7686
rect 8312 7546 8340 7822
rect 8588 7800 8616 8026
rect 8496 7772 8616 7800
rect 8392 7744 8444 7750
rect 8392 7686 8444 7692
rect 8300 7540 8352 7546
rect 8300 7482 8352 7488
rect 8300 7336 8352 7342
rect 8300 7278 8352 7284
rect 8208 7268 8260 7274
rect 8208 7210 8260 7216
rect 8220 7002 8248 7210
rect 8208 6996 8260 7002
rect 8208 6938 8260 6944
rect 8312 6934 8340 7278
rect 8300 6928 8352 6934
rect 8300 6870 8352 6876
rect 8116 6384 8168 6390
rect 8116 6326 8168 6332
rect 8404 6089 8432 7686
rect 8496 6866 8524 7772
rect 8680 7290 8708 14470
rect 8747 13628 9055 13637
rect 8747 13626 8753 13628
rect 8809 13626 8833 13628
rect 8889 13626 8913 13628
rect 8969 13626 8993 13628
rect 9049 13626 9055 13628
rect 8809 13574 8811 13626
rect 8991 13574 8993 13626
rect 8747 13572 8753 13574
rect 8809 13572 8833 13574
rect 8889 13572 8913 13574
rect 8969 13572 8993 13574
rect 9049 13572 9055 13574
rect 8747 13563 9055 13572
rect 9140 13512 9168 14991
rect 9220 13864 9272 13870
rect 9220 13806 9272 13812
rect 9048 13484 9168 13512
rect 8852 12844 8904 12850
rect 8852 12786 8904 12792
rect 8864 12628 8892 12786
rect 9048 12753 9076 13484
rect 9232 13326 9260 13806
rect 9220 13320 9272 13326
rect 9220 13262 9272 13268
rect 9220 13184 9272 13190
rect 9220 13126 9272 13132
rect 9034 12744 9090 12753
rect 9034 12679 9090 12688
rect 8864 12600 9168 12628
rect 8747 12540 9055 12549
rect 8747 12538 8753 12540
rect 8809 12538 8833 12540
rect 8889 12538 8913 12540
rect 8969 12538 8993 12540
rect 9049 12538 9055 12540
rect 8809 12486 8811 12538
rect 8991 12486 8993 12538
rect 8747 12484 8753 12486
rect 8809 12484 8833 12486
rect 8889 12484 8913 12486
rect 8969 12484 8993 12486
rect 9049 12484 9055 12486
rect 8747 12475 9055 12484
rect 8747 11452 9055 11461
rect 8747 11450 8753 11452
rect 8809 11450 8833 11452
rect 8889 11450 8913 11452
rect 8969 11450 8993 11452
rect 9049 11450 9055 11452
rect 8809 11398 8811 11450
rect 8991 11398 8993 11450
rect 8747 11396 8753 11398
rect 8809 11396 8833 11398
rect 8889 11396 8913 11398
rect 8969 11396 8993 11398
rect 9049 11396 9055 11398
rect 8747 11387 9055 11396
rect 9036 11348 9088 11354
rect 9036 11290 9088 11296
rect 9048 11150 9076 11290
rect 9036 11144 9088 11150
rect 9036 11086 9088 11092
rect 9048 10470 9076 11086
rect 9140 10742 9168 12600
rect 9128 10736 9180 10742
rect 9128 10678 9180 10684
rect 9036 10464 9088 10470
rect 9036 10406 9088 10412
rect 8747 10364 9055 10373
rect 8747 10362 8753 10364
rect 8809 10362 8833 10364
rect 8889 10362 8913 10364
rect 8969 10362 8993 10364
rect 9049 10362 9055 10364
rect 8809 10310 8811 10362
rect 8991 10310 8993 10362
rect 8747 10308 8753 10310
rect 8809 10308 8833 10310
rect 8889 10308 8913 10310
rect 8969 10308 8993 10310
rect 9049 10308 9055 10310
rect 8747 10299 9055 10308
rect 8760 10056 8812 10062
rect 8760 9998 8812 10004
rect 8772 9761 8800 9998
rect 9128 9920 9180 9926
rect 9128 9862 9180 9868
rect 8758 9752 8814 9761
rect 8758 9687 8814 9696
rect 9140 9586 9168 9862
rect 9128 9580 9180 9586
rect 9128 9522 9180 9528
rect 8747 9276 9055 9285
rect 8747 9274 8753 9276
rect 8809 9274 8833 9276
rect 8889 9274 8913 9276
rect 8969 9274 8993 9276
rect 9049 9274 9055 9276
rect 8809 9222 8811 9274
rect 8991 9222 8993 9274
rect 8747 9220 8753 9222
rect 8809 9220 8833 9222
rect 8889 9220 8913 9222
rect 8969 9220 8993 9222
rect 9049 9220 9055 9222
rect 8747 9211 9055 9220
rect 9140 9160 9168 9522
rect 8956 9132 9168 9160
rect 8956 8294 8984 9132
rect 9232 8922 9260 13126
rect 9324 12918 9352 15370
rect 9312 12912 9364 12918
rect 9312 12854 9364 12860
rect 9312 12232 9364 12238
rect 9312 12174 9364 12180
rect 9140 8894 9260 8922
rect 8944 8288 8996 8294
rect 8944 8230 8996 8236
rect 8747 8188 9055 8197
rect 8747 8186 8753 8188
rect 8809 8186 8833 8188
rect 8889 8186 8913 8188
rect 8969 8186 8993 8188
rect 9049 8186 9055 8188
rect 8809 8134 8811 8186
rect 8991 8134 8993 8186
rect 8747 8132 8753 8134
rect 8809 8132 8833 8134
rect 8889 8132 8913 8134
rect 8969 8132 8993 8134
rect 9049 8132 9055 8134
rect 8747 8123 9055 8132
rect 8852 8084 8904 8090
rect 8852 8026 8904 8032
rect 8864 7857 8892 8026
rect 8850 7848 8906 7857
rect 8760 7812 8812 7818
rect 8850 7783 8906 7792
rect 8760 7754 8812 7760
rect 8772 7721 8800 7754
rect 8758 7712 8814 7721
rect 8758 7647 8814 7656
rect 8760 7404 8812 7410
rect 8760 7346 8812 7352
rect 8588 7262 8708 7290
rect 8484 6860 8536 6866
rect 8484 6802 8536 6808
rect 8390 6080 8446 6089
rect 8390 6015 8446 6024
rect 8024 5704 8076 5710
rect 8024 5646 8076 5652
rect 8208 5704 8260 5710
rect 8208 5646 8260 5652
rect 7840 4072 7892 4078
rect 7470 4040 7526 4049
rect 7840 4014 7892 4020
rect 7470 3975 7526 3984
rect 7286 3904 7342 3913
rect 7286 3839 7342 3848
rect 7196 3596 7248 3602
rect 7196 3538 7248 3544
rect 7300 3482 7328 3839
rect 7656 3528 7708 3534
rect 7208 3454 7328 3482
rect 7484 3476 7656 3482
rect 7484 3470 7708 3476
rect 7748 3528 7800 3534
rect 7748 3470 7800 3476
rect 7484 3454 7696 3470
rect 7208 3058 7236 3454
rect 7196 3052 7248 3058
rect 7380 3052 7432 3058
rect 7196 2994 7248 3000
rect 7300 3012 7380 3040
rect 7104 2916 7156 2922
rect 7104 2858 7156 2864
rect 7024 2746 7144 2774
rect 6920 2440 6972 2446
rect 6920 2382 6972 2388
rect 6920 2304 6972 2310
rect 6920 2246 6972 2252
rect 7012 2304 7064 2310
rect 7012 2246 7064 2252
rect 6828 1964 6880 1970
rect 6828 1906 6880 1912
rect 6828 1352 6880 1358
rect 6828 1294 6880 1300
rect 6736 1012 6788 1018
rect 6736 954 6788 960
rect 6840 160 6868 1294
rect 6932 1018 6960 2246
rect 7024 1873 7052 2246
rect 7010 1864 7066 1873
rect 7010 1799 7066 1808
rect 7116 1562 7144 2746
rect 7194 2680 7250 2689
rect 7194 2615 7196 2624
rect 7248 2615 7250 2624
rect 7196 2586 7248 2592
rect 7196 2304 7248 2310
rect 7196 2246 7248 2252
rect 7208 2106 7236 2246
rect 7196 2100 7248 2106
rect 7196 2042 7248 2048
rect 7196 1760 7248 1766
rect 7196 1702 7248 1708
rect 7104 1556 7156 1562
rect 7104 1498 7156 1504
rect 7208 1465 7236 1702
rect 7194 1456 7250 1465
rect 7194 1391 7250 1400
rect 7104 1352 7156 1358
rect 7104 1294 7156 1300
rect 6920 1012 6972 1018
rect 6920 954 6972 960
rect 6274 82 6330 160
rect 6196 54 6330 82
rect 6274 -300 6330 54
rect 6458 -300 6514 160
rect 6642 -300 6698 160
rect 6826 -300 6882 160
rect 7010 82 7066 160
rect 7116 82 7144 1294
rect 7300 1290 7328 3012
rect 7380 2994 7432 3000
rect 7380 2848 7432 2854
rect 7380 2790 7432 2796
rect 7392 2038 7420 2790
rect 7380 2032 7432 2038
rect 7380 1974 7432 1980
rect 7380 1352 7432 1358
rect 7378 1320 7380 1329
rect 7432 1320 7434 1329
rect 7288 1284 7340 1290
rect 7378 1255 7434 1264
rect 7288 1226 7340 1232
rect 7196 1216 7248 1222
rect 7196 1158 7248 1164
rect 7208 160 7236 1158
rect 7010 54 7144 82
rect 7010 -300 7066 54
rect 7194 -300 7250 160
rect 7378 82 7434 160
rect 7484 82 7512 3454
rect 7564 3392 7616 3398
rect 7564 3334 7616 3340
rect 7576 2446 7604 3334
rect 7760 2938 7788 3470
rect 7840 3052 7892 3058
rect 7892 3012 8156 3040
rect 7840 2994 7892 3000
rect 7760 2910 7880 2938
rect 7656 2848 7708 2854
rect 7656 2790 7708 2796
rect 7748 2848 7800 2854
rect 7748 2790 7800 2796
rect 7668 2446 7696 2790
rect 7564 2440 7616 2446
rect 7564 2382 7616 2388
rect 7656 2440 7708 2446
rect 7760 2428 7788 2790
rect 7852 2496 7880 2910
rect 7932 2848 7984 2854
rect 7984 2808 8064 2836
rect 7932 2790 7984 2796
rect 7930 2680 7986 2689
rect 7930 2615 7932 2624
rect 7984 2615 7986 2624
rect 7932 2586 7984 2592
rect 7852 2468 7972 2496
rect 7760 2400 7880 2428
rect 7656 2382 7708 2388
rect 7852 2038 7880 2400
rect 7840 2032 7892 2038
rect 7840 1974 7892 1980
rect 7654 1864 7710 1873
rect 7944 1816 7972 2468
rect 8036 2106 8064 2808
rect 8024 2100 8076 2106
rect 8024 2042 8076 2048
rect 8024 1896 8076 1902
rect 8024 1838 8076 1844
rect 7654 1799 7710 1808
rect 7668 1766 7696 1799
rect 7760 1788 7972 1816
rect 7656 1760 7708 1766
rect 7656 1702 7708 1708
rect 7564 1556 7616 1562
rect 7564 1498 7616 1504
rect 7576 160 7604 1498
rect 7760 160 7788 1788
rect 8036 1562 8064 1838
rect 8024 1556 8076 1562
rect 8024 1498 8076 1504
rect 7840 1284 7892 1290
rect 7840 1226 7892 1232
rect 7378 54 7512 82
rect 7378 -300 7434 54
rect 7562 -300 7618 160
rect 7746 -300 7802 160
rect 7852 82 7880 1226
rect 8128 160 8156 3012
rect 8220 2961 8248 5646
rect 8496 5370 8524 6802
rect 8484 5364 8536 5370
rect 8484 5306 8536 5312
rect 8588 3584 8616 7262
rect 8772 7188 8800 7346
rect 8680 7160 8800 7188
rect 8680 7002 8708 7160
rect 8747 7100 9055 7109
rect 8747 7098 8753 7100
rect 8809 7098 8833 7100
rect 8889 7098 8913 7100
rect 8969 7098 8993 7100
rect 9049 7098 9055 7100
rect 8809 7046 8811 7098
rect 8991 7046 8993 7098
rect 8747 7044 8753 7046
rect 8809 7044 8833 7046
rect 8889 7044 8913 7046
rect 8969 7044 8993 7046
rect 9049 7044 9055 7046
rect 8747 7035 9055 7044
rect 8668 6996 8720 7002
rect 8668 6938 8720 6944
rect 8747 6012 9055 6021
rect 8747 6010 8753 6012
rect 8809 6010 8833 6012
rect 8889 6010 8913 6012
rect 8969 6010 8993 6012
rect 9049 6010 9055 6012
rect 8809 5958 8811 6010
rect 8991 5958 8993 6010
rect 8747 5956 8753 5958
rect 8809 5956 8833 5958
rect 8889 5956 8913 5958
rect 8969 5956 8993 5958
rect 9049 5956 9055 5958
rect 8747 5947 9055 5956
rect 8942 5672 8998 5681
rect 9140 5658 9168 8894
rect 9220 8832 9272 8838
rect 9220 8774 9272 8780
rect 8998 5630 9168 5658
rect 8942 5607 8998 5616
rect 8747 4924 9055 4933
rect 8747 4922 8753 4924
rect 8809 4922 8833 4924
rect 8889 4922 8913 4924
rect 8969 4922 8993 4924
rect 9049 4922 9055 4924
rect 8809 4870 8811 4922
rect 8991 4870 8993 4922
rect 8747 4868 8753 4870
rect 8809 4868 8833 4870
rect 8889 4868 8913 4870
rect 8969 4868 8993 4870
rect 9049 4868 9055 4870
rect 8747 4859 9055 4868
rect 9232 4729 9260 8774
rect 9324 8634 9352 12174
rect 9312 8628 9364 8634
rect 9312 8570 9364 8576
rect 9312 8288 9364 8294
rect 9312 8230 9364 8236
rect 9324 7274 9352 8230
rect 9312 7268 9364 7274
rect 9312 7210 9364 7216
rect 9312 6860 9364 6866
rect 9312 6802 9364 6808
rect 9324 6322 9352 6802
rect 9312 6316 9364 6322
rect 9312 6258 9364 6264
rect 9218 4720 9274 4729
rect 9218 4655 9274 4664
rect 8747 3836 9055 3845
rect 8747 3834 8753 3836
rect 8809 3834 8833 3836
rect 8889 3834 8913 3836
rect 8969 3834 8993 3836
rect 9049 3834 9055 3836
rect 8809 3782 8811 3834
rect 8991 3782 8993 3834
rect 8747 3780 8753 3782
rect 8809 3780 8833 3782
rect 8889 3780 8913 3782
rect 8969 3780 8993 3782
rect 9049 3780 9055 3782
rect 8747 3771 9055 3780
rect 8668 3596 8720 3602
rect 8588 3556 8668 3584
rect 8668 3538 8720 3544
rect 9416 3534 9444 17190
rect 9496 16992 9548 16998
rect 9496 16934 9548 16940
rect 9508 15162 9536 16934
rect 9600 15881 9628 17711
rect 9784 17270 9812 18906
rect 9772 17264 9824 17270
rect 9772 17206 9824 17212
rect 9678 16552 9734 16561
rect 9678 16487 9734 16496
rect 9692 16182 9720 16487
rect 9680 16176 9732 16182
rect 9680 16118 9732 16124
rect 9680 16040 9732 16046
rect 9680 15982 9732 15988
rect 9586 15872 9642 15881
rect 9586 15807 9642 15816
rect 9496 15156 9548 15162
rect 9496 15098 9548 15104
rect 9496 13796 9548 13802
rect 9496 13738 9548 13744
rect 9508 13530 9536 13738
rect 9586 13560 9642 13569
rect 9496 13524 9548 13530
rect 9586 13495 9642 13504
rect 9496 13466 9548 13472
rect 9600 12424 9628 13495
rect 9692 13326 9720 15982
rect 9784 14618 9812 17206
rect 9876 17134 9904 19314
rect 9968 18698 9996 20318
rect 10060 20233 10088 20946
rect 10046 20224 10102 20233
rect 10046 20159 10102 20168
rect 9956 18692 10008 18698
rect 9956 18634 10008 18640
rect 9968 18601 9996 18634
rect 9954 18592 10010 18601
rect 9954 18527 10010 18536
rect 10060 18306 10088 20159
rect 10152 19854 10180 24006
rect 10244 21690 10272 24364
rect 10322 24304 10378 24313
rect 10322 24239 10378 24248
rect 10336 24206 10364 24239
rect 10324 24200 10376 24206
rect 10324 24142 10376 24148
rect 10336 23905 10364 24142
rect 10322 23896 10378 23905
rect 10322 23831 10378 23840
rect 10324 23044 10376 23050
rect 10324 22986 10376 22992
rect 10336 22778 10364 22986
rect 10324 22772 10376 22778
rect 10324 22714 10376 22720
rect 10336 22642 10364 22714
rect 10324 22636 10376 22642
rect 10324 22578 10376 22584
rect 10322 22400 10378 22409
rect 10322 22335 10378 22344
rect 10336 22030 10364 22335
rect 10324 22024 10376 22030
rect 10324 21966 10376 21972
rect 10232 21684 10284 21690
rect 10232 21626 10284 21632
rect 10140 19848 10192 19854
rect 10140 19790 10192 19796
rect 10152 18834 10180 19790
rect 10244 18873 10272 21626
rect 10324 21344 10376 21350
rect 10322 21312 10324 21321
rect 10376 21312 10378 21321
rect 10322 21247 10378 21256
rect 10324 20800 10376 20806
rect 10324 20742 10376 20748
rect 10336 20466 10364 20742
rect 10324 20460 10376 20466
rect 10324 20402 10376 20408
rect 10428 20074 10456 28358
rect 10520 26246 10548 34886
rect 10692 34604 10744 34610
rect 10692 34546 10744 34552
rect 10600 34468 10652 34474
rect 10600 34410 10652 34416
rect 10612 29714 10640 34410
rect 10704 34066 10732 34546
rect 10692 34060 10744 34066
rect 10692 34002 10744 34008
rect 10796 33522 10824 42588
rect 11152 42560 11204 42566
rect 10874 42528 10930 42537
rect 11152 42502 11204 42508
rect 11244 42560 11296 42566
rect 11244 42502 11296 42508
rect 10874 42463 10930 42472
rect 10888 37262 10916 42463
rect 11164 42265 11192 42502
rect 11256 42294 11284 42502
rect 11346 42460 11654 42469
rect 11346 42458 11352 42460
rect 11408 42458 11432 42460
rect 11488 42458 11512 42460
rect 11568 42458 11592 42460
rect 11648 42458 11654 42460
rect 11408 42406 11410 42458
rect 11590 42406 11592 42458
rect 11346 42404 11352 42406
rect 11408 42404 11432 42406
rect 11488 42404 11512 42406
rect 11568 42404 11592 42406
rect 11648 42404 11654 42406
rect 11346 42395 11654 42404
rect 11244 42288 11296 42294
rect 11150 42256 11206 42265
rect 11244 42230 11296 42236
rect 11150 42191 11206 42200
rect 11716 42090 11744 43046
rect 11808 42684 11836 44540
rect 11888 43308 11940 43314
rect 11992 43296 12020 44540
rect 12176 43790 12204 44540
rect 12360 43874 12388 44540
rect 12268 43846 12388 43874
rect 12164 43784 12216 43790
rect 12164 43726 12216 43732
rect 11940 43268 12020 43296
rect 12072 43308 12124 43314
rect 11888 43250 11940 43256
rect 12268 43296 12296 43846
rect 12348 43784 12400 43790
rect 12348 43726 12400 43732
rect 12360 43382 12388 43726
rect 12440 43648 12492 43654
rect 12440 43590 12492 43596
rect 12544 43602 12572 44540
rect 12452 43450 12480 43590
rect 12544 43574 12664 43602
rect 12440 43444 12492 43450
rect 12440 43386 12492 43392
rect 12348 43376 12400 43382
rect 12348 43318 12400 43324
rect 12124 43268 12296 43296
rect 12072 43250 12124 43256
rect 12070 43208 12126 43217
rect 12070 43143 12126 43152
rect 11888 42696 11940 42702
rect 11808 42656 11888 42684
rect 12084 42650 12112 43143
rect 12164 42900 12216 42906
rect 12164 42842 12216 42848
rect 11888 42638 11940 42644
rect 11992 42622 12112 42650
rect 11992 42242 12020 42622
rect 12072 42560 12124 42566
rect 12072 42502 12124 42508
rect 11808 42214 12020 42242
rect 11704 42084 11756 42090
rect 11704 42026 11756 42032
rect 11808 41414 11836 42214
rect 11980 42084 12032 42090
rect 11980 42026 12032 42032
rect 11716 41386 11836 41414
rect 11346 41372 11654 41381
rect 11346 41370 11352 41372
rect 11408 41370 11432 41372
rect 11488 41370 11512 41372
rect 11568 41370 11592 41372
rect 11648 41370 11654 41372
rect 11408 41318 11410 41370
rect 11590 41318 11592 41370
rect 11346 41316 11352 41318
rect 11408 41316 11432 41318
rect 11488 41316 11512 41318
rect 11568 41316 11592 41318
rect 11648 41316 11654 41318
rect 11346 41307 11654 41316
rect 11152 41132 11204 41138
rect 11152 41074 11204 41080
rect 11060 40996 11112 41002
rect 11060 40938 11112 40944
rect 11072 38457 11100 40938
rect 11058 38448 11114 38457
rect 11058 38383 11114 38392
rect 11164 38298 11192 41074
rect 11346 40284 11654 40293
rect 11346 40282 11352 40284
rect 11408 40282 11432 40284
rect 11488 40282 11512 40284
rect 11568 40282 11592 40284
rect 11648 40282 11654 40284
rect 11408 40230 11410 40282
rect 11590 40230 11592 40282
rect 11346 40228 11352 40230
rect 11408 40228 11432 40230
rect 11488 40228 11512 40230
rect 11568 40228 11592 40230
rect 11648 40228 11654 40230
rect 11346 40219 11654 40228
rect 11346 39196 11654 39205
rect 11346 39194 11352 39196
rect 11408 39194 11432 39196
rect 11488 39194 11512 39196
rect 11568 39194 11592 39196
rect 11648 39194 11654 39196
rect 11408 39142 11410 39194
rect 11590 39142 11592 39194
rect 11346 39140 11352 39142
rect 11408 39140 11432 39142
rect 11488 39140 11512 39142
rect 11568 39140 11592 39142
rect 11648 39140 11654 39142
rect 11346 39131 11654 39140
rect 11072 38270 11192 38298
rect 11716 38282 11744 41386
rect 11888 38820 11940 38826
rect 11888 38762 11940 38768
rect 11704 38276 11756 38282
rect 10876 37256 10928 37262
rect 10876 37198 10928 37204
rect 10968 37188 11020 37194
rect 10968 37130 11020 37136
rect 10980 36378 11008 37130
rect 10968 36372 11020 36378
rect 10968 36314 11020 36320
rect 10980 36009 11008 36314
rect 10966 36000 11022 36009
rect 10966 35935 11022 35944
rect 10968 35624 11020 35630
rect 10968 35566 11020 35572
rect 10874 35184 10930 35193
rect 10874 35119 10930 35128
rect 10888 35018 10916 35119
rect 10876 35012 10928 35018
rect 10876 34954 10928 34960
rect 10876 34740 10928 34746
rect 10876 34682 10928 34688
rect 10888 34513 10916 34682
rect 10874 34504 10930 34513
rect 10874 34439 10930 34448
rect 10980 33946 11008 35566
rect 11072 35476 11100 38270
rect 11704 38218 11756 38224
rect 11346 38108 11654 38117
rect 11346 38106 11352 38108
rect 11408 38106 11432 38108
rect 11488 38106 11512 38108
rect 11568 38106 11592 38108
rect 11648 38106 11654 38108
rect 11408 38054 11410 38106
rect 11590 38054 11592 38106
rect 11346 38052 11352 38054
rect 11408 38052 11432 38054
rect 11488 38052 11512 38054
rect 11568 38052 11592 38054
rect 11648 38052 11654 38054
rect 11346 38043 11654 38052
rect 11244 37868 11296 37874
rect 11244 37810 11296 37816
rect 11152 37664 11204 37670
rect 11152 37606 11204 37612
rect 11164 35630 11192 37606
rect 11256 36156 11284 37810
rect 11716 37262 11744 38218
rect 11704 37256 11756 37262
rect 11334 37224 11390 37233
rect 11704 37198 11756 37204
rect 11334 37159 11390 37168
rect 11348 37126 11376 37159
rect 11336 37120 11388 37126
rect 11336 37062 11388 37068
rect 11346 37020 11654 37029
rect 11346 37018 11352 37020
rect 11408 37018 11432 37020
rect 11488 37018 11512 37020
rect 11568 37018 11592 37020
rect 11648 37018 11654 37020
rect 11408 36966 11410 37018
rect 11590 36966 11592 37018
rect 11346 36964 11352 36966
rect 11408 36964 11432 36966
rect 11488 36964 11512 36966
rect 11568 36964 11592 36966
rect 11648 36964 11654 36966
rect 11346 36955 11654 36964
rect 11704 36780 11756 36786
rect 11704 36722 11756 36728
rect 11428 36168 11480 36174
rect 11256 36128 11428 36156
rect 11428 36110 11480 36116
rect 11346 35932 11654 35941
rect 11346 35930 11352 35932
rect 11408 35930 11432 35932
rect 11488 35930 11512 35932
rect 11568 35930 11592 35932
rect 11648 35930 11654 35932
rect 11408 35878 11410 35930
rect 11590 35878 11592 35930
rect 11346 35876 11352 35878
rect 11408 35876 11432 35878
rect 11488 35876 11512 35878
rect 11568 35876 11592 35878
rect 11648 35876 11654 35878
rect 11346 35867 11654 35876
rect 11610 35728 11666 35737
rect 11716 35698 11744 36722
rect 11796 36644 11848 36650
rect 11796 36586 11848 36592
rect 11610 35663 11666 35672
rect 11704 35692 11756 35698
rect 11152 35624 11204 35630
rect 11152 35566 11204 35572
rect 11072 35448 11192 35476
rect 11060 34400 11112 34406
rect 11060 34342 11112 34348
rect 11072 34202 11100 34342
rect 11060 34196 11112 34202
rect 11060 34138 11112 34144
rect 10888 33918 11008 33946
rect 10888 33590 10916 33918
rect 10968 33856 11020 33862
rect 10968 33798 11020 33804
rect 10876 33584 10928 33590
rect 10876 33526 10928 33532
rect 10784 33516 10836 33522
rect 10784 33458 10836 33464
rect 10782 33416 10838 33425
rect 10782 33351 10838 33360
rect 10796 33318 10824 33351
rect 10784 33312 10836 33318
rect 10784 33254 10836 33260
rect 10980 32978 11008 33798
rect 11072 33590 11100 34138
rect 11060 33584 11112 33590
rect 11164 33572 11192 35448
rect 11624 35086 11652 35663
rect 11704 35634 11756 35640
rect 11808 35290 11836 36586
rect 11796 35284 11848 35290
rect 11796 35226 11848 35232
rect 11612 35080 11664 35086
rect 11612 35022 11664 35028
rect 11796 35080 11848 35086
rect 11796 35022 11848 35028
rect 11244 35012 11296 35018
rect 11244 34954 11296 34960
rect 11256 33969 11284 34954
rect 11346 34844 11654 34853
rect 11346 34842 11352 34844
rect 11408 34842 11432 34844
rect 11488 34842 11512 34844
rect 11568 34842 11592 34844
rect 11648 34842 11654 34844
rect 11408 34790 11410 34842
rect 11590 34790 11592 34842
rect 11346 34788 11352 34790
rect 11408 34788 11432 34790
rect 11488 34788 11512 34790
rect 11568 34788 11592 34790
rect 11648 34788 11654 34790
rect 11346 34779 11654 34788
rect 11336 34672 11388 34678
rect 11808 34649 11836 35022
rect 11336 34614 11388 34620
rect 11794 34640 11850 34649
rect 11242 33960 11298 33969
rect 11242 33895 11298 33904
rect 11348 33844 11376 34614
rect 11794 34575 11850 34584
rect 11900 34105 11928 38762
rect 11702 34096 11758 34105
rect 11702 34031 11758 34040
rect 11886 34096 11942 34105
rect 11886 34031 11942 34040
rect 11256 33816 11376 33844
rect 11256 33640 11284 33816
rect 11346 33756 11654 33765
rect 11346 33754 11352 33756
rect 11408 33754 11432 33756
rect 11488 33754 11512 33756
rect 11568 33754 11592 33756
rect 11648 33754 11654 33756
rect 11408 33702 11410 33754
rect 11590 33702 11592 33754
rect 11346 33700 11352 33702
rect 11408 33700 11432 33702
rect 11488 33700 11512 33702
rect 11568 33700 11592 33702
rect 11648 33700 11654 33702
rect 11346 33691 11654 33700
rect 11716 33674 11744 34031
rect 11794 33688 11850 33697
rect 11716 33646 11794 33674
rect 11256 33612 11468 33640
rect 11794 33623 11850 33632
rect 11164 33544 11376 33572
rect 11060 33526 11112 33532
rect 11152 33448 11204 33454
rect 11058 33416 11114 33425
rect 11152 33390 11204 33396
rect 11058 33351 11114 33360
rect 10968 32972 11020 32978
rect 10968 32914 11020 32920
rect 10876 32904 10928 32910
rect 10876 32846 10928 32852
rect 10784 32768 10836 32774
rect 10784 32710 10836 32716
rect 10690 32464 10746 32473
rect 10690 32399 10692 32408
rect 10744 32399 10746 32408
rect 10692 32370 10744 32376
rect 10692 32224 10744 32230
rect 10692 32166 10744 32172
rect 10704 31890 10732 32166
rect 10692 31884 10744 31890
rect 10692 31826 10744 31832
rect 10796 31686 10824 32710
rect 10888 32026 10916 32846
rect 11072 32745 11100 33351
rect 11058 32736 11114 32745
rect 11058 32671 11114 32680
rect 10968 32564 11020 32570
rect 10968 32506 11020 32512
rect 10980 32337 11008 32506
rect 11060 32428 11112 32434
rect 11060 32370 11112 32376
rect 10966 32328 11022 32337
rect 10966 32263 11022 32272
rect 10876 32020 10928 32026
rect 10876 31962 10928 31968
rect 10968 31816 11020 31822
rect 10968 31758 11020 31764
rect 10784 31680 10836 31686
rect 10784 31622 10836 31628
rect 10980 31482 11008 31758
rect 10968 31476 11020 31482
rect 10968 31418 11020 31424
rect 10876 31272 10928 31278
rect 10876 31214 10928 31220
rect 10692 30320 10744 30326
rect 10692 30262 10744 30268
rect 10600 29708 10652 29714
rect 10600 29650 10652 29656
rect 10612 29102 10640 29650
rect 10600 29096 10652 29102
rect 10600 29038 10652 29044
rect 10704 28966 10732 30262
rect 10888 29646 10916 31214
rect 11072 30938 11100 32370
rect 11164 31890 11192 33390
rect 11244 33312 11296 33318
rect 11244 33254 11296 33260
rect 11256 32910 11284 33254
rect 11244 32904 11296 32910
rect 11244 32846 11296 32852
rect 11348 32756 11376 33544
rect 11440 33454 11468 33612
rect 11428 33448 11480 33454
rect 11428 33390 11480 33396
rect 11794 33144 11850 33153
rect 11794 33079 11850 33088
rect 11704 32904 11756 32910
rect 11704 32846 11756 32852
rect 11256 32728 11376 32756
rect 11256 32298 11284 32728
rect 11346 32668 11654 32677
rect 11346 32666 11352 32668
rect 11408 32666 11432 32668
rect 11488 32666 11512 32668
rect 11568 32666 11592 32668
rect 11648 32666 11654 32668
rect 11408 32614 11410 32666
rect 11590 32614 11592 32666
rect 11346 32612 11352 32614
rect 11408 32612 11432 32614
rect 11488 32612 11512 32614
rect 11568 32612 11592 32614
rect 11648 32612 11654 32614
rect 11346 32603 11654 32612
rect 11336 32428 11388 32434
rect 11336 32370 11388 32376
rect 11244 32292 11296 32298
rect 11244 32234 11296 32240
rect 11152 31884 11204 31890
rect 11152 31826 11204 31832
rect 11060 30932 11112 30938
rect 11060 30874 11112 30880
rect 10966 30424 11022 30433
rect 10966 30359 11022 30368
rect 10980 30274 11008 30359
rect 10980 30246 11100 30274
rect 10968 29844 11020 29850
rect 10968 29786 11020 29792
rect 10876 29640 10928 29646
rect 10782 29608 10838 29617
rect 10876 29582 10928 29588
rect 10782 29543 10838 29552
rect 10796 29034 10824 29543
rect 10888 29170 10916 29582
rect 10980 29238 11008 29786
rect 10968 29232 11020 29238
rect 10968 29174 11020 29180
rect 10876 29164 10928 29170
rect 10876 29106 10928 29112
rect 10784 29028 10836 29034
rect 10784 28970 10836 28976
rect 10692 28960 10744 28966
rect 10692 28902 10744 28908
rect 10704 27962 10732 28902
rect 10888 28257 10916 29106
rect 10874 28248 10930 28257
rect 10980 28218 11008 29174
rect 11072 28801 11100 30246
rect 11058 28792 11114 28801
rect 11058 28727 11114 28736
rect 11060 28552 11112 28558
rect 11060 28494 11112 28500
rect 10874 28183 10930 28192
rect 10968 28212 11020 28218
rect 10968 28154 11020 28160
rect 11072 28014 11100 28494
rect 11060 28008 11112 28014
rect 10704 27934 11008 27962
rect 11060 27950 11112 27956
rect 10600 27396 10652 27402
rect 10600 27338 10652 27344
rect 10508 26240 10560 26246
rect 10508 26182 10560 26188
rect 10612 25906 10640 27338
rect 10784 27328 10836 27334
rect 10784 27270 10836 27276
rect 10692 27124 10744 27130
rect 10692 27066 10744 27072
rect 10704 26994 10732 27066
rect 10796 27062 10824 27270
rect 10784 27056 10836 27062
rect 10784 26998 10836 27004
rect 10692 26988 10744 26994
rect 10692 26930 10744 26936
rect 10600 25900 10652 25906
rect 10600 25842 10652 25848
rect 10508 24812 10560 24818
rect 10508 24754 10560 24760
rect 10520 23905 10548 24754
rect 10598 24712 10654 24721
rect 10598 24647 10654 24656
rect 10506 23896 10562 23905
rect 10506 23831 10562 23840
rect 10508 23588 10560 23594
rect 10508 23530 10560 23536
rect 10520 22778 10548 23530
rect 10508 22772 10560 22778
rect 10508 22714 10560 22720
rect 10508 22636 10560 22642
rect 10508 22578 10560 22584
rect 10520 21010 10548 22578
rect 10612 22556 10640 24647
rect 10704 23322 10732 26930
rect 10784 26376 10836 26382
rect 10876 26376 10928 26382
rect 10784 26318 10836 26324
rect 10874 26344 10876 26353
rect 10928 26344 10930 26353
rect 10796 25945 10824 26318
rect 10874 26279 10930 26288
rect 10876 26036 10928 26042
rect 10876 25978 10928 25984
rect 10782 25936 10838 25945
rect 10782 25871 10838 25880
rect 10784 25696 10836 25702
rect 10784 25638 10836 25644
rect 10796 25498 10824 25638
rect 10784 25492 10836 25498
rect 10784 25434 10836 25440
rect 10784 24880 10836 24886
rect 10784 24822 10836 24828
rect 10692 23316 10744 23322
rect 10692 23258 10744 23264
rect 10692 22976 10744 22982
rect 10692 22918 10744 22924
rect 10704 22710 10732 22918
rect 10692 22704 10744 22710
rect 10692 22646 10744 22652
rect 10612 22528 10732 22556
rect 10600 22092 10652 22098
rect 10600 22034 10652 22040
rect 10508 21004 10560 21010
rect 10508 20946 10560 20952
rect 10612 20942 10640 22034
rect 10600 20936 10652 20942
rect 10600 20878 10652 20884
rect 10704 20788 10732 22528
rect 10336 20046 10456 20074
rect 10520 20760 10732 20788
rect 10230 18864 10286 18873
rect 10140 18828 10192 18834
rect 10230 18799 10286 18808
rect 10140 18770 10192 18776
rect 10336 18408 10364 20046
rect 10416 19916 10468 19922
rect 10416 19858 10468 19864
rect 10428 18970 10456 19858
rect 10416 18964 10468 18970
rect 10416 18906 10468 18912
rect 10336 18380 10456 18408
rect 10060 18290 10272 18306
rect 9956 18284 10008 18290
rect 10060 18284 10284 18290
rect 10060 18278 10232 18284
rect 9956 18226 10008 18232
rect 10284 18244 10364 18272
rect 10232 18226 10284 18232
rect 9968 17882 9996 18226
rect 10048 18216 10100 18222
rect 10048 18158 10100 18164
rect 10060 17882 10088 18158
rect 9956 17876 10008 17882
rect 9956 17818 10008 17824
rect 10048 17876 10100 17882
rect 10048 17818 10100 17824
rect 9954 17504 10010 17513
rect 9954 17439 10010 17448
rect 9864 17128 9916 17134
rect 9864 17070 9916 17076
rect 9968 16402 9996 17439
rect 10232 17332 10284 17338
rect 10232 17274 10284 17280
rect 10140 16584 10192 16590
rect 10140 16526 10192 16532
rect 9876 16374 9996 16402
rect 10048 16448 10100 16454
rect 10048 16390 10100 16396
rect 9772 14612 9824 14618
rect 9772 14554 9824 14560
rect 9876 14498 9904 16374
rect 9956 16244 10008 16250
rect 9956 16186 10008 16192
rect 9784 14470 9904 14498
rect 9784 13841 9812 14470
rect 9864 14408 9916 14414
rect 9864 14350 9916 14356
rect 9770 13832 9826 13841
rect 9770 13767 9826 13776
rect 9772 13728 9824 13734
rect 9772 13670 9824 13676
rect 9680 13320 9732 13326
rect 9680 13262 9732 13268
rect 9784 13002 9812 13670
rect 9876 13394 9904 14350
rect 9968 13938 9996 16186
rect 10060 16046 10088 16390
rect 10048 16040 10100 16046
rect 10048 15982 10100 15988
rect 10048 14816 10100 14822
rect 10048 14758 10100 14764
rect 10060 13938 10088 14758
rect 10152 14482 10180 16526
rect 10244 16046 10272 17274
rect 10232 16040 10284 16046
rect 10232 15982 10284 15988
rect 10232 15360 10284 15366
rect 10232 15302 10284 15308
rect 10244 14550 10272 15302
rect 10336 15094 10364 18244
rect 10428 17610 10456 18380
rect 10416 17604 10468 17610
rect 10416 17546 10468 17552
rect 10416 16992 10468 16998
rect 10416 16934 10468 16940
rect 10428 16436 10456 16934
rect 10520 16697 10548 20760
rect 10690 20360 10746 20369
rect 10690 20295 10746 20304
rect 10704 19786 10732 20295
rect 10692 19780 10744 19786
rect 10692 19722 10744 19728
rect 10704 19378 10732 19722
rect 10692 19372 10744 19378
rect 10692 19314 10744 19320
rect 10600 18420 10652 18426
rect 10600 18362 10652 18368
rect 10612 17678 10640 18362
rect 10692 18352 10744 18358
rect 10692 18294 10744 18300
rect 10704 18057 10732 18294
rect 10690 18048 10746 18057
rect 10690 17983 10746 17992
rect 10600 17672 10652 17678
rect 10600 17614 10652 17620
rect 10692 17672 10744 17678
rect 10692 17614 10744 17620
rect 10600 17196 10652 17202
rect 10600 17138 10652 17144
rect 10506 16688 10562 16697
rect 10506 16623 10562 16632
rect 10520 16590 10548 16623
rect 10508 16584 10560 16590
rect 10508 16526 10560 16532
rect 10428 16408 10548 16436
rect 10416 16040 10468 16046
rect 10416 15982 10468 15988
rect 10324 15088 10376 15094
rect 10324 15030 10376 15036
rect 10232 14544 10284 14550
rect 10232 14486 10284 14492
rect 10140 14476 10192 14482
rect 10140 14418 10192 14424
rect 9956 13932 10008 13938
rect 9956 13874 10008 13880
rect 10048 13932 10100 13938
rect 10048 13874 10100 13880
rect 10048 13524 10100 13530
rect 10048 13466 10100 13472
rect 9864 13388 9916 13394
rect 9864 13330 9916 13336
rect 9876 13025 9904 13330
rect 9956 13320 10008 13326
rect 9956 13262 10008 13268
rect 9692 12974 9812 13002
rect 9862 13016 9918 13025
rect 9692 12434 9720 12974
rect 9862 12951 9918 12960
rect 9968 12866 9996 13262
rect 9508 12396 9628 12424
rect 9690 12396 9720 12434
rect 9508 12102 9536 12396
rect 9692 12322 9720 12396
rect 9600 12294 9720 12322
rect 9784 12838 9996 12866
rect 9496 12096 9548 12102
rect 9494 12064 9496 12073
rect 9548 12064 9550 12073
rect 9494 11999 9550 12008
rect 9600 11880 9628 12294
rect 9680 12232 9732 12238
rect 9680 12174 9732 12180
rect 9508 11852 9628 11880
rect 9508 10577 9536 11852
rect 9588 11756 9640 11762
rect 9588 11698 9640 11704
rect 9600 10674 9628 11698
rect 9692 11354 9720 12174
rect 9784 11694 9812 12838
rect 9862 12744 9918 12753
rect 10060 12730 10088 13466
rect 9862 12679 9918 12688
rect 9968 12702 10088 12730
rect 9876 12238 9904 12679
rect 9864 12232 9916 12238
rect 9864 12174 9916 12180
rect 9772 11688 9824 11694
rect 9772 11630 9824 11636
rect 9680 11348 9732 11354
rect 9680 11290 9732 11296
rect 9784 11234 9812 11630
rect 9862 11248 9918 11257
rect 9784 11218 9862 11234
rect 9772 11212 9862 11218
rect 9824 11206 9862 11212
rect 9862 11183 9918 11192
rect 9772 11154 9824 11160
rect 9588 10668 9640 10674
rect 9588 10610 9640 10616
rect 9680 10668 9732 10674
rect 9680 10610 9732 10616
rect 9494 10568 9550 10577
rect 9494 10503 9550 10512
rect 9692 10248 9720 10610
rect 9968 10588 9996 12702
rect 10048 12640 10100 12646
rect 10048 12582 10100 12588
rect 10060 11762 10088 12582
rect 10152 12306 10180 14418
rect 10232 13864 10284 13870
rect 10232 13806 10284 13812
rect 10244 13025 10272 13806
rect 10230 13016 10286 13025
rect 10230 12951 10286 12960
rect 10230 12880 10286 12889
rect 10336 12850 10364 15030
rect 10428 13530 10456 15982
rect 10416 13524 10468 13530
rect 10416 13466 10468 13472
rect 10416 13388 10468 13394
rect 10416 13330 10468 13336
rect 10428 12918 10456 13330
rect 10416 12912 10468 12918
rect 10416 12854 10468 12860
rect 10230 12815 10286 12824
rect 10324 12844 10376 12850
rect 10244 12442 10272 12815
rect 10324 12786 10376 12792
rect 10520 12764 10548 16408
rect 10612 16114 10640 17138
rect 10704 16998 10732 17614
rect 10692 16992 10744 16998
rect 10692 16934 10744 16940
rect 10690 16824 10746 16833
rect 10690 16759 10746 16768
rect 10704 16726 10732 16759
rect 10692 16720 10744 16726
rect 10692 16662 10744 16668
rect 10600 16108 10652 16114
rect 10600 16050 10652 16056
rect 10612 14482 10640 16050
rect 10692 15904 10744 15910
rect 10692 15846 10744 15852
rect 10600 14476 10652 14482
rect 10600 14418 10652 14424
rect 10704 14362 10732 15846
rect 10796 15638 10824 24822
rect 10888 24070 10916 25978
rect 10876 24064 10928 24070
rect 10876 24006 10928 24012
rect 10980 23866 11008 27934
rect 11072 25906 11100 27950
rect 11164 27334 11192 31826
rect 11348 31668 11376 32370
rect 11256 31640 11376 31668
rect 11256 31346 11284 31640
rect 11346 31580 11654 31589
rect 11346 31578 11352 31580
rect 11408 31578 11432 31580
rect 11488 31578 11512 31580
rect 11568 31578 11592 31580
rect 11648 31578 11654 31580
rect 11408 31526 11410 31578
rect 11590 31526 11592 31578
rect 11346 31524 11352 31526
rect 11408 31524 11432 31526
rect 11488 31524 11512 31526
rect 11568 31524 11592 31526
rect 11648 31524 11654 31526
rect 11346 31515 11654 31524
rect 11716 31385 11744 32846
rect 11808 32570 11836 33079
rect 11886 32736 11942 32745
rect 11886 32671 11942 32680
rect 11796 32564 11848 32570
rect 11796 32506 11848 32512
rect 11900 32337 11928 32671
rect 11886 32328 11942 32337
rect 11796 32292 11848 32298
rect 11886 32263 11942 32272
rect 11796 32234 11848 32240
rect 11702 31376 11758 31385
rect 11244 31340 11296 31346
rect 11702 31311 11758 31320
rect 11244 31282 11296 31288
rect 11346 30492 11654 30501
rect 11346 30490 11352 30492
rect 11408 30490 11432 30492
rect 11488 30490 11512 30492
rect 11568 30490 11592 30492
rect 11648 30490 11654 30492
rect 11408 30438 11410 30490
rect 11590 30438 11592 30490
rect 11346 30436 11352 30438
rect 11408 30436 11432 30438
rect 11488 30436 11512 30438
rect 11568 30436 11592 30438
rect 11648 30436 11654 30438
rect 11346 30427 11654 30436
rect 11610 30288 11666 30297
rect 11610 30223 11612 30232
rect 11664 30223 11666 30232
rect 11612 30194 11664 30200
rect 11716 30190 11744 31311
rect 11808 31113 11836 32234
rect 11888 31136 11940 31142
rect 11794 31104 11850 31113
rect 11888 31078 11940 31084
rect 11794 31039 11850 31048
rect 11900 30802 11928 31078
rect 11888 30796 11940 30802
rect 11888 30738 11940 30744
rect 11244 30184 11296 30190
rect 11244 30126 11296 30132
rect 11704 30184 11756 30190
rect 11704 30126 11756 30132
rect 11888 30184 11940 30190
rect 11888 30126 11940 30132
rect 11256 28422 11284 30126
rect 11612 30116 11664 30122
rect 11612 30058 11664 30064
rect 11334 29880 11390 29889
rect 11334 29815 11390 29824
rect 11348 29714 11376 29815
rect 11624 29782 11652 30058
rect 11612 29776 11664 29782
rect 11612 29718 11664 29724
rect 11336 29708 11388 29714
rect 11336 29650 11388 29656
rect 11794 29472 11850 29481
rect 11346 29404 11654 29413
rect 11794 29407 11850 29416
rect 11346 29402 11352 29404
rect 11408 29402 11432 29404
rect 11488 29402 11512 29404
rect 11568 29402 11592 29404
rect 11648 29402 11654 29404
rect 11408 29350 11410 29402
rect 11590 29350 11592 29402
rect 11346 29348 11352 29350
rect 11408 29348 11432 29350
rect 11488 29348 11512 29350
rect 11568 29348 11592 29350
rect 11648 29348 11654 29350
rect 11346 29339 11654 29348
rect 11702 29200 11758 29209
rect 11702 29135 11758 29144
rect 11520 28960 11572 28966
rect 11520 28902 11572 28908
rect 11532 28540 11560 28902
rect 11612 28552 11664 28558
rect 11532 28512 11612 28540
rect 11612 28494 11664 28500
rect 11244 28416 11296 28422
rect 11244 28358 11296 28364
rect 11256 27878 11284 28358
rect 11346 28316 11654 28325
rect 11346 28314 11352 28316
rect 11408 28314 11432 28316
rect 11488 28314 11512 28316
rect 11568 28314 11592 28316
rect 11648 28314 11654 28316
rect 11408 28262 11410 28314
rect 11590 28262 11592 28314
rect 11346 28260 11352 28262
rect 11408 28260 11432 28262
rect 11488 28260 11512 28262
rect 11568 28260 11592 28262
rect 11648 28260 11654 28262
rect 11346 28251 11654 28260
rect 11610 27976 11666 27985
rect 11610 27911 11666 27920
rect 11244 27872 11296 27878
rect 11244 27814 11296 27820
rect 11624 27470 11652 27911
rect 11612 27464 11664 27470
rect 11612 27406 11664 27412
rect 11152 27328 11204 27334
rect 11152 27270 11204 27276
rect 11164 27130 11192 27270
rect 11346 27228 11654 27237
rect 11346 27226 11352 27228
rect 11408 27226 11432 27228
rect 11488 27226 11512 27228
rect 11568 27226 11592 27228
rect 11648 27226 11654 27228
rect 11408 27174 11410 27226
rect 11590 27174 11592 27226
rect 11346 27172 11352 27174
rect 11408 27172 11432 27174
rect 11488 27172 11512 27174
rect 11568 27172 11592 27174
rect 11648 27172 11654 27174
rect 11346 27163 11654 27172
rect 11152 27124 11204 27130
rect 11152 27066 11204 27072
rect 11164 26246 11192 27066
rect 11152 26240 11204 26246
rect 11152 26182 11204 26188
rect 11060 25900 11112 25906
rect 11060 25842 11112 25848
rect 11164 25158 11192 26182
rect 11346 26140 11654 26149
rect 11346 26138 11352 26140
rect 11408 26138 11432 26140
rect 11488 26138 11512 26140
rect 11568 26138 11592 26140
rect 11648 26138 11654 26140
rect 11408 26086 11410 26138
rect 11590 26086 11592 26138
rect 11346 26084 11352 26086
rect 11408 26084 11432 26086
rect 11488 26084 11512 26086
rect 11568 26084 11592 26086
rect 11648 26084 11654 26086
rect 11346 26075 11654 26084
rect 11244 25900 11296 25906
rect 11244 25842 11296 25848
rect 11152 25152 11204 25158
rect 11152 25094 11204 25100
rect 11256 24818 11284 25842
rect 11346 25052 11654 25061
rect 11346 25050 11352 25052
rect 11408 25050 11432 25052
rect 11488 25050 11512 25052
rect 11568 25050 11592 25052
rect 11648 25050 11654 25052
rect 11408 24998 11410 25050
rect 11590 24998 11592 25050
rect 11346 24996 11352 24998
rect 11408 24996 11432 24998
rect 11488 24996 11512 24998
rect 11568 24996 11592 24998
rect 11648 24996 11654 24998
rect 11346 24987 11654 24996
rect 11716 24857 11744 29135
rect 11808 27146 11836 29407
rect 11900 29306 11928 30126
rect 11888 29300 11940 29306
rect 11888 29242 11940 29248
rect 11888 27872 11940 27878
rect 11888 27814 11940 27820
rect 11900 27402 11928 27814
rect 11992 27402 12020 42026
rect 12084 37670 12112 42502
rect 12072 37664 12124 37670
rect 12072 37606 12124 37612
rect 12176 37233 12204 42842
rect 12256 42764 12308 42770
rect 12256 42706 12308 42712
rect 12268 41818 12296 42706
rect 12636 42702 12664 43574
rect 12728 43364 12756 44540
rect 12912 43874 12940 44540
rect 12912 43846 13032 43874
rect 12900 43376 12952 43382
rect 12728 43336 12900 43364
rect 13004 43364 13032 43846
rect 13096 43602 13124 44540
rect 13096 43574 13216 43602
rect 13084 43376 13136 43382
rect 13004 43336 13084 43364
rect 12900 43318 12952 43324
rect 13084 43318 13136 43324
rect 13084 43172 13136 43178
rect 13084 43114 13136 43120
rect 13096 42945 13124 43114
rect 13082 42936 13138 42945
rect 13082 42871 13138 42880
rect 13188 42702 13216 43574
rect 13280 43246 13308 44540
rect 13360 43920 13412 43926
rect 13360 43862 13412 43868
rect 13372 43314 13400 43862
rect 13464 43602 13492 44540
rect 13648 43874 13676 44540
rect 13648 43846 13768 43874
rect 13464 43574 13676 43602
rect 13360 43308 13412 43314
rect 13360 43250 13412 43256
rect 13268 43240 13320 43246
rect 13268 43182 13320 43188
rect 13450 43208 13506 43217
rect 13450 43143 13452 43152
rect 13504 43143 13506 43152
rect 13544 43172 13596 43178
rect 13452 43114 13504 43120
rect 13544 43114 13596 43120
rect 13360 43104 13412 43110
rect 13360 43046 13412 43052
rect 12624 42696 12676 42702
rect 12624 42638 12676 42644
rect 13176 42696 13228 42702
rect 13176 42638 13228 42644
rect 12348 42560 12400 42566
rect 12348 42502 12400 42508
rect 12900 42560 12952 42566
rect 12900 42502 12952 42508
rect 12992 42560 13044 42566
rect 12992 42502 13044 42508
rect 12256 41812 12308 41818
rect 12256 41754 12308 41760
rect 12254 41576 12310 41585
rect 12254 41511 12310 41520
rect 12268 38826 12296 41511
rect 12256 38820 12308 38826
rect 12256 38762 12308 38768
rect 12256 37868 12308 37874
rect 12256 37810 12308 37816
rect 12268 37330 12296 37810
rect 12256 37324 12308 37330
rect 12256 37266 12308 37272
rect 12162 37224 12218 37233
rect 12162 37159 12218 37168
rect 12072 37120 12124 37126
rect 12072 37062 12124 37068
rect 12084 33674 12112 37062
rect 12268 36394 12296 37266
rect 12176 36366 12296 36394
rect 12176 36174 12204 36366
rect 12256 36304 12308 36310
rect 12256 36246 12308 36252
rect 12164 36168 12216 36174
rect 12164 36110 12216 36116
rect 12176 35494 12204 36110
rect 12164 35488 12216 35494
rect 12164 35430 12216 35436
rect 12176 34202 12204 35430
rect 12268 35222 12296 36246
rect 12256 35216 12308 35222
rect 12256 35158 12308 35164
rect 12256 34944 12308 34950
rect 12256 34886 12308 34892
rect 12164 34196 12216 34202
rect 12164 34138 12216 34144
rect 12084 33646 12204 33674
rect 12072 33584 12124 33590
rect 12072 33526 12124 33532
rect 12084 32609 12112 33526
rect 12070 32600 12126 32609
rect 12070 32535 12126 32544
rect 12176 32473 12204 33646
rect 12162 32464 12218 32473
rect 12162 32399 12218 32408
rect 12268 32314 12296 34886
rect 12176 32286 12296 32314
rect 12176 31754 12204 32286
rect 12084 31726 12204 31754
rect 11888 27396 11940 27402
rect 11888 27338 11940 27344
rect 11980 27396 12032 27402
rect 11980 27338 12032 27344
rect 11808 27118 11928 27146
rect 11796 27056 11848 27062
rect 11796 26998 11848 27004
rect 11702 24848 11758 24857
rect 11244 24812 11296 24818
rect 11702 24783 11758 24792
rect 11244 24754 11296 24760
rect 11244 24132 11296 24138
rect 11244 24074 11296 24080
rect 11152 24064 11204 24070
rect 11152 24006 11204 24012
rect 10968 23860 11020 23866
rect 10968 23802 11020 23808
rect 11164 23712 11192 24006
rect 11256 23848 11284 24074
rect 11704 24064 11756 24070
rect 11704 24006 11756 24012
rect 11346 23964 11654 23973
rect 11346 23962 11352 23964
rect 11408 23962 11432 23964
rect 11488 23962 11512 23964
rect 11568 23962 11592 23964
rect 11648 23962 11654 23964
rect 11408 23910 11410 23962
rect 11590 23910 11592 23962
rect 11346 23908 11352 23910
rect 11408 23908 11432 23910
rect 11488 23908 11512 23910
rect 11568 23908 11592 23910
rect 11648 23908 11654 23910
rect 11346 23899 11654 23908
rect 11716 23866 11744 24006
rect 11612 23860 11664 23866
rect 11256 23820 11376 23848
rect 11244 23724 11296 23730
rect 11164 23684 11244 23712
rect 11244 23666 11296 23672
rect 10968 23588 11020 23594
rect 10968 23530 11020 23536
rect 10874 23488 10930 23497
rect 10874 23423 10930 23432
rect 10888 22710 10916 23423
rect 10980 22710 11008 23530
rect 11152 23520 11204 23526
rect 11348 23508 11376 23820
rect 11612 23802 11664 23808
rect 11704 23860 11756 23866
rect 11704 23802 11756 23808
rect 11426 23624 11482 23633
rect 11624 23594 11652 23802
rect 11704 23724 11756 23730
rect 11704 23666 11756 23672
rect 11426 23559 11482 23568
rect 11612 23588 11664 23594
rect 11440 23526 11468 23559
rect 11612 23530 11664 23536
rect 11204 23480 11376 23508
rect 11428 23520 11480 23526
rect 11152 23462 11204 23468
rect 11428 23462 11480 23468
rect 11520 23316 11572 23322
rect 11520 23258 11572 23264
rect 11244 23112 11296 23118
rect 11072 23072 11244 23100
rect 10876 22704 10928 22710
rect 10968 22704 11020 22710
rect 10876 22646 10928 22652
rect 10966 22672 10968 22681
rect 11020 22672 11022 22681
rect 10966 22607 11022 22616
rect 11072 22488 11100 23072
rect 11244 23054 11296 23060
rect 11532 22982 11560 23258
rect 11520 22976 11572 22982
rect 11150 22944 11206 22953
rect 11206 22902 11284 22930
rect 11520 22918 11572 22924
rect 11150 22879 11206 22888
rect 11150 22808 11206 22817
rect 11150 22743 11206 22752
rect 11164 22574 11192 22743
rect 11256 22642 11284 22902
rect 11346 22876 11654 22885
rect 11346 22874 11352 22876
rect 11408 22874 11432 22876
rect 11488 22874 11512 22876
rect 11568 22874 11592 22876
rect 11648 22874 11654 22876
rect 11408 22822 11410 22874
rect 11590 22822 11592 22874
rect 11346 22820 11352 22822
rect 11408 22820 11432 22822
rect 11488 22820 11512 22822
rect 11568 22820 11592 22822
rect 11648 22820 11654 22822
rect 11346 22811 11654 22820
rect 11244 22636 11296 22642
rect 11244 22578 11296 22584
rect 11152 22568 11204 22574
rect 11152 22510 11204 22516
rect 10888 22460 11100 22488
rect 10888 22234 10916 22460
rect 11152 22432 11204 22438
rect 10966 22400 11022 22409
rect 11152 22374 11204 22380
rect 10966 22335 11022 22344
rect 10876 22228 10928 22234
rect 10876 22170 10928 22176
rect 10980 20913 11008 22335
rect 11164 22273 11192 22374
rect 11150 22264 11206 22273
rect 11060 22228 11112 22234
rect 11150 22199 11206 22208
rect 11060 22170 11112 22176
rect 11072 21622 11100 22170
rect 11716 22098 11744 23666
rect 11808 22710 11836 26998
rect 11900 25401 11928 27118
rect 11992 27062 12020 27338
rect 11980 27056 12032 27062
rect 11980 26998 12032 27004
rect 11992 26314 12020 26998
rect 11980 26308 12032 26314
rect 11980 26250 12032 26256
rect 11886 25392 11942 25401
rect 11886 25327 11942 25336
rect 11992 25294 12020 26250
rect 11980 25288 12032 25294
rect 11980 25230 12032 25236
rect 11888 25220 11940 25226
rect 11888 25162 11940 25168
rect 11900 24954 11928 25162
rect 11888 24948 11940 24954
rect 11888 24890 11940 24896
rect 11888 23860 11940 23866
rect 11888 23802 11940 23808
rect 11796 22704 11848 22710
rect 11796 22646 11848 22652
rect 11704 22092 11756 22098
rect 11704 22034 11756 22040
rect 11704 21888 11756 21894
rect 11704 21830 11756 21836
rect 11346 21788 11654 21797
rect 11346 21786 11352 21788
rect 11408 21786 11432 21788
rect 11488 21786 11512 21788
rect 11568 21786 11592 21788
rect 11648 21786 11654 21788
rect 11408 21734 11410 21786
rect 11590 21734 11592 21786
rect 11346 21732 11352 21734
rect 11408 21732 11432 21734
rect 11488 21732 11512 21734
rect 11568 21732 11592 21734
rect 11648 21732 11654 21734
rect 11346 21723 11654 21732
rect 11716 21672 11744 21830
rect 11624 21644 11744 21672
rect 11060 21616 11112 21622
rect 11060 21558 11112 21564
rect 10966 20904 11022 20913
rect 10966 20839 11022 20848
rect 10980 20330 11008 20839
rect 11072 20777 11100 21558
rect 11244 21548 11296 21554
rect 11244 21490 11296 21496
rect 11256 21146 11284 21490
rect 11624 21486 11652 21644
rect 11612 21480 11664 21486
rect 11426 21448 11482 21457
rect 11612 21422 11664 21428
rect 11426 21383 11482 21392
rect 11244 21140 11296 21146
rect 11244 21082 11296 21088
rect 11058 20768 11114 20777
rect 11058 20703 11114 20712
rect 11058 20632 11114 20641
rect 11114 20590 11192 20618
rect 11058 20567 11114 20576
rect 10968 20324 11020 20330
rect 10968 20266 11020 20272
rect 11060 20256 11112 20262
rect 11060 20198 11112 20204
rect 11072 19922 11100 20198
rect 11164 20058 11192 20590
rect 11256 20262 11284 21082
rect 11440 20942 11468 21383
rect 11794 21176 11850 21185
rect 11794 21111 11850 21120
rect 11428 20936 11480 20942
rect 11428 20878 11480 20884
rect 11808 20874 11836 21111
rect 11796 20868 11848 20874
rect 11796 20810 11848 20816
rect 11346 20700 11654 20709
rect 11346 20698 11352 20700
rect 11408 20698 11432 20700
rect 11488 20698 11512 20700
rect 11568 20698 11592 20700
rect 11648 20698 11654 20700
rect 11408 20646 11410 20698
rect 11590 20646 11592 20698
rect 11346 20644 11352 20646
rect 11408 20644 11432 20646
rect 11488 20644 11512 20646
rect 11568 20644 11592 20646
rect 11648 20644 11654 20646
rect 11346 20635 11654 20644
rect 11428 20460 11480 20466
rect 11428 20402 11480 20408
rect 11440 20369 11468 20402
rect 11520 20392 11572 20398
rect 11426 20360 11482 20369
rect 11336 20324 11388 20330
rect 11520 20334 11572 20340
rect 11426 20295 11482 20304
rect 11336 20266 11388 20272
rect 11244 20256 11296 20262
rect 11244 20198 11296 20204
rect 11152 20052 11204 20058
rect 11152 19994 11204 20000
rect 11256 19938 11284 20198
rect 11348 20058 11376 20266
rect 11532 20058 11560 20334
rect 11336 20052 11388 20058
rect 11336 19994 11388 20000
rect 11520 20052 11572 20058
rect 11520 19994 11572 20000
rect 11060 19916 11112 19922
rect 11060 19858 11112 19864
rect 11164 19910 11284 19938
rect 11164 19802 11192 19910
rect 10980 19774 11192 19802
rect 11242 19816 11298 19825
rect 10874 18728 10930 18737
rect 10874 18663 10930 18672
rect 10888 18358 10916 18663
rect 10876 18352 10928 18358
rect 10876 18294 10928 18300
rect 10980 17270 11008 19774
rect 11242 19751 11298 19760
rect 11704 19780 11756 19786
rect 11060 19712 11112 19718
rect 11060 19654 11112 19660
rect 11152 19712 11204 19718
rect 11152 19654 11204 19660
rect 11072 19553 11100 19654
rect 11058 19544 11114 19553
rect 11058 19479 11114 19488
rect 11072 19446 11100 19479
rect 11060 19440 11112 19446
rect 11060 19382 11112 19388
rect 11072 18834 11100 19382
rect 11060 18828 11112 18834
rect 11060 18770 11112 18776
rect 11164 18630 11192 19654
rect 11152 18624 11204 18630
rect 11152 18566 11204 18572
rect 11150 18184 11206 18193
rect 11150 18119 11206 18128
rect 11164 18086 11192 18119
rect 11060 18080 11112 18086
rect 11060 18022 11112 18028
rect 11152 18080 11204 18086
rect 11152 18022 11204 18028
rect 10968 17264 11020 17270
rect 10968 17206 11020 17212
rect 10876 17128 10928 17134
rect 10876 17070 10928 17076
rect 10888 16658 10916 17070
rect 10968 16992 11020 16998
rect 10968 16934 11020 16940
rect 10980 16833 11008 16934
rect 10966 16824 11022 16833
rect 10966 16759 11022 16768
rect 11072 16674 11100 18022
rect 11256 17649 11284 19751
rect 11704 19722 11756 19728
rect 11346 19612 11654 19621
rect 11346 19610 11352 19612
rect 11408 19610 11432 19612
rect 11488 19610 11512 19612
rect 11568 19610 11592 19612
rect 11648 19610 11654 19612
rect 11408 19558 11410 19610
rect 11590 19558 11592 19610
rect 11346 19556 11352 19558
rect 11408 19556 11432 19558
rect 11488 19556 11512 19558
rect 11568 19556 11592 19558
rect 11648 19556 11654 19558
rect 11346 19547 11654 19556
rect 11428 19508 11480 19514
rect 11428 19450 11480 19456
rect 11440 18766 11468 19450
rect 11716 19417 11744 19722
rect 11796 19712 11848 19718
rect 11796 19654 11848 19660
rect 11702 19408 11758 19417
rect 11702 19343 11758 19352
rect 11808 19242 11836 19654
rect 11900 19514 11928 23802
rect 11992 23730 12020 25230
rect 11980 23724 12032 23730
rect 11980 23666 12032 23672
rect 11980 23588 12032 23594
rect 11980 23530 12032 23536
rect 11888 19508 11940 19514
rect 11888 19450 11940 19456
rect 11888 19372 11940 19378
rect 11888 19314 11940 19320
rect 11796 19236 11848 19242
rect 11796 19178 11848 19184
rect 11612 18828 11664 18834
rect 11612 18770 11664 18776
rect 11428 18760 11480 18766
rect 11624 18737 11652 18770
rect 11428 18702 11480 18708
rect 11610 18728 11666 18737
rect 11610 18663 11666 18672
rect 11346 18524 11654 18533
rect 11346 18522 11352 18524
rect 11408 18522 11432 18524
rect 11488 18522 11512 18524
rect 11568 18522 11592 18524
rect 11648 18522 11654 18524
rect 11408 18470 11410 18522
rect 11590 18470 11592 18522
rect 11346 18468 11352 18470
rect 11408 18468 11432 18470
rect 11488 18468 11512 18470
rect 11568 18468 11592 18470
rect 11648 18468 11654 18470
rect 11346 18459 11654 18468
rect 11808 18222 11836 19178
rect 11900 18873 11928 19314
rect 11886 18864 11942 18873
rect 11886 18799 11942 18808
rect 11886 18456 11942 18465
rect 11886 18391 11942 18400
rect 11796 18216 11848 18222
rect 11796 18158 11848 18164
rect 11796 17740 11848 17746
rect 11796 17682 11848 17688
rect 11242 17640 11298 17649
rect 11242 17575 11298 17584
rect 11704 17536 11756 17542
rect 11704 17478 11756 17484
rect 11346 17436 11654 17445
rect 11346 17434 11352 17436
rect 11408 17434 11432 17436
rect 11488 17434 11512 17436
rect 11568 17434 11592 17436
rect 11648 17434 11654 17436
rect 11408 17382 11410 17434
rect 11590 17382 11592 17434
rect 11346 17380 11352 17382
rect 11408 17380 11432 17382
rect 11488 17380 11512 17382
rect 11568 17380 11592 17382
rect 11648 17380 11654 17382
rect 11150 17368 11206 17377
rect 11346 17371 11654 17380
rect 11206 17312 11376 17320
rect 11150 17303 11376 17312
rect 11164 17292 11376 17303
rect 11244 17196 11296 17202
rect 11244 17138 11296 17144
rect 11150 17096 11206 17105
rect 11150 17031 11206 17040
rect 11164 16998 11192 17031
rect 11152 16992 11204 16998
rect 11152 16934 11204 16940
rect 10876 16652 10928 16658
rect 10876 16594 10928 16600
rect 10980 16646 11100 16674
rect 10876 16040 10928 16046
rect 10980 15994 11008 16646
rect 11060 16448 11112 16454
rect 11060 16390 11112 16396
rect 11072 16289 11100 16390
rect 11058 16280 11114 16289
rect 11256 16250 11284 17138
rect 11348 16590 11376 17292
rect 11716 16658 11744 17478
rect 11704 16652 11756 16658
rect 11704 16594 11756 16600
rect 11336 16584 11388 16590
rect 11808 16538 11836 17682
rect 11900 17626 11928 18391
rect 11992 17746 12020 23530
rect 12084 22234 12112 31726
rect 12164 31680 12216 31686
rect 12164 31622 12216 31628
rect 12176 29714 12204 31622
rect 12256 31272 12308 31278
rect 12256 31214 12308 31220
rect 12268 30870 12296 31214
rect 12256 30864 12308 30870
rect 12256 30806 12308 30812
rect 12268 30569 12296 30806
rect 12254 30560 12310 30569
rect 12254 30495 12310 30504
rect 12254 29880 12310 29889
rect 12254 29815 12256 29824
rect 12308 29815 12310 29824
rect 12256 29786 12308 29792
rect 12164 29708 12216 29714
rect 12164 29650 12216 29656
rect 12176 28694 12204 29650
rect 12360 29481 12388 42502
rect 12912 42362 12940 42502
rect 12900 42356 12952 42362
rect 12900 42298 12952 42304
rect 12438 42120 12494 42129
rect 12438 42055 12494 42064
rect 12452 30841 12480 42055
rect 12532 41472 12584 41478
rect 12532 41414 12584 41420
rect 12544 36281 12572 41414
rect 12624 38752 12676 38758
rect 12624 38694 12676 38700
rect 12636 37194 12664 38694
rect 12716 38412 12768 38418
rect 12716 38354 12768 38360
rect 12624 37188 12676 37194
rect 12624 37130 12676 37136
rect 12530 36272 12586 36281
rect 12530 36207 12586 36216
rect 12532 35556 12584 35562
rect 12532 35498 12584 35504
rect 12544 35154 12572 35498
rect 12532 35148 12584 35154
rect 12532 35090 12584 35096
rect 12624 35080 12676 35086
rect 12624 35022 12676 35028
rect 12636 34610 12664 35022
rect 12624 34604 12676 34610
rect 12624 34546 12676 34552
rect 12624 33312 12676 33318
rect 12624 33254 12676 33260
rect 12636 32978 12664 33254
rect 12624 32972 12676 32978
rect 12624 32914 12676 32920
rect 12532 32904 12584 32910
rect 12530 32872 12532 32881
rect 12584 32872 12586 32881
rect 12530 32807 12586 32816
rect 12532 32768 12584 32774
rect 12532 32710 12584 32716
rect 12624 32768 12676 32774
rect 12624 32710 12676 32716
rect 12544 32570 12572 32710
rect 12532 32564 12584 32570
rect 12532 32506 12584 32512
rect 12636 31822 12664 32710
rect 12624 31816 12676 31822
rect 12624 31758 12676 31764
rect 12728 31754 12756 38354
rect 13004 36854 13032 42502
rect 13176 38548 13228 38554
rect 13176 38490 13228 38496
rect 13188 37874 13216 38490
rect 13176 37868 13228 37874
rect 13176 37810 13228 37816
rect 13082 37360 13138 37369
rect 13082 37295 13084 37304
rect 13136 37295 13138 37304
rect 13084 37266 13136 37272
rect 12992 36848 13044 36854
rect 12992 36790 13044 36796
rect 13176 36712 13228 36718
rect 13176 36654 13228 36660
rect 13084 35828 13136 35834
rect 13084 35770 13136 35776
rect 13096 35601 13124 35770
rect 13082 35592 13138 35601
rect 13082 35527 13138 35536
rect 12808 35488 12860 35494
rect 12808 35430 12860 35436
rect 12820 35154 12848 35430
rect 12808 35148 12860 35154
rect 12808 35090 12860 35096
rect 13096 34678 13124 35527
rect 13084 34672 13136 34678
rect 13084 34614 13136 34620
rect 13188 34066 13216 36654
rect 13372 36530 13400 43046
rect 13556 42702 13584 43114
rect 13648 42702 13676 43574
rect 13740 43450 13768 43846
rect 13728 43444 13780 43450
rect 13728 43386 13780 43392
rect 13832 42702 13860 44540
rect 14016 43897 14044 44540
rect 14002 43888 14058 43897
rect 14200 43874 14228 44540
rect 14200 43846 14320 43874
rect 14002 43823 14058 43832
rect 14292 43450 14320 43846
rect 13912 43444 13964 43450
rect 13912 43386 13964 43392
rect 14280 43444 14332 43450
rect 14280 43386 14332 43392
rect 13924 43353 13952 43386
rect 13910 43344 13966 43353
rect 13910 43279 13966 43288
rect 14280 43240 14332 43246
rect 14280 43182 14332 43188
rect 13945 43004 14253 43013
rect 13945 43002 13951 43004
rect 14007 43002 14031 43004
rect 14087 43002 14111 43004
rect 14167 43002 14191 43004
rect 14247 43002 14253 43004
rect 14007 42950 14009 43002
rect 14189 42950 14191 43002
rect 13945 42948 13951 42950
rect 14007 42948 14031 42950
rect 14087 42948 14111 42950
rect 14167 42948 14191 42950
rect 14247 42948 14253 42950
rect 13945 42939 14253 42948
rect 13544 42696 13596 42702
rect 13544 42638 13596 42644
rect 13636 42696 13688 42702
rect 13636 42638 13688 42644
rect 13820 42696 13872 42702
rect 13820 42638 13872 42644
rect 14096 42628 14148 42634
rect 14096 42570 14148 42576
rect 13820 42560 13872 42566
rect 13820 42502 13872 42508
rect 13728 42220 13780 42226
rect 13728 42162 13780 42168
rect 13544 42016 13596 42022
rect 13544 41958 13596 41964
rect 13556 39914 13584 41958
rect 13740 41818 13768 42162
rect 13832 42090 13860 42502
rect 14108 42226 14136 42570
rect 14096 42220 14148 42226
rect 14096 42162 14148 42168
rect 14002 42120 14058 42129
rect 13820 42084 13872 42090
rect 14002 42055 14058 42064
rect 13820 42026 13872 42032
rect 14016 42022 14044 42055
rect 14004 42016 14056 42022
rect 14004 41958 14056 41964
rect 13945 41916 14253 41925
rect 13945 41914 13951 41916
rect 14007 41914 14031 41916
rect 14087 41914 14111 41916
rect 14167 41914 14191 41916
rect 14247 41914 14253 41916
rect 14007 41862 14009 41914
rect 14189 41862 14191 41914
rect 13945 41860 13951 41862
rect 14007 41860 14031 41862
rect 14087 41860 14111 41862
rect 14167 41860 14191 41862
rect 14247 41860 14253 41862
rect 13945 41851 14253 41860
rect 13728 41812 13780 41818
rect 13728 41754 13780 41760
rect 14186 41712 14242 41721
rect 13912 41676 13964 41682
rect 14186 41647 14242 41656
rect 13912 41618 13964 41624
rect 13924 41414 13952 41618
rect 14200 41478 14228 41647
rect 14188 41472 14240 41478
rect 14188 41414 14240 41420
rect 13740 41386 13952 41414
rect 13544 39908 13596 39914
rect 13544 39850 13596 39856
rect 13544 38344 13596 38350
rect 13544 38286 13596 38292
rect 13556 37942 13584 38286
rect 13544 37936 13596 37942
rect 13544 37878 13596 37884
rect 13452 37120 13504 37126
rect 13452 37062 13504 37068
rect 13464 36718 13492 37062
rect 13452 36712 13504 36718
rect 13452 36654 13504 36660
rect 13636 36712 13688 36718
rect 13636 36654 13688 36660
rect 13372 36502 13492 36530
rect 13464 35698 13492 36502
rect 13452 35692 13504 35698
rect 13452 35634 13504 35640
rect 13176 34060 13228 34066
rect 13176 34002 13228 34008
rect 12900 33924 12952 33930
rect 12900 33866 12952 33872
rect 12808 33312 12860 33318
rect 12808 33254 12860 33260
rect 12820 32434 12848 33254
rect 12808 32428 12860 32434
rect 12808 32370 12860 32376
rect 12912 31754 12940 33866
rect 13544 33856 13596 33862
rect 13544 33798 13596 33804
rect 13084 33584 13136 33590
rect 12990 33552 13046 33561
rect 13360 33584 13412 33590
rect 13084 33526 13136 33532
rect 13280 33544 13360 33572
rect 12990 33487 13046 33496
rect 13004 33318 13032 33487
rect 12992 33312 13044 33318
rect 12992 33254 13044 33260
rect 13096 32570 13124 33526
rect 13084 32564 13136 32570
rect 13084 32506 13136 32512
rect 13096 32178 13124 32506
rect 13174 32328 13230 32337
rect 13280 32314 13308 33544
rect 13360 33526 13412 33532
rect 13360 32768 13412 32774
rect 13360 32710 13412 32716
rect 13230 32286 13308 32314
rect 13174 32263 13230 32272
rect 13096 32150 13308 32178
rect 13174 32056 13230 32065
rect 13174 31991 13230 32000
rect 12728 31726 12848 31754
rect 12912 31726 13032 31754
rect 12438 30832 12494 30841
rect 12438 30767 12494 30776
rect 12624 30728 12676 30734
rect 12624 30670 12676 30676
rect 12636 30394 12664 30670
rect 12624 30388 12676 30394
rect 12624 30330 12676 30336
rect 12440 30252 12492 30258
rect 12440 30194 12492 30200
rect 12452 29866 12480 30194
rect 12716 30184 12768 30190
rect 12716 30126 12768 30132
rect 12452 29838 12664 29866
rect 12346 29472 12402 29481
rect 12346 29407 12402 29416
rect 12348 29300 12400 29306
rect 12348 29242 12400 29248
rect 12256 29096 12308 29102
rect 12256 29038 12308 29044
rect 12164 28688 12216 28694
rect 12164 28630 12216 28636
rect 12268 28422 12296 29038
rect 12256 28416 12308 28422
rect 12256 28358 12308 28364
rect 12256 27396 12308 27402
rect 12256 27338 12308 27344
rect 12162 27296 12218 27305
rect 12162 27231 12218 27240
rect 12176 27062 12204 27231
rect 12268 27062 12296 27338
rect 12164 27056 12216 27062
rect 12164 26998 12216 27004
rect 12256 27056 12308 27062
rect 12256 26998 12308 27004
rect 12268 26314 12296 26998
rect 12256 26308 12308 26314
rect 12256 26250 12308 26256
rect 12164 26240 12216 26246
rect 12164 26182 12216 26188
rect 12176 25906 12204 26182
rect 12164 25900 12216 25906
rect 12164 25842 12216 25848
rect 12176 23322 12204 25842
rect 12268 25226 12296 26250
rect 12360 25294 12388 29242
rect 12636 29186 12664 29838
rect 12728 29714 12756 30126
rect 12716 29708 12768 29714
rect 12716 29650 12768 29656
rect 12728 29306 12756 29650
rect 12716 29300 12768 29306
rect 12716 29242 12768 29248
rect 12636 29158 12756 29186
rect 12440 28960 12492 28966
rect 12440 28902 12492 28908
rect 12348 25288 12400 25294
rect 12348 25230 12400 25236
rect 12256 25220 12308 25226
rect 12256 25162 12308 25168
rect 12164 23316 12216 23322
rect 12164 23258 12216 23264
rect 12164 23180 12216 23186
rect 12164 23122 12216 23128
rect 12072 22228 12124 22234
rect 12072 22170 12124 22176
rect 12072 21548 12124 21554
rect 12072 21490 12124 21496
rect 12084 21146 12112 21490
rect 12072 21140 12124 21146
rect 12072 21082 12124 21088
rect 12072 19848 12124 19854
rect 12072 19790 12124 19796
rect 12084 19378 12112 19790
rect 12072 19372 12124 19378
rect 12072 19314 12124 19320
rect 12072 19236 12124 19242
rect 12072 19178 12124 19184
rect 12084 18834 12112 19178
rect 12072 18828 12124 18834
rect 12072 18770 12124 18776
rect 12070 18728 12126 18737
rect 12070 18663 12126 18672
rect 12084 17882 12112 18663
rect 12072 17876 12124 17882
rect 12072 17818 12124 17824
rect 11980 17740 12032 17746
rect 11980 17682 12032 17688
rect 11900 17598 12020 17626
rect 11888 17536 11940 17542
rect 11888 17478 11940 17484
rect 11336 16526 11388 16532
rect 11348 16454 11376 16526
rect 11716 16510 11836 16538
rect 11336 16448 11388 16454
rect 11336 16390 11388 16396
rect 11346 16348 11654 16357
rect 11346 16346 11352 16348
rect 11408 16346 11432 16348
rect 11488 16346 11512 16348
rect 11568 16346 11592 16348
rect 11648 16346 11654 16348
rect 11408 16294 11410 16346
rect 11590 16294 11592 16346
rect 11346 16292 11352 16294
rect 11408 16292 11432 16294
rect 11488 16292 11512 16294
rect 11568 16292 11592 16294
rect 11648 16292 11654 16294
rect 11346 16283 11654 16292
rect 11058 16215 11114 16224
rect 11244 16244 11296 16250
rect 11244 16186 11296 16192
rect 10928 15988 11008 15994
rect 10876 15982 11008 15988
rect 10888 15966 11008 15982
rect 10784 15632 10836 15638
rect 10784 15574 10836 15580
rect 10796 14600 10824 15574
rect 11716 15366 11744 16510
rect 11900 15722 11928 17478
rect 11808 15694 11928 15722
rect 11704 15360 11756 15366
rect 11704 15302 11756 15308
rect 11346 15260 11654 15269
rect 11346 15258 11352 15260
rect 11408 15258 11432 15260
rect 11488 15258 11512 15260
rect 11568 15258 11592 15260
rect 11648 15258 11654 15260
rect 11408 15206 11410 15258
rect 11590 15206 11592 15258
rect 11346 15204 11352 15206
rect 11408 15204 11432 15206
rect 11488 15204 11512 15206
rect 11568 15204 11592 15206
rect 11648 15204 11654 15206
rect 11346 15195 11654 15204
rect 11060 14816 11112 14822
rect 11060 14758 11112 14764
rect 10968 14612 11020 14618
rect 10796 14572 10916 14600
rect 10782 14512 10838 14521
rect 10782 14447 10838 14456
rect 10796 14414 10824 14447
rect 10612 14334 10732 14362
rect 10784 14408 10836 14414
rect 10784 14350 10836 14356
rect 10612 13274 10640 14334
rect 10692 13388 10744 13394
rect 10796 13376 10824 14350
rect 10888 13938 10916 14572
rect 10968 14554 11020 14560
rect 10980 14278 11008 14554
rect 11072 14414 11100 14758
rect 11612 14612 11664 14618
rect 11612 14554 11664 14560
rect 11624 14482 11652 14554
rect 11612 14476 11664 14482
rect 11612 14418 11664 14424
rect 11060 14408 11112 14414
rect 11060 14350 11112 14356
rect 10968 14272 11020 14278
rect 10968 14214 11020 14220
rect 11704 14272 11756 14278
rect 11704 14214 11756 14220
rect 10876 13932 10928 13938
rect 10876 13874 10928 13880
rect 10980 13530 11008 14214
rect 11346 14172 11654 14181
rect 11346 14170 11352 14172
rect 11408 14170 11432 14172
rect 11488 14170 11512 14172
rect 11568 14170 11592 14172
rect 11648 14170 11654 14172
rect 11408 14118 11410 14170
rect 11590 14118 11592 14170
rect 11346 14116 11352 14118
rect 11408 14116 11432 14118
rect 11488 14116 11512 14118
rect 11568 14116 11592 14118
rect 11648 14116 11654 14118
rect 11346 14107 11654 14116
rect 11716 14074 11744 14214
rect 11060 14068 11112 14074
rect 11060 14010 11112 14016
rect 11704 14068 11756 14074
rect 11704 14010 11756 14016
rect 10968 13524 11020 13530
rect 10968 13466 11020 13472
rect 10744 13348 10824 13376
rect 10692 13330 10744 13336
rect 10612 13246 10732 13274
rect 10598 13016 10654 13025
rect 10598 12951 10654 12960
rect 10322 12744 10378 12753
rect 10322 12679 10378 12688
rect 10428 12736 10548 12764
rect 10336 12646 10364 12679
rect 10324 12640 10376 12646
rect 10324 12582 10376 12588
rect 10232 12436 10284 12442
rect 10232 12378 10284 12384
rect 10140 12300 10192 12306
rect 10140 12242 10192 12248
rect 10048 11756 10100 11762
rect 10048 11698 10100 11704
rect 10060 10674 10088 11698
rect 10048 10668 10100 10674
rect 10048 10610 10100 10616
rect 9508 10220 9720 10248
rect 9784 10560 9996 10588
rect 9508 9178 9536 10220
rect 9784 10146 9812 10560
rect 9600 10118 9812 10146
rect 9600 9364 9628 10118
rect 9680 10056 9732 10062
rect 9680 9998 9732 10004
rect 9692 9466 9720 9998
rect 10152 9738 10180 12242
rect 10244 10962 10272 12378
rect 10322 11928 10378 11937
rect 10428 11914 10456 12736
rect 10612 12306 10640 12951
rect 10508 12300 10560 12306
rect 10508 12242 10560 12248
rect 10600 12300 10652 12306
rect 10600 12242 10652 12248
rect 10378 11886 10456 11914
rect 10322 11863 10378 11872
rect 10416 11144 10468 11150
rect 10416 11086 10468 11092
rect 10244 10934 10364 10962
rect 10336 10674 10364 10934
rect 10428 10810 10456 11086
rect 10416 10804 10468 10810
rect 10416 10746 10468 10752
rect 10232 10668 10284 10674
rect 10232 10610 10284 10616
rect 10324 10668 10376 10674
rect 10324 10610 10376 10616
rect 10060 9710 10180 9738
rect 9956 9580 10008 9586
rect 9956 9522 10008 9528
rect 10060 9552 10088 9710
rect 10060 9524 10180 9552
rect 9692 9438 9812 9466
rect 9680 9376 9732 9382
rect 9600 9336 9680 9364
rect 9680 9318 9732 9324
rect 9496 9172 9548 9178
rect 9496 9114 9548 9120
rect 9692 8838 9720 9318
rect 9680 8832 9732 8838
rect 9680 8774 9732 8780
rect 9496 8492 9548 8498
rect 9496 8434 9548 8440
rect 9508 8294 9536 8434
rect 9680 8424 9732 8430
rect 9586 8392 9642 8401
rect 9680 8366 9732 8372
rect 9586 8327 9642 8336
rect 9496 8288 9548 8294
rect 9496 8230 9548 8236
rect 9494 7848 9550 7857
rect 9494 7783 9550 7792
rect 8760 3528 8812 3534
rect 8760 3470 8812 3476
rect 9404 3528 9456 3534
rect 9404 3470 9456 3476
rect 8300 3392 8352 3398
rect 8300 3334 8352 3340
rect 8576 3392 8628 3398
rect 8576 3334 8628 3340
rect 8312 3176 8340 3334
rect 8312 3148 8524 3176
rect 8300 3052 8352 3058
rect 8300 2994 8352 3000
rect 8392 3052 8444 3058
rect 8392 2994 8444 3000
rect 8206 2952 8262 2961
rect 8206 2887 8262 2896
rect 8208 2848 8260 2854
rect 8208 2790 8260 2796
rect 8220 2446 8248 2790
rect 8208 2440 8260 2446
rect 8208 2382 8260 2388
rect 8206 2272 8262 2281
rect 8206 2207 8262 2216
rect 8220 2038 8248 2207
rect 8208 2032 8260 2038
rect 8208 1974 8260 1980
rect 8206 1456 8262 1465
rect 8206 1391 8262 1400
rect 8220 1358 8248 1391
rect 8208 1352 8260 1358
rect 8208 1294 8260 1300
rect 8312 160 8340 2994
rect 8404 1442 8432 2994
rect 8496 2990 8524 3148
rect 8588 3097 8616 3334
rect 8772 3233 8800 3470
rect 9312 3460 9364 3466
rect 9312 3402 9364 3408
rect 9220 3392 9272 3398
rect 9220 3334 9272 3340
rect 9232 3233 9260 3334
rect 8758 3224 8814 3233
rect 8758 3159 8814 3168
rect 9218 3224 9274 3233
rect 9218 3159 9274 3168
rect 8574 3088 8630 3097
rect 8944 3052 8996 3058
rect 8574 3023 8630 3032
rect 8680 3012 8944 3040
rect 8484 2984 8536 2990
rect 8484 2926 8536 2932
rect 8484 2848 8536 2854
rect 8484 2790 8536 2796
rect 8576 2848 8628 2854
rect 8576 2790 8628 2796
rect 8496 2292 8524 2790
rect 8588 2446 8616 2790
rect 8576 2440 8628 2446
rect 8576 2382 8628 2388
rect 8496 2264 8616 2292
rect 8404 1414 8524 1442
rect 8392 1284 8444 1290
rect 8392 1226 8444 1232
rect 8404 950 8432 1226
rect 8392 944 8444 950
rect 8392 886 8444 892
rect 8496 160 8524 1414
rect 8588 1358 8616 2264
rect 8680 1544 8708 3012
rect 8944 2994 8996 3000
rect 9220 3052 9272 3058
rect 9220 2994 9272 3000
rect 9128 2848 9180 2854
rect 9128 2790 9180 2796
rect 8747 2748 9055 2757
rect 8747 2746 8753 2748
rect 8809 2746 8833 2748
rect 8889 2746 8913 2748
rect 8969 2746 8993 2748
rect 9049 2746 9055 2748
rect 8809 2694 8811 2746
rect 8991 2694 8993 2746
rect 8747 2692 8753 2694
rect 8809 2692 8833 2694
rect 8889 2692 8913 2694
rect 8969 2692 8993 2694
rect 9049 2692 9055 2694
rect 8747 2683 9055 2692
rect 8758 2544 8814 2553
rect 8758 2479 8814 2488
rect 8772 1766 8800 2479
rect 9140 2038 9168 2790
rect 9128 2032 9180 2038
rect 9128 1974 9180 1980
rect 8760 1760 8812 1766
rect 8760 1702 8812 1708
rect 8747 1660 9055 1669
rect 8747 1658 8753 1660
rect 8809 1658 8833 1660
rect 8889 1658 8913 1660
rect 8969 1658 8993 1660
rect 9049 1658 9055 1660
rect 8809 1606 8811 1658
rect 8991 1606 8993 1658
rect 8747 1604 8753 1606
rect 8809 1604 8833 1606
rect 8889 1604 8913 1606
rect 8969 1604 8993 1606
rect 9049 1604 9055 1606
rect 8747 1595 9055 1604
rect 9036 1556 9088 1562
rect 8680 1516 8892 1544
rect 8576 1352 8628 1358
rect 8576 1294 8628 1300
rect 8668 1284 8720 1290
rect 8668 1226 8720 1232
rect 8680 160 8708 1226
rect 8864 160 8892 1516
rect 9036 1498 9088 1504
rect 9048 1290 9076 1498
rect 9036 1284 9088 1290
rect 9036 1226 9088 1232
rect 8956 190 9076 218
rect 7930 82 7986 160
rect 7852 54 7986 82
rect 7930 -300 7986 54
rect 8114 -300 8170 160
rect 8298 -300 8354 160
rect 8482 -300 8538 160
rect 8666 -300 8722 160
rect 8850 -300 8906 160
rect 8956 105 8984 190
rect 9048 160 9076 190
rect 9232 160 9260 2994
rect 9324 1562 9352 3402
rect 9508 3346 9536 7783
rect 9416 3318 9536 3346
rect 9416 2106 9444 3318
rect 9494 3088 9550 3097
rect 9494 3023 9496 3032
rect 9548 3023 9550 3032
rect 9496 2994 9548 3000
rect 9496 2916 9548 2922
rect 9496 2858 9548 2864
rect 9404 2100 9456 2106
rect 9404 2042 9456 2048
rect 9312 1556 9364 1562
rect 9312 1498 9364 1504
rect 9402 1456 9458 1465
rect 9324 1414 9402 1442
rect 9324 762 9352 1414
rect 9402 1391 9458 1400
rect 9404 1352 9456 1358
rect 9508 1340 9536 2858
rect 9600 2446 9628 8327
rect 9692 7342 9720 8366
rect 9680 7336 9732 7342
rect 9680 7278 9732 7284
rect 9784 6390 9812 9438
rect 9864 9376 9916 9382
rect 9864 9318 9916 9324
rect 9772 6384 9824 6390
rect 9772 6326 9824 6332
rect 9680 6112 9732 6118
rect 9680 6054 9732 6060
rect 9770 6080 9826 6089
rect 9692 3942 9720 6054
rect 9770 6015 9826 6024
rect 9784 5710 9812 6015
rect 9876 5914 9904 9318
rect 9968 9160 9996 9522
rect 10048 9172 10100 9178
rect 9968 9132 10048 9160
rect 10048 9114 10100 9120
rect 10046 9072 10102 9081
rect 10046 9007 10102 9016
rect 10060 8673 10088 9007
rect 10046 8664 10102 8673
rect 9956 8628 10008 8634
rect 10046 8599 10102 8608
rect 9956 8570 10008 8576
rect 9968 6798 9996 8570
rect 10060 7750 10088 8599
rect 10152 8430 10180 9524
rect 10140 8424 10192 8430
rect 10140 8366 10192 8372
rect 10048 7744 10100 7750
rect 10048 7686 10100 7692
rect 10244 7528 10272 10610
rect 10324 10464 10376 10470
rect 10324 10406 10376 10412
rect 10336 9382 10364 10406
rect 10520 10266 10548 12242
rect 10508 10260 10560 10266
rect 10508 10202 10560 10208
rect 10416 10124 10468 10130
rect 10416 10066 10468 10072
rect 10324 9376 10376 9382
rect 10324 9318 10376 9324
rect 10324 8900 10376 8906
rect 10324 8842 10376 8848
rect 10336 8634 10364 8842
rect 10428 8838 10456 10066
rect 10506 9752 10562 9761
rect 10506 9687 10508 9696
rect 10560 9687 10562 9696
rect 10508 9658 10560 9664
rect 10612 9586 10640 12242
rect 10704 10062 10732 13246
rect 10796 11354 10824 13348
rect 10876 13388 10928 13394
rect 10876 13330 10928 13336
rect 10784 11348 10836 11354
rect 10784 11290 10836 11296
rect 10888 11286 10916 13330
rect 10968 13320 11020 13326
rect 10968 13262 11020 13268
rect 10980 12782 11008 13262
rect 10968 12776 11020 12782
rect 10968 12718 11020 12724
rect 10968 12232 11020 12238
rect 11072 12209 11100 14010
rect 11152 13864 11204 13870
rect 11152 13806 11204 13812
rect 11164 13138 11192 13806
rect 11336 13728 11388 13734
rect 11336 13670 11388 13676
rect 11348 13394 11376 13670
rect 11336 13388 11388 13394
rect 11336 13330 11388 13336
rect 11704 13252 11756 13258
rect 11704 13194 11756 13200
rect 11164 13110 11284 13138
rect 11150 13016 11206 13025
rect 11150 12951 11206 12960
rect 11164 12918 11192 12951
rect 11152 12912 11204 12918
rect 11152 12854 11204 12860
rect 11152 12776 11204 12782
rect 11152 12718 11204 12724
rect 10968 12174 11020 12180
rect 11058 12200 11114 12209
rect 10980 12084 11008 12174
rect 11058 12135 11114 12144
rect 11164 12084 11192 12718
rect 10980 12056 11192 12084
rect 10876 11280 10928 11286
rect 10876 11222 10928 11228
rect 11256 11150 11284 13110
rect 11346 13084 11654 13093
rect 11346 13082 11352 13084
rect 11408 13082 11432 13084
rect 11488 13082 11512 13084
rect 11568 13082 11592 13084
rect 11648 13082 11654 13084
rect 11408 13030 11410 13082
rect 11590 13030 11592 13082
rect 11346 13028 11352 13030
rect 11408 13028 11432 13030
rect 11488 13028 11512 13030
rect 11568 13028 11592 13030
rect 11648 13028 11654 13030
rect 11346 13019 11654 13028
rect 11716 12782 11744 13194
rect 11704 12776 11756 12782
rect 11704 12718 11756 12724
rect 11704 12096 11756 12102
rect 11704 12038 11756 12044
rect 11346 11996 11654 12005
rect 11346 11994 11352 11996
rect 11408 11994 11432 11996
rect 11488 11994 11512 11996
rect 11568 11994 11592 11996
rect 11648 11994 11654 11996
rect 11408 11942 11410 11994
rect 11590 11942 11592 11994
rect 11346 11940 11352 11942
rect 11408 11940 11432 11942
rect 11488 11940 11512 11942
rect 11568 11940 11592 11942
rect 11648 11940 11654 11942
rect 11346 11931 11654 11940
rect 11612 11688 11664 11694
rect 11612 11630 11664 11636
rect 11334 11248 11390 11257
rect 11334 11183 11336 11192
rect 11388 11183 11390 11192
rect 11336 11154 11388 11160
rect 11244 11144 11296 11150
rect 11164 11104 11244 11132
rect 11060 11076 11112 11082
rect 11060 11018 11112 11024
rect 10968 11008 11020 11014
rect 10966 10976 10968 10985
rect 11020 10976 11022 10985
rect 10966 10911 11022 10920
rect 10874 10840 10930 10849
rect 10874 10775 10930 10784
rect 10782 10568 10838 10577
rect 10782 10503 10838 10512
rect 10692 10056 10744 10062
rect 10692 9998 10744 10004
rect 10600 9580 10652 9586
rect 10600 9522 10652 9528
rect 10416 8832 10468 8838
rect 10416 8774 10468 8780
rect 10324 8628 10376 8634
rect 10324 8570 10376 8576
rect 10324 8492 10376 8498
rect 10428 8480 10456 8774
rect 10612 8548 10640 9522
rect 10692 9376 10744 9382
rect 10692 9318 10744 9324
rect 10566 8520 10640 8548
rect 10566 8514 10594 8520
rect 10376 8452 10456 8480
rect 10324 8434 10376 8440
rect 10244 7500 10364 7528
rect 10230 7440 10286 7449
rect 10230 7375 10286 7384
rect 10048 7336 10100 7342
rect 10048 7278 10100 7284
rect 9956 6792 10008 6798
rect 9956 6734 10008 6740
rect 10060 6254 10088 7278
rect 10140 7268 10192 7274
rect 10140 7210 10192 7216
rect 10152 6458 10180 7210
rect 10140 6452 10192 6458
rect 10140 6394 10192 6400
rect 10048 6248 10100 6254
rect 10048 6190 10100 6196
rect 9864 5908 9916 5914
rect 9864 5850 9916 5856
rect 9772 5704 9824 5710
rect 9772 5646 9824 5652
rect 10048 5296 10100 5302
rect 10048 5238 10100 5244
rect 9680 3936 9732 3942
rect 9680 3878 9732 3884
rect 9772 3596 9824 3602
rect 9772 3538 9824 3544
rect 9784 3194 9812 3538
rect 9864 3392 9916 3398
rect 9864 3334 9916 3340
rect 9772 3188 9824 3194
rect 9772 3130 9824 3136
rect 9680 2848 9732 2854
rect 9680 2790 9732 2796
rect 9588 2440 9640 2446
rect 9588 2382 9640 2388
rect 9692 2038 9720 2790
rect 9772 2372 9824 2378
rect 9772 2314 9824 2320
rect 9680 2032 9732 2038
rect 9784 2009 9812 2314
rect 9680 1974 9732 1980
rect 9770 2000 9826 2009
rect 9770 1935 9826 1944
rect 9588 1760 9640 1766
rect 9588 1702 9640 1708
rect 9456 1312 9536 1340
rect 9404 1294 9456 1300
rect 9404 1216 9456 1222
rect 9404 1158 9456 1164
rect 9416 950 9444 1158
rect 9404 944 9456 950
rect 9404 886 9456 892
rect 9324 734 9444 762
rect 9416 160 9444 734
rect 9600 160 9628 1702
rect 9876 1442 9904 3334
rect 9956 2304 10008 2310
rect 9956 2246 10008 2252
rect 9968 2106 9996 2246
rect 9956 2100 10008 2106
rect 9956 2042 10008 2048
rect 10060 1834 10088 5238
rect 10244 3058 10272 7375
rect 10336 5030 10364 7500
rect 10428 7410 10456 8452
rect 10520 8486 10594 8514
rect 10520 8430 10548 8486
rect 10508 8424 10560 8430
rect 10508 8366 10560 8372
rect 10600 8424 10652 8430
rect 10600 8366 10652 8372
rect 10520 7546 10548 8366
rect 10612 8090 10640 8366
rect 10600 8084 10652 8090
rect 10600 8026 10652 8032
rect 10508 7540 10560 7546
rect 10508 7482 10560 7488
rect 10520 7410 10548 7482
rect 10704 7426 10732 9318
rect 10796 8974 10824 10503
rect 10784 8968 10836 8974
rect 10784 8910 10836 8916
rect 10796 8265 10824 8910
rect 10888 8548 10916 10775
rect 10980 10305 11008 10911
rect 10966 10296 11022 10305
rect 10966 10231 11022 10240
rect 10888 8520 10962 8548
rect 10934 8294 10962 8520
rect 10888 8266 10962 8294
rect 10782 8256 10838 8265
rect 10782 8191 10838 8200
rect 10796 7818 10824 8191
rect 10784 7812 10836 7818
rect 10784 7754 10836 7760
rect 10416 7404 10468 7410
rect 10416 7346 10468 7352
rect 10508 7404 10560 7410
rect 10508 7346 10560 7352
rect 10612 7398 10732 7426
rect 10428 7002 10456 7346
rect 10416 6996 10468 7002
rect 10416 6938 10468 6944
rect 10416 5568 10468 5574
rect 10416 5510 10468 5516
rect 10324 5024 10376 5030
rect 10324 4966 10376 4972
rect 10428 3194 10456 5510
rect 10612 4570 10640 7398
rect 10692 7336 10744 7342
rect 10692 7278 10744 7284
rect 10704 7002 10732 7278
rect 10692 6996 10744 7002
rect 10692 6938 10744 6944
rect 10784 6792 10836 6798
rect 10784 6734 10836 6740
rect 10796 6225 10824 6734
rect 10782 6216 10838 6225
rect 10782 6151 10838 6160
rect 10692 5568 10744 5574
rect 10692 5510 10744 5516
rect 10520 4542 10640 4570
rect 10520 3505 10548 4542
rect 10600 4480 10652 4486
rect 10600 4422 10652 4428
rect 10506 3496 10562 3505
rect 10506 3431 10562 3440
rect 10416 3188 10468 3194
rect 10416 3130 10468 3136
rect 10232 3052 10284 3058
rect 10232 2994 10284 3000
rect 10324 2916 10376 2922
rect 10324 2858 10376 2864
rect 10232 2304 10284 2310
rect 10232 2246 10284 2252
rect 10138 2000 10194 2009
rect 10138 1935 10194 1944
rect 10152 1902 10180 1935
rect 10140 1896 10192 1902
rect 10140 1838 10192 1844
rect 10048 1828 10100 1834
rect 10048 1770 10100 1776
rect 10244 1766 10272 2246
rect 10140 1760 10192 1766
rect 10140 1702 10192 1708
rect 10232 1760 10284 1766
rect 10232 1702 10284 1708
rect 9784 1414 9904 1442
rect 10048 1420 10100 1426
rect 9784 1222 9812 1414
rect 10048 1362 10100 1368
rect 9864 1352 9916 1358
rect 9862 1320 9864 1329
rect 9916 1320 9918 1329
rect 9862 1255 9918 1264
rect 9772 1216 9824 1222
rect 9772 1158 9824 1164
rect 9864 1216 9916 1222
rect 9864 1158 9916 1164
rect 9876 1018 9904 1158
rect 9864 1012 9916 1018
rect 9864 954 9916 960
rect 9956 672 10008 678
rect 9956 614 10008 620
rect 9968 490 9996 614
rect 9876 462 9996 490
rect 8942 96 8998 105
rect 8942 31 8998 40
rect 9034 -300 9090 160
rect 9218 -300 9274 160
rect 9402 -300 9458 160
rect 9586 -300 9642 160
rect 9770 82 9826 160
rect 9876 82 9904 462
rect 9770 54 9904 82
rect 9954 82 10010 160
rect 10060 82 10088 1362
rect 10152 160 10180 1702
rect 10336 160 10364 2858
rect 10508 2848 10560 2854
rect 10428 2808 10508 2836
rect 10428 2038 10456 2808
rect 10508 2790 10560 2796
rect 10612 2446 10640 4422
rect 10704 2650 10732 5510
rect 10784 3052 10836 3058
rect 10888 3040 10916 8266
rect 10968 7744 11020 7750
rect 10968 7686 11020 7692
rect 10980 7041 11008 7686
rect 10966 7032 11022 7041
rect 10966 6967 11022 6976
rect 10968 6860 11020 6866
rect 10968 6802 11020 6808
rect 10980 6662 11008 6802
rect 10968 6656 11020 6662
rect 10968 6598 11020 6604
rect 11072 6458 11100 11018
rect 11164 8294 11192 11104
rect 11244 11086 11296 11092
rect 11624 10996 11652 11630
rect 11716 11064 11744 12038
rect 11808 11642 11836 15694
rect 11888 15496 11940 15502
rect 11888 15438 11940 15444
rect 11900 14414 11928 15438
rect 11888 14408 11940 14414
rect 11888 14350 11940 14356
rect 11900 11762 11928 14350
rect 11992 14006 12020 17598
rect 12072 17536 12124 17542
rect 12072 17478 12124 17484
rect 12084 16114 12112 17478
rect 12176 16794 12204 23122
rect 12268 22030 12296 25162
rect 12348 25152 12400 25158
rect 12348 25094 12400 25100
rect 12360 23186 12388 25094
rect 12452 24886 12480 28902
rect 12532 28688 12584 28694
rect 12532 28630 12584 28636
rect 12544 26586 12572 28630
rect 12624 28416 12676 28422
rect 12624 28358 12676 28364
rect 12636 27305 12664 28358
rect 12728 27334 12756 29158
rect 12820 28121 12848 31726
rect 12898 31648 12954 31657
rect 12898 31583 12954 31592
rect 12912 30818 12940 31583
rect 13004 31498 13032 31726
rect 13082 31512 13138 31521
rect 13004 31470 13082 31498
rect 13082 31447 13138 31456
rect 13084 31340 13136 31346
rect 13084 31282 13136 31288
rect 12992 31136 13044 31142
rect 12992 31078 13044 31084
rect 13004 30938 13032 31078
rect 13096 30938 13124 31282
rect 12992 30932 13044 30938
rect 12992 30874 13044 30880
rect 13084 30932 13136 30938
rect 13084 30874 13136 30880
rect 12912 30790 13032 30818
rect 12900 30728 12952 30734
rect 12900 30670 12952 30676
rect 12912 29850 12940 30670
rect 12900 29844 12952 29850
rect 12900 29786 12952 29792
rect 12900 29708 12952 29714
rect 12900 29650 12952 29656
rect 12806 28112 12862 28121
rect 12806 28047 12862 28056
rect 12716 27328 12768 27334
rect 12622 27296 12678 27305
rect 12716 27270 12768 27276
rect 12622 27231 12678 27240
rect 12624 27056 12676 27062
rect 12624 26998 12676 27004
rect 12532 26580 12584 26586
rect 12532 26522 12584 26528
rect 12636 26314 12664 26998
rect 12728 26450 12756 27270
rect 12912 26772 12940 29650
rect 13004 27470 13032 30790
rect 13084 30184 13136 30190
rect 13084 30126 13136 30132
rect 13096 27470 13124 30126
rect 12992 27464 13044 27470
rect 12992 27406 13044 27412
rect 13084 27464 13136 27470
rect 13084 27406 13136 27412
rect 13004 27062 13032 27406
rect 12992 27056 13044 27062
rect 12992 26998 13044 27004
rect 12992 26784 13044 26790
rect 12912 26752 12992 26772
rect 13044 26752 13046 26761
rect 12912 26744 12990 26752
rect 12990 26687 13046 26696
rect 12716 26444 12768 26450
rect 12716 26386 12768 26392
rect 12624 26308 12676 26314
rect 12624 26250 12676 26256
rect 12532 25696 12584 25702
rect 12532 25638 12584 25644
rect 12544 25362 12572 25638
rect 12532 25356 12584 25362
rect 12532 25298 12584 25304
rect 12636 25158 12664 26250
rect 12624 25152 12676 25158
rect 12624 25094 12676 25100
rect 12440 24880 12492 24886
rect 12440 24822 12492 24828
rect 12530 24848 12586 24857
rect 12530 24783 12532 24792
rect 12584 24783 12586 24792
rect 12532 24754 12584 24760
rect 12440 24404 12492 24410
rect 12440 24346 12492 24352
rect 12348 23180 12400 23186
rect 12348 23122 12400 23128
rect 12348 22704 12400 22710
rect 12348 22646 12400 22652
rect 12256 22024 12308 22030
rect 12256 21966 12308 21972
rect 12164 16788 12216 16794
rect 12164 16730 12216 16736
rect 12164 16448 12216 16454
rect 12164 16390 12216 16396
rect 12072 16108 12124 16114
rect 12072 16050 12124 16056
rect 12072 15360 12124 15366
rect 12072 15302 12124 15308
rect 12084 14074 12112 15302
rect 12072 14068 12124 14074
rect 12072 14010 12124 14016
rect 11980 14000 12032 14006
rect 11980 13942 12032 13948
rect 11992 13530 12020 13942
rect 11980 13524 12032 13530
rect 11980 13466 12032 13472
rect 11992 12753 12020 13466
rect 11978 12744 12034 12753
rect 11978 12679 12034 12688
rect 11992 12170 12020 12679
rect 11980 12164 12032 12170
rect 11980 12106 12032 12112
rect 11888 11756 11940 11762
rect 11888 11698 11940 11704
rect 11808 11614 12020 11642
rect 11796 11280 11848 11286
rect 11848 11240 11928 11268
rect 11796 11222 11848 11228
rect 11716 11036 11836 11064
rect 11624 10968 11744 10996
rect 11346 10908 11654 10917
rect 11346 10906 11352 10908
rect 11408 10906 11432 10908
rect 11488 10906 11512 10908
rect 11568 10906 11592 10908
rect 11648 10906 11654 10908
rect 11408 10854 11410 10906
rect 11590 10854 11592 10906
rect 11346 10852 11352 10854
rect 11408 10852 11432 10854
rect 11488 10852 11512 10854
rect 11568 10852 11592 10854
rect 11648 10852 11654 10854
rect 11346 10843 11654 10852
rect 11242 10432 11298 10441
rect 11242 10367 11298 10376
rect 11152 8288 11204 8294
rect 11152 8230 11204 8236
rect 11256 8106 11284 10367
rect 11716 10062 11744 10968
rect 11808 10713 11836 11036
rect 11900 10810 11928 11240
rect 11888 10804 11940 10810
rect 11888 10746 11940 10752
rect 11794 10704 11850 10713
rect 11794 10639 11850 10648
rect 11888 10600 11940 10606
rect 11888 10542 11940 10548
rect 11900 10130 11928 10542
rect 11888 10124 11940 10130
rect 11888 10066 11940 10072
rect 11704 10056 11756 10062
rect 11704 9998 11756 10004
rect 11796 9988 11848 9994
rect 11796 9930 11848 9936
rect 11346 9820 11654 9829
rect 11346 9818 11352 9820
rect 11408 9818 11432 9820
rect 11488 9818 11512 9820
rect 11568 9818 11592 9820
rect 11648 9818 11654 9820
rect 11408 9766 11410 9818
rect 11590 9766 11592 9818
rect 11346 9764 11352 9766
rect 11408 9764 11432 9766
rect 11488 9764 11512 9766
rect 11568 9764 11592 9766
rect 11648 9764 11654 9766
rect 11346 9755 11654 9764
rect 11704 9580 11756 9586
rect 11704 9522 11756 9528
rect 11336 9376 11388 9382
rect 11336 9318 11388 9324
rect 11348 8838 11376 9318
rect 11336 8832 11388 8838
rect 11336 8774 11388 8780
rect 11346 8732 11654 8741
rect 11346 8730 11352 8732
rect 11408 8730 11432 8732
rect 11488 8730 11512 8732
rect 11568 8730 11592 8732
rect 11648 8730 11654 8732
rect 11408 8678 11410 8730
rect 11590 8678 11592 8730
rect 11346 8676 11352 8678
rect 11408 8676 11432 8678
rect 11488 8676 11512 8678
rect 11568 8676 11592 8678
rect 11648 8676 11654 8678
rect 11346 8667 11654 8676
rect 11716 8634 11744 9522
rect 11808 9489 11836 9930
rect 11992 9625 12020 11614
rect 12070 11384 12126 11393
rect 12070 11319 12072 11328
rect 12124 11319 12126 11328
rect 12072 11290 12124 11296
rect 12072 11212 12124 11218
rect 12072 11154 12124 11160
rect 12084 11014 12112 11154
rect 12072 11008 12124 11014
rect 12072 10950 12124 10956
rect 12072 10192 12124 10198
rect 12072 10134 12124 10140
rect 11978 9616 12034 9625
rect 11978 9551 12034 9560
rect 11888 9512 11940 9518
rect 11794 9480 11850 9489
rect 11888 9454 11940 9460
rect 11794 9415 11850 9424
rect 11808 9042 11836 9415
rect 11900 9353 11928 9454
rect 11886 9344 11942 9353
rect 11886 9279 11942 9288
rect 11796 9036 11848 9042
rect 11796 8978 11848 8984
rect 11704 8628 11756 8634
rect 11704 8570 11756 8576
rect 11704 8492 11756 8498
rect 11808 8480 11836 8978
rect 11756 8452 11836 8480
rect 11888 8492 11940 8498
rect 11704 8434 11756 8440
rect 11992 8480 12020 9551
rect 12084 9450 12112 10134
rect 12072 9444 12124 9450
rect 12072 9386 12124 9392
rect 12090 8492 12142 8498
rect 11940 8452 12020 8480
rect 11888 8434 11940 8440
rect 12084 8440 12090 8480
rect 12084 8434 12142 8440
rect 11612 8288 11664 8294
rect 11612 8230 11664 8236
rect 11796 8288 11848 8294
rect 11796 8230 11848 8236
rect 11164 8078 11284 8106
rect 11060 6452 11112 6458
rect 11060 6394 11112 6400
rect 10968 6112 11020 6118
rect 10968 6054 11020 6060
rect 10980 5681 11008 6054
rect 10966 5672 11022 5681
rect 10966 5607 11022 5616
rect 11164 5166 11192 8078
rect 11624 7834 11652 8230
rect 11808 8106 11836 8230
rect 11716 8078 11836 8106
rect 11716 8022 11744 8078
rect 12084 8072 12112 8434
rect 11992 8044 12112 8072
rect 12176 8072 12204 16390
rect 12268 11937 12296 21966
rect 12360 13841 12388 22646
rect 12452 22273 12480 24346
rect 12544 23100 12572 24754
rect 12636 24721 12664 25094
rect 12622 24712 12678 24721
rect 12622 24647 12678 24656
rect 12728 23798 12756 26386
rect 12992 26308 13044 26314
rect 12992 26250 13044 26256
rect 12898 25936 12954 25945
rect 12898 25871 12954 25880
rect 12912 25838 12940 25871
rect 12900 25832 12952 25838
rect 12900 25774 12952 25780
rect 12808 25764 12860 25770
rect 12808 25706 12860 25712
rect 12820 25498 12848 25706
rect 12808 25492 12860 25498
rect 12808 25434 12860 25440
rect 12808 25288 12860 25294
rect 13004 25276 13032 26250
rect 12860 25248 13032 25276
rect 12808 25230 12860 25236
rect 12820 23866 12848 25230
rect 12992 24812 13044 24818
rect 12992 24754 13044 24760
rect 12808 23860 12860 23866
rect 12808 23802 12860 23808
rect 12716 23792 12768 23798
rect 12716 23734 12768 23740
rect 12900 23792 12952 23798
rect 12900 23734 12952 23740
rect 12624 23724 12676 23730
rect 12624 23666 12676 23672
rect 12636 23361 12664 23666
rect 12912 23662 12940 23734
rect 12900 23656 12952 23662
rect 12900 23598 12952 23604
rect 12716 23588 12768 23594
rect 12716 23530 12768 23536
rect 12622 23352 12678 23361
rect 12622 23287 12678 23296
rect 12624 23112 12676 23118
rect 12544 23072 12624 23100
rect 12438 22264 12494 22273
rect 12438 22199 12494 22208
rect 12544 22148 12572 23072
rect 12624 23054 12676 23060
rect 12624 22976 12676 22982
rect 12624 22918 12676 22924
rect 12636 22166 12664 22918
rect 12452 22120 12572 22148
rect 12624 22160 12676 22166
rect 12452 20369 12480 22120
rect 12624 22102 12676 22108
rect 12622 21992 12678 22001
rect 12544 21950 12622 21978
rect 12438 20360 12494 20369
rect 12438 20295 12494 20304
rect 12440 19712 12492 19718
rect 12440 19654 12492 19660
rect 12452 19514 12480 19654
rect 12440 19508 12492 19514
rect 12440 19450 12492 19456
rect 12440 19168 12492 19174
rect 12440 19110 12492 19116
rect 12452 18834 12480 19110
rect 12440 18828 12492 18834
rect 12440 18770 12492 18776
rect 12544 18408 12572 21950
rect 12622 21927 12678 21936
rect 12728 21690 12756 23530
rect 12808 23112 12860 23118
rect 12912 23089 12940 23598
rect 12808 23054 12860 23060
rect 12898 23080 12954 23089
rect 12820 22778 12848 23054
rect 12898 23015 12954 23024
rect 12808 22772 12860 22778
rect 12808 22714 12860 22720
rect 12808 22636 12860 22642
rect 12808 22578 12860 22584
rect 12624 21684 12676 21690
rect 12624 21626 12676 21632
rect 12716 21684 12768 21690
rect 12716 21626 12768 21632
rect 12820 21672 12848 22578
rect 12900 21684 12952 21690
rect 12820 21644 12900 21672
rect 12636 21146 12664 21626
rect 12624 21140 12676 21146
rect 12624 21082 12676 21088
rect 12624 20936 12676 20942
rect 12624 20878 12676 20884
rect 12636 20505 12664 20878
rect 12622 20496 12678 20505
rect 12622 20431 12678 20440
rect 12624 20256 12676 20262
rect 12624 20198 12676 20204
rect 12636 18970 12664 20198
rect 12728 19718 12756 21626
rect 12820 20466 12848 21644
rect 12900 21626 12952 21632
rect 13004 21434 13032 24754
rect 13188 24698 13216 31991
rect 13280 30938 13308 32150
rect 13372 31890 13400 32710
rect 13452 32564 13504 32570
rect 13452 32506 13504 32512
rect 13360 31884 13412 31890
rect 13360 31826 13412 31832
rect 13360 31748 13412 31754
rect 13360 31690 13412 31696
rect 13268 30932 13320 30938
rect 13268 30874 13320 30880
rect 13280 30569 13308 30874
rect 13266 30560 13322 30569
rect 13266 30495 13322 30504
rect 13266 30288 13322 30297
rect 13266 30223 13322 30232
rect 13280 29646 13308 30223
rect 13372 30054 13400 31690
rect 13464 30802 13492 32506
rect 13556 32366 13584 33798
rect 13648 33572 13676 36654
rect 13740 34513 13768 41386
rect 14292 41206 14320 43182
rect 14384 41614 14412 44540
rect 14464 42560 14516 42566
rect 14464 42502 14516 42508
rect 14476 42362 14504 42502
rect 14464 42356 14516 42362
rect 14464 42298 14516 42304
rect 14464 42016 14516 42022
rect 14464 41958 14516 41964
rect 14372 41608 14424 41614
rect 14372 41550 14424 41556
rect 14280 41200 14332 41206
rect 14280 41142 14332 41148
rect 13945 40828 14253 40837
rect 13945 40826 13951 40828
rect 14007 40826 14031 40828
rect 14087 40826 14111 40828
rect 14167 40826 14191 40828
rect 14247 40826 14253 40828
rect 14007 40774 14009 40826
rect 14189 40774 14191 40826
rect 13945 40772 13951 40774
rect 14007 40772 14031 40774
rect 14087 40772 14111 40774
rect 14167 40772 14191 40774
rect 14247 40772 14253 40774
rect 13945 40763 14253 40772
rect 13945 39740 14253 39749
rect 13945 39738 13951 39740
rect 14007 39738 14031 39740
rect 14087 39738 14111 39740
rect 14167 39738 14191 39740
rect 14247 39738 14253 39740
rect 14007 39686 14009 39738
rect 14189 39686 14191 39738
rect 13945 39684 13951 39686
rect 14007 39684 14031 39686
rect 14087 39684 14111 39686
rect 14167 39684 14191 39686
rect 14247 39684 14253 39686
rect 13945 39675 14253 39684
rect 14476 39545 14504 41958
rect 14568 41138 14596 44540
rect 14752 43466 14780 44540
rect 14660 43438 14780 43466
rect 14660 43246 14688 43438
rect 14740 43308 14792 43314
rect 14740 43250 14792 43256
rect 14648 43240 14700 43246
rect 14648 43182 14700 43188
rect 14648 43104 14700 43110
rect 14648 43046 14700 43052
rect 14660 42906 14688 43046
rect 14648 42900 14700 42906
rect 14648 42842 14700 42848
rect 14752 42650 14780 43250
rect 14832 43104 14884 43110
rect 14832 43046 14884 43052
rect 14660 42622 14780 42650
rect 14660 41274 14688 42622
rect 14740 42560 14792 42566
rect 14740 42502 14792 42508
rect 14752 42362 14780 42502
rect 14740 42356 14792 42362
rect 14740 42298 14792 42304
rect 14844 42294 14872 43046
rect 14832 42288 14884 42294
rect 14738 42256 14794 42265
rect 14832 42230 14884 42236
rect 14738 42191 14794 42200
rect 14648 41268 14700 41274
rect 14648 41210 14700 41216
rect 14646 41168 14702 41177
rect 14556 41132 14608 41138
rect 14646 41103 14702 41112
rect 14556 41074 14608 41080
rect 14660 40882 14688 41103
rect 14752 41070 14780 42191
rect 14936 42106 14964 44540
rect 15014 42936 15070 42945
rect 15120 42922 15148 44540
rect 15304 44010 15332 44540
rect 15212 43982 15332 44010
rect 15212 43926 15240 43982
rect 15200 43920 15252 43926
rect 15200 43862 15252 43868
rect 15292 43308 15344 43314
rect 15070 42894 15148 42922
rect 15212 43268 15292 43296
rect 15014 42871 15070 42880
rect 15212 42786 15240 43268
rect 15292 43250 15344 43256
rect 15292 43104 15344 43110
rect 15292 43046 15344 43052
rect 15384 43104 15436 43110
rect 15384 43046 15436 43052
rect 14844 42078 14964 42106
rect 15028 42758 15240 42786
rect 14844 41478 14872 42078
rect 14924 42016 14976 42022
rect 14924 41958 14976 41964
rect 14832 41472 14884 41478
rect 14832 41414 14884 41420
rect 14740 41064 14792 41070
rect 14740 41006 14792 41012
rect 14660 40854 14780 40882
rect 14462 39536 14518 39545
rect 14462 39471 14518 39480
rect 14462 39400 14518 39409
rect 14462 39335 14518 39344
rect 13945 38652 14253 38661
rect 13945 38650 13951 38652
rect 14007 38650 14031 38652
rect 14087 38650 14111 38652
rect 14167 38650 14191 38652
rect 14247 38650 14253 38652
rect 14007 38598 14009 38650
rect 14189 38598 14191 38650
rect 13945 38596 13951 38598
rect 14007 38596 14031 38598
rect 14087 38596 14111 38598
rect 14167 38596 14191 38598
rect 14247 38596 14253 38598
rect 13945 38587 14253 38596
rect 14188 37936 14240 37942
rect 14186 37904 14188 37913
rect 14240 37904 14242 37913
rect 14186 37839 14242 37848
rect 14280 37664 14332 37670
rect 14280 37606 14332 37612
rect 13945 37564 14253 37573
rect 13945 37562 13951 37564
rect 14007 37562 14031 37564
rect 14087 37562 14111 37564
rect 14167 37562 14191 37564
rect 14247 37562 14253 37564
rect 14007 37510 14009 37562
rect 14189 37510 14191 37562
rect 13945 37508 13951 37510
rect 14007 37508 14031 37510
rect 14087 37508 14111 37510
rect 14167 37508 14191 37510
rect 14247 37508 14253 37510
rect 13945 37499 14253 37508
rect 14004 37460 14056 37466
rect 14004 37402 14056 37408
rect 14016 37126 14044 37402
rect 13912 37120 13964 37126
rect 13912 37062 13964 37068
rect 14004 37120 14056 37126
rect 14004 37062 14056 37068
rect 13820 36712 13872 36718
rect 13924 36689 13952 37062
rect 14016 36786 14044 37062
rect 14004 36780 14056 36786
rect 14004 36722 14056 36728
rect 14292 36718 14320 37606
rect 14372 37120 14424 37126
rect 14372 37062 14424 37068
rect 14280 36712 14332 36718
rect 13820 36654 13872 36660
rect 13910 36680 13966 36689
rect 13832 36378 13860 36654
rect 14280 36654 14332 36660
rect 13910 36615 13966 36624
rect 13945 36476 14253 36485
rect 13945 36474 13951 36476
rect 14007 36474 14031 36476
rect 14087 36474 14111 36476
rect 14167 36474 14191 36476
rect 14247 36474 14253 36476
rect 14007 36422 14009 36474
rect 14189 36422 14191 36474
rect 13945 36420 13951 36422
rect 14007 36420 14031 36422
rect 14087 36420 14111 36422
rect 14167 36420 14191 36422
rect 14247 36420 14253 36422
rect 13945 36411 14253 36420
rect 13820 36372 13872 36378
rect 13820 36314 13872 36320
rect 13820 36032 13872 36038
rect 13820 35974 13872 35980
rect 13832 35737 13860 35974
rect 13818 35728 13874 35737
rect 13818 35663 13874 35672
rect 13832 34678 13860 35663
rect 14280 35556 14332 35562
rect 14280 35498 14332 35504
rect 13945 35388 14253 35397
rect 13945 35386 13951 35388
rect 14007 35386 14031 35388
rect 14087 35386 14111 35388
rect 14167 35386 14191 35388
rect 14247 35386 14253 35388
rect 14007 35334 14009 35386
rect 14189 35334 14191 35386
rect 13945 35332 13951 35334
rect 14007 35332 14031 35334
rect 14087 35332 14111 35334
rect 14167 35332 14191 35334
rect 14247 35332 14253 35334
rect 13945 35323 14253 35332
rect 13820 34672 13872 34678
rect 13820 34614 13872 34620
rect 14292 34610 14320 35498
rect 14280 34604 14332 34610
rect 14280 34546 14332 34552
rect 13726 34504 13782 34513
rect 13726 34439 13782 34448
rect 13820 34400 13872 34406
rect 13820 34342 13872 34348
rect 13728 33584 13780 33590
rect 13648 33544 13728 33572
rect 13728 33526 13780 33532
rect 13634 33008 13690 33017
rect 13634 32943 13690 32952
rect 13648 32434 13676 32943
rect 13636 32428 13688 32434
rect 13636 32370 13688 32376
rect 13544 32360 13596 32366
rect 13544 32302 13596 32308
rect 13636 32224 13688 32230
rect 13636 32166 13688 32172
rect 13648 31890 13676 32166
rect 13636 31884 13688 31890
rect 13636 31826 13688 31832
rect 13544 31748 13596 31754
rect 13596 31708 13676 31736
rect 13544 31690 13596 31696
rect 13648 31385 13676 31708
rect 13634 31376 13690 31385
rect 13544 31340 13596 31346
rect 13634 31311 13690 31320
rect 13544 31282 13596 31288
rect 13452 30796 13504 30802
rect 13452 30738 13504 30744
rect 13464 30258 13492 30738
rect 13556 30598 13584 31282
rect 13544 30592 13596 30598
rect 13544 30534 13596 30540
rect 13452 30252 13504 30258
rect 13636 30252 13688 30258
rect 13452 30194 13504 30200
rect 13556 30212 13636 30240
rect 13360 30048 13412 30054
rect 13360 29990 13412 29996
rect 13268 29640 13320 29646
rect 13268 29582 13320 29588
rect 13372 29458 13400 29990
rect 13280 29430 13400 29458
rect 13280 29306 13308 29430
rect 13268 29300 13320 29306
rect 13556 29288 13584 30212
rect 13636 30194 13688 30200
rect 13634 29608 13690 29617
rect 13634 29543 13690 29552
rect 13268 29242 13320 29248
rect 13372 29260 13584 29288
rect 13268 29096 13320 29102
rect 13268 29038 13320 29044
rect 13280 28937 13308 29038
rect 13266 28928 13322 28937
rect 13266 28863 13322 28872
rect 13280 28490 13308 28863
rect 13268 28484 13320 28490
rect 13268 28426 13320 28432
rect 13268 27464 13320 27470
rect 13268 27406 13320 27412
rect 13280 25974 13308 27406
rect 13372 27010 13400 29260
rect 13648 29220 13676 29543
rect 13740 29345 13768 33526
rect 13832 33454 13860 34342
rect 13945 34300 14253 34309
rect 13945 34298 13951 34300
rect 14007 34298 14031 34300
rect 14087 34298 14111 34300
rect 14167 34298 14191 34300
rect 14247 34298 14253 34300
rect 14007 34246 14009 34298
rect 14189 34246 14191 34298
rect 13945 34244 13951 34246
rect 14007 34244 14031 34246
rect 14087 34244 14111 34246
rect 14167 34244 14191 34246
rect 14247 34244 14253 34246
rect 13945 34235 14253 34244
rect 13912 34196 13964 34202
rect 13912 34138 13964 34144
rect 13820 33448 13872 33454
rect 13820 33390 13872 33396
rect 13924 33300 13952 34138
rect 14280 34060 14332 34066
rect 14280 34002 14332 34008
rect 14292 33590 14320 34002
rect 14280 33584 14332 33590
rect 14280 33526 14332 33532
rect 13832 33272 13952 33300
rect 13832 32552 13860 33272
rect 13945 33212 14253 33221
rect 13945 33210 13951 33212
rect 14007 33210 14031 33212
rect 14087 33210 14111 33212
rect 14167 33210 14191 33212
rect 14247 33210 14253 33212
rect 14007 33158 14009 33210
rect 14189 33158 14191 33210
rect 13945 33156 13951 33158
rect 14007 33156 14031 33158
rect 14087 33156 14111 33158
rect 14167 33156 14191 33158
rect 14247 33156 14253 33158
rect 13945 33147 14253 33156
rect 14292 33096 14320 33526
rect 14384 33266 14412 37062
rect 14476 33454 14504 39335
rect 14646 38720 14702 38729
rect 14646 38655 14702 38664
rect 14556 38412 14608 38418
rect 14556 38354 14608 38360
rect 14568 37806 14596 38354
rect 14556 37800 14608 37806
rect 14556 37742 14608 37748
rect 14556 37188 14608 37194
rect 14556 37130 14608 37136
rect 14568 36922 14596 37130
rect 14556 36916 14608 36922
rect 14556 36858 14608 36864
rect 14556 36576 14608 36582
rect 14556 36518 14608 36524
rect 14568 36310 14596 36518
rect 14556 36304 14608 36310
rect 14556 36246 14608 36252
rect 14556 35828 14608 35834
rect 14556 35770 14608 35776
rect 14568 35290 14596 35770
rect 14556 35284 14608 35290
rect 14556 35226 14608 35232
rect 14556 33992 14608 33998
rect 14556 33934 14608 33940
rect 14568 33590 14596 33934
rect 14556 33584 14608 33590
rect 14556 33526 14608 33532
rect 14464 33448 14516 33454
rect 14568 33425 14596 33526
rect 14464 33390 14516 33396
rect 14554 33416 14610 33425
rect 14554 33351 14610 33360
rect 14554 33280 14610 33289
rect 14384 33238 14504 33266
rect 14016 33068 14320 33096
rect 13912 32564 13964 32570
rect 13832 32524 13912 32552
rect 13912 32506 13964 32512
rect 13820 32428 13872 32434
rect 13820 32370 13872 32376
rect 13832 30394 13860 32370
rect 13924 32366 13952 32506
rect 13912 32360 13964 32366
rect 14016 32337 14044 33068
rect 14372 32904 14424 32910
rect 14372 32846 14424 32852
rect 14280 32836 14332 32842
rect 14280 32778 14332 32784
rect 13912 32302 13964 32308
rect 14002 32328 14058 32337
rect 14002 32263 14058 32272
rect 13945 32124 14253 32133
rect 13945 32122 13951 32124
rect 14007 32122 14031 32124
rect 14087 32122 14111 32124
rect 14167 32122 14191 32124
rect 14247 32122 14253 32124
rect 14007 32070 14009 32122
rect 14189 32070 14191 32122
rect 13945 32068 13951 32070
rect 14007 32068 14031 32070
rect 14087 32068 14111 32070
rect 14167 32068 14191 32070
rect 14247 32068 14253 32070
rect 13945 32059 14253 32068
rect 13912 31952 13964 31958
rect 13910 31920 13912 31929
rect 13964 31920 13966 31929
rect 14292 31890 14320 32778
rect 14384 32230 14412 32846
rect 14372 32224 14424 32230
rect 14372 32166 14424 32172
rect 13910 31855 13966 31864
rect 14280 31884 14332 31890
rect 14280 31826 14332 31832
rect 14096 31816 14148 31822
rect 14148 31764 14228 31770
rect 14096 31758 14228 31764
rect 14108 31742 14228 31758
rect 14200 31226 14228 31742
rect 14200 31198 14320 31226
rect 13945 31036 14253 31045
rect 13945 31034 13951 31036
rect 14007 31034 14031 31036
rect 14087 31034 14111 31036
rect 14167 31034 14191 31036
rect 14247 31034 14253 31036
rect 14007 30982 14009 31034
rect 14189 30982 14191 31034
rect 13945 30980 13951 30982
rect 14007 30980 14031 30982
rect 14087 30980 14111 30982
rect 14167 30980 14191 30982
rect 14247 30980 14253 30982
rect 13945 30971 14253 30980
rect 14186 30696 14242 30705
rect 14186 30631 14188 30640
rect 14240 30631 14242 30640
rect 14188 30602 14240 30608
rect 13820 30388 13872 30394
rect 13820 30330 13872 30336
rect 13820 30048 13872 30054
rect 13820 29990 13872 29996
rect 13832 29594 13860 29990
rect 13945 29948 14253 29957
rect 13945 29946 13951 29948
rect 14007 29946 14031 29948
rect 14087 29946 14111 29948
rect 14167 29946 14191 29948
rect 14247 29946 14253 29948
rect 14007 29894 14009 29946
rect 14189 29894 14191 29946
rect 13945 29892 13951 29894
rect 14007 29892 14031 29894
rect 14087 29892 14111 29894
rect 14167 29892 14191 29894
rect 14247 29892 14253 29894
rect 13945 29883 14253 29892
rect 13910 29744 13966 29753
rect 13910 29679 13912 29688
rect 13964 29679 13966 29688
rect 14188 29708 14240 29714
rect 13912 29650 13964 29656
rect 14292 29696 14320 31198
rect 14240 29668 14320 29696
rect 14188 29650 14240 29656
rect 13832 29566 14136 29594
rect 14004 29504 14056 29510
rect 14004 29446 14056 29452
rect 13726 29336 13782 29345
rect 13726 29271 13782 29280
rect 14016 29220 14044 29446
rect 13556 29192 13676 29220
rect 13740 29192 14044 29220
rect 13452 28960 13504 28966
rect 13452 28902 13504 28908
rect 13464 28626 13492 28902
rect 13452 28620 13504 28626
rect 13452 28562 13504 28568
rect 13372 26982 13492 27010
rect 13360 26920 13412 26926
rect 13360 26862 13412 26868
rect 13268 25968 13320 25974
rect 13268 25910 13320 25916
rect 13268 25696 13320 25702
rect 13268 25638 13320 25644
rect 13096 24670 13216 24698
rect 13096 23526 13124 24670
rect 13176 24608 13228 24614
rect 13176 24550 13228 24556
rect 13188 24410 13216 24550
rect 13176 24404 13228 24410
rect 13176 24346 13228 24352
rect 13280 24290 13308 25638
rect 13372 25158 13400 26862
rect 13464 26353 13492 26982
rect 13450 26344 13506 26353
rect 13450 26279 13506 26288
rect 13464 26058 13492 26279
rect 13556 26246 13584 29192
rect 13740 29050 13768 29192
rect 14016 29102 14044 29192
rect 13648 29022 13768 29050
rect 13912 29096 13964 29102
rect 13912 29038 13964 29044
rect 14004 29096 14056 29102
rect 14004 29038 14056 29044
rect 13648 26926 13676 29022
rect 13924 28994 13952 29038
rect 14108 28994 14136 29566
rect 14188 29504 14240 29510
rect 14188 29446 14240 29452
rect 14200 29050 14228 29446
rect 14280 29300 14332 29306
rect 14280 29242 14332 29248
rect 14292 29170 14320 29242
rect 14280 29164 14332 29170
rect 14280 29106 14332 29112
rect 14200 29022 14320 29050
rect 13924 28966 14136 28994
rect 13945 28860 14253 28869
rect 13945 28858 13951 28860
rect 14007 28858 14031 28860
rect 14087 28858 14111 28860
rect 14167 28858 14191 28860
rect 14247 28858 14253 28860
rect 14007 28806 14009 28858
rect 14189 28806 14191 28858
rect 13945 28804 13951 28806
rect 14007 28804 14031 28806
rect 14087 28804 14111 28806
rect 14167 28804 14191 28806
rect 14247 28804 14253 28806
rect 13726 28792 13782 28801
rect 13945 28795 14253 28804
rect 13726 28727 13782 28736
rect 13636 26920 13688 26926
rect 13636 26862 13688 26868
rect 13636 26784 13688 26790
rect 13636 26726 13688 26732
rect 13648 26586 13676 26726
rect 13636 26580 13688 26586
rect 13636 26522 13688 26528
rect 13544 26240 13596 26246
rect 13544 26182 13596 26188
rect 13464 26030 13584 26058
rect 13360 25152 13412 25158
rect 13360 25094 13412 25100
rect 13188 24262 13308 24290
rect 13084 23520 13136 23526
rect 13084 23462 13136 23468
rect 13082 22808 13138 22817
rect 13082 22743 13138 22752
rect 13096 22642 13124 22743
rect 13084 22636 13136 22642
rect 13084 22578 13136 22584
rect 13084 22500 13136 22506
rect 13084 22442 13136 22448
rect 13096 22137 13124 22442
rect 13082 22128 13138 22137
rect 13082 22063 13138 22072
rect 13084 22024 13136 22030
rect 13084 21966 13136 21972
rect 13096 21690 13124 21966
rect 13188 21876 13216 24262
rect 13268 22976 13320 22982
rect 13268 22918 13320 22924
rect 13280 22098 13308 22918
rect 13268 22092 13320 22098
rect 13268 22034 13320 22040
rect 13188 21848 13308 21876
rect 13174 21720 13230 21729
rect 13084 21684 13136 21690
rect 13174 21655 13230 21664
rect 13084 21626 13136 21632
rect 12912 21406 13032 21434
rect 12912 20602 12940 21406
rect 12992 21344 13044 21350
rect 12992 21286 13044 21292
rect 13004 20913 13032 21286
rect 12990 20904 13046 20913
rect 12990 20839 13046 20848
rect 13188 20788 13216 21655
rect 13280 21418 13308 21848
rect 13268 21412 13320 21418
rect 13268 21354 13320 21360
rect 13372 21298 13400 25094
rect 13452 24812 13504 24818
rect 13452 24754 13504 24760
rect 13464 24585 13492 24754
rect 13450 24576 13506 24585
rect 13450 24511 13506 24520
rect 13452 24064 13504 24070
rect 13452 24006 13504 24012
rect 13464 23662 13492 24006
rect 13452 23656 13504 23662
rect 13452 23598 13504 23604
rect 13464 22574 13492 23598
rect 13556 23338 13584 26030
rect 13636 25900 13688 25906
rect 13636 25842 13688 25848
rect 13648 25265 13676 25842
rect 13634 25256 13690 25265
rect 13634 25191 13690 25200
rect 13648 23508 13676 25191
rect 13740 23633 13768 28727
rect 14004 28552 14056 28558
rect 14002 28520 14004 28529
rect 14056 28520 14058 28529
rect 14002 28455 14058 28464
rect 13912 28212 13964 28218
rect 13912 28154 13964 28160
rect 13924 28082 13952 28154
rect 13912 28076 13964 28082
rect 13912 28018 13964 28024
rect 14188 28076 14240 28082
rect 14188 28018 14240 28024
rect 14094 27976 14150 27985
rect 14200 27962 14228 28018
rect 14150 27934 14228 27962
rect 14094 27911 14150 27920
rect 13945 27772 14253 27781
rect 13945 27770 13951 27772
rect 14007 27770 14031 27772
rect 14087 27770 14111 27772
rect 14167 27770 14191 27772
rect 14247 27770 14253 27772
rect 14007 27718 14009 27770
rect 14189 27718 14191 27770
rect 13945 27716 13951 27718
rect 14007 27716 14031 27718
rect 14087 27716 14111 27718
rect 14167 27716 14191 27718
rect 14247 27716 14253 27718
rect 13945 27707 14253 27716
rect 13945 26684 14253 26693
rect 13945 26682 13951 26684
rect 14007 26682 14031 26684
rect 14087 26682 14111 26684
rect 14167 26682 14191 26684
rect 14247 26682 14253 26684
rect 14007 26630 14009 26682
rect 14189 26630 14191 26682
rect 13945 26628 13951 26630
rect 14007 26628 14031 26630
rect 14087 26628 14111 26630
rect 14167 26628 14191 26630
rect 14247 26628 14253 26630
rect 13945 26619 14253 26628
rect 14292 26466 14320 29022
rect 14384 28694 14412 32166
rect 14476 31754 14504 33238
rect 14554 33215 14610 33224
rect 14568 33046 14596 33215
rect 14556 33040 14608 33046
rect 14556 32982 14608 32988
rect 14476 31726 14596 31754
rect 14464 30592 14516 30598
rect 14464 30534 14516 30540
rect 14476 29170 14504 30534
rect 14464 29164 14516 29170
rect 14464 29106 14516 29112
rect 14372 28688 14424 28694
rect 14372 28630 14424 28636
rect 14568 27962 14596 31726
rect 14660 31113 14688 38655
rect 14752 36378 14780 40854
rect 14832 38208 14884 38214
rect 14832 38150 14884 38156
rect 14740 36372 14792 36378
rect 14740 36314 14792 36320
rect 14740 36100 14792 36106
rect 14740 36042 14792 36048
rect 14752 33998 14780 36042
rect 14844 35329 14872 38150
rect 14830 35320 14886 35329
rect 14830 35255 14886 35264
rect 14830 34504 14886 34513
rect 14830 34439 14886 34448
rect 14740 33992 14792 33998
rect 14740 33934 14792 33940
rect 14844 31793 14872 34439
rect 14936 32881 14964 41958
rect 15028 41274 15056 42758
rect 15108 42628 15160 42634
rect 15108 42570 15160 42576
rect 15016 41268 15068 41274
rect 15016 41210 15068 41216
rect 15120 37262 15148 42570
rect 15200 42288 15252 42294
rect 15200 42230 15252 42236
rect 15212 42106 15240 42230
rect 15304 42226 15332 43046
rect 15292 42220 15344 42226
rect 15292 42162 15344 42168
rect 15212 42078 15332 42106
rect 15200 42016 15252 42022
rect 15200 41958 15252 41964
rect 15212 41721 15240 41958
rect 15198 41712 15254 41721
rect 15198 41647 15254 41656
rect 15304 41664 15332 42078
rect 15396 41818 15424 43046
rect 15488 42770 15516 44540
rect 15672 44010 15700 44540
rect 15672 43982 15792 44010
rect 15658 43888 15714 43897
rect 15658 43823 15714 43832
rect 15672 43314 15700 43823
rect 15568 43308 15620 43314
rect 15568 43250 15620 43256
rect 15660 43308 15712 43314
rect 15660 43250 15712 43256
rect 15476 42764 15528 42770
rect 15476 42706 15528 42712
rect 15476 42628 15528 42634
rect 15476 42570 15528 42576
rect 15384 41812 15436 41818
rect 15384 41754 15436 41760
rect 15488 41682 15516 42570
rect 15384 41676 15436 41682
rect 15304 41636 15384 41664
rect 15384 41618 15436 41624
rect 15476 41676 15528 41682
rect 15476 41618 15528 41624
rect 15382 41576 15438 41585
rect 15382 41511 15438 41520
rect 15396 41478 15424 41511
rect 15200 41472 15252 41478
rect 15200 41414 15252 41420
rect 15384 41472 15436 41478
rect 15476 41472 15528 41478
rect 15384 41414 15436 41420
rect 15474 41440 15476 41449
rect 15528 41440 15530 41449
rect 15212 41138 15240 41414
rect 15474 41375 15530 41384
rect 15580 41274 15608 43250
rect 15660 43104 15712 43110
rect 15660 43046 15712 43052
rect 15672 42906 15700 43046
rect 15660 42900 15712 42906
rect 15660 42842 15712 42848
rect 15764 42838 15792 43982
rect 15752 42832 15804 42838
rect 15752 42774 15804 42780
rect 15660 42152 15712 42158
rect 15660 42094 15712 42100
rect 15568 41268 15620 41274
rect 15568 41210 15620 41216
rect 15476 41200 15528 41206
rect 15476 41142 15528 41148
rect 15200 41132 15252 41138
rect 15200 41074 15252 41080
rect 15200 38208 15252 38214
rect 15200 38150 15252 38156
rect 15212 37874 15240 38150
rect 15200 37868 15252 37874
rect 15200 37810 15252 37816
rect 15108 37256 15160 37262
rect 15108 37198 15160 37204
rect 15120 36786 15148 37198
rect 15108 36780 15160 36786
rect 15108 36722 15160 36728
rect 15016 36372 15068 36378
rect 15016 36314 15068 36320
rect 15028 33590 15056 36314
rect 15120 35290 15148 36722
rect 15200 35692 15252 35698
rect 15200 35634 15252 35640
rect 15108 35284 15160 35290
rect 15108 35226 15160 35232
rect 15120 34184 15148 35226
rect 15212 35018 15240 35634
rect 15292 35488 15344 35494
rect 15292 35430 15344 35436
rect 15200 35012 15252 35018
rect 15200 34954 15252 34960
rect 15304 34746 15332 35430
rect 15292 34740 15344 34746
rect 15292 34682 15344 34688
rect 15488 34490 15516 41142
rect 15672 40186 15700 42094
rect 15752 42016 15804 42022
rect 15752 41958 15804 41964
rect 15660 40180 15712 40186
rect 15660 40122 15712 40128
rect 15764 38758 15792 41958
rect 15856 41138 15884 44540
rect 15936 43104 15988 43110
rect 15936 43046 15988 43052
rect 15948 42226 15976 43046
rect 16040 42906 16068 44540
rect 16120 43308 16172 43314
rect 16120 43250 16172 43256
rect 16028 42900 16080 42906
rect 16028 42842 16080 42848
rect 15936 42220 15988 42226
rect 15936 42162 15988 42168
rect 16028 42220 16080 42226
rect 16028 42162 16080 42168
rect 15936 42016 15988 42022
rect 15936 41958 15988 41964
rect 15948 41721 15976 41958
rect 16040 41818 16068 42162
rect 16028 41812 16080 41818
rect 16028 41754 16080 41760
rect 15934 41712 15990 41721
rect 15934 41647 15990 41656
rect 16026 41576 16082 41585
rect 16026 41511 16082 41520
rect 15844 41132 15896 41138
rect 15844 41074 15896 41080
rect 15936 39908 15988 39914
rect 15936 39850 15988 39856
rect 15844 38956 15896 38962
rect 15844 38898 15896 38904
rect 15752 38752 15804 38758
rect 15752 38694 15804 38700
rect 15856 38010 15884 38898
rect 15844 38004 15896 38010
rect 15844 37946 15896 37952
rect 15568 37664 15620 37670
rect 15568 37606 15620 37612
rect 15580 37330 15608 37606
rect 15660 37392 15712 37398
rect 15660 37334 15712 37340
rect 15568 37324 15620 37330
rect 15568 37266 15620 37272
rect 15580 36650 15608 37266
rect 15568 36644 15620 36650
rect 15568 36586 15620 36592
rect 15672 36394 15700 37334
rect 15752 37256 15804 37262
rect 15752 37198 15804 37204
rect 15764 36922 15792 37198
rect 15844 37120 15896 37126
rect 15844 37062 15896 37068
rect 15856 36922 15884 37062
rect 15752 36916 15804 36922
rect 15752 36858 15804 36864
rect 15844 36916 15896 36922
rect 15844 36858 15896 36864
rect 15304 34462 15516 34490
rect 15580 36366 15700 36394
rect 15200 34196 15252 34202
rect 15120 34156 15200 34184
rect 15200 34138 15252 34144
rect 15304 34048 15332 34462
rect 15384 34400 15436 34406
rect 15384 34342 15436 34348
rect 15212 34020 15332 34048
rect 15016 33584 15068 33590
rect 15016 33526 15068 33532
rect 14922 32872 14978 32881
rect 14922 32807 14978 32816
rect 14922 32600 14978 32609
rect 14922 32535 14978 32544
rect 14830 31784 14886 31793
rect 14830 31719 14886 31728
rect 14832 31680 14884 31686
rect 14832 31622 14884 31628
rect 14740 31136 14792 31142
rect 14646 31104 14702 31113
rect 14740 31078 14792 31084
rect 14646 31039 14702 31048
rect 14648 30388 14700 30394
rect 14648 30330 14700 30336
rect 14660 30297 14688 30330
rect 14646 30288 14702 30297
rect 14646 30223 14702 30232
rect 14660 28082 14688 30223
rect 14752 30190 14780 31078
rect 14740 30184 14792 30190
rect 14740 30126 14792 30132
rect 14752 29306 14780 30126
rect 14740 29300 14792 29306
rect 14740 29242 14792 29248
rect 14738 28792 14794 28801
rect 14738 28727 14794 28736
rect 14752 28626 14780 28727
rect 14740 28620 14792 28626
rect 14740 28562 14792 28568
rect 14648 28076 14700 28082
rect 14648 28018 14700 28024
rect 14568 27934 14688 27962
rect 14372 27872 14424 27878
rect 14372 27814 14424 27820
rect 14462 27840 14518 27849
rect 14384 27674 14412 27814
rect 14462 27775 14518 27784
rect 14372 27668 14424 27674
rect 14372 27610 14424 27616
rect 14476 27418 14504 27775
rect 14556 27668 14608 27674
rect 14556 27610 14608 27616
rect 14200 26438 14320 26466
rect 14384 27390 14504 27418
rect 14200 26382 14228 26438
rect 13912 26376 13964 26382
rect 13912 26318 13964 26324
rect 14188 26376 14240 26382
rect 14188 26318 14240 26324
rect 13924 26042 13952 26318
rect 13912 26036 13964 26042
rect 13912 25978 13964 25984
rect 13945 25596 14253 25605
rect 13945 25594 13951 25596
rect 14007 25594 14031 25596
rect 14087 25594 14111 25596
rect 14167 25594 14191 25596
rect 14247 25594 14253 25596
rect 14007 25542 14009 25594
rect 14189 25542 14191 25594
rect 13945 25540 13951 25542
rect 14007 25540 14031 25542
rect 14087 25540 14111 25542
rect 14167 25540 14191 25542
rect 14247 25540 14253 25542
rect 13945 25531 14253 25540
rect 14280 25152 14332 25158
rect 14280 25094 14332 25100
rect 13820 24880 13872 24886
rect 13820 24822 13872 24828
rect 13832 24206 13860 24822
rect 13945 24508 14253 24517
rect 13945 24506 13951 24508
rect 14007 24506 14031 24508
rect 14087 24506 14111 24508
rect 14167 24506 14191 24508
rect 14247 24506 14253 24508
rect 14007 24454 14009 24506
rect 14189 24454 14191 24506
rect 13945 24452 13951 24454
rect 14007 24452 14031 24454
rect 14087 24452 14111 24454
rect 14167 24452 14191 24454
rect 14247 24452 14253 24454
rect 13945 24443 14253 24452
rect 14292 24206 14320 25094
rect 14384 24954 14412 27390
rect 14464 27328 14516 27334
rect 14464 27270 14516 27276
rect 14476 26926 14504 27270
rect 14464 26920 14516 26926
rect 14464 26862 14516 26868
rect 14476 26586 14504 26862
rect 14464 26580 14516 26586
rect 14464 26522 14516 26528
rect 14372 24948 14424 24954
rect 14372 24890 14424 24896
rect 14372 24676 14424 24682
rect 14372 24618 14424 24624
rect 14384 24410 14412 24618
rect 14372 24404 14424 24410
rect 14372 24346 14424 24352
rect 13820 24200 13872 24206
rect 13820 24142 13872 24148
rect 14280 24200 14332 24206
rect 14280 24142 14332 24148
rect 14372 24132 14424 24138
rect 14568 24120 14596 27610
rect 14660 26994 14688 27934
rect 14844 27130 14872 31622
rect 14936 27713 14964 32535
rect 15016 32224 15068 32230
rect 15016 32166 15068 32172
rect 15028 32026 15056 32166
rect 15016 32020 15068 32026
rect 15016 31962 15068 31968
rect 15108 31816 15160 31822
rect 15028 31764 15108 31770
rect 15028 31758 15160 31764
rect 15028 31742 15148 31758
rect 15028 29510 15056 31742
rect 15212 31278 15240 34020
rect 15292 33924 15344 33930
rect 15292 33866 15344 33872
rect 15304 31414 15332 33866
rect 15396 33658 15424 34342
rect 15384 33652 15436 33658
rect 15384 33594 15436 33600
rect 15382 33144 15438 33153
rect 15382 33079 15438 33088
rect 15396 31754 15424 33079
rect 15476 32904 15528 32910
rect 15476 32846 15528 32852
rect 15488 32434 15516 32846
rect 15476 32428 15528 32434
rect 15476 32370 15528 32376
rect 15396 31726 15516 31754
rect 15382 31648 15438 31657
rect 15382 31583 15438 31592
rect 15292 31408 15344 31414
rect 15292 31350 15344 31356
rect 15200 31272 15252 31278
rect 15200 31214 15252 31220
rect 15198 30968 15254 30977
rect 15108 30932 15160 30938
rect 15198 30903 15254 30912
rect 15108 30874 15160 30880
rect 15120 29646 15148 30874
rect 15212 30326 15240 30903
rect 15304 30734 15332 31350
rect 15292 30728 15344 30734
rect 15292 30670 15344 30676
rect 15200 30320 15252 30326
rect 15200 30262 15252 30268
rect 15108 29640 15160 29646
rect 15212 29617 15240 30262
rect 15108 29582 15160 29588
rect 15198 29608 15254 29617
rect 15016 29504 15068 29510
rect 15016 29446 15068 29452
rect 15016 28552 15068 28558
rect 15016 28494 15068 28500
rect 14922 27704 14978 27713
rect 14922 27639 14978 27648
rect 14832 27124 14884 27130
rect 14832 27066 14884 27072
rect 14648 26988 14700 26994
rect 14648 26930 14700 26936
rect 14660 26042 14688 26930
rect 14740 26920 14792 26926
rect 14740 26862 14792 26868
rect 14752 26790 14780 26862
rect 14740 26784 14792 26790
rect 14740 26726 14792 26732
rect 14648 26036 14700 26042
rect 14648 25978 14700 25984
rect 14752 25922 14780 26726
rect 15028 26586 15056 28494
rect 15120 26602 15148 29582
rect 15198 29543 15254 29552
rect 15200 28756 15252 28762
rect 15200 28698 15252 28704
rect 15292 28756 15344 28762
rect 15292 28698 15344 28704
rect 15212 27946 15240 28698
rect 15304 28558 15332 28698
rect 15292 28552 15344 28558
rect 15292 28494 15344 28500
rect 15200 27940 15252 27946
rect 15200 27882 15252 27888
rect 15292 27872 15344 27878
rect 15292 27814 15344 27820
rect 15304 26926 15332 27814
rect 15292 26920 15344 26926
rect 15292 26862 15344 26868
rect 15016 26580 15068 26586
rect 15120 26574 15240 26602
rect 15016 26522 15068 26528
rect 14922 26480 14978 26489
rect 14978 26438 15148 26466
rect 15212 26450 15240 26574
rect 15304 26450 15332 26862
rect 14922 26415 14978 26424
rect 14660 25894 14780 25922
rect 14924 25900 14976 25906
rect 14660 24721 14688 25894
rect 14924 25842 14976 25848
rect 14832 25288 14884 25294
rect 14832 25230 14884 25236
rect 14740 24812 14792 24818
rect 14740 24754 14792 24760
rect 14646 24712 14702 24721
rect 14646 24647 14702 24656
rect 14648 24608 14700 24614
rect 14648 24550 14700 24556
rect 14660 24410 14688 24550
rect 14648 24404 14700 24410
rect 14648 24346 14700 24352
rect 14424 24092 14596 24120
rect 14372 24074 14424 24080
rect 13820 24064 13872 24070
rect 13820 24006 13872 24012
rect 13832 23730 13860 24006
rect 13820 23724 13872 23730
rect 13820 23666 13872 23672
rect 13912 23656 13964 23662
rect 13726 23624 13782 23633
rect 13726 23559 13782 23568
rect 13832 23604 13912 23610
rect 13832 23598 13964 23604
rect 14280 23656 14332 23662
rect 14280 23598 14332 23604
rect 13832 23582 13952 23598
rect 13648 23480 13768 23508
rect 13556 23310 13676 23338
rect 13452 22568 13504 22574
rect 13452 22510 13504 22516
rect 13450 22128 13506 22137
rect 13506 22086 13584 22114
rect 13450 22063 13506 22072
rect 13450 21856 13506 21865
rect 13450 21791 13506 21800
rect 13464 21554 13492 21791
rect 13452 21548 13504 21554
rect 13452 21490 13504 21496
rect 13452 21412 13504 21418
rect 13452 21354 13504 21360
rect 13004 20760 13216 20788
rect 13280 21270 13400 21298
rect 12900 20596 12952 20602
rect 12900 20538 12952 20544
rect 12808 20460 12860 20466
rect 12808 20402 12860 20408
rect 12900 20460 12952 20466
rect 12900 20402 12952 20408
rect 12716 19712 12768 19718
rect 12716 19654 12768 19660
rect 12624 18964 12676 18970
rect 12624 18906 12676 18912
rect 12728 18426 12756 19654
rect 12806 19136 12862 19145
rect 12806 19071 12862 19080
rect 12820 18970 12848 19071
rect 12808 18964 12860 18970
rect 12808 18906 12860 18912
rect 12452 18380 12572 18408
rect 12716 18420 12768 18426
rect 12452 17542 12480 18380
rect 12716 18362 12768 18368
rect 12530 18320 12586 18329
rect 12912 18306 12940 20402
rect 12530 18255 12586 18264
rect 12728 18278 12940 18306
rect 12440 17536 12492 17542
rect 12440 17478 12492 17484
rect 12440 16992 12492 16998
rect 12440 16934 12492 16940
rect 12452 16590 12480 16934
rect 12440 16584 12492 16590
rect 12440 16526 12492 16532
rect 12452 16182 12480 16526
rect 12440 16176 12492 16182
rect 12440 16118 12492 16124
rect 12452 15473 12480 16118
rect 12438 15464 12494 15473
rect 12438 15399 12494 15408
rect 12452 15094 12480 15399
rect 12440 15088 12492 15094
rect 12440 15030 12492 15036
rect 12440 14476 12492 14482
rect 12440 14418 12492 14424
rect 12346 13832 12402 13841
rect 12346 13767 12402 13776
rect 12452 13530 12480 14418
rect 12544 13705 12572 18255
rect 12624 17740 12676 17746
rect 12624 17682 12676 17688
rect 12636 17610 12664 17682
rect 12624 17604 12676 17610
rect 12624 17546 12676 17552
rect 12636 16998 12664 17546
rect 12624 16992 12676 16998
rect 12624 16934 12676 16940
rect 12728 16794 12756 18278
rect 12808 18080 12860 18086
rect 12808 18022 12860 18028
rect 12820 17785 12848 18022
rect 12900 17876 12952 17882
rect 12900 17818 12952 17824
rect 12806 17776 12862 17785
rect 12806 17711 12862 17720
rect 12808 17060 12860 17066
rect 12808 17002 12860 17008
rect 12716 16788 12768 16794
rect 12716 16730 12768 16736
rect 12624 16584 12676 16590
rect 12624 16526 12676 16532
rect 12636 16153 12664 16526
rect 12622 16144 12678 16153
rect 12622 16079 12678 16088
rect 12728 15994 12756 16730
rect 12820 16250 12848 17002
rect 12808 16244 12860 16250
rect 12808 16186 12860 16192
rect 12636 15966 12756 15994
rect 12636 15570 12664 15966
rect 12624 15564 12676 15570
rect 12624 15506 12676 15512
rect 12716 15564 12768 15570
rect 12716 15506 12768 15512
rect 12530 13696 12586 13705
rect 12530 13631 12586 13640
rect 12440 13524 12492 13530
rect 12440 13466 12492 13472
rect 12440 13184 12492 13190
rect 12440 13126 12492 13132
rect 12254 11928 12310 11937
rect 12254 11863 12310 11872
rect 12348 11552 12400 11558
rect 12348 11494 12400 11500
rect 12360 11150 12388 11494
rect 12348 11144 12400 11150
rect 12348 11086 12400 11092
rect 12452 10996 12480 13126
rect 12532 12912 12584 12918
rect 12532 12854 12584 12860
rect 12544 12442 12572 12854
rect 12532 12436 12584 12442
rect 12532 12378 12584 12384
rect 12636 12220 12664 15506
rect 12728 15162 12756 15506
rect 12716 15156 12768 15162
rect 12716 15098 12768 15104
rect 12912 15042 12940 17818
rect 13004 17338 13032 20760
rect 13174 20632 13230 20641
rect 13084 20596 13136 20602
rect 13174 20567 13176 20576
rect 13084 20538 13136 20544
rect 13228 20567 13230 20576
rect 13176 20538 13228 20544
rect 13096 19786 13124 20538
rect 13176 20392 13228 20398
rect 13176 20334 13228 20340
rect 13084 19780 13136 19786
rect 13084 19722 13136 19728
rect 13084 19236 13136 19242
rect 13084 19178 13136 19184
rect 13096 18426 13124 19178
rect 13084 18420 13136 18426
rect 13084 18362 13136 18368
rect 13084 18216 13136 18222
rect 13084 18158 13136 18164
rect 13096 17610 13124 18158
rect 13084 17604 13136 17610
rect 13084 17546 13136 17552
rect 12992 17332 13044 17338
rect 12992 17274 13044 17280
rect 13084 16108 13136 16114
rect 13084 16050 13136 16056
rect 12728 15014 12940 15042
rect 12728 14521 12756 15014
rect 12900 14952 12952 14958
rect 12900 14894 12952 14900
rect 12808 14884 12860 14890
rect 12808 14826 12860 14832
rect 12714 14512 12770 14521
rect 12714 14447 12716 14456
rect 12768 14447 12770 14456
rect 12716 14418 12768 14424
rect 12820 12850 12848 14826
rect 12912 14618 12940 14894
rect 12900 14612 12952 14618
rect 12900 14554 12952 14560
rect 12912 13938 12940 14554
rect 12992 14408 13044 14414
rect 12992 14350 13044 14356
rect 13004 14074 13032 14350
rect 12992 14068 13044 14074
rect 12992 14010 13044 14016
rect 12900 13932 12952 13938
rect 12900 13874 12952 13880
rect 12808 12844 12860 12850
rect 12808 12786 12860 12792
rect 12898 12744 12954 12753
rect 13096 12730 13124 16050
rect 13188 15502 13216 20334
rect 13280 17134 13308 21270
rect 13360 21004 13412 21010
rect 13360 20946 13412 20952
rect 13372 20058 13400 20946
rect 13360 20052 13412 20058
rect 13360 19994 13412 20000
rect 13360 19304 13412 19310
rect 13360 19246 13412 19252
rect 13372 18970 13400 19246
rect 13360 18964 13412 18970
rect 13360 18906 13412 18912
rect 13358 18320 13414 18329
rect 13358 18255 13414 18264
rect 13372 17678 13400 18255
rect 13360 17672 13412 17678
rect 13360 17614 13412 17620
rect 13268 17128 13320 17134
rect 13268 17070 13320 17076
rect 13360 17128 13412 17134
rect 13360 17070 13412 17076
rect 13280 16674 13308 17070
rect 13372 16794 13400 17070
rect 13360 16788 13412 16794
rect 13360 16730 13412 16736
rect 13280 16646 13400 16674
rect 13268 16040 13320 16046
rect 13268 15982 13320 15988
rect 13176 15496 13228 15502
rect 13280 15473 13308 15982
rect 13176 15438 13228 15444
rect 13266 15464 13322 15473
rect 13188 14074 13216 15438
rect 13266 15399 13322 15408
rect 13372 15348 13400 16646
rect 13464 16250 13492 21354
rect 13556 19378 13584 22086
rect 13648 21622 13676 23310
rect 13636 21616 13688 21622
rect 13636 21558 13688 21564
rect 13740 21468 13768 23480
rect 13832 23254 13860 23582
rect 13945 23420 14253 23429
rect 13945 23418 13951 23420
rect 14007 23418 14031 23420
rect 14087 23418 14111 23420
rect 14167 23418 14191 23420
rect 14247 23418 14253 23420
rect 14007 23366 14009 23418
rect 14189 23366 14191 23418
rect 13945 23364 13951 23366
rect 14007 23364 14031 23366
rect 14087 23364 14111 23366
rect 14167 23364 14191 23366
rect 14247 23364 14253 23366
rect 13945 23355 14253 23364
rect 14292 23322 14320 23598
rect 14280 23316 14332 23322
rect 14280 23258 14332 23264
rect 13820 23248 13872 23254
rect 13820 23190 13872 23196
rect 14292 22574 14320 23258
rect 13912 22568 13964 22574
rect 13832 22516 13912 22522
rect 13832 22510 13964 22516
rect 14280 22568 14332 22574
rect 14280 22510 14332 22516
rect 13832 22494 13952 22510
rect 13832 22234 13860 22494
rect 13945 22332 14253 22341
rect 13945 22330 13951 22332
rect 14007 22330 14031 22332
rect 14087 22330 14111 22332
rect 14167 22330 14191 22332
rect 14247 22330 14253 22332
rect 14007 22278 14009 22330
rect 14189 22278 14191 22330
rect 13945 22276 13951 22278
rect 14007 22276 14031 22278
rect 14087 22276 14111 22278
rect 14167 22276 14191 22278
rect 14247 22276 14253 22278
rect 13945 22267 14253 22276
rect 14384 22234 14412 24074
rect 14648 24064 14700 24070
rect 14462 24032 14518 24041
rect 14648 24006 14700 24012
rect 14462 23967 14518 23976
rect 13820 22228 13872 22234
rect 13820 22170 13872 22176
rect 14188 22228 14240 22234
rect 14188 22170 14240 22176
rect 14372 22228 14424 22234
rect 14372 22170 14424 22176
rect 13820 22092 13872 22098
rect 13820 22034 13872 22040
rect 13648 21440 13768 21468
rect 13544 19372 13596 19378
rect 13544 19314 13596 19320
rect 13556 16998 13584 19314
rect 13544 16992 13596 16998
rect 13544 16934 13596 16940
rect 13452 16244 13504 16250
rect 13452 16186 13504 16192
rect 13280 15320 13400 15348
rect 13176 14068 13228 14074
rect 13176 14010 13228 14016
rect 13176 13932 13228 13938
rect 13176 13874 13228 13880
rect 13188 13172 13216 13874
rect 13280 13326 13308 15320
rect 13556 14890 13584 16934
rect 13648 16182 13676 21440
rect 13728 21344 13780 21350
rect 13728 21286 13780 21292
rect 13740 20890 13768 21286
rect 13832 21010 13860 22034
rect 14200 21332 14228 22170
rect 14476 22094 14504 23967
rect 14556 23520 14608 23526
rect 14556 23462 14608 23468
rect 14568 23322 14596 23462
rect 14556 23316 14608 23322
rect 14556 23258 14608 23264
rect 14556 23044 14608 23050
rect 14556 22986 14608 22992
rect 14384 22066 14504 22094
rect 14384 21978 14412 22066
rect 14292 21950 14412 21978
rect 14292 21457 14320 21950
rect 14372 21888 14424 21894
rect 14372 21830 14424 21836
rect 14278 21448 14334 21457
rect 14278 21383 14334 21392
rect 14280 21344 14332 21350
rect 14200 21304 14280 21332
rect 14280 21286 14332 21292
rect 13945 21244 14253 21253
rect 13945 21242 13951 21244
rect 14007 21242 14031 21244
rect 14087 21242 14111 21244
rect 14167 21242 14191 21244
rect 14247 21242 14253 21244
rect 14007 21190 14009 21242
rect 14189 21190 14191 21242
rect 13945 21188 13951 21190
rect 14007 21188 14031 21190
rect 14087 21188 14111 21190
rect 14167 21188 14191 21190
rect 14247 21188 14253 21190
rect 13945 21179 14253 21188
rect 13820 21004 13872 21010
rect 13820 20946 13872 20952
rect 14096 21004 14148 21010
rect 14096 20946 14148 20952
rect 13910 20904 13966 20913
rect 13740 20862 13860 20890
rect 13728 20324 13780 20330
rect 13728 20266 13780 20272
rect 13740 19990 13768 20266
rect 13728 19984 13780 19990
rect 13728 19926 13780 19932
rect 13728 19780 13780 19786
rect 13728 19722 13780 19728
rect 13740 19009 13768 19722
rect 13726 19000 13782 19009
rect 13726 18935 13782 18944
rect 13728 18420 13780 18426
rect 13728 18362 13780 18368
rect 13740 18057 13768 18362
rect 13832 18290 13860 20862
rect 13910 20839 13966 20848
rect 13924 20806 13952 20839
rect 13912 20800 13964 20806
rect 13912 20742 13964 20748
rect 14108 20602 14136 20946
rect 14096 20596 14148 20602
rect 14096 20538 14148 20544
rect 14142 20392 14194 20398
rect 14292 20380 14320 21286
rect 14194 20352 14320 20380
rect 14142 20334 14194 20340
rect 13945 20156 14253 20165
rect 13945 20154 13951 20156
rect 14007 20154 14031 20156
rect 14087 20154 14111 20156
rect 14167 20154 14191 20156
rect 14247 20154 14253 20156
rect 14007 20102 14009 20154
rect 14189 20102 14191 20154
rect 13945 20100 13951 20102
rect 14007 20100 14031 20102
rect 14087 20100 14111 20102
rect 14167 20100 14191 20102
rect 14247 20100 14253 20102
rect 13945 20091 14253 20100
rect 14094 19952 14150 19961
rect 14094 19887 14150 19896
rect 14278 19952 14334 19961
rect 14278 19887 14334 19896
rect 14108 19689 14136 19887
rect 14292 19854 14320 19887
rect 14280 19848 14332 19854
rect 14280 19790 14332 19796
rect 14094 19680 14150 19689
rect 14094 19615 14150 19624
rect 14280 19168 14332 19174
rect 14280 19110 14332 19116
rect 13945 19068 14253 19077
rect 13945 19066 13951 19068
rect 14007 19066 14031 19068
rect 14087 19066 14111 19068
rect 14167 19066 14191 19068
rect 14247 19066 14253 19068
rect 14007 19014 14009 19066
rect 14189 19014 14191 19066
rect 13945 19012 13951 19014
rect 14007 19012 14031 19014
rect 14087 19012 14111 19014
rect 14167 19012 14191 19014
rect 14247 19012 14253 19014
rect 13945 19003 14253 19012
rect 14292 18630 14320 19110
rect 14280 18624 14332 18630
rect 14280 18566 14332 18572
rect 13820 18284 13872 18290
rect 13820 18226 13872 18232
rect 13726 18048 13782 18057
rect 13726 17983 13782 17992
rect 13636 16176 13688 16182
rect 13636 16118 13688 16124
rect 13832 15688 13860 18226
rect 13945 17980 14253 17989
rect 13945 17978 13951 17980
rect 14007 17978 14031 17980
rect 14087 17978 14111 17980
rect 14167 17978 14191 17980
rect 14247 17978 14253 17980
rect 14007 17926 14009 17978
rect 14189 17926 14191 17978
rect 13945 17924 13951 17926
rect 14007 17924 14031 17926
rect 14087 17924 14111 17926
rect 14167 17924 14191 17926
rect 14247 17924 14253 17926
rect 13945 17915 14253 17924
rect 14280 16992 14332 16998
rect 14280 16934 14332 16940
rect 13945 16892 14253 16901
rect 13945 16890 13951 16892
rect 14007 16890 14031 16892
rect 14087 16890 14111 16892
rect 14167 16890 14191 16892
rect 14247 16890 14253 16892
rect 14007 16838 14009 16890
rect 14189 16838 14191 16890
rect 13945 16836 13951 16838
rect 14007 16836 14031 16838
rect 14087 16836 14111 16838
rect 14167 16836 14191 16838
rect 14247 16836 14253 16838
rect 13945 16827 14253 16836
rect 14292 16590 14320 16934
rect 14280 16584 14332 16590
rect 14280 16526 14332 16532
rect 14280 15904 14332 15910
rect 14280 15846 14332 15852
rect 13945 15804 14253 15813
rect 13945 15802 13951 15804
rect 14007 15802 14031 15804
rect 14087 15802 14111 15804
rect 14167 15802 14191 15804
rect 14247 15802 14253 15804
rect 14007 15750 14009 15802
rect 14189 15750 14191 15802
rect 13945 15748 13951 15750
rect 14007 15748 14031 15750
rect 14087 15748 14111 15750
rect 14167 15748 14191 15750
rect 14247 15748 14253 15750
rect 13945 15739 14253 15748
rect 14292 15706 14320 15846
rect 14280 15700 14332 15706
rect 13832 15660 13952 15688
rect 13820 15360 13872 15366
rect 13740 15308 13820 15314
rect 13740 15302 13872 15308
rect 13740 15286 13860 15302
rect 13544 14884 13596 14890
rect 13544 14826 13596 14832
rect 13556 14482 13584 14826
rect 13636 14816 13688 14822
rect 13636 14758 13688 14764
rect 13648 14618 13676 14758
rect 13636 14612 13688 14618
rect 13636 14554 13688 14560
rect 13360 14476 13412 14482
rect 13360 14418 13412 14424
rect 13544 14476 13596 14482
rect 13544 14418 13596 14424
rect 13372 13734 13400 14418
rect 13544 14068 13596 14074
rect 13544 14010 13596 14016
rect 13360 13728 13412 13734
rect 13360 13670 13412 13676
rect 13268 13320 13320 13326
rect 13268 13262 13320 13268
rect 13188 13144 13308 13172
rect 13174 13016 13230 13025
rect 13174 12951 13230 12960
rect 12898 12679 12900 12688
rect 12952 12679 12954 12688
rect 13004 12702 13124 12730
rect 12900 12650 12952 12656
rect 12806 12472 12862 12481
rect 12806 12407 12862 12416
rect 12900 12436 12952 12442
rect 12636 12192 12756 12220
rect 12622 12064 12678 12073
rect 12622 11999 12678 12008
rect 12532 11688 12584 11694
rect 12532 11630 12584 11636
rect 12268 10968 12480 10996
rect 12268 9382 12296 10968
rect 12544 10606 12572 11630
rect 12532 10600 12584 10606
rect 12532 10542 12584 10548
rect 12360 10130 12572 10146
rect 12348 10124 12572 10130
rect 12400 10118 12572 10124
rect 12348 10066 12400 10072
rect 12544 9874 12572 10118
rect 12452 9846 12572 9874
rect 12348 9512 12400 9518
rect 12348 9454 12400 9460
rect 12256 9376 12308 9382
rect 12360 9353 12388 9454
rect 12256 9318 12308 9324
rect 12346 9344 12402 9353
rect 12268 8974 12296 9318
rect 12346 9279 12402 9288
rect 12346 9072 12402 9081
rect 12346 9007 12402 9016
rect 12256 8968 12308 8974
rect 12256 8910 12308 8916
rect 12360 8906 12388 9007
rect 12348 8900 12400 8906
rect 12348 8842 12400 8848
rect 12256 8832 12308 8838
rect 12256 8774 12308 8780
rect 12268 8430 12296 8774
rect 12452 8634 12480 9846
rect 12530 9752 12586 9761
rect 12530 9687 12586 9696
rect 12440 8628 12492 8634
rect 12440 8570 12492 8576
rect 12256 8424 12308 8430
rect 12256 8366 12308 8372
rect 12438 8392 12494 8401
rect 12438 8327 12494 8336
rect 12176 8044 12294 8072
rect 11704 8016 11756 8022
rect 11704 7958 11756 7964
rect 11796 8016 11848 8022
rect 11796 7958 11848 7964
rect 11992 7970 12020 8044
rect 11244 7812 11296 7818
rect 11624 7806 11744 7834
rect 11244 7754 11296 7760
rect 11256 7478 11284 7754
rect 11346 7644 11654 7653
rect 11346 7642 11352 7644
rect 11408 7642 11432 7644
rect 11488 7642 11512 7644
rect 11568 7642 11592 7644
rect 11648 7642 11654 7644
rect 11408 7590 11410 7642
rect 11590 7590 11592 7642
rect 11346 7588 11352 7590
rect 11408 7588 11432 7590
rect 11488 7588 11512 7590
rect 11568 7588 11592 7590
rect 11648 7588 11654 7590
rect 11346 7579 11654 7588
rect 11716 7546 11744 7806
rect 11704 7540 11756 7546
rect 11704 7482 11756 7488
rect 11244 7472 11296 7478
rect 11244 7414 11296 7420
rect 11704 7404 11756 7410
rect 11704 7346 11756 7352
rect 11244 7200 11296 7206
rect 11244 7142 11296 7148
rect 11256 6458 11284 7142
rect 11716 6934 11744 7346
rect 11808 7002 11836 7958
rect 11992 7954 12112 7970
rect 11992 7948 12124 7954
rect 11992 7942 12072 7948
rect 12072 7890 12124 7896
rect 12164 7880 12216 7886
rect 11900 7828 12164 7834
rect 11900 7822 12216 7828
rect 12266 7834 12294 8044
rect 12348 7948 12400 7954
rect 12348 7890 12400 7896
rect 11900 7806 12202 7822
rect 12266 7806 12296 7834
rect 11900 7206 11928 7806
rect 11980 7744 12032 7750
rect 12268 7732 12296 7806
rect 11980 7686 12032 7692
rect 12176 7704 12296 7732
rect 11888 7200 11940 7206
rect 11888 7142 11940 7148
rect 11796 6996 11848 7002
rect 11796 6938 11848 6944
rect 11704 6928 11756 6934
rect 11704 6870 11756 6876
rect 11888 6656 11940 6662
rect 11888 6598 11940 6604
rect 11346 6556 11654 6565
rect 11346 6554 11352 6556
rect 11408 6554 11432 6556
rect 11488 6554 11512 6556
rect 11568 6554 11592 6556
rect 11648 6554 11654 6556
rect 11408 6502 11410 6554
rect 11590 6502 11592 6554
rect 11346 6500 11352 6502
rect 11408 6500 11432 6502
rect 11488 6500 11512 6502
rect 11568 6500 11592 6502
rect 11648 6500 11654 6502
rect 11346 6491 11654 6500
rect 11244 6452 11296 6458
rect 11244 6394 11296 6400
rect 11900 6186 11928 6598
rect 11888 6180 11940 6186
rect 11888 6122 11940 6128
rect 11796 6112 11848 6118
rect 11796 6054 11848 6060
rect 11704 5908 11756 5914
rect 11704 5850 11756 5856
rect 11346 5468 11654 5477
rect 11346 5466 11352 5468
rect 11408 5466 11432 5468
rect 11488 5466 11512 5468
rect 11568 5466 11592 5468
rect 11648 5466 11654 5468
rect 11408 5414 11410 5466
rect 11590 5414 11592 5466
rect 11346 5412 11352 5414
rect 11408 5412 11432 5414
rect 11488 5412 11512 5414
rect 11568 5412 11592 5414
rect 11648 5412 11654 5414
rect 11346 5403 11654 5412
rect 11152 5160 11204 5166
rect 11152 5102 11204 5108
rect 11346 4380 11654 4389
rect 11346 4378 11352 4380
rect 11408 4378 11432 4380
rect 11488 4378 11512 4380
rect 11568 4378 11592 4380
rect 11648 4378 11654 4380
rect 11408 4326 11410 4378
rect 11590 4326 11592 4378
rect 11346 4324 11352 4326
rect 11408 4324 11432 4326
rect 11488 4324 11512 4326
rect 11568 4324 11592 4326
rect 11648 4324 11654 4326
rect 11346 4315 11654 4324
rect 11612 3732 11664 3738
rect 11612 3674 11664 3680
rect 11624 3398 11652 3674
rect 11612 3392 11664 3398
rect 11612 3334 11664 3340
rect 11346 3292 11654 3301
rect 11346 3290 11352 3292
rect 11408 3290 11432 3292
rect 11488 3290 11512 3292
rect 11568 3290 11592 3292
rect 11648 3290 11654 3292
rect 11408 3238 11410 3290
rect 11590 3238 11592 3290
rect 11346 3236 11352 3238
rect 11408 3236 11432 3238
rect 11488 3236 11512 3238
rect 11568 3236 11592 3238
rect 11648 3236 11654 3238
rect 11346 3227 11654 3236
rect 10836 3012 10916 3040
rect 11060 3052 11112 3058
rect 10784 2994 10836 3000
rect 11060 2994 11112 3000
rect 11072 2774 11100 2994
rect 10980 2746 11100 2774
rect 10980 2650 11008 2746
rect 10692 2644 10744 2650
rect 10692 2586 10744 2592
rect 10968 2644 11020 2650
rect 10968 2586 11020 2592
rect 10876 2576 10928 2582
rect 11060 2576 11112 2582
rect 10876 2518 10928 2524
rect 10980 2524 11060 2530
rect 10980 2518 11112 2524
rect 10784 2508 10836 2514
rect 10784 2450 10836 2456
rect 10600 2440 10652 2446
rect 10600 2382 10652 2388
rect 10508 2304 10560 2310
rect 10508 2246 10560 2252
rect 10416 2032 10468 2038
rect 10416 1974 10468 1980
rect 10520 1902 10548 2246
rect 10508 1896 10560 1902
rect 10508 1838 10560 1844
rect 10796 1834 10824 2450
rect 10888 2378 10916 2518
rect 10980 2502 11100 2518
rect 10876 2372 10928 2378
rect 10876 2314 10928 2320
rect 10600 1828 10652 1834
rect 10600 1770 10652 1776
rect 10784 1828 10836 1834
rect 10784 1770 10836 1776
rect 10508 1760 10560 1766
rect 10508 1702 10560 1708
rect 10416 1420 10468 1426
rect 10416 1362 10468 1368
rect 10428 678 10456 1362
rect 10416 672 10468 678
rect 10416 614 10468 620
rect 10520 160 10548 1702
rect 10612 1358 10640 1770
rect 10980 1562 11008 2502
rect 11612 2440 11664 2446
rect 11716 2428 11744 5850
rect 11808 3738 11836 6054
rect 11992 4282 12020 7686
rect 12070 7576 12126 7585
rect 12070 7511 12126 7520
rect 11980 4276 12032 4282
rect 11980 4218 12032 4224
rect 11796 3732 11848 3738
rect 11796 3674 11848 3680
rect 12084 3058 12112 7511
rect 12176 6322 12204 7704
rect 12360 7546 12388 7890
rect 12348 7540 12400 7546
rect 12348 7482 12400 7488
rect 12452 7410 12480 8327
rect 12440 7404 12492 7410
rect 12440 7346 12492 7352
rect 12544 7313 12572 9687
rect 12530 7304 12586 7313
rect 12440 7268 12492 7274
rect 12530 7239 12586 7248
rect 12440 7210 12492 7216
rect 12346 7168 12402 7177
rect 12346 7103 12402 7112
rect 12254 7032 12310 7041
rect 12254 6967 12310 6976
rect 12268 6798 12296 6967
rect 12256 6792 12308 6798
rect 12256 6734 12308 6740
rect 12164 6316 12216 6322
rect 12164 6258 12216 6264
rect 12360 6066 12388 7103
rect 12268 6038 12388 6066
rect 12164 5636 12216 5642
rect 12164 5578 12216 5584
rect 12176 5545 12204 5578
rect 12162 5536 12218 5545
rect 12162 5471 12218 5480
rect 12268 5273 12296 6038
rect 12452 5302 12480 7210
rect 12530 6896 12586 6905
rect 12530 6831 12586 6840
rect 12544 5778 12572 6831
rect 12532 5772 12584 5778
rect 12532 5714 12584 5720
rect 12440 5296 12492 5302
rect 12254 5264 12310 5273
rect 12440 5238 12492 5244
rect 12254 5199 12310 5208
rect 12636 3602 12664 11999
rect 12728 10130 12756 12192
rect 12716 10124 12768 10130
rect 12716 10066 12768 10072
rect 12716 9444 12768 9450
rect 12716 9386 12768 9392
rect 12728 9178 12756 9386
rect 12716 9172 12768 9178
rect 12716 9114 12768 9120
rect 12714 9072 12770 9081
rect 12714 9007 12770 9016
rect 12728 5574 12756 9007
rect 12820 6089 12848 12407
rect 12900 12378 12952 12384
rect 12912 10146 12940 12378
rect 13004 12238 13032 12702
rect 13084 12640 13136 12646
rect 13084 12582 13136 12588
rect 12992 12232 13044 12238
rect 12992 12174 13044 12180
rect 13096 11626 13124 12582
rect 12992 11620 13044 11626
rect 12992 11562 13044 11568
rect 13084 11620 13136 11626
rect 13084 11562 13136 11568
rect 13004 11150 13032 11562
rect 12992 11144 13044 11150
rect 12992 11086 13044 11092
rect 13084 10464 13136 10470
rect 13084 10406 13136 10412
rect 12912 10118 13032 10146
rect 12900 10056 12952 10062
rect 12900 9998 12952 10004
rect 12912 9178 12940 9998
rect 13004 9897 13032 10118
rect 12990 9888 13046 9897
rect 12990 9823 13046 9832
rect 12990 9616 13046 9625
rect 12990 9551 13046 9560
rect 12900 9172 12952 9178
rect 12900 9114 12952 9120
rect 12900 8424 12952 8430
rect 12900 8366 12952 8372
rect 12912 8022 12940 8366
rect 12900 8016 12952 8022
rect 12900 7958 12952 7964
rect 13004 7834 13032 9551
rect 13096 8906 13124 10406
rect 13084 8900 13136 8906
rect 13084 8842 13136 8848
rect 13096 8498 13124 8842
rect 13084 8492 13136 8498
rect 13084 8434 13136 8440
rect 13004 7806 13124 7834
rect 12900 7744 12952 7750
rect 12900 7686 12952 7692
rect 12992 7744 13044 7750
rect 12992 7686 13044 7692
rect 12912 7546 12940 7686
rect 12900 7540 12952 7546
rect 12900 7482 12952 7488
rect 12898 7304 12954 7313
rect 12898 7239 12954 7248
rect 12912 7002 12940 7239
rect 12900 6996 12952 7002
rect 12900 6938 12952 6944
rect 12900 6384 12952 6390
rect 12900 6326 12952 6332
rect 12806 6080 12862 6089
rect 12806 6015 12862 6024
rect 12716 5568 12768 5574
rect 12716 5510 12768 5516
rect 12912 5166 12940 6326
rect 13004 5370 13032 7686
rect 12992 5364 13044 5370
rect 12992 5306 13044 5312
rect 12900 5160 12952 5166
rect 12900 5102 12952 5108
rect 12808 4820 12860 4826
rect 12808 4762 12860 4768
rect 12624 3596 12676 3602
rect 12624 3538 12676 3544
rect 12820 3058 12848 4762
rect 13096 4214 13124 7806
rect 13188 5273 13216 12951
rect 13280 10810 13308 13144
rect 13372 11762 13400 13670
rect 13452 12640 13504 12646
rect 13452 12582 13504 12588
rect 13464 12442 13492 12582
rect 13452 12436 13504 12442
rect 13452 12378 13504 12384
rect 13452 12164 13504 12170
rect 13452 12106 13504 12112
rect 13360 11756 13412 11762
rect 13360 11698 13412 11704
rect 13372 11558 13400 11698
rect 13360 11552 13412 11558
rect 13360 11494 13412 11500
rect 13360 11348 13412 11354
rect 13360 11290 13412 11296
rect 13268 10804 13320 10810
rect 13268 10746 13320 10752
rect 13280 9722 13308 10746
rect 13372 10606 13400 11290
rect 13464 11218 13492 12106
rect 13556 11801 13584 14010
rect 13740 12986 13768 15286
rect 13924 15178 13952 15660
rect 14280 15642 14332 15648
rect 14384 15502 14412 21830
rect 14464 21412 14516 21418
rect 14464 21354 14516 21360
rect 14476 19922 14504 21354
rect 14464 19916 14516 19922
rect 14464 19858 14516 19864
rect 14464 17672 14516 17678
rect 14464 17614 14516 17620
rect 14372 15496 14424 15502
rect 14372 15438 14424 15444
rect 14476 15314 14504 17614
rect 14568 15570 14596 22986
rect 14660 19922 14688 24006
rect 14752 23322 14780 24754
rect 14844 24410 14872 25230
rect 14936 25158 14964 25842
rect 15016 25288 15068 25294
rect 15016 25230 15068 25236
rect 14924 25152 14976 25158
rect 14924 25094 14976 25100
rect 14936 24818 14964 25094
rect 15028 24868 15056 25230
rect 15120 24970 15148 26438
rect 15200 26444 15252 26450
rect 15200 26386 15252 26392
rect 15292 26444 15344 26450
rect 15292 26386 15344 26392
rect 15292 25900 15344 25906
rect 15292 25842 15344 25848
rect 15304 25809 15332 25842
rect 15290 25800 15346 25809
rect 15290 25735 15346 25744
rect 15396 25294 15424 31583
rect 15488 31498 15516 31726
rect 15580 31686 15608 36366
rect 15844 36032 15896 36038
rect 15844 35974 15896 35980
rect 15856 33833 15884 35974
rect 15948 34626 15976 39850
rect 16040 38554 16068 41511
rect 16132 41002 16160 43250
rect 16120 40996 16172 41002
rect 16120 40938 16172 40944
rect 16224 40730 16252 44540
rect 16408 43330 16436 44540
rect 16592 43738 16620 44540
rect 16776 43858 16804 44540
rect 16960 43926 16988 44540
rect 16948 43920 17000 43926
rect 16948 43862 17000 43868
rect 16764 43852 16816 43858
rect 16764 43794 16816 43800
rect 16592 43710 16988 43738
rect 16544 43548 16852 43557
rect 16544 43546 16550 43548
rect 16606 43546 16630 43548
rect 16686 43546 16710 43548
rect 16766 43546 16790 43548
rect 16846 43546 16852 43548
rect 16606 43494 16608 43546
rect 16788 43494 16790 43546
rect 16544 43492 16550 43494
rect 16606 43492 16630 43494
rect 16686 43492 16710 43494
rect 16766 43492 16790 43494
rect 16846 43492 16852 43494
rect 16544 43483 16852 43492
rect 16960 43450 16988 43710
rect 16580 43444 16632 43450
rect 16580 43386 16632 43392
rect 16948 43444 17000 43450
rect 16948 43386 17000 43392
rect 16592 43330 16620 43386
rect 16408 43302 16620 43330
rect 16304 43240 16356 43246
rect 16304 43182 16356 43188
rect 16316 42158 16344 43182
rect 16396 42900 16448 42906
rect 17144 42888 17172 44540
rect 17328 43382 17356 44540
rect 17408 43920 17460 43926
rect 17408 43862 17460 43868
rect 17316 43376 17368 43382
rect 17316 43318 17368 43324
rect 17316 43240 17368 43246
rect 17316 43182 17368 43188
rect 17224 42900 17276 42906
rect 17144 42860 17224 42888
rect 16396 42842 16448 42848
rect 17224 42842 17276 42848
rect 16304 42152 16356 42158
rect 16304 42094 16356 42100
rect 16302 41848 16358 41857
rect 16302 41783 16358 41792
rect 16316 41614 16344 41783
rect 16304 41608 16356 41614
rect 16304 41550 16356 41556
rect 16408 41206 16436 42842
rect 17132 42764 17184 42770
rect 17132 42706 17184 42712
rect 17040 42628 17092 42634
rect 17040 42570 17092 42576
rect 16544 42460 16852 42469
rect 16544 42458 16550 42460
rect 16606 42458 16630 42460
rect 16686 42458 16710 42460
rect 16766 42458 16790 42460
rect 16846 42458 16852 42460
rect 16606 42406 16608 42458
rect 16788 42406 16790 42458
rect 16544 42404 16550 42406
rect 16606 42404 16630 42406
rect 16686 42404 16710 42406
rect 16766 42404 16790 42406
rect 16846 42404 16852 42406
rect 16544 42395 16852 42404
rect 16764 42220 16816 42226
rect 16764 42162 16816 42168
rect 16776 41818 16804 42162
rect 16856 42016 16908 42022
rect 16856 41958 16908 41964
rect 16948 42016 17000 42022
rect 16948 41958 17000 41964
rect 16764 41812 16816 41818
rect 16764 41754 16816 41760
rect 16868 41721 16896 41958
rect 16960 41818 16988 41958
rect 16948 41812 17000 41818
rect 16948 41754 17000 41760
rect 16854 41712 16910 41721
rect 16854 41647 16910 41656
rect 16672 41608 16724 41614
rect 16670 41576 16672 41585
rect 16948 41608 17000 41614
rect 16724 41576 16726 41585
rect 16670 41511 16726 41520
rect 16854 41576 16910 41585
rect 16948 41550 17000 41556
rect 17052 41562 17080 42570
rect 17144 41750 17172 42706
rect 17328 42362 17356 43182
rect 17420 42362 17448 43862
rect 17512 42906 17540 44540
rect 17696 43178 17724 44540
rect 17776 43852 17828 43858
rect 17776 43794 17828 43800
rect 17788 43450 17816 43794
rect 17776 43444 17828 43450
rect 17776 43386 17828 43392
rect 17776 43308 17828 43314
rect 17776 43250 17828 43256
rect 17684 43172 17736 43178
rect 17684 43114 17736 43120
rect 17500 42900 17552 42906
rect 17500 42842 17552 42848
rect 17788 42684 17816 43250
rect 17880 42786 17908 44540
rect 18064 43296 18092 44540
rect 18064 43268 18184 43296
rect 17880 42770 18092 42786
rect 17880 42764 18104 42770
rect 17880 42758 18052 42764
rect 18052 42706 18104 42712
rect 17788 42656 17908 42684
rect 17500 42628 17552 42634
rect 17500 42570 17552 42576
rect 17592 42628 17644 42634
rect 17592 42570 17644 42576
rect 17512 42537 17540 42570
rect 17498 42528 17554 42537
rect 17498 42463 17554 42472
rect 17316 42356 17368 42362
rect 17316 42298 17368 42304
rect 17408 42356 17460 42362
rect 17408 42298 17460 42304
rect 17500 42220 17552 42226
rect 17500 42162 17552 42168
rect 17408 42152 17460 42158
rect 17408 42094 17460 42100
rect 17132 41744 17184 41750
rect 17132 41686 17184 41692
rect 17420 41682 17448 42094
rect 17316 41676 17368 41682
rect 17316 41618 17368 41624
rect 17408 41676 17460 41682
rect 17408 41618 17460 41624
rect 17224 41608 17276 41614
rect 16854 41511 16910 41520
rect 16868 41478 16896 41511
rect 16856 41472 16908 41478
rect 16856 41414 16908 41420
rect 16544 41372 16852 41381
rect 16544 41370 16550 41372
rect 16606 41370 16630 41372
rect 16686 41370 16710 41372
rect 16766 41370 16790 41372
rect 16846 41370 16852 41372
rect 16606 41318 16608 41370
rect 16788 41318 16790 41370
rect 16544 41316 16550 41318
rect 16606 41316 16630 41318
rect 16686 41316 16710 41318
rect 16766 41316 16790 41318
rect 16846 41316 16852 41318
rect 16544 41307 16852 41316
rect 16960 41256 16988 41550
rect 17052 41534 17172 41562
rect 17224 41550 17276 41556
rect 17040 41472 17092 41478
rect 17040 41414 17092 41420
rect 16776 41228 16988 41256
rect 16396 41200 16448 41206
rect 16396 41142 16448 41148
rect 16580 41064 16632 41070
rect 16578 41032 16580 41041
rect 16632 41032 16634 41041
rect 16578 40967 16634 40976
rect 16776 40934 16804 41228
rect 17052 41177 17080 41414
rect 17038 41168 17094 41177
rect 16856 41132 16908 41138
rect 17038 41103 17094 41112
rect 16856 41074 16908 41080
rect 16764 40928 16816 40934
rect 16764 40870 16816 40876
rect 16212 40724 16264 40730
rect 16212 40666 16264 40672
rect 16868 40474 16896 41074
rect 17144 40662 17172 41534
rect 17236 41002 17264 41550
rect 17328 41274 17356 41618
rect 17408 41540 17460 41546
rect 17408 41482 17460 41488
rect 17316 41268 17368 41274
rect 17316 41210 17368 41216
rect 17316 41132 17368 41138
rect 17316 41074 17368 41080
rect 17224 40996 17276 41002
rect 17224 40938 17276 40944
rect 17132 40656 17184 40662
rect 17132 40598 17184 40604
rect 16868 40446 16988 40474
rect 16544 40284 16852 40293
rect 16544 40282 16550 40284
rect 16606 40282 16630 40284
rect 16686 40282 16710 40284
rect 16766 40282 16790 40284
rect 16846 40282 16852 40284
rect 16606 40230 16608 40282
rect 16788 40230 16790 40282
rect 16544 40228 16550 40230
rect 16606 40228 16630 40230
rect 16686 40228 16710 40230
rect 16766 40228 16790 40230
rect 16846 40228 16852 40230
rect 16544 40219 16852 40228
rect 16304 40044 16356 40050
rect 16304 39986 16356 39992
rect 16212 39840 16264 39846
rect 16212 39782 16264 39788
rect 16120 39432 16172 39438
rect 16120 39374 16172 39380
rect 16132 39098 16160 39374
rect 16120 39092 16172 39098
rect 16120 39034 16172 39040
rect 16224 38894 16252 39782
rect 16316 39642 16344 39986
rect 16304 39636 16356 39642
rect 16304 39578 16356 39584
rect 16544 39196 16852 39205
rect 16544 39194 16550 39196
rect 16606 39194 16630 39196
rect 16686 39194 16710 39196
rect 16766 39194 16790 39196
rect 16846 39194 16852 39196
rect 16606 39142 16608 39194
rect 16788 39142 16790 39194
rect 16544 39140 16550 39142
rect 16606 39140 16630 39142
rect 16686 39140 16710 39142
rect 16766 39140 16790 39142
rect 16846 39140 16852 39142
rect 16544 39131 16852 39140
rect 16486 38992 16542 39001
rect 16408 38950 16486 38978
rect 16212 38888 16264 38894
rect 16212 38830 16264 38836
rect 16212 38752 16264 38758
rect 16212 38694 16264 38700
rect 16028 38548 16080 38554
rect 16028 38490 16080 38496
rect 16028 38412 16080 38418
rect 16028 38354 16080 38360
rect 16040 36242 16068 38354
rect 16120 37120 16172 37126
rect 16120 37062 16172 37068
rect 16132 36922 16160 37062
rect 16120 36916 16172 36922
rect 16120 36858 16172 36864
rect 16224 36802 16252 38694
rect 16408 36922 16436 38950
rect 16486 38927 16542 38936
rect 16544 38108 16852 38117
rect 16544 38106 16550 38108
rect 16606 38106 16630 38108
rect 16686 38106 16710 38108
rect 16766 38106 16790 38108
rect 16846 38106 16852 38108
rect 16606 38054 16608 38106
rect 16788 38054 16790 38106
rect 16544 38052 16550 38054
rect 16606 38052 16630 38054
rect 16686 38052 16710 38054
rect 16766 38052 16790 38054
rect 16846 38052 16852 38054
rect 16544 38043 16852 38052
rect 16960 37398 16988 40446
rect 17224 40384 17276 40390
rect 17224 40326 17276 40332
rect 17236 40225 17264 40326
rect 17222 40216 17278 40225
rect 17222 40151 17278 40160
rect 17040 39296 17092 39302
rect 17040 39238 17092 39244
rect 17052 38962 17080 39238
rect 17040 38956 17092 38962
rect 17040 38898 17092 38904
rect 16948 37392 17000 37398
rect 16948 37334 17000 37340
rect 17052 37274 17080 38898
rect 17222 38720 17278 38729
rect 16960 37246 17080 37274
rect 17144 38678 17222 38706
rect 16544 37020 16852 37029
rect 16544 37018 16550 37020
rect 16606 37018 16630 37020
rect 16686 37018 16710 37020
rect 16766 37018 16790 37020
rect 16846 37018 16852 37020
rect 16606 36966 16608 37018
rect 16788 36966 16790 37018
rect 16544 36964 16550 36966
rect 16606 36964 16630 36966
rect 16686 36964 16710 36966
rect 16766 36964 16790 36966
rect 16846 36964 16852 36966
rect 16544 36955 16852 36964
rect 16396 36916 16448 36922
rect 16396 36858 16448 36864
rect 16580 36916 16632 36922
rect 16580 36858 16632 36864
rect 16132 36774 16252 36802
rect 16304 36780 16356 36786
rect 16028 36236 16080 36242
rect 16028 36178 16080 36184
rect 16028 35692 16080 35698
rect 16028 35634 16080 35640
rect 16040 34746 16068 35634
rect 16028 34740 16080 34746
rect 16028 34682 16080 34688
rect 15948 34598 16068 34626
rect 15936 33856 15988 33862
rect 15842 33824 15898 33833
rect 15936 33798 15988 33804
rect 15842 33759 15898 33768
rect 15844 33516 15896 33522
rect 15844 33458 15896 33464
rect 15660 33312 15712 33318
rect 15660 33254 15712 33260
rect 15672 33114 15700 33254
rect 15660 33108 15712 33114
rect 15660 33050 15712 33056
rect 15752 33108 15804 33114
rect 15752 33050 15804 33056
rect 15764 33017 15792 33050
rect 15750 33008 15806 33017
rect 15750 32943 15806 32952
rect 15660 32292 15712 32298
rect 15660 32234 15712 32240
rect 15672 31890 15700 32234
rect 15752 32224 15804 32230
rect 15752 32166 15804 32172
rect 15660 31884 15712 31890
rect 15660 31826 15712 31832
rect 15764 31754 15792 32166
rect 15672 31726 15792 31754
rect 15568 31680 15620 31686
rect 15568 31622 15620 31628
rect 15488 31470 15608 31498
rect 15476 31136 15528 31142
rect 15476 31078 15528 31084
rect 15488 29714 15516 31078
rect 15476 29708 15528 29714
rect 15476 29650 15528 29656
rect 15474 27432 15530 27441
rect 15474 27367 15530 27376
rect 15488 27334 15516 27367
rect 15476 27328 15528 27334
rect 15476 27270 15528 27276
rect 15384 25288 15436 25294
rect 15384 25230 15436 25236
rect 15120 24942 15332 24970
rect 15028 24840 15148 24868
rect 14924 24812 14976 24818
rect 14924 24754 14976 24760
rect 14922 24712 14978 24721
rect 14922 24647 14978 24656
rect 14832 24404 14884 24410
rect 14832 24346 14884 24352
rect 14936 24290 14964 24647
rect 15016 24608 15068 24614
rect 15016 24550 15068 24556
rect 14844 24262 14964 24290
rect 14844 24138 14872 24262
rect 14924 24200 14976 24206
rect 14924 24142 14976 24148
rect 14832 24132 14884 24138
rect 14832 24074 14884 24080
rect 14936 23866 14964 24142
rect 14924 23860 14976 23866
rect 14924 23802 14976 23808
rect 14832 23656 14884 23662
rect 15028 23644 15056 24550
rect 14884 23616 15056 23644
rect 14832 23598 14884 23604
rect 14740 23316 14792 23322
rect 14740 23258 14792 23264
rect 14832 23112 14884 23118
rect 14832 23054 14884 23060
rect 14844 22778 14872 23054
rect 14832 22772 14884 22778
rect 14832 22714 14884 22720
rect 14740 22568 14792 22574
rect 14740 22510 14792 22516
rect 14752 22234 14780 22510
rect 14830 22264 14886 22273
rect 14740 22228 14792 22234
rect 14830 22199 14886 22208
rect 14740 22170 14792 22176
rect 14648 19916 14700 19922
rect 14648 19858 14700 19864
rect 14648 19372 14700 19378
rect 14648 19314 14700 19320
rect 14660 18902 14688 19314
rect 14648 18896 14700 18902
rect 14646 18864 14648 18873
rect 14700 18864 14702 18873
rect 14646 18799 14702 18808
rect 14752 18086 14780 22170
rect 14844 20074 14872 22199
rect 14936 22114 14964 23616
rect 15120 23066 15148 24840
rect 15304 24206 15332 24942
rect 15200 24200 15252 24206
rect 15200 24142 15252 24148
rect 15292 24200 15344 24206
rect 15292 24142 15344 24148
rect 15212 23798 15240 24142
rect 15200 23792 15252 23798
rect 15200 23734 15252 23740
rect 15212 23186 15240 23734
rect 15200 23180 15252 23186
rect 15200 23122 15252 23128
rect 15304 23118 15332 24142
rect 15396 23361 15424 25230
rect 15488 24410 15516 27270
rect 15476 24404 15528 24410
rect 15476 24346 15528 24352
rect 15382 23352 15438 23361
rect 15382 23287 15438 23296
rect 15474 23216 15530 23225
rect 15474 23151 15530 23160
rect 15292 23112 15344 23118
rect 15120 23038 15240 23066
rect 15292 23054 15344 23060
rect 15382 23080 15438 23089
rect 15014 22536 15070 22545
rect 15014 22471 15070 22480
rect 15028 22438 15056 22471
rect 15016 22432 15068 22438
rect 15016 22374 15068 22380
rect 15212 22234 15240 23038
rect 15382 23015 15438 23024
rect 15200 22228 15252 22234
rect 15200 22170 15252 22176
rect 14936 22086 15332 22114
rect 15396 22098 15424 23015
rect 15200 22024 15252 22030
rect 15200 21966 15252 21972
rect 15212 21690 15240 21966
rect 15200 21684 15252 21690
rect 15200 21626 15252 21632
rect 15200 21548 15252 21554
rect 15200 21490 15252 21496
rect 15016 21072 15068 21078
rect 15016 21014 15068 21020
rect 14924 20800 14976 20806
rect 14924 20742 14976 20748
rect 14936 20398 14964 20742
rect 14924 20392 14976 20398
rect 14924 20334 14976 20340
rect 14844 20046 14964 20074
rect 14832 19916 14884 19922
rect 14832 19858 14884 19864
rect 14740 18080 14792 18086
rect 14740 18022 14792 18028
rect 14738 17640 14794 17649
rect 14660 17598 14738 17626
rect 14660 16658 14688 17598
rect 14738 17575 14794 17584
rect 14844 17542 14872 19858
rect 14832 17536 14884 17542
rect 14832 17478 14884 17484
rect 14740 17128 14792 17134
rect 14738 17096 14740 17105
rect 14792 17096 14794 17105
rect 14738 17031 14794 17040
rect 14738 16688 14794 16697
rect 14648 16652 14700 16658
rect 14738 16623 14740 16632
rect 14648 16594 14700 16600
rect 14792 16623 14794 16632
rect 14740 16594 14792 16600
rect 14648 16040 14700 16046
rect 14648 15982 14700 15988
rect 14556 15564 14608 15570
rect 14556 15506 14608 15512
rect 13832 15150 13952 15178
rect 14292 15286 14504 15314
rect 13832 13258 13860 15150
rect 14292 14958 14320 15286
rect 14280 14952 14332 14958
rect 14280 14894 14332 14900
rect 13945 14716 14253 14725
rect 13945 14714 13951 14716
rect 14007 14714 14031 14716
rect 14087 14714 14111 14716
rect 14167 14714 14191 14716
rect 14247 14714 14253 14716
rect 14007 14662 14009 14714
rect 14189 14662 14191 14714
rect 13945 14660 13951 14662
rect 14007 14660 14031 14662
rect 14087 14660 14111 14662
rect 14167 14660 14191 14662
rect 14247 14660 14253 14662
rect 13945 14651 14253 14660
rect 14292 14498 14320 14894
rect 14372 14884 14424 14890
rect 14372 14826 14424 14832
rect 14384 14618 14412 14826
rect 14372 14612 14424 14618
rect 14372 14554 14424 14560
rect 14292 14470 14412 14498
rect 14096 14408 14148 14414
rect 14096 14350 14148 14356
rect 14108 14278 14136 14350
rect 14096 14272 14148 14278
rect 14096 14214 14148 14220
rect 14280 14000 14332 14006
rect 14280 13942 14332 13948
rect 13945 13628 14253 13637
rect 13945 13626 13951 13628
rect 14007 13626 14031 13628
rect 14087 13626 14111 13628
rect 14167 13626 14191 13628
rect 14247 13626 14253 13628
rect 14007 13574 14009 13626
rect 14189 13574 14191 13626
rect 13945 13572 13951 13574
rect 14007 13572 14031 13574
rect 14087 13572 14111 13574
rect 14167 13572 14191 13574
rect 14247 13572 14253 13574
rect 13945 13563 14253 13572
rect 14188 13388 14240 13394
rect 14292 13376 14320 13942
rect 14240 13348 14320 13376
rect 14188 13330 14240 13336
rect 13820 13252 13872 13258
rect 13820 13194 13872 13200
rect 13728 12980 13780 12986
rect 13728 12922 13780 12928
rect 13818 12880 13874 12889
rect 13818 12815 13820 12824
rect 13872 12815 13874 12824
rect 13820 12786 13872 12792
rect 13728 12436 13780 12442
rect 13728 12378 13780 12384
rect 13636 12368 13688 12374
rect 13636 12310 13688 12316
rect 13542 11792 13598 11801
rect 13648 11762 13676 12310
rect 13542 11727 13544 11736
rect 13596 11727 13598 11736
rect 13636 11756 13688 11762
rect 13544 11698 13596 11704
rect 13636 11698 13688 11704
rect 13740 11642 13768 12378
rect 13832 12238 13860 12786
rect 13945 12540 14253 12549
rect 13945 12538 13951 12540
rect 14007 12538 14031 12540
rect 14087 12538 14111 12540
rect 14167 12538 14191 12540
rect 14247 12538 14253 12540
rect 14007 12486 14009 12538
rect 14189 12486 14191 12538
rect 13945 12484 13951 12486
rect 14007 12484 14031 12486
rect 14087 12484 14111 12486
rect 14167 12484 14191 12486
rect 14247 12484 14253 12486
rect 13945 12475 14253 12484
rect 13820 12232 13872 12238
rect 13820 12174 13872 12180
rect 13910 12200 13966 12209
rect 13910 12135 13966 12144
rect 13556 11614 13768 11642
rect 13556 11286 13584 11614
rect 13636 11552 13688 11558
rect 13924 11540 13952 12135
rect 14292 11762 14320 13348
rect 14280 11756 14332 11762
rect 14280 11698 14332 11704
rect 13636 11494 13688 11500
rect 13832 11512 13952 11540
rect 13544 11280 13596 11286
rect 13544 11222 13596 11228
rect 13452 11212 13504 11218
rect 13452 11154 13504 11160
rect 13544 11076 13596 11082
rect 13544 11018 13596 11024
rect 13452 11008 13504 11014
rect 13452 10950 13504 10956
rect 13464 10810 13492 10950
rect 13452 10804 13504 10810
rect 13452 10746 13504 10752
rect 13556 10674 13584 11018
rect 13648 10674 13676 11494
rect 13832 11200 13860 11512
rect 13945 11452 14253 11461
rect 13945 11450 13951 11452
rect 14007 11450 14031 11452
rect 14087 11450 14111 11452
rect 14167 11450 14191 11452
rect 14247 11450 14253 11452
rect 14007 11398 14009 11450
rect 14189 11398 14191 11450
rect 13945 11396 13951 11398
rect 14007 11396 14031 11398
rect 14087 11396 14111 11398
rect 14167 11396 14191 11398
rect 14247 11396 14253 11398
rect 13945 11387 14253 11396
rect 13740 11172 13860 11200
rect 14096 11212 14148 11218
rect 13544 10668 13596 10674
rect 13544 10610 13596 10616
rect 13636 10668 13688 10674
rect 13636 10610 13688 10616
rect 13360 10600 13412 10606
rect 13740 10554 13768 11172
rect 14096 11154 14148 11160
rect 13910 11112 13966 11121
rect 13360 10542 13412 10548
rect 13648 10526 13768 10554
rect 13832 11070 13910 11098
rect 13542 10160 13598 10169
rect 13542 10095 13544 10104
rect 13596 10095 13598 10104
rect 13544 10066 13596 10072
rect 13358 9752 13414 9761
rect 13268 9716 13320 9722
rect 13358 9687 13414 9696
rect 13268 9658 13320 9664
rect 13268 9580 13320 9586
rect 13268 9522 13320 9528
rect 13280 8634 13308 9522
rect 13268 8628 13320 8634
rect 13268 8570 13320 8576
rect 13268 8492 13320 8498
rect 13268 8434 13320 8440
rect 13280 8401 13308 8434
rect 13266 8392 13322 8401
rect 13266 8327 13322 8336
rect 13280 7410 13308 8327
rect 13268 7404 13320 7410
rect 13268 7346 13320 7352
rect 13280 6730 13308 7346
rect 13268 6724 13320 6730
rect 13268 6666 13320 6672
rect 13268 6452 13320 6458
rect 13268 6394 13320 6400
rect 13174 5264 13230 5273
rect 13174 5199 13230 5208
rect 13084 4208 13136 4214
rect 13084 4150 13136 4156
rect 12992 3936 13044 3942
rect 12992 3878 13044 3884
rect 12900 3392 12952 3398
rect 12900 3334 12952 3340
rect 12072 3052 12124 3058
rect 12072 2994 12124 3000
rect 12808 3052 12860 3058
rect 12808 2994 12860 3000
rect 11888 2916 11940 2922
rect 11888 2858 11940 2864
rect 11664 2400 11744 2428
rect 11612 2382 11664 2388
rect 11244 2304 11296 2310
rect 11244 2246 11296 2252
rect 11704 2304 11756 2310
rect 11704 2246 11756 2252
rect 11796 2304 11848 2310
rect 11796 2246 11848 2252
rect 11256 2038 11284 2246
rect 11346 2204 11654 2213
rect 11346 2202 11352 2204
rect 11408 2202 11432 2204
rect 11488 2202 11512 2204
rect 11568 2202 11592 2204
rect 11648 2202 11654 2204
rect 11408 2150 11410 2202
rect 11590 2150 11592 2202
rect 11346 2148 11352 2150
rect 11408 2148 11432 2150
rect 11488 2148 11512 2150
rect 11568 2148 11592 2150
rect 11648 2148 11654 2150
rect 11346 2139 11654 2148
rect 11244 2032 11296 2038
rect 11244 1974 11296 1980
rect 11060 1760 11112 1766
rect 11060 1702 11112 1708
rect 11244 1760 11296 1766
rect 11244 1702 11296 1708
rect 10968 1556 11020 1562
rect 10968 1498 11020 1504
rect 11072 1408 11100 1702
rect 10980 1380 11100 1408
rect 11152 1420 11204 1426
rect 10600 1352 10652 1358
rect 10600 1294 10652 1300
rect 10692 1284 10744 1290
rect 10692 1226 10744 1232
rect 10704 160 10732 1226
rect 9954 54 10088 82
rect 9770 -300 9826 54
rect 9954 -300 10010 54
rect 10138 -300 10194 160
rect 10322 -300 10378 160
rect 10506 -300 10562 160
rect 10690 -300 10746 160
rect 10874 82 10930 160
rect 10980 82 11008 1380
rect 11152 1362 11204 1368
rect 11060 1284 11112 1290
rect 11060 1226 11112 1232
rect 11072 160 11100 1226
rect 10874 54 11008 82
rect 10874 -300 10930 54
rect 11058 -300 11114 160
rect 11164 82 11192 1362
rect 11256 898 11284 1702
rect 11716 1494 11744 2246
rect 11704 1488 11756 1494
rect 11704 1430 11756 1436
rect 11704 1216 11756 1222
rect 11704 1158 11756 1164
rect 11346 1116 11654 1125
rect 11346 1114 11352 1116
rect 11408 1114 11432 1116
rect 11488 1114 11512 1116
rect 11568 1114 11592 1116
rect 11648 1114 11654 1116
rect 11408 1062 11410 1114
rect 11590 1062 11592 1114
rect 11346 1060 11352 1062
rect 11408 1060 11432 1062
rect 11488 1060 11512 1062
rect 11568 1060 11592 1062
rect 11648 1060 11654 1062
rect 11346 1051 11654 1060
rect 11256 870 11652 898
rect 11520 808 11572 814
rect 11520 750 11572 756
rect 11242 82 11298 160
rect 11164 54 11298 82
rect 11242 -300 11298 54
rect 11426 82 11482 160
rect 11532 82 11560 750
rect 11624 160 11652 870
rect 11426 54 11560 82
rect 11426 -300 11482 54
rect 11610 -300 11666 160
rect 11716 82 11744 1158
rect 11808 950 11836 2246
rect 11796 944 11848 950
rect 11796 886 11848 892
rect 11900 814 11928 2858
rect 12072 2848 12124 2854
rect 12072 2790 12124 2796
rect 12624 2848 12676 2854
rect 12676 2808 12848 2836
rect 12624 2790 12676 2796
rect 11980 2304 12032 2310
rect 11980 2246 12032 2252
rect 11992 2009 12020 2246
rect 11978 2000 12034 2009
rect 11978 1935 12034 1944
rect 11980 1760 12032 1766
rect 11980 1702 12032 1708
rect 11888 808 11940 814
rect 11888 750 11940 756
rect 11992 160 12020 1702
rect 12084 1358 12112 2790
rect 12440 2304 12492 2310
rect 12440 2246 12492 2252
rect 12348 1556 12400 1562
rect 12348 1498 12400 1504
rect 12072 1352 12124 1358
rect 12072 1294 12124 1300
rect 12072 1216 12124 1222
rect 12124 1176 12204 1204
rect 12072 1158 12124 1164
rect 12176 160 12204 1176
rect 12360 160 12388 1498
rect 12452 1426 12480 2246
rect 12714 2000 12770 2009
rect 12714 1935 12716 1944
rect 12768 1935 12770 1944
rect 12716 1906 12768 1912
rect 12440 1420 12492 1426
rect 12440 1362 12492 1368
rect 12820 1358 12848 2808
rect 12912 1970 12940 3334
rect 13004 2106 13032 3878
rect 13176 3664 13228 3670
rect 13176 3606 13228 3612
rect 12992 2100 13044 2106
rect 12992 2042 13044 2048
rect 12900 1964 12952 1970
rect 12900 1906 12952 1912
rect 13084 1760 13136 1766
rect 13084 1702 13136 1708
rect 12808 1352 12860 1358
rect 12808 1294 12860 1300
rect 12716 1284 12768 1290
rect 12716 1226 12768 1232
rect 12532 1216 12584 1222
rect 12532 1158 12584 1164
rect 12544 160 12572 1158
rect 12728 160 12756 1226
rect 12900 672 12952 678
rect 12900 614 12952 620
rect 12912 160 12940 614
rect 13096 160 13124 1702
rect 13188 1358 13216 3606
rect 13280 2972 13308 6394
rect 13372 3126 13400 9687
rect 13452 9376 13504 9382
rect 13450 9344 13452 9353
rect 13504 9344 13506 9353
rect 13450 9279 13506 9288
rect 13452 8832 13504 8838
rect 13452 8774 13504 8780
rect 13464 3534 13492 8774
rect 13544 8016 13596 8022
rect 13544 7958 13596 7964
rect 13556 6458 13584 7958
rect 13544 6452 13596 6458
rect 13544 6394 13596 6400
rect 13648 6338 13676 10526
rect 13728 10464 13780 10470
rect 13728 10406 13780 10412
rect 13740 7886 13768 10406
rect 13832 9654 13860 11070
rect 13910 11047 13966 11056
rect 14108 10810 14136 11154
rect 14096 10804 14148 10810
rect 14096 10746 14148 10752
rect 14278 10704 14334 10713
rect 14278 10639 14334 10648
rect 13945 10364 14253 10373
rect 13945 10362 13951 10364
rect 14007 10362 14031 10364
rect 14087 10362 14111 10364
rect 14167 10362 14191 10364
rect 14247 10362 14253 10364
rect 14007 10310 14009 10362
rect 14189 10310 14191 10362
rect 13945 10308 13951 10310
rect 14007 10308 14031 10310
rect 14087 10308 14111 10310
rect 14167 10308 14191 10310
rect 14247 10308 14253 10310
rect 13945 10299 14253 10308
rect 14292 10010 14320 10639
rect 14384 10112 14412 14470
rect 14568 14346 14596 15506
rect 14556 14340 14608 14346
rect 14556 14282 14608 14288
rect 14464 14068 14516 14074
rect 14464 14010 14516 14016
rect 14476 11830 14504 14010
rect 14568 12850 14596 14282
rect 14556 12844 14608 12850
rect 14556 12786 14608 12792
rect 14660 12730 14688 15982
rect 14752 14074 14780 16594
rect 14844 14958 14872 17478
rect 14832 14952 14884 14958
rect 14832 14894 14884 14900
rect 14844 14822 14872 14894
rect 14832 14816 14884 14822
rect 14832 14758 14884 14764
rect 14740 14068 14792 14074
rect 14740 14010 14792 14016
rect 14740 13456 14792 13462
rect 14740 13398 14792 13404
rect 14752 12986 14780 13398
rect 14936 13308 14964 20046
rect 15028 19904 15056 21014
rect 15212 20466 15240 21490
rect 15304 20913 15332 22086
rect 15384 22092 15436 22098
rect 15384 22034 15436 22040
rect 15396 21418 15424 22034
rect 15384 21412 15436 21418
rect 15384 21354 15436 21360
rect 15290 20904 15346 20913
rect 15290 20839 15346 20848
rect 15200 20460 15252 20466
rect 15200 20402 15252 20408
rect 15106 19952 15162 19961
rect 15028 19896 15106 19904
rect 15028 19876 15108 19896
rect 15160 19887 15162 19896
rect 15108 19858 15160 19864
rect 15198 19680 15254 19689
rect 15198 19615 15254 19624
rect 15212 19310 15240 19615
rect 15200 19304 15252 19310
rect 15200 19246 15252 19252
rect 15108 19236 15160 19242
rect 15108 19178 15160 19184
rect 15120 18834 15148 19178
rect 15212 18970 15240 19246
rect 15200 18964 15252 18970
rect 15200 18906 15252 18912
rect 15108 18828 15160 18834
rect 15108 18770 15160 18776
rect 15200 18760 15252 18766
rect 15200 18702 15252 18708
rect 15212 18154 15240 18702
rect 15304 18204 15332 20839
rect 15384 20256 15436 20262
rect 15384 20198 15436 20204
rect 15396 20058 15424 20198
rect 15384 20052 15436 20058
rect 15384 19994 15436 20000
rect 15384 19372 15436 19378
rect 15384 19314 15436 19320
rect 15396 18970 15424 19314
rect 15384 18964 15436 18970
rect 15384 18906 15436 18912
rect 15384 18216 15436 18222
rect 15304 18176 15384 18204
rect 15384 18158 15436 18164
rect 15200 18148 15252 18154
rect 15200 18090 15252 18096
rect 15292 18080 15344 18086
rect 15292 18022 15344 18028
rect 15304 17746 15332 18022
rect 15292 17740 15344 17746
rect 15292 17682 15344 17688
rect 15108 17672 15160 17678
rect 15160 17632 15240 17660
rect 15108 17614 15160 17620
rect 15106 17368 15162 17377
rect 15016 17332 15068 17338
rect 15106 17303 15162 17312
rect 15016 17274 15068 17280
rect 15028 17241 15056 17274
rect 15014 17232 15070 17241
rect 15014 17167 15070 17176
rect 15016 13320 15068 13326
rect 14936 13280 15016 13308
rect 14740 12980 14792 12986
rect 14740 12922 14792 12928
rect 14568 12702 14688 12730
rect 14464 11824 14516 11830
rect 14464 11766 14516 11772
rect 14568 10554 14596 12702
rect 14936 12442 14964 13280
rect 15016 13262 15068 13268
rect 15016 12844 15068 12850
rect 15016 12786 15068 12792
rect 14924 12436 14976 12442
rect 14924 12378 14976 12384
rect 15028 12322 15056 12786
rect 14740 12300 14792 12306
rect 14740 12242 14792 12248
rect 14936 12294 15056 12322
rect 14648 12096 14700 12102
rect 14648 12038 14700 12044
rect 14660 10810 14688 12038
rect 14648 10804 14700 10810
rect 14648 10746 14700 10752
rect 14752 10674 14780 12242
rect 14832 11824 14884 11830
rect 14832 11766 14884 11772
rect 14740 10668 14792 10674
rect 14740 10610 14792 10616
rect 14568 10526 14780 10554
rect 14556 10260 14608 10266
rect 14556 10202 14608 10208
rect 14568 10169 14596 10202
rect 14554 10160 14610 10169
rect 14384 10084 14504 10112
rect 14554 10095 14610 10104
rect 13924 9982 14320 10010
rect 14372 9988 14424 9994
rect 13820 9648 13872 9654
rect 13820 9590 13872 9596
rect 13924 9364 13952 9982
rect 14372 9930 14424 9936
rect 14280 9920 14332 9926
rect 14280 9862 14332 9868
rect 14292 9654 14320 9862
rect 14280 9648 14332 9654
rect 14280 9590 14332 9596
rect 13832 9336 13952 9364
rect 13728 7880 13780 7886
rect 13728 7822 13780 7828
rect 13832 7834 13860 9336
rect 13945 9276 14253 9285
rect 13945 9274 13951 9276
rect 14007 9274 14031 9276
rect 14087 9274 14111 9276
rect 14167 9274 14191 9276
rect 14247 9274 14253 9276
rect 14007 9222 14009 9274
rect 14189 9222 14191 9274
rect 13945 9220 13951 9222
rect 14007 9220 14031 9222
rect 14087 9220 14111 9222
rect 14167 9220 14191 9222
rect 14247 9220 14253 9222
rect 13945 9211 14253 9220
rect 14186 8664 14242 8673
rect 14186 8599 14242 8608
rect 14200 8498 14228 8599
rect 14188 8492 14240 8498
rect 14188 8434 14240 8440
rect 14292 8294 14320 9590
rect 14384 8294 14412 9930
rect 14476 9674 14504 10084
rect 14646 10024 14702 10033
rect 14646 9959 14702 9968
rect 14476 9646 14596 9674
rect 14568 9450 14596 9646
rect 14556 9444 14608 9450
rect 14556 9386 14608 9392
rect 14464 8492 14516 8498
rect 14464 8434 14516 8440
rect 14280 8288 14332 8294
rect 14280 8230 14332 8236
rect 14372 8288 14424 8294
rect 14372 8230 14424 8236
rect 13945 8188 14253 8197
rect 13945 8186 13951 8188
rect 14007 8186 14031 8188
rect 14087 8186 14111 8188
rect 14167 8186 14191 8188
rect 14247 8186 14253 8188
rect 14007 8134 14009 8186
rect 14189 8134 14191 8186
rect 13945 8132 13951 8134
rect 14007 8132 14031 8134
rect 14087 8132 14111 8134
rect 14167 8132 14191 8134
rect 14247 8132 14253 8134
rect 13945 8123 14253 8132
rect 14004 7880 14056 7886
rect 14002 7848 14004 7857
rect 14096 7880 14148 7886
rect 14056 7848 14058 7857
rect 13832 7806 13952 7834
rect 13820 7744 13872 7750
rect 13820 7686 13872 7692
rect 13728 6792 13780 6798
rect 13728 6734 13780 6740
rect 13740 6458 13768 6734
rect 13728 6452 13780 6458
rect 13728 6394 13780 6400
rect 13648 6310 13768 6338
rect 13544 5568 13596 5574
rect 13544 5510 13596 5516
rect 13452 3528 13504 3534
rect 13452 3470 13504 3476
rect 13452 3392 13504 3398
rect 13452 3334 13504 3340
rect 13360 3120 13412 3126
rect 13360 3062 13412 3068
rect 13280 2944 13400 2972
rect 13268 1556 13320 1562
rect 13268 1498 13320 1504
rect 13176 1352 13228 1358
rect 13176 1294 13228 1300
rect 13280 160 13308 1498
rect 13372 1358 13400 2944
rect 13464 2009 13492 3334
rect 13556 3074 13584 5510
rect 13634 4448 13690 4457
rect 13634 4383 13690 4392
rect 13648 3194 13676 4383
rect 13740 3754 13768 6310
rect 13832 4146 13860 7686
rect 13924 7274 13952 7806
rect 14148 7840 14320 7868
rect 14096 7822 14148 7828
rect 14002 7783 14058 7792
rect 14292 7392 14320 7840
rect 14292 7364 14412 7392
rect 13912 7268 13964 7274
rect 13912 7210 13964 7216
rect 14280 7268 14332 7274
rect 14280 7210 14332 7216
rect 13945 7100 14253 7109
rect 13945 7098 13951 7100
rect 14007 7098 14031 7100
rect 14087 7098 14111 7100
rect 14167 7098 14191 7100
rect 14247 7098 14253 7100
rect 14007 7046 14009 7098
rect 14189 7046 14191 7098
rect 13945 7044 13951 7046
rect 14007 7044 14031 7046
rect 14087 7044 14111 7046
rect 14167 7044 14191 7046
rect 14247 7044 14253 7046
rect 13945 7035 14253 7044
rect 14096 6792 14148 6798
rect 14096 6734 14148 6740
rect 14108 6390 14136 6734
rect 14292 6633 14320 7210
rect 14278 6624 14334 6633
rect 14278 6559 14334 6568
rect 14188 6452 14240 6458
rect 14188 6394 14240 6400
rect 14096 6384 14148 6390
rect 14096 6326 14148 6332
rect 14200 6186 14228 6394
rect 14384 6390 14412 7364
rect 14476 6798 14504 8434
rect 14568 7585 14596 9386
rect 14554 7576 14610 7585
rect 14554 7511 14610 7520
rect 14556 7404 14608 7410
rect 14556 7346 14608 7352
rect 14568 7002 14596 7346
rect 14556 6996 14608 7002
rect 14556 6938 14608 6944
rect 14464 6792 14516 6798
rect 14660 6746 14688 9959
rect 14752 9092 14780 10526
rect 14844 9654 14872 11766
rect 14936 11082 14964 12294
rect 15120 11914 15148 17303
rect 15212 16794 15240 17632
rect 15292 17536 15344 17542
rect 15292 17478 15344 17484
rect 15304 17338 15332 17478
rect 15292 17332 15344 17338
rect 15292 17274 15344 17280
rect 15292 16992 15344 16998
rect 15396 16980 15424 18158
rect 15344 16952 15424 16980
rect 15292 16934 15344 16940
rect 15290 16824 15346 16833
rect 15200 16788 15252 16794
rect 15290 16759 15346 16768
rect 15200 16730 15252 16736
rect 15304 16726 15332 16759
rect 15292 16720 15344 16726
rect 15292 16662 15344 16668
rect 15200 16652 15252 16658
rect 15200 16594 15252 16600
rect 15212 15502 15240 16594
rect 15292 16448 15344 16454
rect 15292 16390 15344 16396
rect 15384 16448 15436 16454
rect 15384 16390 15436 16396
rect 15200 15496 15252 15502
rect 15200 15438 15252 15444
rect 15200 14340 15252 14346
rect 15200 14282 15252 14288
rect 15212 14006 15240 14282
rect 15200 14000 15252 14006
rect 15200 13942 15252 13948
rect 15304 13410 15332 16390
rect 15396 16182 15424 16390
rect 15384 16176 15436 16182
rect 15384 16118 15436 16124
rect 15384 15564 15436 15570
rect 15384 15506 15436 15512
rect 15212 13382 15332 13410
rect 15212 12345 15240 13382
rect 15292 13320 15344 13326
rect 15292 13262 15344 13268
rect 15304 12986 15332 13262
rect 15292 12980 15344 12986
rect 15292 12922 15344 12928
rect 15290 12744 15346 12753
rect 15396 12730 15424 15506
rect 15346 12702 15424 12730
rect 15290 12679 15346 12688
rect 15198 12336 15254 12345
rect 15198 12271 15254 12280
rect 15120 11886 15240 11914
rect 15108 11756 15160 11762
rect 15028 11716 15108 11744
rect 14924 11076 14976 11082
rect 14924 11018 14976 11024
rect 15028 9994 15056 11716
rect 15108 11698 15160 11704
rect 15212 10690 15240 11886
rect 15304 11354 15332 12679
rect 15292 11348 15344 11354
rect 15292 11290 15344 11296
rect 15212 10662 15424 10690
rect 15292 10532 15344 10538
rect 15292 10474 15344 10480
rect 15108 10124 15160 10130
rect 15108 10066 15160 10072
rect 15016 9988 15068 9994
rect 15016 9930 15068 9936
rect 15028 9654 15056 9930
rect 14832 9648 14884 9654
rect 14832 9590 14884 9596
rect 15016 9648 15068 9654
rect 15016 9590 15068 9596
rect 15014 9344 15070 9353
rect 15014 9279 15070 9288
rect 14832 9104 14884 9110
rect 14752 9064 14832 9092
rect 14752 8673 14780 9064
rect 14832 9046 14884 9052
rect 14738 8664 14794 8673
rect 14738 8599 14794 8608
rect 14738 8392 14794 8401
rect 15028 8378 15056 9279
rect 15120 9178 15148 10066
rect 15304 9994 15332 10474
rect 15292 9988 15344 9994
rect 15292 9930 15344 9936
rect 15304 9654 15332 9930
rect 15292 9648 15344 9654
rect 15290 9616 15292 9625
rect 15344 9616 15346 9625
rect 15200 9580 15252 9586
rect 15290 9551 15346 9560
rect 15200 9522 15252 9528
rect 15212 9178 15240 9522
rect 15292 9512 15344 9518
rect 15292 9454 15344 9460
rect 15108 9172 15160 9178
rect 15108 9114 15160 9120
rect 15200 9172 15252 9178
rect 15200 9114 15252 9120
rect 15108 8900 15160 8906
rect 15108 8842 15160 8848
rect 14738 8327 14794 8336
rect 14936 8350 15056 8378
rect 14464 6734 14516 6740
rect 14568 6718 14688 6746
rect 14568 6474 14596 6718
rect 14648 6656 14700 6662
rect 14648 6598 14700 6604
rect 14476 6446 14596 6474
rect 14372 6384 14424 6390
rect 14372 6326 14424 6332
rect 14280 6248 14332 6254
rect 14280 6190 14332 6196
rect 14188 6180 14240 6186
rect 14188 6122 14240 6128
rect 13945 6012 14253 6021
rect 13945 6010 13951 6012
rect 14007 6010 14031 6012
rect 14087 6010 14111 6012
rect 14167 6010 14191 6012
rect 14247 6010 14253 6012
rect 14007 5958 14009 6010
rect 14189 5958 14191 6010
rect 13945 5956 13951 5958
rect 14007 5956 14031 5958
rect 14087 5956 14111 5958
rect 14167 5956 14191 5958
rect 14247 5956 14253 5958
rect 13945 5947 14253 5956
rect 14292 5234 14320 6190
rect 14280 5228 14332 5234
rect 14280 5170 14332 5176
rect 13945 4924 14253 4933
rect 13945 4922 13951 4924
rect 14007 4922 14031 4924
rect 14087 4922 14111 4924
rect 14167 4922 14191 4924
rect 14247 4922 14253 4924
rect 14007 4870 14009 4922
rect 14189 4870 14191 4922
rect 13945 4868 13951 4870
rect 14007 4868 14031 4870
rect 14087 4868 14111 4870
rect 14167 4868 14191 4870
rect 14247 4868 14253 4870
rect 13945 4859 14253 4868
rect 14292 4622 14320 5170
rect 14476 5030 14504 6446
rect 14556 6316 14608 6322
rect 14556 6258 14608 6264
rect 14568 6225 14596 6258
rect 14554 6216 14610 6225
rect 14554 6151 14610 6160
rect 14660 6118 14688 6598
rect 14648 6112 14700 6118
rect 14648 6054 14700 6060
rect 14660 5778 14688 6054
rect 14648 5772 14700 5778
rect 14648 5714 14700 5720
rect 14752 5574 14780 8327
rect 14830 8256 14886 8265
rect 14830 8191 14886 8200
rect 14740 5568 14792 5574
rect 14740 5510 14792 5516
rect 14554 5264 14610 5273
rect 14554 5199 14610 5208
rect 14464 5024 14516 5030
rect 14464 4966 14516 4972
rect 14280 4616 14332 4622
rect 14280 4558 14332 4564
rect 14464 4616 14516 4622
rect 14464 4558 14516 4564
rect 13820 4140 13872 4146
rect 13820 4082 13872 4088
rect 14372 4140 14424 4146
rect 14372 4082 14424 4088
rect 13945 3836 14253 3845
rect 13945 3834 13951 3836
rect 14007 3834 14031 3836
rect 14087 3834 14111 3836
rect 14167 3834 14191 3836
rect 14247 3834 14253 3836
rect 14007 3782 14009 3834
rect 14189 3782 14191 3834
rect 13945 3780 13951 3782
rect 14007 3780 14031 3782
rect 14087 3780 14111 3782
rect 14167 3780 14191 3782
rect 14247 3780 14253 3782
rect 13945 3771 14253 3780
rect 14384 3777 14412 4082
rect 14476 4078 14504 4558
rect 14464 4072 14516 4078
rect 14464 4014 14516 4020
rect 14568 3890 14596 5199
rect 14648 5024 14700 5030
rect 14648 4966 14700 4972
rect 14660 4282 14688 4966
rect 14740 4480 14792 4486
rect 14844 4468 14872 8191
rect 14936 7290 14964 8350
rect 15120 8022 15148 8842
rect 15304 8634 15332 9454
rect 15292 8628 15344 8634
rect 15292 8570 15344 8576
rect 15396 8514 15424 10662
rect 15212 8486 15424 8514
rect 15108 8016 15160 8022
rect 15108 7958 15160 7964
rect 15016 7744 15068 7750
rect 15016 7686 15068 7692
rect 15028 7410 15056 7686
rect 15016 7404 15068 7410
rect 15016 7346 15068 7352
rect 14936 7262 15056 7290
rect 14924 5704 14976 5710
rect 14924 5646 14976 5652
rect 14936 5370 14964 5646
rect 14924 5364 14976 5370
rect 14924 5306 14976 5312
rect 14922 4856 14978 4865
rect 14922 4791 14978 4800
rect 14792 4440 14872 4468
rect 14740 4422 14792 4428
rect 14648 4276 14700 4282
rect 14648 4218 14700 4224
rect 14832 4276 14884 4282
rect 14832 4218 14884 4224
rect 14738 4176 14794 4185
rect 14738 4111 14794 4120
rect 14476 3862 14596 3890
rect 14646 3904 14702 3913
rect 14370 3768 14426 3777
rect 13740 3726 13860 3754
rect 13728 3664 13780 3670
rect 13728 3606 13780 3612
rect 13636 3188 13688 3194
rect 13636 3130 13688 3136
rect 13556 3046 13676 3074
rect 13648 2922 13676 3046
rect 13636 2916 13688 2922
rect 13636 2858 13688 2864
rect 13636 2304 13688 2310
rect 13636 2246 13688 2252
rect 13648 2038 13676 2246
rect 13636 2032 13688 2038
rect 13450 2000 13506 2009
rect 13636 1974 13688 1980
rect 13450 1935 13506 1944
rect 13452 1760 13504 1766
rect 13452 1702 13504 1708
rect 13360 1352 13412 1358
rect 13360 1294 13412 1300
rect 13464 160 13492 1702
rect 13636 1488 13688 1494
rect 13636 1430 13688 1436
rect 13648 160 13676 1430
rect 13740 1340 13768 3606
rect 13832 3534 13860 3726
rect 14370 3703 14426 3712
rect 14094 3632 14150 3641
rect 14094 3567 14150 3576
rect 13820 3528 13872 3534
rect 13820 3470 13872 3476
rect 14108 3194 14136 3567
rect 14476 3534 14504 3862
rect 14646 3839 14702 3848
rect 14464 3528 14516 3534
rect 14464 3470 14516 3476
rect 14660 3466 14688 3839
rect 14752 3534 14780 4111
rect 14844 3534 14872 4218
rect 14936 4146 14964 4791
rect 15028 4162 15056 7262
rect 15106 6896 15162 6905
rect 15106 6831 15162 6840
rect 15120 5914 15148 6831
rect 15108 5908 15160 5914
rect 15108 5850 15160 5856
rect 15106 5808 15162 5817
rect 15106 5743 15162 5752
rect 15120 4282 15148 5743
rect 15212 4826 15240 8486
rect 15384 8424 15436 8430
rect 15384 8366 15436 8372
rect 15488 8378 15516 23151
rect 15580 23089 15608 31470
rect 15672 28218 15700 31726
rect 15856 30394 15884 33458
rect 15948 32978 15976 33798
rect 15936 32972 15988 32978
rect 15936 32914 15988 32920
rect 15936 32564 15988 32570
rect 15936 32506 15988 32512
rect 15948 31958 15976 32506
rect 15936 31952 15988 31958
rect 15936 31894 15988 31900
rect 16040 31754 16068 34598
rect 15948 31726 16068 31754
rect 15844 30388 15896 30394
rect 15844 30330 15896 30336
rect 15948 30138 15976 31726
rect 16132 31668 16160 36774
rect 16304 36722 16356 36728
rect 16396 36780 16448 36786
rect 16396 36722 16448 36728
rect 16488 36780 16540 36786
rect 16488 36722 16540 36728
rect 16212 36236 16264 36242
rect 16212 36178 16264 36184
rect 16224 35154 16252 36178
rect 16212 35148 16264 35154
rect 16212 35090 16264 35096
rect 16212 34944 16264 34950
rect 16212 34886 16264 34892
rect 16224 34746 16252 34886
rect 16212 34740 16264 34746
rect 16212 34682 16264 34688
rect 16316 34626 16344 36722
rect 16408 36378 16436 36722
rect 16500 36582 16528 36722
rect 16488 36576 16540 36582
rect 16488 36518 16540 36524
rect 16396 36372 16448 36378
rect 16396 36314 16448 36320
rect 16500 36174 16528 36518
rect 16592 36378 16620 36858
rect 16580 36372 16632 36378
rect 16580 36314 16632 36320
rect 16488 36168 16540 36174
rect 16488 36110 16540 36116
rect 16544 35932 16852 35941
rect 16544 35930 16550 35932
rect 16606 35930 16630 35932
rect 16686 35930 16710 35932
rect 16766 35930 16790 35932
rect 16846 35930 16852 35932
rect 16606 35878 16608 35930
rect 16788 35878 16790 35930
rect 16544 35876 16550 35878
rect 16606 35876 16630 35878
rect 16686 35876 16710 35878
rect 16766 35876 16790 35878
rect 16846 35876 16852 35878
rect 16544 35867 16852 35876
rect 16960 35086 16988 37246
rect 17040 35624 17092 35630
rect 17040 35566 17092 35572
rect 17052 35290 17080 35566
rect 17040 35284 17092 35290
rect 17040 35226 17092 35232
rect 16948 35080 17000 35086
rect 16948 35022 17000 35028
rect 16396 35012 16448 35018
rect 16396 34954 16448 34960
rect 16408 34746 16436 34954
rect 17040 34944 17092 34950
rect 17040 34886 17092 34892
rect 16544 34844 16852 34853
rect 16544 34842 16550 34844
rect 16606 34842 16630 34844
rect 16686 34842 16710 34844
rect 16766 34842 16790 34844
rect 16846 34842 16852 34844
rect 16606 34790 16608 34842
rect 16788 34790 16790 34842
rect 16544 34788 16550 34790
rect 16606 34788 16630 34790
rect 16686 34788 16710 34790
rect 16766 34788 16790 34790
rect 16846 34788 16852 34790
rect 16544 34779 16852 34788
rect 16396 34740 16448 34746
rect 16396 34682 16448 34688
rect 16316 34598 16436 34626
rect 17052 34610 17080 34886
rect 16212 34400 16264 34406
rect 16212 34342 16264 34348
rect 16224 32230 16252 34342
rect 16304 34060 16356 34066
rect 16304 34002 16356 34008
rect 16316 32978 16344 34002
rect 16304 32972 16356 32978
rect 16304 32914 16356 32920
rect 16212 32224 16264 32230
rect 16212 32166 16264 32172
rect 16224 31822 16252 32166
rect 16212 31816 16264 31822
rect 16212 31758 16264 31764
rect 16040 31640 16160 31668
rect 16040 30938 16068 31640
rect 16120 31476 16172 31482
rect 16120 31418 16172 31424
rect 16028 30932 16080 30938
rect 16028 30874 16080 30880
rect 16028 30592 16080 30598
rect 16028 30534 16080 30540
rect 16040 30326 16068 30534
rect 16028 30320 16080 30326
rect 16028 30262 16080 30268
rect 15764 30110 15976 30138
rect 15660 28212 15712 28218
rect 15660 28154 15712 28160
rect 15672 27062 15700 28154
rect 15764 27962 15792 30110
rect 15844 30048 15896 30054
rect 15844 29990 15896 29996
rect 15934 30016 15990 30025
rect 15856 29850 15884 29990
rect 15934 29951 15990 29960
rect 15844 29844 15896 29850
rect 15844 29786 15896 29792
rect 15948 29345 15976 29951
rect 15934 29336 15990 29345
rect 15934 29271 15990 29280
rect 15948 29170 15976 29271
rect 16028 29232 16080 29238
rect 16028 29174 16080 29180
rect 15936 29164 15988 29170
rect 15936 29106 15988 29112
rect 15844 28620 15896 28626
rect 15844 28562 15896 28568
rect 15856 28506 15884 28562
rect 16040 28558 16068 29174
rect 16028 28552 16080 28558
rect 15856 28478 15976 28506
rect 16028 28494 16080 28500
rect 15844 28416 15896 28422
rect 15844 28358 15896 28364
rect 15856 28150 15884 28358
rect 15948 28150 15976 28478
rect 15844 28144 15896 28150
rect 15844 28086 15896 28092
rect 15936 28144 15988 28150
rect 15936 28086 15988 28092
rect 15764 27934 15884 27962
rect 15660 27056 15712 27062
rect 15660 26998 15712 27004
rect 15660 26784 15712 26790
rect 15660 26726 15712 26732
rect 15752 26784 15804 26790
rect 15752 26726 15804 26732
rect 15672 26042 15700 26726
rect 15660 26036 15712 26042
rect 15660 25978 15712 25984
rect 15764 25906 15792 26726
rect 15856 26330 15884 27934
rect 15948 27402 15976 28086
rect 15936 27396 15988 27402
rect 15936 27338 15988 27344
rect 15934 26344 15990 26353
rect 15856 26302 15934 26330
rect 15934 26279 15990 26288
rect 15752 25900 15804 25906
rect 15752 25842 15804 25848
rect 15936 25696 15988 25702
rect 15936 25638 15988 25644
rect 15948 25401 15976 25638
rect 15934 25392 15990 25401
rect 15934 25327 15990 25336
rect 16040 25226 16068 28494
rect 16132 27130 16160 31418
rect 16316 31346 16344 32914
rect 16304 31340 16356 31346
rect 16304 31282 16356 31288
rect 16316 30734 16344 31282
rect 16304 30728 16356 30734
rect 16302 30696 16304 30705
rect 16356 30696 16358 30705
rect 16212 30660 16264 30666
rect 16302 30631 16358 30640
rect 16212 30602 16264 30608
rect 16224 29646 16252 30602
rect 16212 29640 16264 29646
rect 16212 29582 16264 29588
rect 16224 29306 16252 29582
rect 16212 29300 16264 29306
rect 16212 29242 16264 29248
rect 16316 29170 16344 30631
rect 16408 30138 16436 34598
rect 16948 34604 17000 34610
rect 16948 34546 17000 34552
rect 17040 34604 17092 34610
rect 17040 34546 17092 34552
rect 16960 33930 16988 34546
rect 16948 33924 17000 33930
rect 16948 33866 17000 33872
rect 16544 33756 16852 33765
rect 16544 33754 16550 33756
rect 16606 33754 16630 33756
rect 16686 33754 16710 33756
rect 16766 33754 16790 33756
rect 16846 33754 16852 33756
rect 16606 33702 16608 33754
rect 16788 33702 16790 33754
rect 16544 33700 16550 33702
rect 16606 33700 16630 33702
rect 16686 33700 16710 33702
rect 16766 33700 16790 33702
rect 16846 33700 16852 33702
rect 16544 33691 16852 33700
rect 16580 33584 16632 33590
rect 16580 33526 16632 33532
rect 16592 33386 16620 33526
rect 16764 33448 16816 33454
rect 16764 33390 16816 33396
rect 16580 33380 16632 33386
rect 16580 33322 16632 33328
rect 16776 32842 16804 33390
rect 16764 32836 16816 32842
rect 16764 32778 16816 32784
rect 16544 32668 16852 32677
rect 16544 32666 16550 32668
rect 16606 32666 16630 32668
rect 16686 32666 16710 32668
rect 16766 32666 16790 32668
rect 16846 32666 16852 32668
rect 16606 32614 16608 32666
rect 16788 32614 16790 32666
rect 16544 32612 16550 32614
rect 16606 32612 16630 32614
rect 16686 32612 16710 32614
rect 16766 32612 16790 32614
rect 16846 32612 16852 32614
rect 16544 32603 16852 32612
rect 16488 32224 16540 32230
rect 16488 32166 16540 32172
rect 16856 32224 16908 32230
rect 16856 32166 16908 32172
rect 16500 32026 16528 32166
rect 16488 32020 16540 32026
rect 16488 31962 16540 31968
rect 16868 31668 16896 32166
rect 16960 31822 16988 33866
rect 17052 32212 17080 34546
rect 17144 33658 17172 38678
rect 17222 38655 17278 38664
rect 17224 37256 17276 37262
rect 17224 37198 17276 37204
rect 17328 37210 17356 41074
rect 17420 40066 17448 41482
rect 17512 41070 17540 42162
rect 17604 41834 17632 42570
rect 17880 42514 17908 42656
rect 18052 42628 18104 42634
rect 18052 42570 18104 42576
rect 17880 42486 18000 42514
rect 17776 42220 17828 42226
rect 17776 42162 17828 42168
rect 17788 42022 17816 42162
rect 17776 42016 17828 42022
rect 17776 41958 17828 41964
rect 17866 41848 17922 41857
rect 17604 41806 17724 41834
rect 17592 41744 17644 41750
rect 17592 41686 17644 41692
rect 17604 41274 17632 41686
rect 17592 41268 17644 41274
rect 17592 41210 17644 41216
rect 17592 41132 17644 41138
rect 17592 41074 17644 41080
rect 17500 41064 17552 41070
rect 17500 41006 17552 41012
rect 17498 40896 17554 40905
rect 17498 40831 17554 40840
rect 17512 40662 17540 40831
rect 17500 40656 17552 40662
rect 17500 40598 17552 40604
rect 17604 40186 17632 41074
rect 17696 41070 17724 41806
rect 17866 41783 17922 41792
rect 17880 41750 17908 41783
rect 17868 41744 17920 41750
rect 17868 41686 17920 41692
rect 17776 41608 17828 41614
rect 17774 41576 17776 41585
rect 17828 41576 17830 41585
rect 17774 41511 17830 41520
rect 17972 41274 18000 42486
rect 17868 41268 17920 41274
rect 17868 41210 17920 41216
rect 17960 41268 18012 41274
rect 17960 41210 18012 41216
rect 17880 41154 17908 41210
rect 18064 41154 18092 42570
rect 18156 42362 18184 43268
rect 18248 42838 18276 44540
rect 18432 43450 18460 44540
rect 18616 43874 18644 44540
rect 18800 44010 18828 44540
rect 18800 43982 18920 44010
rect 18616 43846 18828 43874
rect 18420 43444 18472 43450
rect 18420 43386 18472 43392
rect 18420 43308 18472 43314
rect 18420 43250 18472 43256
rect 18604 43308 18656 43314
rect 18604 43250 18656 43256
rect 18326 43208 18382 43217
rect 18326 43143 18382 43152
rect 18236 42832 18288 42838
rect 18236 42774 18288 42780
rect 18340 42702 18368 43143
rect 18328 42696 18380 42702
rect 18328 42638 18380 42644
rect 18144 42356 18196 42362
rect 18144 42298 18196 42304
rect 18328 42152 18380 42158
rect 18328 42094 18380 42100
rect 18340 41698 18368 42094
rect 18432 41818 18460 43250
rect 18512 43240 18564 43246
rect 18512 43182 18564 43188
rect 18420 41812 18472 41818
rect 18420 41754 18472 41760
rect 18340 41682 18460 41698
rect 18340 41676 18472 41682
rect 18340 41670 18420 41676
rect 18420 41618 18472 41624
rect 18328 41608 18380 41614
rect 17880 41126 18092 41154
rect 18156 41534 18276 41562
rect 18328 41550 18380 41556
rect 17684 41064 17736 41070
rect 17684 41006 17736 41012
rect 17958 41032 18014 41041
rect 17868 40996 17920 41002
rect 17958 40967 18014 40976
rect 17868 40938 17920 40944
rect 17880 40662 17908 40938
rect 17868 40656 17920 40662
rect 17774 40624 17830 40633
rect 17868 40598 17920 40604
rect 17774 40559 17830 40568
rect 17684 40520 17736 40526
rect 17684 40462 17736 40468
rect 17696 40186 17724 40462
rect 17788 40186 17816 40559
rect 17972 40526 18000 40967
rect 17960 40520 18012 40526
rect 17960 40462 18012 40468
rect 18050 40352 18106 40361
rect 18050 40287 18106 40296
rect 18064 40186 18092 40287
rect 17592 40180 17644 40186
rect 17592 40122 17644 40128
rect 17684 40180 17736 40186
rect 17684 40122 17736 40128
rect 17776 40180 17828 40186
rect 17776 40122 17828 40128
rect 18052 40180 18104 40186
rect 18052 40122 18104 40128
rect 18156 40118 18184 41534
rect 18248 41478 18276 41534
rect 18236 41472 18288 41478
rect 18236 41414 18288 41420
rect 18340 41313 18368 41550
rect 18420 41472 18472 41478
rect 18420 41414 18472 41420
rect 18524 41414 18552 43182
rect 18616 42945 18644 43250
rect 18800 43110 18828 43846
rect 18788 43104 18840 43110
rect 18788 43046 18840 43052
rect 18602 42936 18658 42945
rect 18602 42871 18658 42880
rect 18788 42900 18840 42906
rect 18788 42842 18840 42848
rect 18604 42220 18656 42226
rect 18800 42208 18828 42842
rect 18892 42786 18920 43982
rect 18984 43654 19012 44540
rect 18972 43648 19024 43654
rect 18972 43590 19024 43596
rect 19168 43296 19196 44540
rect 19352 43874 19380 44540
rect 19352 43846 19472 43874
rect 19076 43268 19196 43296
rect 19076 42888 19104 43268
rect 19444 43178 19472 43846
rect 19432 43172 19484 43178
rect 19432 43114 19484 43120
rect 19143 43004 19451 43013
rect 19143 43002 19149 43004
rect 19205 43002 19229 43004
rect 19285 43002 19309 43004
rect 19365 43002 19389 43004
rect 19445 43002 19451 43004
rect 19205 42950 19207 43002
rect 19387 42950 19389 43002
rect 19143 42948 19149 42950
rect 19205 42948 19229 42950
rect 19285 42948 19309 42950
rect 19365 42948 19389 42950
rect 19445 42948 19451 42950
rect 19143 42939 19451 42948
rect 19536 42888 19564 44540
rect 19720 43296 19748 44540
rect 19904 43602 19932 44540
rect 20812 43648 20864 43654
rect 19904 43574 20024 43602
rect 20812 43590 20864 43596
rect 22374 43616 22430 43625
rect 19720 43268 19840 43296
rect 19708 42900 19760 42906
rect 19076 42860 19196 42888
rect 19536 42860 19708 42888
rect 18892 42758 19104 42786
rect 19076 42702 19104 42758
rect 19064 42696 19116 42702
rect 19064 42638 19116 42644
rect 18970 42528 19026 42537
rect 19026 42486 19104 42514
rect 18970 42463 19026 42472
rect 19076 42294 19104 42486
rect 19168 42362 19196 42860
rect 19708 42842 19760 42848
rect 19812 42786 19840 43268
rect 19720 42758 19840 42786
rect 19996 42770 20024 43574
rect 20824 43382 20852 43590
rect 21742 43548 22050 43557
rect 22374 43551 22430 43560
rect 21742 43546 21748 43548
rect 21804 43546 21828 43548
rect 21884 43546 21908 43548
rect 21964 43546 21988 43548
rect 22044 43546 22050 43548
rect 21804 43494 21806 43546
rect 21986 43494 21988 43546
rect 21742 43492 21748 43494
rect 21804 43492 21828 43494
rect 21884 43492 21908 43494
rect 21964 43492 21988 43494
rect 22044 43492 22050 43494
rect 21742 43483 22050 43492
rect 20720 43376 20772 43382
rect 20720 43318 20772 43324
rect 20812 43376 20864 43382
rect 20812 43318 20864 43324
rect 20534 43072 20590 43081
rect 20534 43007 20590 43016
rect 19984 42764 20036 42770
rect 19340 42628 19392 42634
rect 19340 42570 19392 42576
rect 19616 42628 19668 42634
rect 19616 42570 19668 42576
rect 19156 42356 19208 42362
rect 19156 42298 19208 42304
rect 19064 42288 19116 42294
rect 19064 42230 19116 42236
rect 18880 42220 18932 42226
rect 18800 42180 18880 42208
rect 18604 42162 18656 42168
rect 18880 42162 18932 42168
rect 18972 42220 19024 42226
rect 18972 42162 19024 42168
rect 18616 41562 18644 42162
rect 18880 42084 18932 42090
rect 18880 42026 18932 42032
rect 18892 41750 18920 42026
rect 18984 41857 19012 42162
rect 19352 42072 19380 42570
rect 19524 42220 19576 42226
rect 19524 42162 19576 42168
rect 19536 42129 19564 42162
rect 19076 42044 19380 42072
rect 19522 42120 19578 42129
rect 19522 42055 19578 42064
rect 18970 41848 19026 41857
rect 18970 41783 19026 41792
rect 18880 41744 18932 41750
rect 18880 41686 18932 41692
rect 18616 41534 19012 41562
rect 18326 41304 18382 41313
rect 18326 41239 18382 41248
rect 18234 41168 18290 41177
rect 18234 41103 18236 41112
rect 18288 41103 18290 41112
rect 18236 41074 18288 41080
rect 18432 41018 18460 41414
rect 18524 41386 18736 41414
rect 18708 41274 18736 41386
rect 18696 41268 18748 41274
rect 18696 41210 18748 41216
rect 18788 41268 18840 41274
rect 18788 41210 18840 41216
rect 18800 41154 18828 41210
rect 18248 40990 18460 41018
rect 18524 41126 18828 41154
rect 18878 41168 18934 41177
rect 18248 40526 18276 40990
rect 18236 40520 18288 40526
rect 18236 40462 18288 40468
rect 18328 40520 18380 40526
rect 18328 40462 18380 40468
rect 18418 40488 18474 40497
rect 18144 40112 18196 40118
rect 17420 40038 17632 40066
rect 18144 40054 18196 40060
rect 17500 39432 17552 39438
rect 17500 39374 17552 39380
rect 17236 36922 17264 37198
rect 17328 37182 17448 37210
rect 17316 37120 17368 37126
rect 17316 37062 17368 37068
rect 17328 36922 17356 37062
rect 17224 36916 17276 36922
rect 17224 36858 17276 36864
rect 17316 36916 17368 36922
rect 17316 36858 17368 36864
rect 17314 35320 17370 35329
rect 17314 35255 17370 35264
rect 17132 33652 17184 33658
rect 17132 33594 17184 33600
rect 17224 33516 17276 33522
rect 17224 33458 17276 33464
rect 17236 33425 17264 33458
rect 17222 33416 17278 33425
rect 17132 33380 17184 33386
rect 17222 33351 17278 33360
rect 17132 33322 17184 33328
rect 17144 32722 17172 33322
rect 17144 32694 17264 32722
rect 17132 32224 17184 32230
rect 17052 32184 17132 32212
rect 17132 32166 17184 32172
rect 17236 32042 17264 32694
rect 17144 32014 17264 32042
rect 16948 31816 17000 31822
rect 16948 31758 17000 31764
rect 17144 31754 17172 32014
rect 17224 31884 17276 31890
rect 17224 31826 17276 31832
rect 17052 31726 17172 31754
rect 16868 31640 16988 31668
rect 16544 31580 16852 31589
rect 16544 31578 16550 31580
rect 16606 31578 16630 31580
rect 16686 31578 16710 31580
rect 16766 31578 16790 31580
rect 16846 31578 16852 31580
rect 16606 31526 16608 31578
rect 16788 31526 16790 31578
rect 16544 31524 16550 31526
rect 16606 31524 16630 31526
rect 16686 31524 16710 31526
rect 16766 31524 16790 31526
rect 16846 31524 16852 31526
rect 16544 31515 16852 31524
rect 16544 30492 16852 30501
rect 16544 30490 16550 30492
rect 16606 30490 16630 30492
rect 16686 30490 16710 30492
rect 16766 30490 16790 30492
rect 16846 30490 16852 30492
rect 16606 30438 16608 30490
rect 16788 30438 16790 30490
rect 16544 30436 16550 30438
rect 16606 30436 16630 30438
rect 16686 30436 16710 30438
rect 16766 30436 16790 30438
rect 16846 30436 16852 30438
rect 16544 30427 16852 30436
rect 16960 30274 16988 31640
rect 16868 30258 16988 30274
rect 16856 30252 16988 30258
rect 16908 30246 16988 30252
rect 17052 30274 17080 31726
rect 17236 31482 17264 31826
rect 17224 31476 17276 31482
rect 17224 31418 17276 31424
rect 17224 31340 17276 31346
rect 17224 31282 17276 31288
rect 17236 30666 17264 31282
rect 17224 30660 17276 30666
rect 17224 30602 17276 30608
rect 17052 30246 17172 30274
rect 16856 30194 16908 30200
rect 16408 30110 16528 30138
rect 16396 30048 16448 30054
rect 16396 29990 16448 29996
rect 16408 29850 16436 29990
rect 16396 29844 16448 29850
rect 16396 29786 16448 29792
rect 16500 29730 16528 30110
rect 16764 30048 16816 30054
rect 16764 29990 16816 29996
rect 16408 29702 16528 29730
rect 16304 29164 16356 29170
rect 16304 29106 16356 29112
rect 16212 28960 16264 28966
rect 16212 28902 16264 28908
rect 16224 28801 16252 28902
rect 16210 28792 16266 28801
rect 16210 28727 16266 28736
rect 16212 28552 16264 28558
rect 16210 28520 16212 28529
rect 16264 28520 16266 28529
rect 16210 28455 16266 28464
rect 16212 28008 16264 28014
rect 16212 27950 16264 27956
rect 16408 27962 16436 29702
rect 16776 29646 16804 29990
rect 16764 29640 16816 29646
rect 16764 29582 16816 29588
rect 17040 29504 17092 29510
rect 17040 29446 17092 29452
rect 16544 29404 16852 29413
rect 16544 29402 16550 29404
rect 16606 29402 16630 29404
rect 16686 29402 16710 29404
rect 16766 29402 16790 29404
rect 16846 29402 16852 29404
rect 16606 29350 16608 29402
rect 16788 29350 16790 29402
rect 16544 29348 16550 29350
rect 16606 29348 16630 29350
rect 16686 29348 16710 29350
rect 16766 29348 16790 29350
rect 16846 29348 16852 29350
rect 16544 29339 16852 29348
rect 17052 29306 17080 29446
rect 17040 29300 17092 29306
rect 17040 29242 17092 29248
rect 16672 29164 16724 29170
rect 16672 29106 16724 29112
rect 16684 28994 16712 29106
rect 16684 28966 16988 28994
rect 16960 28694 16988 28966
rect 17038 28928 17094 28937
rect 17038 28863 17094 28872
rect 16948 28688 17000 28694
rect 16948 28630 17000 28636
rect 16544 28316 16852 28325
rect 16544 28314 16550 28316
rect 16606 28314 16630 28316
rect 16686 28314 16710 28316
rect 16766 28314 16790 28316
rect 16846 28314 16852 28316
rect 16606 28262 16608 28314
rect 16788 28262 16790 28314
rect 16544 28260 16550 28262
rect 16606 28260 16630 28262
rect 16686 28260 16710 28262
rect 16766 28260 16790 28262
rect 16846 28260 16852 28262
rect 16544 28251 16852 28260
rect 17052 28218 17080 28863
rect 17040 28212 17092 28218
rect 17040 28154 17092 28160
rect 17040 28008 17092 28014
rect 16224 27674 16252 27950
rect 16408 27934 16528 27962
rect 17144 27985 17172 30246
rect 17224 29504 17276 29510
rect 17224 29446 17276 29452
rect 17236 28558 17264 29446
rect 17224 28552 17276 28558
rect 17224 28494 17276 28500
rect 17040 27950 17092 27956
rect 17130 27976 17186 27985
rect 16396 27872 16448 27878
rect 16396 27814 16448 27820
rect 16212 27668 16264 27674
rect 16212 27610 16264 27616
rect 16120 27124 16172 27130
rect 16120 27066 16172 27072
rect 16120 26988 16172 26994
rect 16120 26930 16172 26936
rect 16132 26586 16160 26930
rect 16120 26580 16172 26586
rect 16120 26522 16172 26528
rect 16224 26466 16252 27610
rect 16304 27056 16356 27062
rect 16304 26998 16356 27004
rect 16132 26438 16252 26466
rect 16132 26314 16160 26438
rect 16316 26314 16344 26998
rect 16408 26382 16436 27814
rect 16500 27554 16528 27934
rect 17052 27674 17080 27950
rect 17130 27911 17186 27920
rect 17328 27690 17356 35255
rect 17040 27668 17092 27674
rect 17040 27610 17092 27616
rect 17144 27662 17356 27690
rect 16500 27526 16620 27554
rect 16592 27418 16620 27526
rect 16592 27390 16988 27418
rect 16544 27228 16852 27237
rect 16544 27226 16550 27228
rect 16606 27226 16630 27228
rect 16686 27226 16710 27228
rect 16766 27226 16790 27228
rect 16846 27226 16852 27228
rect 16606 27174 16608 27226
rect 16788 27174 16790 27226
rect 16544 27172 16550 27174
rect 16606 27172 16630 27174
rect 16686 27172 16710 27174
rect 16766 27172 16790 27174
rect 16846 27172 16852 27174
rect 16544 27163 16852 27172
rect 16856 27124 16908 27130
rect 16856 27066 16908 27072
rect 16868 26994 16896 27066
rect 16856 26988 16908 26994
rect 16856 26930 16908 26936
rect 16396 26376 16448 26382
rect 16396 26318 16448 26324
rect 16120 26308 16172 26314
rect 16120 26250 16172 26256
rect 16304 26308 16356 26314
rect 16304 26250 16356 26256
rect 16212 26240 16264 26246
rect 16212 26182 16264 26188
rect 16224 25906 16252 26182
rect 16212 25900 16264 25906
rect 16212 25842 16264 25848
rect 16316 25786 16344 26250
rect 16544 26140 16852 26149
rect 16544 26138 16550 26140
rect 16606 26138 16630 26140
rect 16686 26138 16710 26140
rect 16766 26138 16790 26140
rect 16846 26138 16852 26140
rect 16606 26086 16608 26138
rect 16788 26086 16790 26138
rect 16544 26084 16550 26086
rect 16606 26084 16630 26086
rect 16686 26084 16710 26086
rect 16766 26084 16790 26086
rect 16846 26084 16852 26086
rect 16544 26075 16852 26084
rect 16224 25758 16344 25786
rect 16028 25220 16080 25226
rect 16028 25162 16080 25168
rect 15844 25152 15896 25158
rect 15844 25094 15896 25100
rect 16120 25152 16172 25158
rect 16120 25094 16172 25100
rect 15658 24984 15714 24993
rect 15658 24919 15714 24928
rect 15566 23080 15622 23089
rect 15566 23015 15622 23024
rect 15566 22944 15622 22953
rect 15566 22879 15622 22888
rect 15580 22166 15608 22879
rect 15568 22160 15620 22166
rect 15568 22102 15620 22108
rect 15580 21078 15608 22102
rect 15672 21185 15700 24919
rect 15856 23662 15884 25094
rect 16028 24608 16080 24614
rect 16028 24550 16080 24556
rect 15844 23656 15896 23662
rect 15844 23598 15896 23604
rect 16040 23254 16068 24550
rect 16132 24342 16160 25094
rect 16120 24336 16172 24342
rect 16120 24278 16172 24284
rect 16120 23656 16172 23662
rect 16120 23598 16172 23604
rect 16028 23248 16080 23254
rect 16028 23190 16080 23196
rect 15752 23180 15804 23186
rect 15752 23122 15804 23128
rect 15764 22778 15792 23122
rect 15752 22772 15804 22778
rect 15752 22714 15804 22720
rect 15936 22432 15988 22438
rect 15936 22374 15988 22380
rect 15948 22166 15976 22374
rect 15936 22160 15988 22166
rect 15936 22102 15988 22108
rect 15752 21344 15804 21350
rect 15752 21286 15804 21292
rect 15658 21176 15714 21185
rect 15658 21111 15714 21120
rect 15568 21072 15620 21078
rect 15568 21014 15620 21020
rect 15568 20596 15620 20602
rect 15568 20538 15620 20544
rect 15580 15570 15608 20538
rect 15660 20528 15712 20534
rect 15660 20470 15712 20476
rect 15672 18358 15700 20470
rect 15764 19718 15792 21286
rect 16132 21078 16160 23598
rect 16224 21486 16252 25758
rect 16544 25052 16852 25061
rect 16544 25050 16550 25052
rect 16606 25050 16630 25052
rect 16686 25050 16710 25052
rect 16766 25050 16790 25052
rect 16846 25050 16852 25052
rect 16606 24998 16608 25050
rect 16788 24998 16790 25050
rect 16544 24996 16550 24998
rect 16606 24996 16630 24998
rect 16686 24996 16710 24998
rect 16766 24996 16790 24998
rect 16846 24996 16852 24998
rect 16544 24987 16852 24996
rect 16960 24857 16988 27390
rect 17052 26790 17080 27610
rect 17040 26784 17092 26790
rect 17040 26726 17092 26732
rect 17040 26036 17092 26042
rect 17040 25978 17092 25984
rect 17052 25158 17080 25978
rect 17040 25152 17092 25158
rect 17040 25094 17092 25100
rect 16946 24848 17002 24857
rect 16946 24783 17002 24792
rect 16394 24440 16450 24449
rect 16394 24375 16450 24384
rect 16948 24404 17000 24410
rect 16408 24206 16436 24375
rect 16948 24346 17000 24352
rect 16304 24200 16356 24206
rect 16304 24142 16356 24148
rect 16396 24200 16448 24206
rect 16396 24142 16448 24148
rect 16316 24070 16344 24142
rect 16304 24064 16356 24070
rect 16304 24006 16356 24012
rect 16544 23964 16852 23973
rect 16544 23962 16550 23964
rect 16606 23962 16630 23964
rect 16686 23962 16710 23964
rect 16766 23962 16790 23964
rect 16846 23962 16852 23964
rect 16606 23910 16608 23962
rect 16788 23910 16790 23962
rect 16544 23908 16550 23910
rect 16606 23908 16630 23910
rect 16686 23908 16710 23910
rect 16766 23908 16790 23910
rect 16846 23908 16852 23910
rect 16544 23899 16852 23908
rect 16396 23316 16448 23322
rect 16396 23258 16448 23264
rect 16408 23118 16436 23258
rect 16396 23112 16448 23118
rect 16396 23054 16448 23060
rect 16302 22808 16358 22817
rect 16408 22778 16436 23054
rect 16544 22876 16852 22885
rect 16544 22874 16550 22876
rect 16606 22874 16630 22876
rect 16686 22874 16710 22876
rect 16766 22874 16790 22876
rect 16846 22874 16852 22876
rect 16606 22822 16608 22874
rect 16788 22822 16790 22874
rect 16544 22820 16550 22822
rect 16606 22820 16630 22822
rect 16686 22820 16710 22822
rect 16766 22820 16790 22822
rect 16846 22820 16852 22822
rect 16544 22811 16852 22820
rect 16302 22743 16358 22752
rect 16396 22772 16448 22778
rect 16316 22030 16344 22743
rect 16396 22714 16448 22720
rect 16960 22642 16988 24346
rect 17052 23338 17080 25094
rect 17144 23497 17172 27662
rect 17420 27554 17448 37182
rect 17512 35562 17540 39374
rect 17604 35578 17632 40038
rect 17684 40044 17736 40050
rect 17684 39986 17736 39992
rect 17696 39642 17724 39986
rect 18052 39976 18104 39982
rect 18052 39918 18104 39924
rect 18064 39642 18092 39918
rect 17684 39636 17736 39642
rect 17684 39578 17736 39584
rect 18052 39636 18104 39642
rect 18052 39578 18104 39584
rect 17774 39536 17830 39545
rect 17774 39471 17830 39480
rect 17684 39432 17736 39438
rect 17684 39374 17736 39380
rect 17696 38554 17724 39374
rect 17684 38548 17736 38554
rect 17684 38490 17736 38496
rect 17788 35680 17816 39471
rect 18340 37738 18368 40462
rect 18418 40423 18474 40432
rect 18432 40186 18460 40423
rect 18524 40390 18552 41126
rect 18878 41103 18934 41112
rect 18892 41018 18920 41103
rect 18696 40996 18748 41002
rect 18696 40938 18748 40944
rect 18800 40990 18920 41018
rect 18602 40624 18658 40633
rect 18602 40559 18658 40568
rect 18616 40390 18644 40559
rect 18512 40384 18564 40390
rect 18512 40326 18564 40332
rect 18604 40384 18656 40390
rect 18604 40326 18656 40332
rect 18420 40180 18472 40186
rect 18420 40122 18472 40128
rect 18708 40050 18736 40938
rect 18800 40934 18828 40990
rect 18788 40928 18840 40934
rect 18788 40870 18840 40876
rect 18880 40928 18932 40934
rect 18880 40870 18932 40876
rect 18788 40520 18840 40526
rect 18788 40462 18840 40468
rect 18800 40186 18828 40462
rect 18892 40186 18920 40870
rect 18984 40186 19012 41534
rect 19076 41274 19104 42044
rect 19143 41916 19451 41925
rect 19143 41914 19149 41916
rect 19205 41914 19229 41916
rect 19285 41914 19309 41916
rect 19365 41914 19389 41916
rect 19445 41914 19451 41916
rect 19205 41862 19207 41914
rect 19387 41862 19389 41914
rect 19143 41860 19149 41862
rect 19205 41860 19229 41862
rect 19285 41860 19309 41862
rect 19365 41860 19389 41862
rect 19445 41860 19451 41862
rect 19143 41851 19451 41860
rect 19340 41744 19392 41750
rect 19340 41686 19392 41692
rect 19352 41414 19380 41686
rect 19628 41562 19656 42570
rect 19720 42294 19748 42758
rect 19984 42706 20036 42712
rect 20444 42628 20496 42634
rect 20444 42570 20496 42576
rect 20456 42401 20484 42570
rect 20442 42392 20498 42401
rect 20442 42327 20498 42336
rect 19708 42288 19760 42294
rect 19708 42230 19760 42236
rect 19984 42220 20036 42226
rect 19984 42162 20036 42168
rect 20444 42220 20496 42226
rect 20444 42162 20496 42168
rect 19708 42016 19760 42022
rect 19708 41958 19760 41964
rect 19260 41386 19380 41414
rect 19444 41534 19656 41562
rect 19064 41268 19116 41274
rect 19064 41210 19116 41216
rect 19064 41132 19116 41138
rect 19064 41074 19116 41080
rect 18788 40180 18840 40186
rect 18788 40122 18840 40128
rect 18880 40180 18932 40186
rect 18880 40122 18932 40128
rect 18972 40180 19024 40186
rect 18972 40122 19024 40128
rect 19076 40089 19104 41074
rect 19260 41041 19288 41386
rect 19246 41032 19302 41041
rect 19246 40967 19302 40976
rect 19340 40996 19392 41002
rect 19444 40984 19472 41534
rect 19720 41274 19748 41958
rect 19800 41608 19852 41614
rect 19800 41550 19852 41556
rect 19708 41268 19760 41274
rect 19708 41210 19760 41216
rect 19524 41132 19576 41138
rect 19524 41074 19576 41080
rect 19392 40956 19472 40984
rect 19340 40938 19392 40944
rect 19143 40828 19451 40837
rect 19143 40826 19149 40828
rect 19205 40826 19229 40828
rect 19285 40826 19309 40828
rect 19365 40826 19389 40828
rect 19445 40826 19451 40828
rect 19205 40774 19207 40826
rect 19387 40774 19389 40826
rect 19143 40772 19149 40774
rect 19205 40772 19229 40774
rect 19285 40772 19309 40774
rect 19365 40772 19389 40774
rect 19445 40772 19451 40774
rect 19143 40763 19451 40772
rect 19432 40656 19484 40662
rect 19536 40644 19564 41074
rect 19812 40769 19840 41550
rect 19892 41132 19944 41138
rect 19892 41074 19944 41080
rect 19798 40760 19854 40769
rect 19798 40695 19854 40704
rect 19484 40616 19564 40644
rect 19800 40656 19852 40662
rect 19432 40598 19484 40604
rect 19800 40598 19852 40604
rect 19616 40520 19668 40526
rect 19616 40462 19668 40468
rect 19156 40452 19208 40458
rect 19156 40394 19208 40400
rect 19168 40186 19196 40394
rect 19432 40384 19484 40390
rect 19432 40326 19484 40332
rect 19156 40180 19208 40186
rect 19156 40122 19208 40128
rect 19062 40080 19118 40089
rect 18696 40044 18748 40050
rect 18696 39986 18748 39992
rect 18788 40044 18840 40050
rect 18788 39986 18840 39992
rect 18972 40044 19024 40050
rect 19062 40015 19118 40024
rect 18972 39986 19024 39992
rect 18800 39522 18828 39986
rect 18984 39574 19012 39986
rect 19444 39982 19472 40326
rect 19432 39976 19484 39982
rect 19432 39918 19484 39924
rect 19522 39944 19578 39953
rect 19522 39879 19578 39888
rect 19143 39740 19451 39749
rect 19143 39738 19149 39740
rect 19205 39738 19229 39740
rect 19285 39738 19309 39740
rect 19365 39738 19389 39740
rect 19445 39738 19451 39740
rect 19205 39686 19207 39738
rect 19387 39686 19389 39738
rect 19143 39684 19149 39686
rect 19205 39684 19229 39686
rect 19285 39684 19309 39686
rect 19365 39684 19389 39686
rect 19445 39684 19451 39686
rect 19143 39675 19451 39684
rect 18708 39494 18828 39522
rect 18972 39568 19024 39574
rect 18972 39510 19024 39516
rect 19340 39568 19392 39574
rect 19340 39510 19392 39516
rect 18604 38344 18656 38350
rect 18604 38286 18656 38292
rect 18616 38010 18644 38286
rect 18604 38004 18656 38010
rect 18604 37946 18656 37952
rect 18328 37732 18380 37738
rect 18328 37674 18380 37680
rect 17868 37256 17920 37262
rect 17868 37198 17920 37204
rect 18052 37256 18104 37262
rect 18052 37198 18104 37204
rect 18236 37256 18288 37262
rect 18236 37198 18288 37204
rect 17880 36922 17908 37198
rect 17868 36916 17920 36922
rect 17868 36858 17920 36864
rect 18064 36802 18092 37198
rect 18144 37120 18196 37126
rect 18144 37062 18196 37068
rect 18156 36922 18184 37062
rect 18144 36916 18196 36922
rect 18144 36858 18196 36864
rect 18064 36774 18184 36802
rect 18156 36582 18184 36774
rect 17960 36576 18012 36582
rect 17960 36518 18012 36524
rect 18144 36576 18196 36582
rect 18144 36518 18196 36524
rect 17972 35698 18000 36518
rect 18156 36378 18184 36518
rect 18144 36372 18196 36378
rect 18144 36314 18196 36320
rect 18052 36236 18104 36242
rect 18052 36178 18104 36184
rect 17960 35692 18012 35698
rect 17788 35652 17908 35680
rect 17500 35556 17552 35562
rect 17604 35550 17724 35578
rect 17500 35498 17552 35504
rect 17512 35290 17540 35498
rect 17592 35488 17644 35494
rect 17592 35430 17644 35436
rect 17500 35284 17552 35290
rect 17500 35226 17552 35232
rect 17500 33108 17552 33114
rect 17500 33050 17552 33056
rect 17512 30258 17540 33050
rect 17604 30394 17632 35430
rect 17696 35136 17724 35550
rect 17776 35556 17828 35562
rect 17776 35498 17828 35504
rect 17788 35290 17816 35498
rect 17776 35284 17828 35290
rect 17776 35226 17828 35232
rect 17696 35108 17816 35136
rect 17684 32496 17736 32502
rect 17684 32438 17736 32444
rect 17592 30388 17644 30394
rect 17592 30330 17644 30336
rect 17500 30252 17552 30258
rect 17500 30194 17552 30200
rect 17500 29164 17552 29170
rect 17500 29106 17552 29112
rect 17512 28994 17540 29106
rect 17512 28966 17632 28994
rect 17500 28416 17552 28422
rect 17500 28358 17552 28364
rect 17512 28218 17540 28358
rect 17500 28212 17552 28218
rect 17500 28154 17552 28160
rect 17604 27826 17632 28966
rect 17696 27849 17724 32438
rect 17512 27798 17632 27826
rect 17682 27840 17738 27849
rect 17512 27674 17540 27798
rect 17682 27775 17738 27784
rect 17788 27690 17816 35108
rect 17880 32994 17908 35652
rect 17960 35634 18012 35640
rect 18064 35601 18092 36178
rect 18248 35850 18276 37198
rect 18340 36174 18368 37674
rect 18512 36712 18564 36718
rect 18512 36654 18564 36660
rect 18328 36168 18380 36174
rect 18328 36110 18380 36116
rect 18420 36100 18472 36106
rect 18420 36042 18472 36048
rect 18156 35822 18276 35850
rect 18050 35592 18106 35601
rect 17960 35556 18012 35562
rect 18050 35527 18106 35536
rect 17960 35498 18012 35504
rect 17972 34610 18000 35498
rect 18052 34740 18104 34746
rect 18052 34682 18104 34688
rect 17960 34604 18012 34610
rect 17960 34546 18012 34552
rect 17960 34400 18012 34406
rect 17960 34342 18012 34348
rect 17972 33998 18000 34342
rect 18064 34066 18092 34682
rect 18052 34060 18104 34066
rect 18052 34002 18104 34008
rect 17960 33992 18012 33998
rect 18156 33946 18184 35822
rect 18326 35728 18382 35737
rect 18236 35692 18288 35698
rect 18326 35663 18328 35672
rect 18236 35634 18288 35640
rect 18380 35663 18382 35672
rect 18328 35634 18380 35640
rect 18248 35057 18276 35634
rect 18432 35562 18460 36042
rect 18524 36038 18552 36654
rect 18512 36032 18564 36038
rect 18512 35974 18564 35980
rect 18512 35692 18564 35698
rect 18512 35634 18564 35640
rect 18420 35556 18472 35562
rect 18420 35498 18472 35504
rect 18418 35184 18474 35193
rect 18418 35119 18474 35128
rect 18234 35048 18290 35057
rect 18234 34983 18290 34992
rect 18328 34944 18380 34950
rect 18328 34886 18380 34892
rect 18236 34196 18288 34202
rect 18236 34138 18288 34144
rect 17960 33934 18012 33940
rect 18064 33918 18184 33946
rect 18064 33402 18092 33918
rect 17972 33374 18092 33402
rect 17972 33114 18000 33374
rect 18052 33312 18104 33318
rect 18052 33254 18104 33260
rect 18064 33114 18092 33254
rect 17960 33108 18012 33114
rect 17960 33050 18012 33056
rect 18052 33108 18104 33114
rect 18052 33050 18104 33056
rect 18144 33108 18196 33114
rect 18144 33050 18196 33056
rect 17880 32966 18000 32994
rect 18156 32978 18184 33050
rect 17868 32768 17920 32774
rect 17868 32710 17920 32716
rect 17880 32570 17908 32710
rect 17868 32564 17920 32570
rect 17868 32506 17920 32512
rect 17972 32502 18000 32966
rect 18144 32972 18196 32978
rect 18144 32914 18196 32920
rect 18248 32858 18276 34138
rect 18340 33289 18368 34886
rect 18326 33280 18382 33289
rect 18326 33215 18382 33224
rect 18328 33040 18380 33046
rect 18328 32982 18380 32988
rect 18340 32910 18368 32982
rect 18064 32830 18276 32858
rect 18328 32904 18380 32910
rect 18328 32846 18380 32852
rect 17960 32496 18012 32502
rect 17866 32464 17922 32473
rect 17960 32438 18012 32444
rect 17866 32399 17922 32408
rect 17500 27668 17552 27674
rect 17500 27610 17552 27616
rect 17604 27662 17816 27690
rect 17236 27526 17448 27554
rect 17130 23488 17186 23497
rect 17130 23423 17186 23432
rect 17052 23310 17172 23338
rect 16396 22636 16448 22642
rect 16396 22578 16448 22584
rect 16948 22636 17000 22642
rect 16948 22578 17000 22584
rect 16304 22024 16356 22030
rect 16304 21966 16356 21972
rect 16212 21480 16264 21486
rect 16212 21422 16264 21428
rect 16120 21072 16172 21078
rect 16120 21014 16172 21020
rect 16028 20936 16080 20942
rect 16028 20878 16080 20884
rect 16212 20936 16264 20942
rect 16212 20878 16264 20884
rect 15844 20800 15896 20806
rect 15844 20742 15896 20748
rect 15752 19712 15804 19718
rect 15752 19654 15804 19660
rect 15764 18850 15792 19654
rect 15856 19242 15884 20742
rect 15936 20528 15988 20534
rect 15936 20470 15988 20476
rect 15948 20369 15976 20470
rect 15934 20360 15990 20369
rect 15934 20295 15990 20304
rect 15948 19514 15976 20295
rect 16040 20058 16068 20878
rect 16120 20800 16172 20806
rect 16120 20742 16172 20748
rect 16132 20262 16160 20742
rect 16120 20256 16172 20262
rect 16120 20198 16172 20204
rect 16028 20052 16080 20058
rect 16028 19994 16080 20000
rect 16028 19780 16080 19786
rect 16028 19722 16080 19728
rect 15936 19508 15988 19514
rect 15936 19450 15988 19456
rect 15844 19236 15896 19242
rect 15844 19178 15896 19184
rect 15764 18822 15976 18850
rect 15660 18352 15712 18358
rect 15660 18294 15712 18300
rect 15752 18080 15804 18086
rect 15752 18022 15804 18028
rect 15658 17640 15714 17649
rect 15658 17575 15714 17584
rect 15672 17270 15700 17575
rect 15660 17264 15712 17270
rect 15660 17206 15712 17212
rect 15764 16130 15792 18022
rect 15948 17882 15976 18822
rect 15936 17876 15988 17882
rect 15936 17818 15988 17824
rect 16040 17610 16068 19722
rect 16132 19378 16160 20198
rect 16120 19372 16172 19378
rect 16120 19314 16172 19320
rect 16120 18964 16172 18970
rect 16120 18906 16172 18912
rect 16132 18465 16160 18906
rect 16118 18456 16174 18465
rect 16224 18426 16252 20878
rect 16304 20800 16356 20806
rect 16304 20742 16356 20748
rect 16316 19446 16344 20742
rect 16304 19440 16356 19446
rect 16304 19382 16356 19388
rect 16304 19168 16356 19174
rect 16304 19110 16356 19116
rect 16118 18391 16174 18400
rect 16212 18420 16264 18426
rect 16212 18362 16264 18368
rect 16210 18184 16266 18193
rect 16210 18119 16266 18128
rect 16224 18086 16252 18119
rect 16212 18080 16264 18086
rect 16212 18022 16264 18028
rect 16120 17876 16172 17882
rect 16120 17818 16172 17824
rect 16028 17604 16080 17610
rect 16028 17546 16080 17552
rect 16040 16794 16068 17546
rect 16132 17542 16160 17818
rect 16212 17740 16264 17746
rect 16212 17682 16264 17688
rect 16120 17536 16172 17542
rect 16120 17478 16172 17484
rect 15936 16788 15988 16794
rect 15936 16730 15988 16736
rect 16028 16788 16080 16794
rect 16028 16730 16080 16736
rect 15844 16584 15896 16590
rect 15844 16526 15896 16532
rect 15672 16102 15792 16130
rect 15856 16114 15884 16526
rect 15948 16250 15976 16730
rect 16132 16674 16160 17478
rect 16224 17338 16252 17682
rect 16212 17332 16264 17338
rect 16212 17274 16264 17280
rect 16212 16992 16264 16998
rect 16212 16934 16264 16940
rect 16040 16646 16160 16674
rect 15936 16244 15988 16250
rect 15936 16186 15988 16192
rect 15844 16108 15896 16114
rect 15568 15564 15620 15570
rect 15568 15506 15620 15512
rect 15568 15360 15620 15366
rect 15568 15302 15620 15308
rect 15580 15026 15608 15302
rect 15568 15020 15620 15026
rect 15568 14962 15620 14968
rect 15568 14816 15620 14822
rect 15568 14758 15620 14764
rect 15580 14618 15608 14758
rect 15568 14612 15620 14618
rect 15568 14554 15620 14560
rect 15672 14498 15700 16102
rect 15844 16050 15896 16056
rect 15752 16040 15804 16046
rect 15752 15982 15804 15988
rect 15764 15162 15792 15982
rect 15752 15156 15804 15162
rect 15752 15098 15804 15104
rect 15580 14470 15700 14498
rect 15580 13025 15608 14470
rect 15660 14408 15712 14414
rect 15660 14350 15712 14356
rect 15752 14408 15804 14414
rect 15752 14350 15804 14356
rect 15672 13433 15700 14350
rect 15764 13530 15792 14350
rect 15936 14272 15988 14278
rect 15936 14214 15988 14220
rect 15948 13977 15976 14214
rect 15934 13968 15990 13977
rect 15844 13932 15896 13938
rect 15934 13903 15990 13912
rect 15844 13874 15896 13880
rect 15752 13524 15804 13530
rect 15752 13466 15804 13472
rect 15658 13424 15714 13433
rect 15856 13394 15884 13874
rect 15658 13359 15714 13368
rect 15844 13388 15896 13394
rect 15844 13330 15896 13336
rect 15566 13016 15622 13025
rect 15566 12951 15622 12960
rect 15856 12434 15884 13330
rect 15764 12406 15884 12434
rect 15660 12096 15712 12102
rect 15660 12038 15712 12044
rect 15568 11212 15620 11218
rect 15672 11200 15700 12038
rect 15764 11762 15792 12406
rect 15936 12232 15988 12238
rect 15936 12174 15988 12180
rect 15752 11756 15804 11762
rect 15752 11698 15804 11704
rect 15620 11172 15700 11200
rect 15568 11154 15620 11160
rect 15580 9722 15608 11154
rect 15658 10976 15714 10985
rect 15658 10911 15714 10920
rect 15568 9716 15620 9722
rect 15568 9658 15620 9664
rect 15580 8906 15608 9658
rect 15568 8900 15620 8906
rect 15568 8842 15620 8848
rect 15292 8084 15344 8090
rect 15292 8026 15344 8032
rect 15304 7721 15332 8026
rect 15290 7712 15346 7721
rect 15290 7647 15346 7656
rect 15292 6112 15344 6118
rect 15292 6054 15344 6060
rect 15304 5914 15332 6054
rect 15292 5908 15344 5914
rect 15292 5850 15344 5856
rect 15396 5794 15424 8366
rect 15488 8350 15608 8378
rect 15476 8288 15528 8294
rect 15476 8230 15528 8236
rect 15488 5914 15516 8230
rect 15580 7274 15608 8350
rect 15568 7268 15620 7274
rect 15568 7210 15620 7216
rect 15672 6984 15700 10911
rect 15764 10538 15792 11698
rect 15948 11150 15976 12174
rect 16040 11914 16068 16646
rect 16120 16176 16172 16182
rect 16120 16118 16172 16124
rect 16132 15910 16160 16118
rect 16224 15978 16252 16934
rect 16212 15972 16264 15978
rect 16212 15914 16264 15920
rect 16316 15910 16344 19110
rect 16408 18290 16436 22578
rect 17040 21888 17092 21894
rect 17038 21856 17040 21865
rect 17092 21856 17094 21865
rect 16544 21788 16852 21797
rect 17038 21791 17094 21800
rect 16544 21786 16550 21788
rect 16606 21786 16630 21788
rect 16686 21786 16710 21788
rect 16766 21786 16790 21788
rect 16846 21786 16852 21788
rect 16606 21734 16608 21786
rect 16788 21734 16790 21786
rect 16544 21732 16550 21734
rect 16606 21732 16630 21734
rect 16686 21732 16710 21734
rect 16766 21732 16790 21734
rect 16846 21732 16852 21734
rect 16544 21723 16852 21732
rect 16856 21480 16908 21486
rect 16856 21422 16908 21428
rect 16868 20890 16896 21422
rect 17040 20936 17092 20942
rect 16868 20862 16988 20890
rect 17040 20878 17092 20884
rect 16544 20700 16852 20709
rect 16544 20698 16550 20700
rect 16606 20698 16630 20700
rect 16686 20698 16710 20700
rect 16766 20698 16790 20700
rect 16846 20698 16852 20700
rect 16606 20646 16608 20698
rect 16788 20646 16790 20698
rect 16544 20644 16550 20646
rect 16606 20644 16630 20646
rect 16686 20644 16710 20646
rect 16766 20644 16790 20646
rect 16846 20644 16852 20646
rect 16544 20635 16852 20644
rect 16960 20097 16988 20862
rect 16946 20088 17002 20097
rect 16946 20023 17002 20032
rect 16762 19952 16818 19961
rect 16762 19887 16818 19896
rect 16948 19916 17000 19922
rect 16776 19854 16804 19887
rect 16948 19858 17000 19864
rect 16764 19848 16816 19854
rect 16764 19790 16816 19796
rect 16544 19612 16852 19621
rect 16544 19610 16550 19612
rect 16606 19610 16630 19612
rect 16686 19610 16710 19612
rect 16766 19610 16790 19612
rect 16846 19610 16852 19612
rect 16606 19558 16608 19610
rect 16788 19558 16790 19610
rect 16544 19556 16550 19558
rect 16606 19556 16630 19558
rect 16686 19556 16710 19558
rect 16766 19556 16790 19558
rect 16846 19556 16852 19558
rect 16544 19547 16852 19556
rect 16856 19508 16908 19514
rect 16856 19450 16908 19456
rect 16868 19378 16896 19450
rect 16856 19372 16908 19378
rect 16856 19314 16908 19320
rect 16960 18970 16988 19858
rect 16948 18964 17000 18970
rect 16948 18906 17000 18912
rect 16948 18760 17000 18766
rect 17052 18748 17080 20878
rect 17144 20369 17172 23310
rect 17236 20992 17264 27526
rect 17316 27464 17368 27470
rect 17316 27406 17368 27412
rect 17408 27464 17460 27470
rect 17408 27406 17460 27412
rect 17328 27130 17356 27406
rect 17316 27124 17368 27130
rect 17316 27066 17368 27072
rect 17420 26586 17448 27406
rect 17408 26580 17460 26586
rect 17408 26522 17460 26528
rect 17408 25152 17460 25158
rect 17408 25094 17460 25100
rect 17500 25152 17552 25158
rect 17500 25094 17552 25100
rect 17420 24818 17448 25094
rect 17408 24812 17460 24818
rect 17408 24754 17460 24760
rect 17420 24410 17448 24754
rect 17408 24404 17460 24410
rect 17408 24346 17460 24352
rect 17512 24274 17540 25094
rect 17500 24268 17552 24274
rect 17500 24210 17552 24216
rect 17500 24132 17552 24138
rect 17500 24074 17552 24080
rect 17316 24064 17368 24070
rect 17316 24006 17368 24012
rect 17328 23730 17356 24006
rect 17316 23724 17368 23730
rect 17316 23666 17368 23672
rect 17406 23352 17462 23361
rect 17406 23287 17462 23296
rect 17420 22234 17448 23287
rect 17512 23050 17540 24074
rect 17500 23044 17552 23050
rect 17500 22986 17552 22992
rect 17408 22228 17460 22234
rect 17408 22170 17460 22176
rect 17604 21672 17632 27662
rect 17776 27600 17828 27606
rect 17776 27542 17828 27548
rect 17788 25906 17816 27542
rect 17776 25900 17828 25906
rect 17776 25842 17828 25848
rect 17684 25696 17736 25702
rect 17684 25638 17736 25644
rect 17696 24138 17724 25638
rect 17788 24886 17816 25842
rect 17880 25650 17908 32399
rect 17960 32224 18012 32230
rect 17960 32166 18012 32172
rect 17972 31346 18000 32166
rect 17960 31340 18012 31346
rect 17960 31282 18012 31288
rect 17972 29594 18000 31282
rect 18064 29714 18092 32830
rect 18236 32768 18288 32774
rect 18236 32710 18288 32716
rect 18144 31680 18196 31686
rect 18144 31622 18196 31628
rect 18156 31210 18184 31622
rect 18144 31204 18196 31210
rect 18144 31146 18196 31152
rect 18156 30734 18184 31146
rect 18144 30728 18196 30734
rect 18144 30670 18196 30676
rect 18052 29708 18104 29714
rect 18052 29650 18104 29656
rect 18144 29640 18196 29646
rect 17972 29566 18092 29594
rect 18144 29582 18196 29588
rect 17960 29504 18012 29510
rect 17960 29446 18012 29452
rect 17972 28218 18000 29446
rect 18064 29170 18092 29566
rect 18156 29306 18184 29582
rect 18144 29300 18196 29306
rect 18144 29242 18196 29248
rect 18052 29164 18104 29170
rect 18052 29106 18104 29112
rect 18052 28756 18104 28762
rect 18104 28716 18184 28744
rect 18052 28698 18104 28704
rect 17960 28212 18012 28218
rect 17960 28154 18012 28160
rect 18156 27674 18184 28716
rect 18052 27668 18104 27674
rect 18052 27610 18104 27616
rect 18144 27668 18196 27674
rect 18144 27610 18196 27616
rect 18064 27130 18092 27610
rect 18144 27532 18196 27538
rect 18144 27474 18196 27480
rect 18156 27130 18184 27474
rect 18052 27124 18104 27130
rect 18052 27066 18104 27072
rect 18144 27124 18196 27130
rect 18144 27066 18196 27072
rect 18050 27024 18106 27033
rect 18050 26959 18106 26968
rect 17880 25622 18000 25650
rect 17776 24880 17828 24886
rect 17776 24822 17828 24828
rect 17684 24132 17736 24138
rect 17684 24074 17736 24080
rect 17868 24132 17920 24138
rect 17868 24074 17920 24080
rect 17684 23520 17736 23526
rect 17684 23462 17736 23468
rect 17696 23186 17724 23462
rect 17684 23180 17736 23186
rect 17684 23122 17736 23128
rect 17684 23044 17736 23050
rect 17684 22986 17736 22992
rect 17696 22148 17724 22986
rect 17776 22636 17828 22642
rect 17776 22578 17828 22584
rect 17788 22438 17816 22578
rect 17776 22432 17828 22438
rect 17776 22374 17828 22380
rect 17696 22120 17816 22148
rect 17684 21956 17736 21962
rect 17684 21898 17736 21904
rect 17512 21644 17632 21672
rect 17408 21412 17460 21418
rect 17408 21354 17460 21360
rect 17420 21146 17448 21354
rect 17408 21140 17460 21146
rect 17408 21082 17460 21088
rect 17512 21026 17540 21644
rect 17592 21548 17644 21554
rect 17592 21490 17644 21496
rect 17604 21350 17632 21490
rect 17592 21344 17644 21350
rect 17592 21286 17644 21292
rect 17696 21049 17724 21898
rect 17420 20998 17540 21026
rect 17682 21040 17738 21049
rect 17236 20964 17356 20992
rect 17224 20868 17276 20874
rect 17224 20810 17276 20816
rect 17130 20360 17186 20369
rect 17130 20295 17186 20304
rect 17130 20088 17186 20097
rect 17130 20023 17186 20032
rect 17144 19854 17172 20023
rect 17132 19848 17184 19854
rect 17132 19790 17184 19796
rect 17132 19712 17184 19718
rect 17132 19654 17184 19660
rect 17144 19514 17172 19654
rect 17132 19508 17184 19514
rect 17132 19450 17184 19456
rect 17130 19272 17186 19281
rect 17130 19207 17186 19216
rect 17000 18720 17080 18748
rect 16948 18702 17000 18708
rect 16544 18524 16852 18533
rect 16544 18522 16550 18524
rect 16606 18522 16630 18524
rect 16686 18522 16710 18524
rect 16766 18522 16790 18524
rect 16846 18522 16852 18524
rect 16606 18470 16608 18522
rect 16788 18470 16790 18522
rect 16544 18468 16550 18470
rect 16606 18468 16630 18470
rect 16686 18468 16710 18470
rect 16766 18468 16790 18470
rect 16846 18468 16852 18470
rect 16544 18459 16852 18468
rect 16396 18284 16448 18290
rect 16396 18226 16448 18232
rect 16672 18216 16724 18222
rect 16672 18158 16724 18164
rect 16396 18148 16448 18154
rect 16396 18090 16448 18096
rect 16120 15904 16172 15910
rect 16120 15846 16172 15852
rect 16304 15904 16356 15910
rect 16304 15846 16356 15852
rect 16302 15600 16358 15609
rect 16302 15535 16358 15544
rect 16212 15496 16264 15502
rect 16212 15438 16264 15444
rect 16120 15156 16172 15162
rect 16120 15098 16172 15104
rect 16132 14006 16160 15098
rect 16224 14006 16252 15438
rect 16316 14414 16344 15535
rect 16408 15162 16436 18090
rect 16580 18080 16632 18086
rect 16580 18022 16632 18028
rect 16592 17610 16620 18022
rect 16580 17604 16632 17610
rect 16580 17546 16632 17552
rect 16684 17542 16712 18158
rect 16672 17536 16724 17542
rect 16672 17478 16724 17484
rect 16544 17436 16852 17445
rect 16544 17434 16550 17436
rect 16606 17434 16630 17436
rect 16686 17434 16710 17436
rect 16766 17434 16790 17436
rect 16846 17434 16852 17436
rect 16606 17382 16608 17434
rect 16788 17382 16790 17434
rect 16544 17380 16550 17382
rect 16606 17380 16630 17382
rect 16686 17380 16710 17382
rect 16766 17380 16790 17382
rect 16846 17380 16852 17382
rect 16544 17371 16852 17380
rect 16856 17332 16908 17338
rect 16856 17274 16908 17280
rect 16868 17134 16896 17274
rect 16856 17128 16908 17134
rect 16856 17070 16908 17076
rect 16762 16960 16818 16969
rect 16762 16895 16818 16904
rect 16776 16794 16804 16895
rect 16764 16788 16816 16794
rect 16764 16730 16816 16736
rect 16544 16348 16852 16357
rect 16544 16346 16550 16348
rect 16606 16346 16630 16348
rect 16686 16346 16710 16348
rect 16766 16346 16790 16348
rect 16846 16346 16852 16348
rect 16606 16294 16608 16346
rect 16788 16294 16790 16346
rect 16544 16292 16550 16294
rect 16606 16292 16630 16294
rect 16686 16292 16710 16294
rect 16766 16292 16790 16294
rect 16846 16292 16852 16294
rect 16544 16283 16852 16292
rect 16856 16108 16908 16114
rect 16856 16050 16908 16056
rect 16868 15366 16896 16050
rect 16856 15360 16908 15366
rect 16856 15302 16908 15308
rect 16544 15260 16852 15269
rect 16544 15258 16550 15260
rect 16606 15258 16630 15260
rect 16686 15258 16710 15260
rect 16766 15258 16790 15260
rect 16846 15258 16852 15260
rect 16606 15206 16608 15258
rect 16788 15206 16790 15258
rect 16544 15204 16550 15206
rect 16606 15204 16630 15206
rect 16686 15204 16710 15206
rect 16766 15204 16790 15206
rect 16846 15204 16852 15206
rect 16544 15195 16852 15204
rect 16396 15156 16448 15162
rect 16396 15098 16448 15104
rect 16396 14816 16448 14822
rect 16396 14758 16448 14764
rect 16304 14408 16356 14414
rect 16304 14350 16356 14356
rect 16120 14000 16172 14006
rect 16120 13942 16172 13948
rect 16212 14000 16264 14006
rect 16212 13942 16264 13948
rect 16132 13394 16160 13942
rect 16120 13388 16172 13394
rect 16120 13330 16172 13336
rect 16132 12442 16160 13330
rect 16120 12436 16172 12442
rect 16120 12378 16172 12384
rect 16132 12102 16160 12378
rect 16120 12096 16172 12102
rect 16120 12038 16172 12044
rect 16040 11886 16160 11914
rect 15936 11144 15988 11150
rect 15842 11112 15898 11121
rect 15936 11086 15988 11092
rect 15842 11047 15898 11056
rect 15752 10532 15804 10538
rect 15752 10474 15804 10480
rect 15752 9920 15804 9926
rect 15752 9862 15804 9868
rect 15764 9654 15792 9862
rect 15752 9648 15804 9654
rect 15752 9590 15804 9596
rect 15764 7546 15792 9590
rect 15856 9081 15884 11047
rect 15936 10260 15988 10266
rect 15936 10202 15988 10208
rect 15842 9072 15898 9081
rect 15842 9007 15898 9016
rect 15844 8968 15896 8974
rect 15844 8910 15896 8916
rect 15752 7540 15804 7546
rect 15752 7482 15804 7488
rect 15856 7426 15884 8910
rect 15948 8786 15976 10202
rect 16028 10056 16080 10062
rect 16028 9998 16080 10004
rect 16040 9722 16068 9998
rect 16028 9716 16080 9722
rect 16028 9658 16080 9664
rect 16040 9625 16068 9658
rect 16026 9616 16082 9625
rect 16132 9586 16160 11886
rect 16224 11762 16252 13942
rect 16408 13802 16436 14758
rect 16544 14172 16852 14181
rect 16544 14170 16550 14172
rect 16606 14170 16630 14172
rect 16686 14170 16710 14172
rect 16766 14170 16790 14172
rect 16846 14170 16852 14172
rect 16606 14118 16608 14170
rect 16788 14118 16790 14170
rect 16544 14116 16550 14118
rect 16606 14116 16630 14118
rect 16686 14116 16710 14118
rect 16766 14116 16790 14118
rect 16846 14116 16852 14118
rect 16544 14107 16852 14116
rect 16580 14068 16632 14074
rect 16580 14010 16632 14016
rect 16396 13796 16448 13802
rect 16396 13738 16448 13744
rect 16592 13530 16620 14010
rect 16960 13938 16988 18702
rect 17040 17672 17092 17678
rect 17040 17614 17092 17620
rect 17052 16998 17080 17614
rect 17040 16992 17092 16998
rect 17040 16934 17092 16940
rect 17040 16448 17092 16454
rect 17040 16390 17092 16396
rect 17052 15348 17080 16390
rect 17144 15502 17172 19207
rect 17236 18329 17264 20810
rect 17328 19922 17356 20964
rect 17316 19916 17368 19922
rect 17316 19858 17368 19864
rect 17316 19780 17368 19786
rect 17316 19722 17368 19728
rect 17222 18320 17278 18329
rect 17222 18255 17278 18264
rect 17328 17542 17356 19722
rect 17420 18834 17448 20998
rect 17682 20975 17738 20984
rect 17592 20800 17644 20806
rect 17592 20742 17644 20748
rect 17604 20398 17632 20742
rect 17592 20392 17644 20398
rect 17592 20334 17644 20340
rect 17604 19446 17632 20334
rect 17592 19440 17644 19446
rect 17592 19382 17644 19388
rect 17408 18828 17460 18834
rect 17408 18770 17460 18776
rect 17604 17864 17632 19382
rect 17420 17836 17632 17864
rect 17224 17536 17276 17542
rect 17224 17478 17276 17484
rect 17316 17536 17368 17542
rect 17316 17478 17368 17484
rect 17236 16130 17264 17478
rect 17328 17338 17356 17478
rect 17316 17332 17368 17338
rect 17316 17274 17368 17280
rect 17316 17060 17368 17066
rect 17316 17002 17368 17008
rect 17328 16250 17356 17002
rect 17316 16244 17368 16250
rect 17316 16186 17368 16192
rect 17236 16102 17356 16130
rect 17132 15496 17184 15502
rect 17132 15438 17184 15444
rect 17052 15320 17264 15348
rect 17132 15156 17184 15162
rect 17132 15098 17184 15104
rect 16948 13932 17000 13938
rect 16948 13874 17000 13880
rect 16580 13524 16632 13530
rect 16580 13466 16632 13472
rect 17040 13320 17092 13326
rect 17040 13262 17092 13268
rect 16396 13252 16448 13258
rect 16396 13194 16448 13200
rect 16408 12986 16436 13194
rect 16544 13084 16852 13093
rect 16544 13082 16550 13084
rect 16606 13082 16630 13084
rect 16686 13082 16710 13084
rect 16766 13082 16790 13084
rect 16846 13082 16852 13084
rect 16606 13030 16608 13082
rect 16788 13030 16790 13082
rect 16544 13028 16550 13030
rect 16606 13028 16630 13030
rect 16686 13028 16710 13030
rect 16766 13028 16790 13030
rect 16846 13028 16852 13030
rect 16544 13019 16852 13028
rect 16396 12980 16448 12986
rect 16396 12922 16448 12928
rect 16856 12844 16908 12850
rect 16856 12786 16908 12792
rect 16396 12368 16448 12374
rect 16396 12310 16448 12316
rect 16212 11756 16264 11762
rect 16212 11698 16264 11704
rect 16224 9654 16252 11698
rect 16408 11626 16436 12310
rect 16868 12306 16896 12786
rect 16948 12436 17000 12442
rect 16948 12378 17000 12384
rect 16856 12300 16908 12306
rect 16856 12242 16908 12248
rect 16544 11996 16852 12005
rect 16544 11994 16550 11996
rect 16606 11994 16630 11996
rect 16686 11994 16710 11996
rect 16766 11994 16790 11996
rect 16846 11994 16852 11996
rect 16606 11942 16608 11994
rect 16788 11942 16790 11994
rect 16544 11940 16550 11942
rect 16606 11940 16630 11942
rect 16686 11940 16710 11942
rect 16766 11940 16790 11942
rect 16846 11940 16852 11942
rect 16544 11931 16852 11940
rect 16580 11824 16632 11830
rect 16486 11792 16542 11801
rect 16580 11766 16632 11772
rect 16486 11727 16542 11736
rect 16396 11620 16448 11626
rect 16396 11562 16448 11568
rect 16500 11558 16528 11727
rect 16488 11552 16540 11558
rect 16488 11494 16540 11500
rect 16302 11384 16358 11393
rect 16358 11342 16436 11370
rect 16592 11354 16620 11766
rect 16302 11319 16358 11328
rect 16304 11076 16356 11082
rect 16304 11018 16356 11024
rect 16316 10305 16344 11018
rect 16302 10296 16358 10305
rect 16302 10231 16358 10240
rect 16408 10062 16436 11342
rect 16580 11348 16632 11354
rect 16580 11290 16632 11296
rect 16544 10908 16852 10917
rect 16544 10906 16550 10908
rect 16606 10906 16630 10908
rect 16686 10906 16710 10908
rect 16766 10906 16790 10908
rect 16846 10906 16852 10908
rect 16606 10854 16608 10906
rect 16788 10854 16790 10906
rect 16544 10852 16550 10854
rect 16606 10852 16630 10854
rect 16686 10852 16710 10854
rect 16766 10852 16790 10854
rect 16846 10852 16852 10854
rect 16544 10843 16852 10852
rect 16762 10160 16818 10169
rect 16762 10095 16764 10104
rect 16816 10095 16818 10104
rect 16764 10066 16816 10072
rect 16396 10056 16448 10062
rect 16396 9998 16448 10004
rect 16212 9648 16264 9654
rect 16212 9590 16264 9596
rect 16026 9551 16082 9560
rect 16120 9580 16172 9586
rect 16120 9522 16172 9528
rect 16304 9580 16356 9586
rect 16304 9522 16356 9528
rect 16212 9444 16264 9450
rect 16212 9386 16264 9392
rect 16224 8906 16252 9386
rect 16212 8900 16264 8906
rect 16212 8842 16264 8848
rect 15948 8758 16068 8786
rect 16040 7857 16068 8758
rect 16316 8430 16344 9522
rect 16408 8809 16436 9998
rect 16544 9820 16852 9829
rect 16544 9818 16550 9820
rect 16606 9818 16630 9820
rect 16686 9818 16710 9820
rect 16766 9818 16790 9820
rect 16846 9818 16852 9820
rect 16606 9766 16608 9818
rect 16788 9766 16790 9818
rect 16544 9764 16550 9766
rect 16606 9764 16630 9766
rect 16686 9764 16710 9766
rect 16766 9764 16790 9766
rect 16846 9764 16852 9766
rect 16544 9755 16852 9764
rect 16960 8922 16988 12378
rect 17052 11762 17080 13262
rect 17040 11756 17092 11762
rect 17040 11698 17092 11704
rect 17040 10804 17092 10810
rect 17040 10746 17092 10752
rect 17052 9058 17080 10746
rect 17144 9178 17172 15098
rect 17236 12238 17264 15320
rect 17328 14822 17356 16102
rect 17420 16046 17448 17836
rect 17500 17536 17552 17542
rect 17500 17478 17552 17484
rect 17696 17490 17724 20975
rect 17788 18766 17816 22120
rect 17880 21570 17908 24074
rect 17972 23254 18000 25622
rect 18064 24138 18092 26959
rect 18144 26920 18196 26926
rect 18144 26862 18196 26868
rect 18156 24954 18184 26862
rect 18248 26586 18276 32710
rect 18328 31816 18380 31822
rect 18328 31758 18380 31764
rect 18340 31482 18368 31758
rect 18328 31476 18380 31482
rect 18328 31418 18380 31424
rect 18328 30932 18380 30938
rect 18328 30874 18380 30880
rect 18340 29850 18368 30874
rect 18328 29844 18380 29850
rect 18328 29786 18380 29792
rect 18328 29708 18380 29714
rect 18328 29650 18380 29656
rect 18236 26580 18288 26586
rect 18236 26522 18288 26528
rect 18234 26208 18290 26217
rect 18234 26143 18290 26152
rect 18144 24948 18196 24954
rect 18144 24890 18196 24896
rect 18052 24132 18104 24138
rect 18052 24074 18104 24080
rect 17960 23248 18012 23254
rect 17960 23190 18012 23196
rect 18144 22976 18196 22982
rect 18144 22918 18196 22924
rect 18052 22772 18104 22778
rect 18052 22714 18104 22720
rect 17880 21542 18000 21570
rect 17868 21480 17920 21486
rect 17868 21422 17920 21428
rect 17880 20602 17908 21422
rect 17972 20942 18000 21542
rect 17960 20936 18012 20942
rect 17960 20878 18012 20884
rect 17868 20596 17920 20602
rect 17868 20538 17920 20544
rect 18064 19334 18092 22714
rect 18156 22642 18184 22918
rect 18144 22636 18196 22642
rect 18144 22578 18196 22584
rect 18156 21865 18184 22578
rect 18142 21856 18198 21865
rect 18142 21791 18198 21800
rect 18142 19408 18198 19417
rect 18142 19343 18198 19352
rect 17880 19306 18092 19334
rect 17776 18760 17828 18766
rect 17776 18702 17828 18708
rect 17880 17626 17908 19306
rect 17960 18692 18012 18698
rect 17960 18634 18012 18640
rect 17972 18358 18000 18634
rect 17960 18352 18012 18358
rect 17960 18294 18012 18300
rect 17788 17610 17908 17626
rect 17960 17672 18012 17678
rect 17960 17614 18012 17620
rect 17776 17604 17908 17610
rect 17828 17598 17908 17604
rect 17776 17546 17828 17552
rect 17868 17536 17920 17542
rect 17408 16040 17460 16046
rect 17408 15982 17460 15988
rect 17408 15904 17460 15910
rect 17408 15846 17460 15852
rect 17316 14816 17368 14822
rect 17316 14758 17368 14764
rect 17420 12356 17448 15846
rect 17512 14872 17540 17478
rect 17696 17462 17816 17490
rect 17868 17478 17920 17484
rect 17684 17332 17736 17338
rect 17684 17274 17736 17280
rect 17696 17218 17724 17274
rect 17604 17202 17724 17218
rect 17592 17196 17724 17202
rect 17644 17190 17724 17196
rect 17592 17138 17644 17144
rect 17684 17128 17736 17134
rect 17684 17070 17736 17076
rect 17696 16969 17724 17070
rect 17682 16960 17738 16969
rect 17682 16895 17738 16904
rect 17592 16584 17644 16590
rect 17788 16574 17816 17462
rect 17880 17134 17908 17478
rect 17866 17128 17918 17134
rect 17866 17070 17918 17076
rect 17972 16969 18000 17614
rect 17958 16960 18014 16969
rect 17958 16895 18014 16904
rect 17644 16546 17816 16574
rect 17592 16526 17644 16532
rect 17960 16244 18012 16250
rect 17960 16186 18012 16192
rect 17868 16040 17920 16046
rect 17868 15982 17920 15988
rect 17684 14952 17736 14958
rect 17684 14894 17736 14900
rect 17512 14844 17632 14872
rect 17604 12442 17632 14844
rect 17696 14482 17724 14894
rect 17684 14476 17736 14482
rect 17684 14418 17736 14424
rect 17592 12436 17644 12442
rect 17592 12378 17644 12384
rect 17328 12328 17448 12356
rect 17224 12232 17276 12238
rect 17224 12174 17276 12180
rect 17328 12152 17356 12328
rect 17696 12186 17724 14418
rect 17776 12844 17828 12850
rect 17776 12786 17828 12792
rect 17788 12374 17816 12786
rect 17776 12368 17828 12374
rect 17776 12310 17828 12316
rect 17880 12220 17908 15982
rect 17972 14278 18000 16186
rect 18052 15020 18104 15026
rect 18052 14962 18104 14968
rect 18064 14929 18092 14962
rect 18050 14920 18106 14929
rect 18050 14855 18106 14864
rect 18050 14376 18106 14385
rect 18050 14311 18106 14320
rect 17960 14272 18012 14278
rect 17960 14214 18012 14220
rect 17958 13696 18014 13705
rect 17958 13631 18014 13640
rect 17972 12782 18000 13631
rect 17960 12776 18012 12782
rect 17960 12718 18012 12724
rect 18064 12434 18092 14311
rect 17604 12158 17724 12186
rect 17788 12192 17908 12220
rect 17972 12406 18092 12434
rect 17328 12124 17448 12152
rect 17224 12096 17276 12102
rect 17224 12038 17276 12044
rect 17236 10606 17264 12038
rect 17316 11756 17368 11762
rect 17316 11698 17368 11704
rect 17328 10810 17356 11698
rect 17316 10804 17368 10810
rect 17316 10746 17368 10752
rect 17224 10600 17276 10606
rect 17224 10542 17276 10548
rect 17224 9376 17276 9382
rect 17224 9318 17276 9324
rect 17236 9178 17264 9318
rect 17132 9172 17184 9178
rect 17132 9114 17184 9120
rect 17224 9172 17276 9178
rect 17224 9114 17276 9120
rect 17052 9030 17264 9058
rect 17236 8974 17264 9030
rect 17132 8968 17184 8974
rect 17130 8936 17132 8945
rect 17224 8968 17276 8974
rect 17184 8936 17186 8945
rect 16960 8894 17080 8922
rect 16948 8832 17000 8838
rect 16394 8800 16450 8809
rect 16948 8774 17000 8780
rect 16394 8735 16450 8744
rect 16544 8732 16852 8741
rect 16544 8730 16550 8732
rect 16606 8730 16630 8732
rect 16686 8730 16710 8732
rect 16766 8730 16790 8732
rect 16846 8730 16852 8732
rect 16606 8678 16608 8730
rect 16788 8678 16790 8730
rect 16544 8676 16550 8678
rect 16606 8676 16630 8678
rect 16686 8676 16710 8678
rect 16766 8676 16790 8678
rect 16846 8676 16852 8678
rect 16544 8667 16852 8676
rect 16304 8424 16356 8430
rect 16304 8366 16356 8372
rect 16764 8424 16816 8430
rect 16816 8384 16896 8412
rect 16764 8366 16816 8372
rect 16304 8288 16356 8294
rect 16304 8230 16356 8236
rect 16672 8288 16724 8294
rect 16672 8230 16724 8236
rect 16316 7954 16344 8230
rect 16304 7948 16356 7954
rect 16304 7890 16356 7896
rect 16026 7848 16082 7857
rect 15936 7812 15988 7818
rect 16026 7783 16082 7792
rect 16212 7812 16264 7818
rect 15936 7754 15988 7760
rect 16212 7754 16264 7760
rect 15580 6956 15700 6984
rect 15764 7398 15884 7426
rect 15476 5908 15528 5914
rect 15476 5850 15528 5856
rect 15396 5766 15516 5794
rect 15292 5636 15344 5642
rect 15292 5578 15344 5584
rect 15304 5030 15332 5578
rect 15382 5128 15438 5137
rect 15382 5063 15438 5072
rect 15292 5024 15344 5030
rect 15292 4966 15344 4972
rect 15200 4820 15252 4826
rect 15200 4762 15252 4768
rect 15108 4276 15160 4282
rect 15108 4218 15160 4224
rect 14924 4140 14976 4146
rect 15028 4134 15148 4162
rect 14924 4082 14976 4088
rect 15016 4072 15068 4078
rect 15016 4014 15068 4020
rect 14740 3528 14792 3534
rect 14740 3470 14792 3476
rect 14832 3528 14884 3534
rect 14832 3470 14884 3476
rect 14648 3460 14700 3466
rect 14648 3402 14700 3408
rect 14464 3392 14516 3398
rect 14464 3334 14516 3340
rect 14556 3392 14608 3398
rect 14556 3334 14608 3340
rect 14924 3392 14976 3398
rect 14924 3334 14976 3340
rect 14096 3188 14148 3194
rect 14096 3130 14148 3136
rect 14370 3088 14426 3097
rect 14476 3074 14504 3334
rect 14568 3194 14596 3334
rect 14556 3188 14608 3194
rect 14556 3130 14608 3136
rect 14476 3046 14596 3074
rect 14370 3023 14372 3032
rect 14424 3023 14426 3032
rect 14372 2994 14424 3000
rect 14464 2984 14516 2990
rect 13818 2952 13874 2961
rect 14464 2926 14516 2932
rect 13818 2887 13874 2896
rect 13832 2854 13860 2887
rect 13820 2848 13872 2854
rect 13820 2790 13872 2796
rect 14372 2848 14424 2854
rect 14372 2790 14424 2796
rect 13945 2748 14253 2757
rect 13945 2746 13951 2748
rect 14007 2746 14031 2748
rect 14087 2746 14111 2748
rect 14167 2746 14191 2748
rect 14247 2746 14253 2748
rect 14007 2694 14009 2746
rect 14189 2694 14191 2746
rect 13945 2692 13951 2694
rect 14007 2692 14031 2694
rect 14087 2692 14111 2694
rect 14167 2692 14191 2694
rect 14247 2692 14253 2694
rect 13945 2683 14253 2692
rect 14384 2417 14412 2790
rect 14370 2408 14426 2417
rect 14370 2343 14426 2352
rect 14476 1986 14504 2926
rect 14568 2689 14596 3046
rect 14740 3052 14792 3058
rect 14740 2994 14792 3000
rect 14832 3052 14884 3058
rect 14832 2994 14884 3000
rect 14752 2961 14780 2994
rect 14738 2952 14794 2961
rect 14738 2887 14794 2896
rect 14740 2848 14792 2854
rect 14740 2790 14792 2796
rect 14554 2680 14610 2689
rect 14554 2615 14610 2624
rect 14476 1958 14596 1986
rect 14464 1896 14516 1902
rect 14464 1838 14516 1844
rect 14372 1828 14424 1834
rect 14372 1770 14424 1776
rect 14096 1760 14148 1766
rect 13832 1720 14096 1748
rect 13832 1442 13860 1720
rect 14096 1702 14148 1708
rect 13945 1660 14253 1669
rect 13945 1658 13951 1660
rect 14007 1658 14031 1660
rect 14087 1658 14111 1660
rect 14167 1658 14191 1660
rect 14247 1658 14253 1660
rect 14007 1606 14009 1658
rect 14189 1606 14191 1658
rect 13945 1604 13951 1606
rect 14007 1604 14031 1606
rect 14087 1604 14111 1606
rect 14167 1604 14191 1606
rect 14247 1604 14253 1606
rect 13945 1595 14253 1604
rect 14384 1544 14412 1770
rect 14292 1516 14412 1544
rect 13832 1414 13952 1442
rect 13820 1352 13872 1358
rect 13740 1312 13820 1340
rect 13820 1294 13872 1300
rect 13728 1216 13780 1222
rect 13728 1158 13780 1164
rect 13740 678 13768 1158
rect 13924 898 13952 1414
rect 14004 1420 14056 1426
rect 14004 1362 14056 1368
rect 13832 870 13952 898
rect 13728 672 13780 678
rect 13728 614 13780 620
rect 13832 160 13860 870
rect 14016 160 14044 1362
rect 11794 82 11850 160
rect 11716 54 11850 82
rect 11794 -300 11850 54
rect 11978 -300 12034 160
rect 12162 -300 12218 160
rect 12346 -300 12402 160
rect 12530 -300 12586 160
rect 12714 -300 12770 160
rect 12898 -300 12954 160
rect 13082 -300 13138 160
rect 13266 -300 13322 160
rect 13450 -300 13506 160
rect 13634 -300 13690 160
rect 13818 -300 13874 160
rect 14002 -300 14058 160
rect 14186 82 14242 160
rect 14292 82 14320 1516
rect 14370 1456 14426 1465
rect 14370 1391 14426 1400
rect 14384 160 14412 1391
rect 14476 1018 14504 1838
rect 14568 1737 14596 1958
rect 14648 1828 14700 1834
rect 14648 1770 14700 1776
rect 14554 1728 14610 1737
rect 14554 1663 14610 1672
rect 14660 1306 14688 1770
rect 14752 1358 14780 2790
rect 14844 2650 14872 2994
rect 14832 2644 14884 2650
rect 14832 2586 14884 2592
rect 14936 1970 14964 3334
rect 15028 3194 15056 4014
rect 15120 3534 15148 4134
rect 15200 4140 15252 4146
rect 15200 4082 15252 4088
rect 15212 3738 15240 4082
rect 15200 3732 15252 3738
rect 15200 3674 15252 3680
rect 15396 3618 15424 5063
rect 15488 4026 15516 5766
rect 15580 5710 15608 6956
rect 15660 6792 15712 6798
rect 15660 6734 15712 6740
rect 15672 6458 15700 6734
rect 15660 6452 15712 6458
rect 15660 6394 15712 6400
rect 15660 6316 15712 6322
rect 15660 6258 15712 6264
rect 15672 6186 15700 6258
rect 15660 6180 15712 6186
rect 15660 6122 15712 6128
rect 15764 5953 15792 7398
rect 15844 7336 15896 7342
rect 15948 7324 15976 7754
rect 16028 7744 16080 7750
rect 16224 7698 16252 7754
rect 16028 7686 16080 7692
rect 16040 7546 16068 7686
rect 16132 7670 16252 7698
rect 16132 7546 16160 7670
rect 16028 7540 16080 7546
rect 16028 7482 16080 7488
rect 16120 7540 16172 7546
rect 16316 7528 16344 7890
rect 16684 7886 16712 8230
rect 16868 8106 16896 8384
rect 16960 8294 16988 8774
rect 16948 8288 17000 8294
rect 16948 8230 17000 8236
rect 16868 8078 16988 8106
rect 16672 7880 16724 7886
rect 16672 7822 16724 7828
rect 16960 7818 16988 8078
rect 16948 7812 17000 7818
rect 16948 7754 17000 7760
rect 16544 7644 16852 7653
rect 16544 7642 16550 7644
rect 16606 7642 16630 7644
rect 16686 7642 16710 7644
rect 16766 7642 16790 7644
rect 16846 7642 16852 7644
rect 16606 7590 16608 7642
rect 16788 7590 16790 7642
rect 16544 7588 16550 7590
rect 16606 7588 16630 7590
rect 16686 7588 16710 7590
rect 16766 7588 16790 7590
rect 16846 7588 16852 7590
rect 16120 7482 16172 7488
rect 16224 7500 16344 7528
rect 16394 7576 16450 7585
rect 16544 7579 16852 7588
rect 16394 7511 16450 7520
rect 15896 7296 15976 7324
rect 15844 7278 15896 7284
rect 16028 7268 16080 7274
rect 16028 7210 16080 7216
rect 15844 7200 15896 7206
rect 15844 7142 15896 7148
rect 15856 7002 15884 7142
rect 15844 6996 15896 7002
rect 15844 6938 15896 6944
rect 16040 6934 16068 7210
rect 16028 6928 16080 6934
rect 16028 6870 16080 6876
rect 16028 6452 16080 6458
rect 16028 6394 16080 6400
rect 15844 6316 15896 6322
rect 15844 6258 15896 6264
rect 15750 5944 15806 5953
rect 15856 5914 15884 6258
rect 15750 5879 15806 5888
rect 15844 5908 15896 5914
rect 15844 5850 15896 5856
rect 15568 5704 15620 5710
rect 15568 5646 15620 5652
rect 15752 5704 15804 5710
rect 15752 5646 15804 5652
rect 15580 5545 15608 5646
rect 15660 5636 15712 5642
rect 15660 5578 15712 5584
rect 15566 5536 15622 5545
rect 15566 5471 15622 5480
rect 15568 5364 15620 5370
rect 15568 5306 15620 5312
rect 15580 5114 15608 5306
rect 15672 5250 15700 5578
rect 15764 5370 15792 5646
rect 15752 5364 15804 5370
rect 15752 5306 15804 5312
rect 15844 5364 15896 5370
rect 15844 5306 15896 5312
rect 15856 5250 15884 5306
rect 15672 5222 15884 5250
rect 15936 5228 15988 5234
rect 15936 5170 15988 5176
rect 15580 5086 15884 5114
rect 15856 5030 15884 5086
rect 15844 5024 15896 5030
rect 15948 5001 15976 5170
rect 15844 4966 15896 4972
rect 15934 4992 15990 5001
rect 15934 4927 15990 4936
rect 16040 4842 16068 6394
rect 16120 5772 16172 5778
rect 16224 5760 16252 7500
rect 16304 7404 16356 7410
rect 16304 7346 16356 7352
rect 16316 6730 16344 7346
rect 16408 7274 16436 7511
rect 16396 7268 16448 7274
rect 16396 7210 16448 7216
rect 16304 6724 16356 6730
rect 16304 6666 16356 6672
rect 16172 5732 16252 5760
rect 16120 5714 16172 5720
rect 16120 5568 16172 5574
rect 16120 5510 16172 5516
rect 16212 5568 16264 5574
rect 16212 5510 16264 5516
rect 16132 5166 16160 5510
rect 16120 5160 16172 5166
rect 16120 5102 16172 5108
rect 16224 4842 16252 5510
rect 16316 5284 16344 6666
rect 16960 6662 16988 7754
rect 17052 7449 17080 8894
rect 17224 8910 17276 8916
rect 17130 8871 17186 8880
rect 17132 8832 17184 8838
rect 17132 8774 17184 8780
rect 17038 7440 17094 7449
rect 17144 7410 17172 8774
rect 17420 7970 17448 12124
rect 17604 12102 17632 12158
rect 17592 12096 17644 12102
rect 17498 12064 17554 12073
rect 17592 12038 17644 12044
rect 17684 12096 17736 12102
rect 17684 12038 17736 12044
rect 17498 11999 17554 12008
rect 17328 7942 17448 7970
rect 17224 7744 17276 7750
rect 17224 7686 17276 7692
rect 17236 7546 17264 7686
rect 17224 7540 17276 7546
rect 17224 7482 17276 7488
rect 17038 7375 17094 7384
rect 17132 7404 17184 7410
rect 17132 7346 17184 7352
rect 16948 6656 17000 6662
rect 16948 6598 17000 6604
rect 16544 6556 16852 6565
rect 16544 6554 16550 6556
rect 16606 6554 16630 6556
rect 16686 6554 16710 6556
rect 16766 6554 16790 6556
rect 16846 6554 16852 6556
rect 16606 6502 16608 6554
rect 16788 6502 16790 6554
rect 16544 6500 16550 6502
rect 16606 6500 16630 6502
rect 16686 6500 16710 6502
rect 16766 6500 16790 6502
rect 16846 6500 16852 6502
rect 16544 6491 16852 6500
rect 16544 5468 16852 5477
rect 16544 5466 16550 5468
rect 16606 5466 16630 5468
rect 16686 5466 16710 5468
rect 16766 5466 16790 5468
rect 16846 5466 16852 5468
rect 16606 5414 16608 5466
rect 16788 5414 16790 5466
rect 16544 5412 16550 5414
rect 16606 5412 16630 5414
rect 16686 5412 16710 5414
rect 16766 5412 16790 5414
rect 16846 5412 16852 5414
rect 16544 5403 16852 5412
rect 16580 5364 16632 5370
rect 16960 5352 16988 6598
rect 17040 6316 17092 6322
rect 17040 6258 17092 6264
rect 17052 5914 17080 6258
rect 17132 6248 17184 6254
rect 17132 6190 17184 6196
rect 17144 5914 17172 6190
rect 17040 5908 17092 5914
rect 17040 5850 17092 5856
rect 17132 5908 17184 5914
rect 17132 5850 17184 5856
rect 17040 5636 17092 5642
rect 17040 5578 17092 5584
rect 16580 5306 16632 5312
rect 16684 5324 16988 5352
rect 16316 5256 16528 5284
rect 16396 5160 16448 5166
rect 16396 5102 16448 5108
rect 15948 4814 16068 4842
rect 16132 4814 16252 4842
rect 16304 4820 16356 4826
rect 15566 4720 15622 4729
rect 15566 4655 15622 4664
rect 15580 4146 15608 4655
rect 15948 4622 15976 4814
rect 16132 4706 16160 4814
rect 16408 4808 16436 5102
rect 16356 4780 16436 4808
rect 16304 4762 16356 4768
rect 16500 4758 16528 5256
rect 16040 4678 16160 4706
rect 16488 4752 16540 4758
rect 16488 4694 16540 4700
rect 15936 4616 15988 4622
rect 15936 4558 15988 4564
rect 16040 4282 16068 4678
rect 16212 4616 16264 4622
rect 16118 4584 16174 4593
rect 16212 4558 16264 4564
rect 16396 4616 16448 4622
rect 16592 4604 16620 5306
rect 16684 5166 16712 5324
rect 16764 5228 16816 5234
rect 16764 5170 16816 5176
rect 16672 5160 16724 5166
rect 16672 5102 16724 5108
rect 16684 4690 16712 5102
rect 16672 4684 16724 4690
rect 16672 4626 16724 4632
rect 16776 4622 16804 5170
rect 16856 4820 16908 4826
rect 16856 4762 16908 4768
rect 16448 4576 16620 4604
rect 16764 4616 16816 4622
rect 16396 4558 16448 4564
rect 16764 4558 16816 4564
rect 16118 4519 16174 4528
rect 16028 4276 16080 4282
rect 16028 4218 16080 4224
rect 16132 4146 16160 4519
rect 15568 4140 15620 4146
rect 15568 4082 15620 4088
rect 16028 4140 16080 4146
rect 16028 4082 16080 4088
rect 16120 4140 16172 4146
rect 16120 4082 16172 4088
rect 15658 4040 15714 4049
rect 15488 3998 15608 4026
rect 15212 3590 15424 3618
rect 15474 3632 15530 3641
rect 15212 3534 15240 3590
rect 15474 3567 15530 3576
rect 15108 3528 15160 3534
rect 15108 3470 15160 3476
rect 15200 3528 15252 3534
rect 15200 3470 15252 3476
rect 15292 3460 15344 3466
rect 15292 3402 15344 3408
rect 15200 3392 15252 3398
rect 15200 3334 15252 3340
rect 15106 3224 15162 3233
rect 15016 3188 15068 3194
rect 15106 3159 15162 3168
rect 15016 3130 15068 3136
rect 15016 2916 15068 2922
rect 15016 2858 15068 2864
rect 14924 1964 14976 1970
rect 14924 1906 14976 1912
rect 14922 1592 14978 1601
rect 14844 1550 14922 1578
rect 14568 1278 14688 1306
rect 14740 1352 14792 1358
rect 14740 1294 14792 1300
rect 14464 1012 14516 1018
rect 14464 954 14516 960
rect 14568 160 14596 1278
rect 14186 54 14320 82
rect 14186 -300 14242 54
rect 14370 -300 14426 160
rect 14554 -300 14610 160
rect 14738 82 14794 160
rect 14844 82 14872 1550
rect 14922 1527 14978 1536
rect 14924 1488 14976 1494
rect 14924 1430 14976 1436
rect 14936 160 14964 1430
rect 14738 54 14872 82
rect 14738 -300 14794 54
rect 14922 -300 14978 160
rect 15028 82 15056 2858
rect 15120 2514 15148 3159
rect 15212 3058 15240 3334
rect 15200 3052 15252 3058
rect 15200 2994 15252 3000
rect 15108 2508 15160 2514
rect 15108 2450 15160 2456
rect 15108 2304 15160 2310
rect 15108 2246 15160 2252
rect 15120 1426 15148 2246
rect 15200 2032 15252 2038
rect 15200 1974 15252 1980
rect 15212 1562 15240 1974
rect 15200 1556 15252 1562
rect 15200 1498 15252 1504
rect 15108 1420 15160 1426
rect 15108 1362 15160 1368
rect 15304 160 15332 3402
rect 15384 3188 15436 3194
rect 15384 3130 15436 3136
rect 15396 2446 15424 3130
rect 15488 3058 15516 3567
rect 15580 3534 15608 3998
rect 15658 3975 15714 3984
rect 15672 3534 15700 3975
rect 15752 3936 15804 3942
rect 16040 3913 16068 4082
rect 15752 3878 15804 3884
rect 16026 3904 16082 3913
rect 15764 3641 15792 3878
rect 16026 3839 16082 3848
rect 15844 3664 15896 3670
rect 15750 3632 15806 3641
rect 15844 3606 15896 3612
rect 15750 3567 15806 3576
rect 15568 3528 15620 3534
rect 15568 3470 15620 3476
rect 15660 3528 15712 3534
rect 15660 3470 15712 3476
rect 15752 3392 15804 3398
rect 15752 3334 15804 3340
rect 15476 3052 15528 3058
rect 15476 2994 15528 3000
rect 15476 2848 15528 2854
rect 15476 2790 15528 2796
rect 15384 2440 15436 2446
rect 15384 2382 15436 2388
rect 15488 2038 15516 2790
rect 15568 2644 15620 2650
rect 15568 2586 15620 2592
rect 15660 2644 15712 2650
rect 15660 2586 15712 2592
rect 15476 2032 15528 2038
rect 15476 1974 15528 1980
rect 15384 1352 15436 1358
rect 15384 1294 15436 1300
rect 15396 921 15424 1294
rect 15382 912 15438 921
rect 15382 847 15438 856
rect 15106 82 15162 160
rect 15028 54 15162 82
rect 15106 -300 15162 54
rect 15290 -300 15346 160
rect 15474 82 15530 160
rect 15580 82 15608 2586
rect 15672 160 15700 2586
rect 15764 2038 15792 3334
rect 15856 3233 15884 3606
rect 15936 3528 15988 3534
rect 15936 3470 15988 3476
rect 15842 3224 15898 3233
rect 15842 3159 15898 3168
rect 15948 3126 15976 3470
rect 15936 3120 15988 3126
rect 15936 3062 15988 3068
rect 15844 2916 15896 2922
rect 15844 2858 15896 2864
rect 15948 2910 16160 2938
rect 15752 2032 15804 2038
rect 15752 1974 15804 1980
rect 15752 1760 15804 1766
rect 15752 1702 15804 1708
rect 15764 1601 15792 1702
rect 15750 1592 15806 1601
rect 15750 1527 15806 1536
rect 15856 160 15884 2858
rect 15948 1426 15976 2910
rect 16028 2848 16080 2854
rect 16132 2825 16160 2910
rect 16028 2790 16080 2796
rect 16118 2816 16174 2825
rect 15936 1420 15988 1426
rect 15936 1362 15988 1368
rect 16040 160 16068 2790
rect 16118 2751 16174 2760
rect 16118 2680 16174 2689
rect 16118 2615 16174 2624
rect 16132 2514 16160 2615
rect 16120 2508 16172 2514
rect 16120 2450 16172 2456
rect 16120 2304 16172 2310
rect 16120 2246 16172 2252
rect 16132 1494 16160 2246
rect 16120 1488 16172 1494
rect 16120 1430 16172 1436
rect 16224 160 16252 4558
rect 16672 4548 16724 4554
rect 16592 4508 16672 4536
rect 16304 4480 16356 4486
rect 16302 4448 16304 4457
rect 16592 4468 16620 4508
rect 16672 4490 16724 4496
rect 16868 4486 16896 4762
rect 17052 4758 17080 5578
rect 17040 4752 17092 4758
rect 17040 4694 17092 4700
rect 17040 4616 17092 4622
rect 17040 4558 17092 4564
rect 16356 4448 16358 4457
rect 16302 4383 16358 4392
rect 16408 4440 16620 4468
rect 16856 4480 16908 4486
rect 16304 3936 16356 3942
rect 16304 3878 16356 3884
rect 16316 3505 16344 3878
rect 16408 3738 16436 4440
rect 16856 4422 16908 4428
rect 16544 4380 16852 4389
rect 16544 4378 16550 4380
rect 16606 4378 16630 4380
rect 16686 4378 16710 4380
rect 16766 4378 16790 4380
rect 16846 4378 16852 4380
rect 16606 4326 16608 4378
rect 16788 4326 16790 4378
rect 16544 4324 16550 4326
rect 16606 4324 16630 4326
rect 16686 4324 16710 4326
rect 16766 4324 16790 4326
rect 16846 4324 16852 4326
rect 16544 4315 16852 4324
rect 17052 4298 17080 4558
rect 17144 4554 17172 5850
rect 17224 5636 17276 5642
rect 17224 5578 17276 5584
rect 17236 4622 17264 5578
rect 17224 4616 17276 4622
rect 17224 4558 17276 4564
rect 17132 4548 17184 4554
rect 17132 4490 17184 4496
rect 17222 4448 17278 4457
rect 17222 4383 17278 4392
rect 16960 4270 17080 4298
rect 17236 4282 17264 4383
rect 17224 4276 17276 4282
rect 16500 4236 16712 4264
rect 16500 4146 16528 4236
rect 16488 4140 16540 4146
rect 16488 4082 16540 4088
rect 16580 4140 16632 4146
rect 16580 4082 16632 4088
rect 16396 3732 16448 3738
rect 16396 3674 16448 3680
rect 16592 3602 16620 4082
rect 16684 3720 16712 4236
rect 16764 4072 16816 4078
rect 16816 4032 16896 4060
rect 16764 4014 16816 4020
rect 16868 3890 16896 4032
rect 16960 4010 16988 4270
rect 17224 4218 17276 4224
rect 17224 4140 17276 4146
rect 17224 4082 17276 4088
rect 16948 4004 17000 4010
rect 16948 3946 17000 3952
rect 16868 3862 17172 3890
rect 16684 3692 17080 3720
rect 16580 3596 16632 3602
rect 16580 3538 16632 3544
rect 16488 3528 16540 3534
rect 16302 3496 16358 3505
rect 16540 3476 16804 3482
rect 16488 3470 16804 3476
rect 16500 3454 16804 3470
rect 16302 3431 16358 3440
rect 16776 3398 16804 3454
rect 16396 3392 16448 3398
rect 16302 3360 16358 3369
rect 16396 3334 16448 3340
rect 16764 3392 16816 3398
rect 16764 3334 16816 3340
rect 16302 3295 16358 3304
rect 16316 3058 16344 3295
rect 16304 3052 16356 3058
rect 16304 2994 16356 3000
rect 16304 1420 16356 1426
rect 16304 1362 16356 1368
rect 15474 54 15608 82
rect 15474 -300 15530 54
rect 15658 -300 15714 160
rect 15842 -300 15898 160
rect 16026 -300 16082 160
rect 16210 -300 16266 160
rect 16316 82 16344 1362
rect 16408 1358 16436 3334
rect 16544 3292 16852 3301
rect 16544 3290 16550 3292
rect 16606 3290 16630 3292
rect 16686 3290 16710 3292
rect 16766 3290 16790 3292
rect 16846 3290 16852 3292
rect 16606 3238 16608 3290
rect 16788 3238 16790 3290
rect 16544 3236 16550 3238
rect 16606 3236 16630 3238
rect 16686 3236 16710 3238
rect 16766 3236 16790 3238
rect 16846 3236 16852 3238
rect 16544 3227 16852 3236
rect 16578 2680 16634 2689
rect 16578 2615 16634 2624
rect 16592 2582 16620 2615
rect 16580 2576 16632 2582
rect 16580 2518 16632 2524
rect 16544 2204 16852 2213
rect 16544 2202 16550 2204
rect 16606 2202 16630 2204
rect 16686 2202 16710 2204
rect 16766 2202 16790 2204
rect 16846 2202 16852 2204
rect 16606 2150 16608 2202
rect 16788 2150 16790 2202
rect 16544 2148 16550 2150
rect 16606 2148 16630 2150
rect 16686 2148 16710 2150
rect 16766 2148 16790 2150
rect 16846 2148 16852 2150
rect 16544 2139 16852 2148
rect 17052 2038 17080 3692
rect 17144 2106 17172 3862
rect 17236 2922 17264 4082
rect 17328 3602 17356 7942
rect 17512 7834 17540 11999
rect 17590 11928 17646 11937
rect 17590 11863 17646 11872
rect 17420 7806 17540 7834
rect 17420 3670 17448 7806
rect 17500 7744 17552 7750
rect 17500 7686 17552 7692
rect 17512 7546 17540 7686
rect 17500 7540 17552 7546
rect 17500 7482 17552 7488
rect 17498 6624 17554 6633
rect 17604 6610 17632 11863
rect 17696 11354 17724 12038
rect 17684 11348 17736 11354
rect 17684 11290 17736 11296
rect 17788 11234 17816 12192
rect 17868 11552 17920 11558
rect 17868 11494 17920 11500
rect 17696 11206 17816 11234
rect 17696 10033 17724 11206
rect 17880 11150 17908 11494
rect 17776 11144 17828 11150
rect 17776 11086 17828 11092
rect 17868 11144 17920 11150
rect 17868 11086 17920 11092
rect 17788 10810 17816 11086
rect 17972 10996 18000 12406
rect 18156 11098 18184 19343
rect 17880 10968 18000 10996
rect 18064 11070 18184 11098
rect 17776 10804 17828 10810
rect 17776 10746 17828 10752
rect 17682 10024 17738 10033
rect 17682 9959 17738 9968
rect 17684 9920 17736 9926
rect 17684 9862 17736 9868
rect 17696 8566 17724 9862
rect 17788 9518 17816 10746
rect 17776 9512 17828 9518
rect 17776 9454 17828 9460
rect 17684 8560 17736 8566
rect 17684 8502 17736 8508
rect 17684 8016 17736 8022
rect 17684 7958 17736 7964
rect 17696 6746 17724 7958
rect 17788 7886 17816 9454
rect 17880 8022 17908 10968
rect 18064 10266 18092 11070
rect 18144 11008 18196 11014
rect 18144 10950 18196 10956
rect 18052 10260 18104 10266
rect 18052 10202 18104 10208
rect 18156 10198 18184 10950
rect 18144 10192 18196 10198
rect 18144 10134 18196 10140
rect 18144 10056 18196 10062
rect 18144 9998 18196 10004
rect 18052 9580 18104 9586
rect 18052 9522 18104 9528
rect 17960 9172 18012 9178
rect 17960 9114 18012 9120
rect 17972 8974 18000 9114
rect 18064 9058 18092 9522
rect 18156 9178 18184 9998
rect 18144 9172 18196 9178
rect 18144 9114 18196 9120
rect 18064 9030 18184 9058
rect 17960 8968 18012 8974
rect 17960 8910 18012 8916
rect 17958 8528 18014 8537
rect 17958 8463 17960 8472
rect 18012 8463 18014 8472
rect 17960 8434 18012 8440
rect 17960 8084 18012 8090
rect 17960 8026 18012 8032
rect 17868 8016 17920 8022
rect 17868 7958 17920 7964
rect 17776 7880 17828 7886
rect 17776 7822 17828 7828
rect 17972 7546 18000 8026
rect 18052 8016 18104 8022
rect 18052 7958 18104 7964
rect 18064 7857 18092 7958
rect 18050 7848 18106 7857
rect 18050 7783 18106 7792
rect 17960 7540 18012 7546
rect 17960 7482 18012 7488
rect 18052 7540 18104 7546
rect 18052 7482 18104 7488
rect 18064 7426 18092 7482
rect 17880 7398 18092 7426
rect 17774 7304 17830 7313
rect 17774 7239 17830 7248
rect 17788 7206 17816 7239
rect 17776 7200 17828 7206
rect 17776 7142 17828 7148
rect 17696 6718 17816 6746
rect 17604 6582 17724 6610
rect 17498 6559 17554 6568
rect 17512 6458 17540 6559
rect 17500 6452 17552 6458
rect 17500 6394 17552 6400
rect 17500 6316 17552 6322
rect 17500 6258 17552 6264
rect 17512 4826 17540 6258
rect 17592 5772 17644 5778
rect 17592 5714 17644 5720
rect 17604 5370 17632 5714
rect 17696 5370 17724 6582
rect 17592 5364 17644 5370
rect 17592 5306 17644 5312
rect 17684 5364 17736 5370
rect 17684 5306 17736 5312
rect 17684 5024 17736 5030
rect 17684 4966 17736 4972
rect 17500 4820 17552 4826
rect 17500 4762 17552 4768
rect 17500 4548 17552 4554
rect 17500 4490 17552 4496
rect 17408 3664 17460 3670
rect 17408 3606 17460 3612
rect 17316 3596 17368 3602
rect 17316 3538 17368 3544
rect 17408 3528 17460 3534
rect 17408 3470 17460 3476
rect 17420 3369 17448 3470
rect 17406 3360 17462 3369
rect 17406 3295 17462 3304
rect 17224 2916 17276 2922
rect 17224 2858 17276 2864
rect 17224 2440 17276 2446
rect 17224 2382 17276 2388
rect 17132 2100 17184 2106
rect 17132 2042 17184 2048
rect 17040 2032 17092 2038
rect 16868 1970 16988 1986
rect 17040 1974 17092 1980
rect 16856 1964 16988 1970
rect 16908 1958 16988 1964
rect 16856 1906 16908 1912
rect 16856 1556 16908 1562
rect 16856 1498 16908 1504
rect 16868 1465 16896 1498
rect 16854 1456 16910 1465
rect 16854 1391 16910 1400
rect 16396 1352 16448 1358
rect 16396 1294 16448 1300
rect 16544 1116 16852 1125
rect 16544 1114 16550 1116
rect 16606 1114 16630 1116
rect 16686 1114 16710 1116
rect 16766 1114 16790 1116
rect 16846 1114 16852 1116
rect 16606 1062 16608 1114
rect 16788 1062 16790 1114
rect 16544 1060 16550 1062
rect 16606 1060 16630 1062
rect 16686 1060 16710 1062
rect 16766 1060 16790 1062
rect 16846 1060 16852 1062
rect 16544 1051 16852 1060
rect 16960 490 16988 1958
rect 17132 1964 17184 1970
rect 17132 1906 17184 1912
rect 17040 1896 17092 1902
rect 17040 1838 17092 1844
rect 17052 1737 17080 1838
rect 17038 1728 17094 1737
rect 17038 1663 17094 1672
rect 17040 1284 17092 1290
rect 17040 1226 17092 1232
rect 16684 462 16988 490
rect 16394 82 16450 160
rect 16316 54 16450 82
rect 16394 -300 16450 54
rect 16578 82 16634 160
rect 16684 82 16712 462
rect 17052 354 17080 1226
rect 16868 326 17080 354
rect 16578 54 16712 82
rect 16762 82 16818 160
rect 16868 82 16896 326
rect 17144 218 17172 1906
rect 16960 190 17172 218
rect 16960 160 16988 190
rect 16762 54 16896 82
rect 16578 -300 16634 54
rect 16762 -300 16818 54
rect 16946 -300 17002 160
rect 17130 82 17186 160
rect 17236 82 17264 2382
rect 17408 1216 17460 1222
rect 17328 1176 17408 1204
rect 17328 160 17356 1176
rect 17408 1158 17460 1164
rect 17512 1018 17540 4490
rect 17592 4480 17644 4486
rect 17592 4422 17644 4428
rect 17604 4214 17632 4422
rect 17696 4282 17724 4966
rect 17684 4276 17736 4282
rect 17684 4218 17736 4224
rect 17592 4208 17644 4214
rect 17592 4150 17644 4156
rect 17604 3482 17632 4150
rect 17788 3602 17816 6718
rect 17880 5522 17908 7398
rect 18052 7336 18104 7342
rect 18052 7278 18104 7284
rect 18064 7002 18092 7278
rect 18052 6996 18104 7002
rect 18052 6938 18104 6944
rect 18052 6656 18104 6662
rect 18052 6598 18104 6604
rect 18064 5914 18092 6598
rect 18052 5908 18104 5914
rect 18052 5850 18104 5856
rect 17880 5494 18000 5522
rect 17868 5364 17920 5370
rect 17868 5306 17920 5312
rect 17880 4554 17908 5306
rect 17868 4548 17920 4554
rect 17868 4490 17920 4496
rect 17868 4140 17920 4146
rect 17868 4082 17920 4088
rect 17880 3738 17908 4082
rect 17868 3732 17920 3738
rect 17868 3674 17920 3680
rect 17776 3596 17828 3602
rect 17776 3538 17828 3544
rect 17868 3596 17920 3602
rect 17868 3538 17920 3544
rect 17880 3482 17908 3538
rect 17604 3454 17908 3482
rect 17972 3058 18000 5494
rect 18156 5370 18184 9030
rect 18248 7546 18276 26143
rect 18340 24596 18368 29650
rect 18432 24721 18460 35119
rect 18524 31754 18552 35634
rect 18708 35578 18736 39494
rect 18880 39432 18932 39438
rect 19352 39409 19380 39510
rect 19536 39438 19564 39879
rect 19628 39642 19656 40462
rect 19708 40044 19760 40050
rect 19708 39986 19760 39992
rect 19616 39636 19668 39642
rect 19616 39578 19668 39584
rect 19720 39522 19748 39986
rect 19812 39896 19840 40598
rect 19904 40089 19932 41074
rect 19996 41070 20024 42162
rect 20456 41834 20484 42162
rect 20272 41806 20484 41834
rect 20548 41818 20576 43007
rect 20536 41812 20588 41818
rect 20168 41132 20220 41138
rect 20168 41074 20220 41080
rect 19984 41064 20036 41070
rect 19984 41006 20036 41012
rect 20076 40520 20128 40526
rect 20076 40462 20128 40468
rect 20088 40168 20116 40462
rect 19996 40140 20116 40168
rect 19890 40080 19946 40089
rect 19890 40015 19946 40024
rect 19892 39908 19944 39914
rect 19812 39868 19892 39896
rect 19892 39850 19944 39856
rect 19628 39506 19748 39522
rect 19616 39500 19748 39506
rect 19668 39494 19748 39500
rect 19616 39442 19668 39448
rect 19524 39432 19576 39438
rect 18880 39374 18932 39380
rect 19338 39400 19394 39409
rect 18788 39364 18840 39370
rect 18788 39306 18840 39312
rect 18800 39098 18828 39306
rect 18788 39092 18840 39098
rect 18788 39034 18840 39040
rect 18788 37868 18840 37874
rect 18788 37810 18840 37816
rect 18616 35550 18736 35578
rect 18616 34513 18644 35550
rect 18800 34746 18828 37810
rect 18788 34740 18840 34746
rect 18788 34682 18840 34688
rect 18602 34504 18658 34513
rect 18602 34439 18658 34448
rect 18604 34400 18656 34406
rect 18604 34342 18656 34348
rect 18616 34066 18644 34342
rect 18604 34060 18656 34066
rect 18604 34002 18656 34008
rect 18892 33538 18920 39374
rect 19524 39374 19576 39380
rect 19708 39432 19760 39438
rect 19708 39374 19760 39380
rect 19800 39432 19852 39438
rect 19800 39374 19852 39380
rect 19338 39335 19394 39344
rect 19720 39273 19748 39374
rect 19706 39264 19762 39273
rect 19706 39199 19762 39208
rect 19812 38962 19840 39374
rect 18972 38956 19024 38962
rect 18972 38898 19024 38904
rect 19800 38956 19852 38962
rect 19800 38898 19852 38904
rect 18984 38554 19012 38898
rect 19143 38652 19451 38661
rect 19996 38654 20024 40140
rect 20180 39098 20208 41074
rect 20272 40633 20300 41806
rect 20536 41754 20588 41760
rect 20626 41712 20682 41721
rect 20626 41647 20682 41656
rect 20352 41608 20404 41614
rect 20352 41550 20404 41556
rect 20258 40624 20314 40633
rect 20258 40559 20314 40568
rect 20260 40384 20312 40390
rect 20260 40326 20312 40332
rect 20272 40186 20300 40326
rect 20364 40186 20392 41550
rect 20442 41304 20498 41313
rect 20442 41239 20498 41248
rect 20456 41138 20484 41239
rect 20444 41132 20496 41138
rect 20444 41074 20496 41080
rect 20444 40724 20496 40730
rect 20444 40666 20496 40672
rect 20260 40180 20312 40186
rect 20260 40122 20312 40128
rect 20352 40180 20404 40186
rect 20352 40122 20404 40128
rect 20352 39432 20404 39438
rect 20352 39374 20404 39380
rect 20364 39098 20392 39374
rect 20456 39370 20484 40666
rect 20536 40384 20588 40390
rect 20536 40326 20588 40332
rect 20444 39364 20496 39370
rect 20444 39306 20496 39312
rect 20548 39273 20576 40326
rect 20534 39264 20590 39273
rect 20534 39199 20590 39208
rect 20168 39092 20220 39098
rect 20168 39034 20220 39040
rect 20352 39092 20404 39098
rect 20352 39034 20404 39040
rect 20260 38956 20312 38962
rect 20260 38898 20312 38904
rect 20272 38729 20300 38898
rect 20258 38720 20314 38729
rect 20258 38655 20314 38664
rect 19143 38650 19149 38652
rect 19205 38650 19229 38652
rect 19285 38650 19309 38652
rect 19365 38650 19389 38652
rect 19445 38650 19451 38652
rect 19205 38598 19207 38650
rect 19387 38598 19389 38650
rect 19143 38596 19149 38598
rect 19205 38596 19229 38598
rect 19285 38596 19309 38598
rect 19365 38596 19389 38598
rect 19445 38596 19451 38598
rect 19143 38587 19451 38596
rect 19904 38626 20024 38654
rect 18972 38548 19024 38554
rect 18972 38490 19024 38496
rect 19708 37800 19760 37806
rect 19708 37742 19760 37748
rect 19143 37564 19451 37573
rect 19143 37562 19149 37564
rect 19205 37562 19229 37564
rect 19285 37562 19309 37564
rect 19365 37562 19389 37564
rect 19445 37562 19451 37564
rect 19205 37510 19207 37562
rect 19387 37510 19389 37562
rect 19143 37508 19149 37510
rect 19205 37508 19229 37510
rect 19285 37508 19309 37510
rect 19365 37508 19389 37510
rect 19445 37508 19451 37510
rect 19143 37499 19451 37508
rect 19720 37466 19748 37742
rect 19708 37460 19760 37466
rect 19708 37402 19760 37408
rect 19708 37256 19760 37262
rect 19708 37198 19760 37204
rect 19616 36780 19668 36786
rect 19616 36722 19668 36728
rect 19143 36476 19451 36485
rect 19143 36474 19149 36476
rect 19205 36474 19229 36476
rect 19285 36474 19309 36476
rect 19365 36474 19389 36476
rect 19445 36474 19451 36476
rect 19205 36422 19207 36474
rect 19387 36422 19389 36474
rect 19143 36420 19149 36422
rect 19205 36420 19229 36422
rect 19285 36420 19309 36422
rect 19365 36420 19389 36422
rect 19445 36420 19451 36422
rect 19143 36411 19451 36420
rect 19430 36272 19486 36281
rect 19352 36242 19430 36258
rect 19340 36236 19430 36242
rect 19392 36230 19430 36236
rect 19430 36207 19486 36216
rect 19340 36178 19392 36184
rect 18972 36168 19024 36174
rect 18972 36110 19024 36116
rect 18984 35766 19012 36110
rect 19064 36032 19116 36038
rect 19064 35974 19116 35980
rect 18972 35760 19024 35766
rect 18972 35702 19024 35708
rect 19076 35086 19104 35974
rect 19524 35692 19576 35698
rect 19524 35634 19576 35640
rect 19143 35388 19451 35397
rect 19143 35386 19149 35388
rect 19205 35386 19229 35388
rect 19285 35386 19309 35388
rect 19365 35386 19389 35388
rect 19445 35386 19451 35388
rect 19205 35334 19207 35386
rect 19387 35334 19389 35386
rect 19143 35332 19149 35334
rect 19205 35332 19229 35334
rect 19285 35332 19309 35334
rect 19365 35332 19389 35334
rect 19445 35332 19451 35334
rect 19143 35323 19451 35332
rect 19064 35080 19116 35086
rect 19064 35022 19116 35028
rect 19536 34746 19564 35634
rect 19628 34950 19656 36722
rect 19720 36582 19748 37198
rect 19904 36666 19932 38626
rect 19982 38584 20038 38593
rect 19982 38519 20038 38528
rect 19996 38486 20024 38519
rect 19984 38480 20036 38486
rect 19984 38422 20036 38428
rect 20168 38344 20220 38350
rect 20444 38344 20496 38350
rect 20168 38286 20220 38292
rect 20258 38312 20314 38321
rect 20180 38010 20208 38286
rect 20444 38286 20496 38292
rect 20258 38247 20314 38256
rect 20168 38004 20220 38010
rect 20168 37946 20220 37952
rect 20076 37868 20128 37874
rect 20076 37810 20128 37816
rect 20168 37868 20220 37874
rect 20168 37810 20220 37816
rect 20088 37777 20116 37810
rect 20074 37768 20130 37777
rect 20074 37703 20130 37712
rect 20180 37466 20208 37810
rect 20168 37460 20220 37466
rect 20168 37402 20220 37408
rect 20074 36816 20130 36825
rect 20074 36751 20130 36760
rect 19982 36680 20038 36689
rect 19800 36644 19852 36650
rect 19904 36638 19982 36666
rect 19982 36615 20038 36624
rect 19800 36586 19852 36592
rect 19708 36576 19760 36582
rect 19708 36518 19760 36524
rect 19720 36310 19748 36518
rect 19708 36304 19760 36310
rect 19708 36246 19760 36252
rect 19708 36168 19760 36174
rect 19708 36110 19760 36116
rect 19720 35834 19748 36110
rect 19708 35828 19760 35834
rect 19708 35770 19760 35776
rect 19708 35284 19760 35290
rect 19708 35226 19760 35232
rect 19616 34944 19668 34950
rect 19616 34886 19668 34892
rect 19524 34740 19576 34746
rect 19524 34682 19576 34688
rect 19143 34300 19451 34309
rect 19143 34298 19149 34300
rect 19205 34298 19229 34300
rect 19285 34298 19309 34300
rect 19365 34298 19389 34300
rect 19445 34298 19451 34300
rect 19205 34246 19207 34298
rect 19387 34246 19389 34298
rect 19143 34244 19149 34246
rect 19205 34244 19229 34246
rect 19285 34244 19309 34246
rect 19365 34244 19389 34246
rect 19445 34244 19451 34246
rect 19143 34235 19451 34244
rect 19432 33992 19484 33998
rect 19720 33946 19748 35226
rect 19432 33934 19484 33940
rect 19156 33924 19208 33930
rect 19156 33866 19208 33872
rect 19168 33658 19196 33866
rect 19156 33652 19208 33658
rect 19156 33594 19208 33600
rect 19338 33552 19394 33561
rect 18892 33510 19012 33538
rect 18880 33448 18932 33454
rect 18880 33390 18932 33396
rect 18892 33114 18920 33390
rect 18880 33108 18932 33114
rect 18880 33050 18932 33056
rect 18880 32904 18932 32910
rect 18984 32881 19012 33510
rect 19338 33487 19340 33496
rect 19392 33487 19394 33496
rect 19340 33458 19392 33464
rect 19444 33402 19472 33934
rect 19628 33918 19748 33946
rect 19444 33374 19564 33402
rect 19143 33212 19451 33221
rect 19143 33210 19149 33212
rect 19205 33210 19229 33212
rect 19285 33210 19309 33212
rect 19365 33210 19389 33212
rect 19445 33210 19451 33212
rect 19205 33158 19207 33210
rect 19387 33158 19389 33210
rect 19143 33156 19149 33158
rect 19205 33156 19229 33158
rect 19285 33156 19309 33158
rect 19365 33156 19389 33158
rect 19445 33156 19451 33158
rect 19143 33147 19451 33156
rect 19156 32904 19208 32910
rect 18880 32846 18932 32852
rect 18970 32872 19026 32881
rect 18788 32768 18840 32774
rect 18708 32728 18788 32756
rect 18524 31726 18644 31754
rect 18512 31680 18564 31686
rect 18512 31622 18564 31628
rect 18524 30938 18552 31622
rect 18616 31414 18644 31726
rect 18604 31408 18656 31414
rect 18604 31350 18656 31356
rect 18512 30932 18564 30938
rect 18512 30874 18564 30880
rect 18512 29844 18564 29850
rect 18512 29786 18564 29792
rect 18524 29306 18552 29786
rect 18512 29300 18564 29306
rect 18512 29242 18564 29248
rect 18512 29164 18564 29170
rect 18512 29106 18564 29112
rect 18524 27441 18552 29106
rect 18510 27432 18566 27441
rect 18510 27367 18566 27376
rect 18512 26240 18564 26246
rect 18512 26182 18564 26188
rect 18524 25906 18552 26182
rect 18616 26042 18644 31350
rect 18604 26036 18656 26042
rect 18604 25978 18656 25984
rect 18512 25900 18564 25906
rect 18512 25842 18564 25848
rect 18708 25702 18736 32728
rect 18788 32710 18840 32716
rect 18788 32360 18840 32366
rect 18788 32302 18840 32308
rect 18800 30666 18828 32302
rect 18892 32026 18920 32846
rect 18970 32807 19026 32816
rect 19076 32852 19156 32858
rect 19076 32846 19208 32852
rect 19076 32830 19196 32846
rect 18972 32428 19024 32434
rect 18972 32370 19024 32376
rect 18880 32020 18932 32026
rect 18880 31962 18932 31968
rect 18984 31822 19012 32370
rect 18972 31816 19024 31822
rect 18972 31758 19024 31764
rect 18880 31340 18932 31346
rect 18880 31282 18932 31288
rect 18892 30841 18920 31282
rect 18972 31272 19024 31278
rect 18972 31214 19024 31220
rect 18878 30832 18934 30841
rect 18878 30767 18934 30776
rect 18880 30728 18932 30734
rect 18880 30670 18932 30676
rect 18788 30660 18840 30666
rect 18788 30602 18840 30608
rect 18788 30388 18840 30394
rect 18788 30330 18840 30336
rect 18696 25696 18748 25702
rect 18696 25638 18748 25644
rect 18512 25288 18564 25294
rect 18564 25236 18736 25242
rect 18512 25230 18736 25236
rect 18524 25214 18736 25230
rect 18604 25152 18656 25158
rect 18604 25094 18656 25100
rect 18616 24818 18644 25094
rect 18708 24818 18736 25214
rect 18604 24812 18656 24818
rect 18604 24754 18656 24760
rect 18696 24812 18748 24818
rect 18696 24754 18748 24760
rect 18418 24712 18474 24721
rect 18418 24647 18474 24656
rect 18340 24568 18644 24596
rect 18512 23248 18564 23254
rect 18512 23190 18564 23196
rect 18420 23180 18472 23186
rect 18420 23122 18472 23128
rect 18328 22976 18380 22982
rect 18328 22918 18380 22924
rect 18340 22030 18368 22918
rect 18328 22024 18380 22030
rect 18328 21966 18380 21972
rect 18432 19854 18460 23122
rect 18524 22001 18552 23190
rect 18510 21992 18566 22001
rect 18510 21927 18566 21936
rect 18616 21010 18644 24568
rect 18708 24410 18736 24754
rect 18696 24404 18748 24410
rect 18696 24346 18748 24352
rect 18800 22094 18828 30330
rect 18892 27033 18920 30670
rect 18984 30394 19012 31214
rect 19076 30920 19104 32830
rect 19536 32434 19564 33374
rect 19628 32434 19656 33918
rect 19708 33856 19760 33862
rect 19708 33798 19760 33804
rect 19720 33658 19748 33798
rect 19708 33652 19760 33658
rect 19708 33594 19760 33600
rect 19812 33538 19840 36586
rect 19984 36576 20036 36582
rect 19984 36518 20036 36524
rect 19892 36304 19944 36310
rect 19892 36246 19944 36252
rect 19904 34746 19932 36246
rect 19892 34740 19944 34746
rect 19892 34682 19944 34688
rect 19892 33992 19944 33998
rect 19892 33934 19944 33940
rect 19904 33658 19932 33934
rect 19892 33652 19944 33658
rect 19892 33594 19944 33600
rect 19708 33516 19760 33522
rect 19812 33510 19932 33538
rect 19708 33458 19760 33464
rect 19720 32842 19748 33458
rect 19904 33318 19932 33510
rect 19892 33312 19944 33318
rect 19892 33254 19944 33260
rect 19708 32836 19760 32842
rect 19708 32778 19760 32784
rect 19996 32774 20024 36518
rect 19984 32768 20036 32774
rect 19984 32710 20036 32716
rect 20088 32586 20116 36751
rect 20166 35864 20222 35873
rect 20166 35799 20222 35808
rect 20180 34746 20208 35799
rect 20168 34740 20220 34746
rect 20168 34682 20220 34688
rect 20168 34604 20220 34610
rect 20168 34546 20220 34552
rect 20180 33266 20208 34546
rect 20272 33930 20300 38247
rect 20456 37466 20484 38286
rect 20444 37460 20496 37466
rect 20444 37402 20496 37408
rect 20444 37256 20496 37262
rect 20444 37198 20496 37204
rect 20536 37256 20588 37262
rect 20536 37198 20588 37204
rect 20352 36780 20404 36786
rect 20352 36722 20404 36728
rect 20364 35290 20392 36722
rect 20456 36718 20484 37198
rect 20548 36825 20576 37198
rect 20534 36816 20590 36825
rect 20534 36751 20590 36760
rect 20444 36712 20496 36718
rect 20444 36654 20496 36660
rect 20534 36680 20590 36689
rect 20534 36615 20590 36624
rect 20442 36272 20498 36281
rect 20442 36207 20498 36216
rect 20456 36174 20484 36207
rect 20444 36168 20496 36174
rect 20444 36110 20496 36116
rect 20444 36032 20496 36038
rect 20444 35974 20496 35980
rect 20456 35873 20484 35974
rect 20442 35864 20498 35873
rect 20442 35799 20498 35808
rect 20444 35692 20496 35698
rect 20444 35634 20496 35640
rect 20352 35284 20404 35290
rect 20352 35226 20404 35232
rect 20456 34746 20484 35634
rect 20548 35086 20576 36615
rect 20536 35080 20588 35086
rect 20536 35022 20588 35028
rect 20444 34740 20496 34746
rect 20444 34682 20496 34688
rect 20444 34604 20496 34610
rect 20444 34546 20496 34552
rect 20456 34202 20484 34546
rect 20444 34196 20496 34202
rect 20444 34138 20496 34144
rect 20640 34082 20668 41647
rect 20732 40730 20760 43318
rect 20996 43308 21048 43314
rect 20996 43250 21048 43256
rect 20904 42220 20956 42226
rect 20904 42162 20956 42168
rect 20812 42084 20864 42090
rect 20812 42026 20864 42032
rect 20824 41138 20852 42026
rect 20916 41177 20944 42162
rect 20902 41168 20958 41177
rect 20812 41132 20864 41138
rect 20902 41103 20958 41112
rect 20812 41074 20864 41080
rect 21008 41002 21036 43250
rect 21640 43240 21692 43246
rect 21640 43182 21692 43188
rect 21364 42628 21416 42634
rect 21364 42570 21416 42576
rect 21088 41608 21140 41614
rect 21088 41550 21140 41556
rect 20904 40996 20956 41002
rect 20904 40938 20956 40944
rect 20996 40996 21048 41002
rect 20996 40938 21048 40944
rect 20720 40724 20772 40730
rect 20720 40666 20772 40672
rect 20720 40520 20772 40526
rect 20720 40462 20772 40468
rect 20812 40520 20864 40526
rect 20812 40462 20864 40468
rect 20732 39642 20760 40462
rect 20720 39636 20772 39642
rect 20720 39578 20772 39584
rect 20824 39438 20852 40462
rect 20916 40338 20944 40938
rect 20916 40310 21036 40338
rect 20902 40216 20958 40225
rect 20902 40151 20958 40160
rect 20916 40118 20944 40151
rect 20904 40112 20956 40118
rect 20904 40054 20956 40060
rect 21008 39914 21036 40310
rect 21100 40168 21128 41550
rect 21180 41540 21232 41546
rect 21180 41482 21232 41488
rect 21192 40662 21220 41482
rect 21272 41132 21324 41138
rect 21272 41074 21324 41080
rect 21284 40730 21312 41074
rect 21272 40724 21324 40730
rect 21272 40666 21324 40672
rect 21180 40656 21232 40662
rect 21180 40598 21232 40604
rect 21272 40520 21324 40526
rect 21272 40462 21324 40468
rect 21100 40140 21220 40168
rect 21088 40044 21140 40050
rect 21088 39986 21140 39992
rect 20996 39908 21048 39914
rect 20996 39850 21048 39856
rect 20812 39432 20864 39438
rect 20812 39374 20864 39380
rect 20996 39432 21048 39438
rect 20996 39374 21048 39380
rect 20720 39364 20772 39370
rect 20720 39306 20772 39312
rect 20732 39098 20760 39306
rect 20812 39296 20864 39302
rect 20812 39238 20864 39244
rect 20824 39098 20852 39238
rect 20720 39092 20772 39098
rect 20720 39034 20772 39040
rect 20812 39092 20864 39098
rect 20812 39034 20864 39040
rect 20720 38956 20772 38962
rect 20720 38898 20772 38904
rect 20904 38956 20956 38962
rect 20904 38898 20956 38904
rect 20732 38554 20760 38898
rect 20720 38548 20772 38554
rect 20720 38490 20772 38496
rect 20720 38344 20772 38350
rect 20720 38286 20772 38292
rect 20812 38344 20864 38350
rect 20812 38286 20864 38292
rect 20732 38010 20760 38286
rect 20720 38004 20772 38010
rect 20720 37946 20772 37952
rect 20720 37868 20772 37874
rect 20720 37810 20772 37816
rect 20732 37466 20760 37810
rect 20824 37806 20852 38286
rect 20812 37800 20864 37806
rect 20812 37742 20864 37748
rect 20916 37738 20944 38898
rect 21008 38554 21036 39374
rect 21100 38593 21128 39986
rect 21192 39409 21220 40140
rect 21284 39642 21312 40462
rect 21376 39982 21404 42570
rect 21548 42152 21600 42158
rect 21548 42094 21600 42100
rect 21456 41744 21508 41750
rect 21456 41686 21508 41692
rect 21364 39976 21416 39982
rect 21364 39918 21416 39924
rect 21468 39930 21496 41686
rect 21560 41274 21588 42094
rect 21548 41268 21600 41274
rect 21548 41210 21600 41216
rect 21652 41154 21680 43182
rect 22190 42528 22246 42537
rect 21742 42460 22050 42469
rect 22190 42463 22246 42472
rect 21742 42458 21748 42460
rect 21804 42458 21828 42460
rect 21884 42458 21908 42460
rect 21964 42458 21988 42460
rect 22044 42458 22050 42460
rect 21804 42406 21806 42458
rect 21986 42406 21988 42458
rect 21742 42404 21748 42406
rect 21804 42404 21828 42406
rect 21884 42404 21908 42406
rect 21964 42404 21988 42406
rect 22044 42404 22050 42406
rect 21742 42395 22050 42404
rect 22204 42362 22232 42463
rect 22388 42362 22416 43551
rect 22192 42356 22244 42362
rect 22192 42298 22244 42304
rect 22376 42356 22428 42362
rect 22376 42298 22428 42304
rect 21914 41984 21970 41993
rect 21914 41919 21970 41928
rect 21928 41818 21956 41919
rect 21916 41812 21968 41818
rect 21916 41754 21968 41760
rect 22652 41676 22704 41682
rect 22652 41618 22704 41624
rect 22284 41540 22336 41546
rect 22284 41482 22336 41488
rect 22296 41449 22324 41482
rect 22560 41472 22612 41478
rect 22282 41440 22338 41449
rect 22560 41414 22612 41420
rect 21742 41372 22050 41381
rect 22282 41375 22338 41384
rect 21742 41370 21748 41372
rect 21804 41370 21828 41372
rect 21884 41370 21908 41372
rect 21964 41370 21988 41372
rect 22044 41370 22050 41372
rect 21804 41318 21806 41370
rect 21986 41318 21988 41370
rect 21742 41316 21748 41318
rect 21804 41316 21828 41318
rect 21884 41316 21908 41318
rect 21964 41316 21988 41318
rect 22044 41316 22050 41318
rect 21742 41307 22050 41316
rect 21560 41126 21680 41154
rect 21560 40361 21588 41126
rect 21640 41064 21692 41070
rect 21640 41006 21692 41012
rect 21546 40352 21602 40361
rect 21546 40287 21602 40296
rect 21468 39902 21588 39930
rect 21456 39840 21508 39846
rect 21454 39808 21456 39817
rect 21508 39808 21510 39817
rect 21454 39743 21510 39752
rect 21272 39636 21324 39642
rect 21272 39578 21324 39584
rect 21178 39400 21234 39409
rect 21178 39335 21234 39344
rect 21180 38752 21232 38758
rect 21456 38752 21508 38758
rect 21180 38694 21232 38700
rect 21454 38720 21456 38729
rect 21508 38720 21510 38729
rect 21086 38584 21142 38593
rect 20996 38548 21048 38554
rect 21086 38519 21142 38528
rect 20996 38490 21048 38496
rect 21088 38208 21140 38214
rect 21088 38150 21140 38156
rect 20996 37868 21048 37874
rect 20996 37810 21048 37816
rect 20904 37732 20956 37738
rect 20904 37674 20956 37680
rect 20812 37664 20864 37670
rect 20812 37606 20864 37612
rect 20720 37460 20772 37466
rect 20720 37402 20772 37408
rect 20824 36922 20852 37606
rect 20904 37256 20956 37262
rect 20904 37198 20956 37204
rect 20812 36916 20864 36922
rect 20812 36858 20864 36864
rect 20812 36780 20864 36786
rect 20812 36722 20864 36728
rect 20824 36122 20852 36722
rect 20916 36666 20944 37198
rect 21008 36922 21036 37810
rect 21100 37262 21128 38150
rect 21192 37874 21220 38694
rect 21454 38655 21510 38664
rect 21180 37868 21232 37874
rect 21180 37810 21232 37816
rect 21456 37664 21508 37670
rect 21454 37632 21456 37641
rect 21508 37632 21510 37641
rect 21454 37567 21510 37576
rect 21088 37256 21140 37262
rect 21088 37198 21140 37204
rect 21088 37120 21140 37126
rect 21088 37062 21140 37068
rect 20996 36916 21048 36922
rect 20996 36858 21048 36864
rect 20916 36638 21036 36666
rect 20904 36576 20956 36582
rect 20904 36518 20956 36524
rect 20732 36094 20852 36122
rect 20732 35562 20760 36094
rect 20812 36032 20864 36038
rect 20812 35974 20864 35980
rect 20720 35556 20772 35562
rect 20720 35498 20772 35504
rect 20720 34740 20772 34746
rect 20720 34682 20772 34688
rect 20456 34054 20668 34082
rect 20352 33992 20404 33998
rect 20352 33934 20404 33940
rect 20260 33924 20312 33930
rect 20260 33866 20312 33872
rect 20364 33522 20392 33934
rect 20352 33516 20404 33522
rect 20352 33458 20404 33464
rect 20456 33402 20484 34054
rect 20732 33998 20760 34682
rect 20824 34678 20852 35974
rect 20916 35086 20944 36518
rect 21008 36310 21036 36638
rect 20996 36304 21048 36310
rect 20996 36246 21048 36252
rect 21100 35698 21128 37062
rect 21456 36576 21508 36582
rect 21454 36544 21456 36553
rect 21508 36544 21510 36553
rect 21454 36479 21510 36488
rect 21180 36372 21232 36378
rect 21180 36314 21232 36320
rect 20996 35692 21048 35698
rect 20996 35634 21048 35640
rect 21088 35692 21140 35698
rect 21088 35634 21140 35640
rect 21008 35578 21036 35634
rect 21008 35550 21128 35578
rect 20996 35488 21048 35494
rect 20996 35430 21048 35436
rect 20904 35080 20956 35086
rect 20904 35022 20956 35028
rect 20812 34672 20864 34678
rect 20812 34614 20864 34620
rect 20904 34604 20956 34610
rect 20904 34546 20956 34552
rect 20628 33992 20680 33998
rect 20628 33934 20680 33940
rect 20720 33992 20772 33998
rect 20720 33934 20772 33940
rect 20536 33924 20588 33930
rect 20536 33866 20588 33872
rect 20364 33374 20484 33402
rect 20180 33238 20300 33266
rect 19812 32558 20116 32586
rect 19432 32428 19484 32434
rect 19432 32370 19484 32376
rect 19524 32428 19576 32434
rect 19524 32370 19576 32376
rect 19616 32428 19668 32434
rect 19616 32370 19668 32376
rect 19444 32212 19472 32370
rect 19444 32184 19564 32212
rect 19143 32124 19451 32133
rect 19143 32122 19149 32124
rect 19205 32122 19229 32124
rect 19285 32122 19309 32124
rect 19365 32122 19389 32124
rect 19445 32122 19451 32124
rect 19205 32070 19207 32122
rect 19387 32070 19389 32122
rect 19143 32068 19149 32070
rect 19205 32068 19229 32070
rect 19285 32068 19309 32070
rect 19365 32068 19389 32070
rect 19445 32068 19451 32070
rect 19143 32059 19451 32068
rect 19143 31036 19451 31045
rect 19143 31034 19149 31036
rect 19205 31034 19229 31036
rect 19285 31034 19309 31036
rect 19365 31034 19389 31036
rect 19445 31034 19451 31036
rect 19205 30982 19207 31034
rect 19387 30982 19389 31034
rect 19143 30980 19149 30982
rect 19205 30980 19229 30982
rect 19285 30980 19309 30982
rect 19365 30980 19389 30982
rect 19445 30980 19451 30982
rect 19143 30971 19451 30980
rect 19536 30954 19564 32184
rect 19516 30926 19564 30954
rect 19516 30920 19544 30926
rect 19076 30892 19196 30920
rect 19168 30734 19196 30892
rect 19444 30892 19544 30920
rect 19156 30728 19208 30734
rect 19154 30696 19156 30705
rect 19208 30696 19210 30705
rect 19064 30660 19116 30666
rect 19154 30631 19210 30640
rect 19064 30602 19116 30608
rect 18972 30388 19024 30394
rect 18972 30330 19024 30336
rect 19076 30138 19104 30602
rect 18984 30110 19104 30138
rect 18984 29238 19012 30110
rect 19064 30048 19116 30054
rect 19444 30036 19472 30892
rect 19524 30252 19576 30258
rect 19628 30240 19656 32370
rect 19708 32224 19760 32230
rect 19708 32166 19760 32172
rect 19720 31890 19748 32166
rect 19812 31906 19840 32558
rect 19984 32496 20036 32502
rect 19984 32438 20036 32444
rect 20076 32496 20128 32502
rect 20076 32438 20128 32444
rect 19892 32224 19944 32230
rect 19892 32166 19944 32172
rect 19904 32026 19932 32166
rect 19996 32026 20024 32438
rect 19892 32020 19944 32026
rect 19892 31962 19944 31968
rect 19984 32020 20036 32026
rect 19984 31962 20036 31968
rect 20088 31929 20116 32438
rect 20074 31920 20130 31929
rect 19708 31884 19760 31890
rect 19812 31878 19932 31906
rect 19708 31826 19760 31832
rect 19800 31816 19852 31822
rect 19800 31758 19852 31764
rect 19708 31748 19760 31754
rect 19708 31690 19760 31696
rect 19720 31482 19748 31690
rect 19708 31476 19760 31482
rect 19708 31418 19760 31424
rect 19708 31340 19760 31346
rect 19708 31282 19760 31288
rect 19720 30666 19748 31282
rect 19812 30734 19840 31758
rect 19800 30728 19852 30734
rect 19800 30670 19852 30676
rect 19708 30660 19760 30666
rect 19708 30602 19760 30608
rect 19576 30212 19656 30240
rect 19800 30252 19852 30258
rect 19524 30194 19576 30200
rect 19800 30194 19852 30200
rect 19444 30008 19564 30036
rect 19064 29990 19116 29996
rect 19076 29850 19104 29990
rect 19143 29948 19451 29957
rect 19143 29946 19149 29948
rect 19205 29946 19229 29948
rect 19285 29946 19309 29948
rect 19365 29946 19389 29948
rect 19445 29946 19451 29948
rect 19205 29894 19207 29946
rect 19387 29894 19389 29946
rect 19143 29892 19149 29894
rect 19205 29892 19229 29894
rect 19285 29892 19309 29894
rect 19365 29892 19389 29894
rect 19445 29892 19451 29894
rect 19143 29883 19451 29892
rect 19064 29844 19116 29850
rect 19064 29786 19116 29792
rect 18972 29232 19024 29238
rect 18972 29174 19024 29180
rect 19536 29102 19564 30008
rect 19708 29572 19760 29578
rect 19708 29514 19760 29520
rect 19720 29102 19748 29514
rect 19524 29096 19576 29102
rect 19708 29096 19760 29102
rect 19576 29056 19656 29084
rect 19524 29038 19576 29044
rect 19524 28960 19576 28966
rect 18970 28928 19026 28937
rect 19524 28902 19576 28908
rect 19628 28914 19656 29056
rect 19708 29038 19760 29044
rect 18970 28863 19026 28872
rect 18878 27024 18934 27033
rect 18878 26959 18934 26968
rect 18880 26784 18932 26790
rect 18880 26726 18932 26732
rect 18892 25838 18920 26726
rect 18880 25832 18932 25838
rect 18880 25774 18932 25780
rect 18892 25378 18920 25774
rect 18984 25480 19012 28863
rect 19143 28860 19451 28869
rect 19143 28858 19149 28860
rect 19205 28858 19229 28860
rect 19285 28858 19309 28860
rect 19365 28858 19389 28860
rect 19445 28858 19451 28860
rect 19205 28806 19207 28858
rect 19387 28806 19389 28858
rect 19143 28804 19149 28806
rect 19205 28804 19229 28806
rect 19285 28804 19309 28806
rect 19365 28804 19389 28806
rect 19445 28804 19451 28806
rect 19143 28795 19451 28804
rect 19340 28552 19392 28558
rect 19536 28506 19564 28902
rect 19628 28886 19748 28914
rect 19340 28494 19392 28500
rect 19352 28218 19380 28494
rect 19444 28490 19564 28506
rect 19432 28484 19564 28490
rect 19484 28478 19564 28484
rect 19432 28426 19484 28432
rect 19524 28416 19576 28422
rect 19524 28358 19576 28364
rect 19616 28416 19668 28422
rect 19616 28358 19668 28364
rect 19340 28212 19392 28218
rect 19340 28154 19392 28160
rect 19064 27940 19116 27946
rect 19064 27882 19116 27888
rect 19076 27538 19104 27882
rect 19143 27772 19451 27781
rect 19143 27770 19149 27772
rect 19205 27770 19229 27772
rect 19285 27770 19309 27772
rect 19365 27770 19389 27772
rect 19445 27770 19451 27772
rect 19205 27718 19207 27770
rect 19387 27718 19389 27770
rect 19143 27716 19149 27718
rect 19205 27716 19229 27718
rect 19285 27716 19309 27718
rect 19365 27716 19389 27718
rect 19445 27716 19451 27718
rect 19143 27707 19451 27716
rect 19536 27674 19564 28358
rect 19628 28218 19656 28358
rect 19616 28212 19668 28218
rect 19616 28154 19668 28160
rect 19616 28076 19668 28082
rect 19616 28018 19668 28024
rect 19628 27985 19656 28018
rect 19614 27976 19670 27985
rect 19614 27911 19670 27920
rect 19616 27872 19668 27878
rect 19616 27814 19668 27820
rect 19524 27668 19576 27674
rect 19524 27610 19576 27616
rect 19064 27532 19116 27538
rect 19064 27474 19116 27480
rect 19628 27402 19656 27814
rect 19616 27396 19668 27402
rect 19616 27338 19668 27344
rect 19143 26684 19451 26693
rect 19143 26682 19149 26684
rect 19205 26682 19229 26684
rect 19285 26682 19309 26684
rect 19365 26682 19389 26684
rect 19445 26682 19451 26684
rect 19205 26630 19207 26682
rect 19387 26630 19389 26682
rect 19143 26628 19149 26630
rect 19205 26628 19229 26630
rect 19285 26628 19309 26630
rect 19365 26628 19389 26630
rect 19445 26628 19451 26630
rect 19143 26619 19451 26628
rect 19524 26376 19576 26382
rect 19524 26318 19576 26324
rect 19156 26308 19208 26314
rect 19156 26250 19208 26256
rect 19168 26042 19196 26250
rect 19156 26036 19208 26042
rect 19156 25978 19208 25984
rect 19143 25596 19451 25605
rect 19143 25594 19149 25596
rect 19205 25594 19229 25596
rect 19285 25594 19309 25596
rect 19365 25594 19389 25596
rect 19445 25594 19451 25596
rect 19205 25542 19207 25594
rect 19387 25542 19389 25594
rect 19143 25540 19149 25542
rect 19205 25540 19229 25542
rect 19285 25540 19309 25542
rect 19365 25540 19389 25542
rect 19445 25540 19451 25542
rect 19143 25531 19451 25540
rect 19536 25498 19564 26318
rect 19720 26042 19748 28886
rect 19812 28694 19840 30194
rect 19800 28688 19852 28694
rect 19800 28630 19852 28636
rect 19800 27872 19852 27878
rect 19800 27814 19852 27820
rect 19812 26382 19840 27814
rect 19904 27062 19932 31878
rect 20074 31855 20130 31864
rect 20088 31754 20116 31855
rect 20088 31726 20208 31754
rect 20076 31680 20128 31686
rect 20076 31622 20128 31628
rect 19982 31376 20038 31385
rect 19982 31311 20038 31320
rect 19996 29646 20024 31311
rect 19984 29640 20036 29646
rect 19984 29582 20036 29588
rect 19984 29164 20036 29170
rect 19984 29106 20036 29112
rect 19892 27056 19944 27062
rect 19892 26998 19944 27004
rect 19800 26376 19852 26382
rect 19800 26318 19852 26324
rect 19890 26344 19946 26353
rect 19890 26279 19946 26288
rect 19800 26240 19852 26246
rect 19800 26182 19852 26188
rect 19708 26036 19760 26042
rect 19708 25978 19760 25984
rect 19616 25968 19668 25974
rect 19616 25910 19668 25916
rect 19628 25498 19656 25910
rect 19708 25696 19760 25702
rect 19708 25638 19760 25644
rect 19720 25498 19748 25638
rect 19812 25498 19840 26182
rect 19524 25492 19576 25498
rect 18984 25452 19288 25480
rect 18892 25350 19196 25378
rect 18880 25288 18932 25294
rect 18880 25230 18932 25236
rect 18892 24954 18920 25230
rect 18972 25220 19024 25226
rect 18972 25162 19024 25168
rect 18880 24948 18932 24954
rect 18880 24890 18932 24896
rect 18984 24818 19012 25162
rect 18880 24812 18932 24818
rect 18880 24754 18932 24760
rect 18972 24812 19024 24818
rect 18972 24754 19024 24760
rect 18892 24410 18920 24754
rect 19168 24698 19196 25350
rect 19260 24834 19288 25452
rect 19524 25434 19576 25440
rect 19616 25492 19668 25498
rect 19616 25434 19668 25440
rect 19708 25492 19760 25498
rect 19708 25434 19760 25440
rect 19800 25492 19852 25498
rect 19800 25434 19852 25440
rect 19904 25378 19932 26279
rect 19812 25350 19932 25378
rect 19708 25152 19760 25158
rect 19708 25094 19760 25100
rect 19524 24948 19576 24954
rect 19524 24890 19576 24896
rect 19260 24806 19380 24834
rect 19352 24750 19380 24806
rect 18984 24670 19196 24698
rect 19340 24744 19392 24750
rect 19340 24686 19392 24692
rect 18880 24404 18932 24410
rect 18880 24346 18932 24352
rect 18984 24274 19012 24670
rect 19143 24508 19451 24517
rect 19143 24506 19149 24508
rect 19205 24506 19229 24508
rect 19285 24506 19309 24508
rect 19365 24506 19389 24508
rect 19445 24506 19451 24508
rect 19205 24454 19207 24506
rect 19387 24454 19389 24506
rect 19143 24452 19149 24454
rect 19205 24452 19229 24454
rect 19285 24452 19309 24454
rect 19365 24452 19389 24454
rect 19445 24452 19451 24454
rect 19143 24443 19451 24452
rect 19536 24290 19564 24890
rect 18972 24268 19024 24274
rect 18972 24210 19024 24216
rect 19064 24268 19116 24274
rect 19064 24210 19116 24216
rect 19260 24262 19564 24290
rect 18880 24200 18932 24206
rect 18880 24142 18932 24148
rect 18708 22066 18828 22094
rect 18604 21004 18656 21010
rect 18604 20946 18656 20952
rect 18708 20777 18736 22066
rect 18788 21072 18840 21078
rect 18788 21014 18840 21020
rect 18694 20768 18750 20777
rect 18694 20703 18750 20712
rect 18420 19848 18472 19854
rect 18420 19790 18472 19796
rect 18326 19680 18382 19689
rect 18326 19615 18382 19624
rect 18340 16250 18368 19615
rect 18432 19446 18460 19790
rect 18420 19440 18472 19446
rect 18420 19382 18472 19388
rect 18694 19408 18750 19417
rect 18604 19372 18656 19378
rect 18694 19343 18750 19352
rect 18604 19314 18656 19320
rect 18512 16992 18564 16998
rect 18512 16934 18564 16940
rect 18328 16244 18380 16250
rect 18328 16186 18380 16192
rect 18328 16108 18380 16114
rect 18328 16050 18380 16056
rect 18340 15706 18368 16050
rect 18420 15904 18472 15910
rect 18420 15846 18472 15852
rect 18432 15706 18460 15846
rect 18328 15700 18380 15706
rect 18328 15642 18380 15648
rect 18420 15700 18472 15706
rect 18420 15642 18472 15648
rect 18420 15360 18472 15366
rect 18420 15302 18472 15308
rect 18326 13288 18382 13297
rect 18326 13223 18382 13232
rect 18340 12209 18368 13223
rect 18432 12832 18460 15302
rect 18524 13326 18552 16934
rect 18512 13320 18564 13326
rect 18512 13262 18564 13268
rect 18616 13258 18644 19314
rect 18708 16402 18736 19343
rect 18800 16561 18828 21014
rect 18892 20874 18920 24142
rect 18984 23526 19012 24210
rect 18972 23520 19024 23526
rect 18972 23462 19024 23468
rect 19076 23338 19104 24210
rect 19260 23730 19288 24262
rect 19720 24138 19748 25094
rect 19340 24132 19392 24138
rect 19340 24074 19392 24080
rect 19708 24132 19760 24138
rect 19708 24074 19760 24080
rect 19352 23769 19380 24074
rect 19338 23760 19394 23769
rect 19248 23724 19300 23730
rect 19338 23695 19340 23704
rect 19248 23666 19300 23672
rect 19392 23695 19394 23704
rect 19340 23666 19392 23672
rect 19524 23588 19576 23594
rect 19524 23530 19576 23536
rect 19536 23497 19564 23530
rect 19616 23520 19668 23526
rect 19522 23488 19578 23497
rect 19616 23462 19668 23468
rect 19143 23420 19451 23429
rect 19522 23423 19578 23432
rect 19143 23418 19149 23420
rect 19205 23418 19229 23420
rect 19285 23418 19309 23420
rect 19365 23418 19389 23420
rect 19445 23418 19451 23420
rect 19205 23366 19207 23418
rect 19387 23366 19389 23418
rect 19143 23364 19149 23366
rect 19205 23364 19229 23366
rect 19285 23364 19309 23366
rect 19365 23364 19389 23366
rect 19445 23364 19451 23366
rect 19143 23355 19451 23364
rect 19522 23352 19578 23361
rect 18984 23310 19104 23338
rect 18984 22438 19012 23310
rect 19518 23296 19522 23338
rect 19628 23322 19656 23462
rect 19518 23276 19524 23296
rect 19576 23287 19578 23296
rect 19616 23316 19668 23322
rect 19524 23258 19576 23264
rect 19616 23258 19668 23264
rect 19628 23202 19656 23258
rect 19594 23174 19656 23202
rect 19340 23112 19392 23118
rect 19321 23080 19340 23100
rect 19392 23080 19394 23089
rect 19321 23038 19338 23080
rect 19594 23066 19622 23174
rect 19338 23015 19394 23024
rect 19536 23038 19622 23066
rect 19064 22976 19116 22982
rect 19064 22918 19116 22924
rect 19156 22976 19208 22982
rect 19156 22918 19208 22924
rect 19294 22976 19346 22982
rect 19432 22976 19484 22982
rect 19346 22944 19394 22953
rect 19294 22918 19338 22924
rect 19076 22778 19104 22918
rect 19064 22772 19116 22778
rect 19064 22714 19116 22720
rect 19168 22642 19196 22918
rect 19306 22902 19338 22918
rect 19432 22918 19484 22924
rect 19338 22879 19394 22888
rect 19338 22808 19394 22817
rect 19444 22778 19472 22918
rect 19338 22743 19394 22752
rect 19432 22772 19484 22778
rect 19352 22710 19380 22743
rect 19432 22714 19484 22720
rect 19340 22704 19392 22710
rect 19536 22652 19564 23038
rect 19340 22646 19392 22652
rect 19493 22646 19564 22652
rect 19156 22636 19208 22642
rect 19545 22594 19564 22646
rect 19493 22588 19564 22594
rect 19156 22578 19208 22584
rect 18972 22432 19024 22438
rect 18972 22374 19024 22380
rect 18984 22030 19012 22374
rect 19143 22332 19451 22341
rect 19143 22330 19149 22332
rect 19205 22330 19229 22332
rect 19285 22330 19309 22332
rect 19365 22330 19389 22332
rect 19445 22330 19451 22332
rect 19205 22278 19207 22330
rect 19387 22278 19389 22330
rect 19143 22276 19149 22278
rect 19205 22276 19229 22278
rect 19285 22276 19309 22278
rect 19365 22276 19389 22278
rect 19445 22276 19451 22278
rect 19143 22267 19451 22276
rect 19432 22228 19484 22234
rect 19432 22170 19484 22176
rect 18972 22024 19024 22030
rect 18972 21966 19024 21972
rect 18880 20868 18932 20874
rect 18880 20810 18932 20816
rect 18984 19854 19012 21966
rect 19444 21554 19472 22170
rect 19432 21548 19484 21554
rect 19432 21490 19484 21496
rect 19536 21486 19564 22588
rect 19812 22137 19840 25350
rect 19892 25220 19944 25226
rect 19892 25162 19944 25168
rect 19904 24886 19932 25162
rect 19892 24880 19944 24886
rect 19892 24822 19944 24828
rect 19892 24132 19944 24138
rect 19892 24074 19944 24080
rect 19904 23730 19932 24074
rect 19892 23724 19944 23730
rect 19892 23666 19944 23672
rect 19890 23488 19946 23497
rect 19890 23423 19946 23432
rect 19904 23322 19932 23423
rect 19892 23316 19944 23322
rect 19892 23258 19944 23264
rect 19892 23112 19944 23118
rect 19892 23054 19944 23060
rect 19904 22953 19932 23054
rect 19890 22944 19946 22953
rect 19890 22879 19946 22888
rect 19798 22128 19854 22137
rect 19996 22094 20024 29106
rect 20088 29073 20116 31622
rect 20180 29170 20208 31726
rect 20272 30297 20300 33238
rect 20258 30288 20314 30297
rect 20258 30223 20314 30232
rect 20364 29866 20392 33374
rect 20444 33312 20496 33318
rect 20444 33254 20496 33260
rect 20456 31929 20484 33254
rect 20442 31920 20498 31929
rect 20442 31855 20498 31864
rect 20444 31816 20496 31822
rect 20444 31758 20496 31764
rect 20456 31482 20484 31758
rect 20444 31476 20496 31482
rect 20444 31418 20496 31424
rect 20548 30433 20576 33866
rect 20640 33046 20668 33934
rect 20720 33856 20772 33862
rect 20720 33798 20772 33804
rect 20812 33856 20864 33862
rect 20812 33798 20864 33804
rect 20628 33040 20680 33046
rect 20628 32982 20680 32988
rect 20640 32570 20668 32982
rect 20732 32892 20760 33798
rect 20824 33114 20852 33798
rect 20812 33108 20864 33114
rect 20812 33050 20864 33056
rect 20916 32910 20944 34546
rect 21008 33590 21036 35430
rect 21100 34490 21128 35550
rect 21192 35290 21220 36314
rect 21364 36168 21416 36174
rect 21364 36110 21416 36116
rect 21272 35828 21324 35834
rect 21272 35770 21324 35776
rect 21180 35284 21232 35290
rect 21180 35226 21232 35232
rect 21100 34462 21220 34490
rect 21088 34400 21140 34406
rect 21088 34342 21140 34348
rect 20996 33584 21048 33590
rect 20996 33526 21048 33532
rect 20812 32904 20864 32910
rect 20732 32864 20812 32892
rect 20812 32846 20864 32852
rect 20904 32904 20956 32910
rect 20904 32846 20956 32852
rect 20628 32564 20680 32570
rect 20628 32506 20680 32512
rect 20812 32564 20864 32570
rect 20812 32506 20864 32512
rect 20720 31884 20772 31890
rect 20720 31826 20772 31832
rect 20628 31340 20680 31346
rect 20628 31282 20680 31288
rect 20534 30424 20590 30433
rect 20444 30388 20496 30394
rect 20534 30359 20590 30368
rect 20444 30330 20496 30336
rect 20272 29838 20392 29866
rect 20168 29164 20220 29170
rect 20168 29106 20220 29112
rect 20074 29064 20130 29073
rect 20074 28999 20130 29008
rect 20168 28688 20220 28694
rect 20168 28630 20220 28636
rect 20180 28082 20208 28630
rect 20168 28076 20220 28082
rect 20168 28018 20220 28024
rect 20076 27056 20128 27062
rect 20076 26998 20128 27004
rect 20088 26586 20116 26998
rect 20076 26580 20128 26586
rect 20076 26522 20128 26528
rect 20076 25832 20128 25838
rect 20076 25774 20128 25780
rect 20088 25498 20116 25774
rect 20076 25492 20128 25498
rect 20076 25434 20128 25440
rect 20076 24880 20128 24886
rect 20076 24822 20128 24828
rect 19798 22063 19854 22072
rect 19904 22066 20024 22094
rect 20088 22094 20116 24822
rect 20180 24070 20208 28018
rect 20272 27538 20300 29838
rect 20456 29696 20484 30330
rect 20534 30288 20590 30297
rect 20534 30223 20590 30232
rect 20548 29730 20576 30223
rect 20640 29850 20668 31282
rect 20732 29850 20760 31826
rect 20824 30938 20852 32506
rect 20904 32224 20956 32230
rect 20904 32166 20956 32172
rect 20996 32224 21048 32230
rect 20996 32166 21048 32172
rect 20916 31958 20944 32166
rect 20904 31952 20956 31958
rect 20904 31894 20956 31900
rect 20812 30932 20864 30938
rect 20812 30874 20864 30880
rect 20904 30728 20956 30734
rect 20904 30670 20956 30676
rect 20812 30592 20864 30598
rect 20812 30534 20864 30540
rect 20628 29844 20680 29850
rect 20628 29786 20680 29792
rect 20720 29844 20772 29850
rect 20720 29786 20772 29792
rect 20548 29702 20760 29730
rect 20364 29668 20484 29696
rect 20260 27532 20312 27538
rect 20260 27474 20312 27480
rect 20260 27124 20312 27130
rect 20260 27066 20312 27072
rect 20272 26382 20300 27066
rect 20260 26376 20312 26382
rect 20260 26318 20312 26324
rect 20258 24304 20314 24313
rect 20258 24239 20314 24248
rect 20168 24064 20220 24070
rect 20168 24006 20220 24012
rect 20272 23882 20300 24239
rect 20180 23854 20300 23882
rect 20180 22642 20208 23854
rect 20364 23497 20392 29668
rect 20536 29640 20588 29646
rect 20536 29582 20588 29588
rect 20444 29572 20496 29578
rect 20444 29514 20496 29520
rect 20456 29306 20484 29514
rect 20548 29306 20576 29582
rect 20444 29300 20496 29306
rect 20444 29242 20496 29248
rect 20536 29300 20588 29306
rect 20536 29242 20588 29248
rect 20732 28778 20760 29702
rect 20824 29238 20852 30534
rect 20916 29782 20944 30670
rect 21008 30326 21036 32166
rect 21100 31822 21128 34342
rect 21192 34202 21220 34462
rect 21180 34196 21232 34202
rect 21180 34138 21232 34144
rect 21284 33998 21312 35770
rect 21376 34542 21404 36110
rect 21456 35488 21508 35494
rect 21454 35456 21456 35465
rect 21508 35456 21510 35465
rect 21454 35391 21510 35400
rect 21364 34536 21416 34542
rect 21364 34478 21416 34484
rect 21456 34400 21508 34406
rect 21454 34368 21456 34377
rect 21508 34368 21510 34377
rect 21454 34303 21510 34312
rect 21456 34060 21508 34066
rect 21456 34002 21508 34008
rect 21272 33992 21324 33998
rect 21272 33934 21324 33940
rect 21272 33856 21324 33862
rect 21272 33798 21324 33804
rect 21284 33402 21312 33798
rect 21284 33374 21404 33402
rect 21180 33312 21232 33318
rect 21272 33312 21324 33318
rect 21180 33254 21232 33260
rect 21270 33280 21272 33289
rect 21324 33280 21326 33289
rect 21192 33017 21220 33254
rect 21270 33215 21326 33224
rect 21178 33008 21234 33017
rect 21178 32943 21234 32952
rect 21180 32904 21232 32910
rect 21376 32858 21404 33374
rect 21180 32846 21232 32852
rect 21192 32570 21220 32846
rect 21284 32830 21404 32858
rect 21180 32564 21232 32570
rect 21180 32506 21232 32512
rect 21180 32428 21232 32434
rect 21180 32370 21232 32376
rect 21088 31816 21140 31822
rect 21088 31758 21140 31764
rect 21192 31482 21220 32370
rect 21180 31476 21232 31482
rect 21180 31418 21232 31424
rect 21284 31346 21312 32830
rect 21364 32768 21416 32774
rect 21364 32710 21416 32716
rect 21272 31340 21324 31346
rect 21272 31282 21324 31288
rect 21376 31226 21404 32710
rect 21468 32366 21496 34002
rect 21560 33697 21588 39902
rect 21546 33688 21602 33697
rect 21546 33623 21602 33632
rect 21652 33266 21680 41006
rect 22192 40928 22244 40934
rect 22190 40896 22192 40905
rect 22244 40896 22246 40905
rect 22190 40831 22246 40840
rect 22192 40384 22244 40390
rect 22190 40352 22192 40361
rect 22244 40352 22246 40361
rect 21742 40284 22050 40293
rect 22190 40287 22246 40296
rect 21742 40282 21748 40284
rect 21804 40282 21828 40284
rect 21884 40282 21908 40284
rect 21964 40282 21988 40284
rect 22044 40282 22050 40284
rect 21804 40230 21806 40282
rect 21986 40230 21988 40282
rect 21742 40228 21748 40230
rect 21804 40228 21828 40230
rect 21884 40228 21908 40230
rect 21964 40228 21988 40230
rect 22044 40228 22050 40230
rect 21742 40219 22050 40228
rect 22468 39908 22520 39914
rect 22468 39850 22520 39856
rect 22192 39296 22244 39302
rect 22190 39264 22192 39273
rect 22244 39264 22246 39273
rect 21742 39196 22050 39205
rect 22190 39199 22246 39208
rect 21742 39194 21748 39196
rect 21804 39194 21828 39196
rect 21884 39194 21908 39196
rect 21964 39194 21988 39196
rect 22044 39194 22050 39196
rect 21804 39142 21806 39194
rect 21986 39142 21988 39194
rect 21742 39140 21748 39142
rect 21804 39140 21828 39142
rect 21884 39140 21908 39142
rect 21964 39140 21988 39142
rect 22044 39140 22050 39142
rect 21742 39131 22050 39140
rect 22192 38208 22244 38214
rect 22190 38176 22192 38185
rect 22244 38176 22246 38185
rect 21742 38108 22050 38117
rect 22190 38111 22246 38120
rect 21742 38106 21748 38108
rect 21804 38106 21828 38108
rect 21884 38106 21908 38108
rect 21964 38106 21988 38108
rect 22044 38106 22050 38108
rect 21804 38054 21806 38106
rect 21986 38054 21988 38106
rect 21742 38052 21748 38054
rect 21804 38052 21828 38054
rect 21884 38052 21908 38054
rect 21964 38052 21988 38054
rect 22044 38052 22050 38054
rect 21742 38043 22050 38052
rect 22284 37188 22336 37194
rect 22284 37130 22336 37136
rect 22296 37097 22324 37130
rect 22282 37088 22338 37097
rect 21742 37020 22050 37029
rect 22282 37023 22338 37032
rect 21742 37018 21748 37020
rect 21804 37018 21828 37020
rect 21884 37018 21908 37020
rect 21964 37018 21988 37020
rect 22044 37018 22050 37020
rect 21804 36966 21806 37018
rect 21986 36966 21988 37018
rect 21742 36964 21748 36966
rect 21804 36964 21828 36966
rect 21884 36964 21908 36966
rect 21964 36964 21988 36966
rect 22044 36964 22050 36966
rect 21742 36955 22050 36964
rect 22284 36100 22336 36106
rect 22284 36042 22336 36048
rect 22296 36009 22324 36042
rect 22282 36000 22338 36009
rect 21742 35932 22050 35941
rect 22282 35935 22338 35944
rect 21742 35930 21748 35932
rect 21804 35930 21828 35932
rect 21884 35930 21908 35932
rect 21964 35930 21988 35932
rect 22044 35930 22050 35932
rect 21804 35878 21806 35930
rect 21986 35878 21988 35930
rect 21742 35876 21748 35878
rect 21804 35876 21828 35878
rect 21884 35876 21908 35878
rect 21964 35876 21988 35878
rect 22044 35876 22050 35878
rect 21742 35867 22050 35876
rect 22020 35018 22140 35034
rect 22008 35012 22140 35018
rect 22060 35006 22140 35012
rect 22008 34954 22060 34960
rect 21742 34844 22050 34853
rect 21742 34842 21748 34844
rect 21804 34842 21828 34844
rect 21884 34842 21908 34844
rect 21964 34842 21988 34844
rect 22044 34842 22050 34844
rect 21804 34790 21806 34842
rect 21986 34790 21988 34842
rect 21742 34788 21748 34790
rect 21804 34788 21828 34790
rect 21884 34788 21908 34790
rect 21964 34788 21988 34790
rect 22044 34788 22050 34790
rect 21742 34779 22050 34788
rect 21742 33756 22050 33765
rect 21742 33754 21748 33756
rect 21804 33754 21828 33756
rect 21884 33754 21908 33756
rect 21964 33754 21988 33756
rect 22044 33754 22050 33756
rect 21804 33702 21806 33754
rect 21986 33702 21988 33754
rect 21742 33700 21748 33702
rect 21804 33700 21828 33702
rect 21884 33700 21908 33702
rect 21964 33700 21988 33702
rect 22044 33700 22050 33702
rect 21742 33691 22050 33700
rect 22112 33402 22140 35006
rect 22192 34944 22244 34950
rect 22190 34912 22192 34921
rect 22244 34912 22246 34921
rect 22190 34847 22246 34856
rect 22284 34604 22336 34610
rect 22284 34546 22336 34552
rect 22192 33856 22244 33862
rect 22190 33824 22192 33833
rect 22244 33824 22246 33833
rect 22190 33759 22246 33768
rect 22112 33374 22232 33402
rect 21652 33238 22140 33266
rect 21640 33040 21692 33046
rect 21640 32982 21692 32988
rect 21548 32904 21600 32910
rect 21548 32846 21600 32852
rect 21456 32360 21508 32366
rect 21456 32302 21508 32308
rect 21456 32224 21508 32230
rect 21454 32192 21456 32201
rect 21508 32192 21510 32201
rect 21454 32127 21510 32136
rect 21560 32026 21588 32846
rect 21548 32020 21600 32026
rect 21548 31962 21600 31968
rect 21546 31920 21602 31929
rect 21546 31855 21602 31864
rect 21192 31198 21404 31226
rect 21088 31136 21140 31142
rect 21088 31078 21140 31084
rect 20996 30320 21048 30326
rect 20996 30262 21048 30268
rect 20996 30048 21048 30054
rect 20996 29990 21048 29996
rect 20904 29776 20956 29782
rect 20904 29718 20956 29724
rect 21008 29646 21036 29990
rect 21100 29646 21128 31078
rect 21192 30734 21220 31198
rect 21456 31136 21508 31142
rect 21454 31104 21456 31113
rect 21508 31104 21510 31113
rect 21454 31039 21510 31048
rect 21270 30968 21326 30977
rect 21270 30903 21326 30912
rect 21180 30728 21232 30734
rect 21180 30670 21232 30676
rect 20996 29640 21048 29646
rect 20996 29582 21048 29588
rect 21088 29640 21140 29646
rect 21088 29582 21140 29588
rect 20996 29504 21048 29510
rect 20996 29446 21048 29452
rect 21180 29504 21232 29510
rect 21180 29446 21232 29452
rect 20812 29232 20864 29238
rect 20812 29174 20864 29180
rect 20456 28750 20760 28778
rect 20456 26874 20484 28750
rect 20536 28620 20588 28626
rect 20536 28562 20588 28568
rect 20548 28218 20576 28562
rect 21008 28558 21036 29446
rect 20628 28552 20680 28558
rect 20628 28494 20680 28500
rect 20996 28552 21048 28558
rect 20996 28494 21048 28500
rect 20640 28218 20668 28494
rect 20720 28416 20772 28422
rect 20720 28358 20772 28364
rect 20996 28416 21048 28422
rect 20996 28358 21048 28364
rect 20732 28218 20760 28358
rect 20536 28212 20588 28218
rect 20536 28154 20588 28160
rect 20628 28212 20680 28218
rect 20628 28154 20680 28160
rect 20720 28212 20772 28218
rect 20720 28154 20772 28160
rect 20812 28076 20864 28082
rect 20812 28018 20864 28024
rect 20824 27674 20852 28018
rect 20904 27872 20956 27878
rect 20904 27814 20956 27820
rect 20720 27668 20772 27674
rect 20720 27610 20772 27616
rect 20812 27668 20864 27674
rect 20812 27610 20864 27616
rect 20732 27418 20760 27610
rect 20732 27390 20852 27418
rect 20720 27328 20772 27334
rect 20720 27270 20772 27276
rect 20456 26846 20576 26874
rect 20444 26784 20496 26790
rect 20444 26726 20496 26732
rect 20456 26586 20484 26726
rect 20444 26580 20496 26586
rect 20444 26522 20496 26528
rect 20548 25362 20576 26846
rect 20628 26852 20680 26858
rect 20628 26794 20680 26800
rect 20640 26586 20668 26794
rect 20732 26586 20760 27270
rect 20628 26580 20680 26586
rect 20628 26522 20680 26528
rect 20720 26580 20772 26586
rect 20720 26522 20772 26528
rect 20720 25696 20772 25702
rect 20720 25638 20772 25644
rect 20732 25498 20760 25638
rect 20720 25492 20772 25498
rect 20720 25434 20772 25440
rect 20536 25356 20588 25362
rect 20536 25298 20588 25304
rect 20444 25288 20496 25294
rect 20444 25230 20496 25236
rect 20456 24290 20484 25230
rect 20536 25220 20588 25226
rect 20536 25162 20588 25168
rect 20548 24410 20576 25162
rect 20628 25152 20680 25158
rect 20628 25094 20680 25100
rect 20720 25152 20772 25158
rect 20720 25094 20772 25100
rect 20640 24410 20668 25094
rect 20732 24954 20760 25094
rect 20720 24948 20772 24954
rect 20720 24890 20772 24896
rect 20536 24404 20588 24410
rect 20536 24346 20588 24352
rect 20628 24404 20680 24410
rect 20628 24346 20680 24352
rect 20456 24262 20668 24290
rect 20640 24206 20668 24262
rect 20628 24200 20680 24206
rect 20628 24142 20680 24148
rect 20640 23866 20668 24142
rect 20628 23860 20680 23866
rect 20628 23802 20680 23808
rect 20536 23724 20588 23730
rect 20536 23666 20588 23672
rect 20350 23488 20406 23497
rect 20350 23423 20406 23432
rect 20548 23322 20576 23666
rect 20720 23520 20772 23526
rect 20720 23462 20772 23468
rect 20626 23352 20682 23361
rect 20536 23316 20588 23322
rect 20626 23287 20682 23296
rect 20536 23258 20588 23264
rect 20444 23248 20496 23254
rect 20444 23190 20496 23196
rect 20350 23080 20406 23089
rect 20350 23015 20406 23024
rect 20364 22778 20392 23015
rect 20352 22772 20404 22778
rect 20352 22714 20404 22720
rect 20258 22672 20314 22681
rect 20168 22636 20220 22642
rect 20258 22607 20314 22616
rect 20168 22578 20220 22584
rect 20088 22066 20208 22094
rect 19524 21480 19576 21486
rect 19524 21422 19576 21428
rect 19064 21344 19116 21350
rect 19064 21286 19116 21292
rect 19076 19854 19104 21286
rect 19143 21244 19451 21253
rect 19143 21242 19149 21244
rect 19205 21242 19229 21244
rect 19285 21242 19309 21244
rect 19365 21242 19389 21244
rect 19445 21242 19451 21244
rect 19205 21190 19207 21242
rect 19387 21190 19389 21242
rect 19143 21188 19149 21190
rect 19205 21188 19229 21190
rect 19285 21188 19309 21190
rect 19365 21188 19389 21190
rect 19445 21188 19451 21190
rect 19143 21179 19451 21188
rect 19536 20398 19564 21422
rect 19524 20392 19576 20398
rect 19524 20334 19576 20340
rect 19143 20156 19451 20165
rect 19143 20154 19149 20156
rect 19205 20154 19229 20156
rect 19285 20154 19309 20156
rect 19365 20154 19389 20156
rect 19445 20154 19451 20156
rect 19205 20102 19207 20154
rect 19387 20102 19389 20154
rect 19143 20100 19149 20102
rect 19205 20100 19229 20102
rect 19285 20100 19309 20102
rect 19365 20100 19389 20102
rect 19445 20100 19451 20102
rect 19143 20091 19451 20100
rect 18972 19848 19024 19854
rect 18972 19790 19024 19796
rect 19064 19848 19116 19854
rect 19064 19790 19116 19796
rect 18880 19712 18932 19718
rect 18880 19654 18932 19660
rect 18892 19378 18920 19654
rect 18880 19372 18932 19378
rect 18880 19314 18932 19320
rect 18984 19310 19012 19790
rect 18972 19304 19024 19310
rect 18972 19246 19024 19252
rect 18984 18086 19012 19246
rect 19143 19068 19451 19077
rect 19143 19066 19149 19068
rect 19205 19066 19229 19068
rect 19285 19066 19309 19068
rect 19365 19066 19389 19068
rect 19445 19066 19451 19068
rect 19205 19014 19207 19066
rect 19387 19014 19389 19066
rect 19143 19012 19149 19014
rect 19205 19012 19229 19014
rect 19285 19012 19309 19014
rect 19365 19012 19389 19014
rect 19445 19012 19451 19014
rect 19143 19003 19451 19012
rect 19536 18970 19564 20334
rect 19616 19780 19668 19786
rect 19616 19722 19668 19728
rect 19524 18964 19576 18970
rect 19524 18906 19576 18912
rect 19628 18766 19656 19722
rect 19708 18964 19760 18970
rect 19708 18906 19760 18912
rect 19616 18760 19668 18766
rect 19616 18702 19668 18708
rect 19524 18624 19576 18630
rect 19720 18578 19748 18906
rect 19524 18566 19576 18572
rect 19064 18352 19116 18358
rect 19064 18294 19116 18300
rect 18972 18080 19024 18086
rect 18972 18022 19024 18028
rect 18984 17134 19012 18022
rect 19076 17678 19104 18294
rect 19143 17980 19451 17989
rect 19143 17978 19149 17980
rect 19205 17978 19229 17980
rect 19285 17978 19309 17980
rect 19365 17978 19389 17980
rect 19445 17978 19451 17980
rect 19205 17926 19207 17978
rect 19387 17926 19389 17978
rect 19143 17924 19149 17926
rect 19205 17924 19229 17926
rect 19285 17924 19309 17926
rect 19365 17924 19389 17926
rect 19445 17924 19451 17926
rect 19143 17915 19451 17924
rect 19536 17678 19564 18566
rect 19628 18550 19748 18578
rect 19064 17672 19116 17678
rect 19064 17614 19116 17620
rect 19524 17672 19576 17678
rect 19524 17614 19576 17620
rect 19536 17202 19564 17614
rect 19524 17196 19576 17202
rect 19524 17138 19576 17144
rect 18972 17128 19024 17134
rect 18972 17070 19024 17076
rect 18786 16552 18842 16561
rect 18786 16487 18842 16496
rect 18708 16374 18828 16402
rect 18696 16108 18748 16114
rect 18696 16050 18748 16056
rect 18708 15638 18736 16050
rect 18696 15632 18748 15638
rect 18696 15574 18748 15580
rect 18694 15464 18750 15473
rect 18694 15399 18750 15408
rect 18604 13252 18656 13258
rect 18604 13194 18656 13200
rect 18616 12986 18644 13194
rect 18604 12980 18656 12986
rect 18604 12922 18656 12928
rect 18512 12844 18564 12850
rect 18432 12804 18512 12832
rect 18512 12786 18564 12792
rect 18604 12368 18656 12374
rect 18604 12310 18656 12316
rect 18708 12322 18736 15399
rect 18800 12442 18828 16374
rect 18880 16040 18932 16046
rect 18880 15982 18932 15988
rect 18892 15570 18920 15982
rect 18880 15564 18932 15570
rect 18880 15506 18932 15512
rect 18892 15162 18920 15506
rect 18984 15434 19012 17070
rect 19524 16992 19576 16998
rect 19524 16934 19576 16940
rect 19143 16892 19451 16901
rect 19143 16890 19149 16892
rect 19205 16890 19229 16892
rect 19285 16890 19309 16892
rect 19365 16890 19389 16892
rect 19445 16890 19451 16892
rect 19205 16838 19207 16890
rect 19387 16838 19389 16890
rect 19143 16836 19149 16838
rect 19205 16836 19229 16838
rect 19285 16836 19309 16838
rect 19365 16836 19389 16838
rect 19445 16836 19451 16838
rect 19143 16827 19451 16836
rect 19246 16008 19302 16017
rect 19246 15943 19248 15952
rect 19300 15943 19302 15952
rect 19248 15914 19300 15920
rect 19064 15904 19116 15910
rect 19064 15846 19116 15852
rect 19076 15706 19104 15846
rect 19143 15804 19451 15813
rect 19143 15802 19149 15804
rect 19205 15802 19229 15804
rect 19285 15802 19309 15804
rect 19365 15802 19389 15804
rect 19445 15802 19451 15804
rect 19205 15750 19207 15802
rect 19387 15750 19389 15802
rect 19143 15748 19149 15750
rect 19205 15748 19229 15750
rect 19285 15748 19309 15750
rect 19365 15748 19389 15750
rect 19445 15748 19451 15750
rect 19143 15739 19451 15748
rect 19536 15706 19564 16934
rect 19628 16454 19656 18550
rect 19706 17776 19762 17785
rect 19706 17711 19762 17720
rect 19616 16448 19668 16454
rect 19616 16390 19668 16396
rect 19628 16046 19656 16390
rect 19616 16040 19668 16046
rect 19616 15982 19668 15988
rect 19064 15700 19116 15706
rect 19064 15642 19116 15648
rect 19524 15700 19576 15706
rect 19524 15642 19576 15648
rect 19156 15496 19208 15502
rect 19156 15438 19208 15444
rect 18972 15428 19024 15434
rect 18972 15370 19024 15376
rect 19168 15178 19196 15438
rect 18880 15156 18932 15162
rect 18880 15098 18932 15104
rect 19076 15150 19564 15178
rect 18972 13932 19024 13938
rect 18972 13874 19024 13880
rect 18880 13728 18932 13734
rect 18880 13670 18932 13676
rect 18788 12436 18840 12442
rect 18788 12378 18840 12384
rect 18420 12232 18472 12238
rect 18326 12200 18382 12209
rect 18420 12174 18472 12180
rect 18326 12135 18382 12144
rect 18328 12096 18380 12102
rect 18328 12038 18380 12044
rect 18340 11150 18368 12038
rect 18432 11354 18460 12174
rect 18512 12096 18564 12102
rect 18512 12038 18564 12044
rect 18524 11898 18552 12038
rect 18512 11892 18564 11898
rect 18512 11834 18564 11840
rect 18616 11778 18644 12310
rect 18708 12294 18828 12322
rect 18696 12096 18748 12102
rect 18696 12038 18748 12044
rect 18524 11750 18644 11778
rect 18708 11762 18736 12038
rect 18800 11801 18828 12294
rect 18786 11792 18842 11801
rect 18696 11756 18748 11762
rect 18524 11694 18552 11750
rect 18786 11727 18842 11736
rect 18696 11698 18748 11704
rect 18512 11688 18564 11694
rect 18512 11630 18564 11636
rect 18420 11348 18472 11354
rect 18420 11290 18472 11296
rect 18328 11144 18380 11150
rect 18328 11086 18380 11092
rect 18420 10600 18472 10606
rect 18420 10542 18472 10548
rect 18328 10464 18380 10470
rect 18328 10406 18380 10412
rect 18340 10062 18368 10406
rect 18432 10198 18460 10542
rect 18420 10192 18472 10198
rect 18420 10134 18472 10140
rect 18328 10056 18380 10062
rect 18328 9998 18380 10004
rect 18418 10024 18474 10033
rect 18418 9959 18474 9968
rect 18328 8424 18380 8430
rect 18328 8366 18380 8372
rect 18236 7540 18288 7546
rect 18236 7482 18288 7488
rect 18340 7274 18368 8366
rect 18432 8242 18460 9959
rect 18524 8430 18552 11630
rect 18604 10260 18656 10266
rect 18604 10202 18656 10208
rect 18616 9722 18644 10202
rect 18604 9716 18656 9722
rect 18604 9658 18656 9664
rect 18604 9580 18656 9586
rect 18604 9522 18656 9528
rect 18616 9081 18644 9522
rect 18602 9072 18658 9081
rect 18602 9007 18658 9016
rect 18604 8832 18656 8838
rect 18604 8774 18656 8780
rect 18512 8424 18564 8430
rect 18512 8366 18564 8372
rect 18432 8214 18552 8242
rect 18524 8090 18552 8214
rect 18512 8084 18564 8090
rect 18512 8026 18564 8032
rect 18512 7880 18564 7886
rect 18418 7848 18474 7857
rect 18512 7822 18564 7828
rect 18418 7783 18474 7792
rect 18328 7268 18380 7274
rect 18328 7210 18380 7216
rect 18236 6792 18288 6798
rect 18236 6734 18288 6740
rect 18248 6497 18276 6734
rect 18234 6488 18290 6497
rect 18234 6423 18290 6432
rect 18234 6352 18290 6361
rect 18234 6287 18236 6296
rect 18288 6287 18290 6296
rect 18236 6258 18288 6264
rect 18340 5930 18368 7210
rect 18432 6322 18460 7783
rect 18524 7002 18552 7822
rect 18616 7546 18644 8774
rect 18604 7540 18656 7546
rect 18604 7482 18656 7488
rect 18512 6996 18564 7002
rect 18512 6938 18564 6944
rect 18708 6662 18736 11698
rect 18788 11552 18840 11558
rect 18788 11494 18840 11500
rect 18800 11150 18828 11494
rect 18788 11144 18840 11150
rect 18788 11086 18840 11092
rect 18788 10056 18840 10062
rect 18788 9998 18840 10004
rect 18800 9382 18828 9998
rect 18892 9761 18920 13670
rect 18984 13530 19012 13874
rect 18972 13524 19024 13530
rect 18972 13466 19024 13472
rect 19076 13462 19104 15150
rect 19143 14716 19451 14725
rect 19143 14714 19149 14716
rect 19205 14714 19229 14716
rect 19285 14714 19309 14716
rect 19365 14714 19389 14716
rect 19445 14714 19451 14716
rect 19205 14662 19207 14714
rect 19387 14662 19389 14714
rect 19143 14660 19149 14662
rect 19205 14660 19229 14662
rect 19285 14660 19309 14662
rect 19365 14660 19389 14662
rect 19445 14660 19451 14662
rect 19143 14651 19451 14660
rect 19536 13938 19564 15150
rect 19628 14618 19656 15982
rect 19616 14612 19668 14618
rect 19616 14554 19668 14560
rect 19524 13932 19576 13938
rect 19524 13874 19576 13880
rect 19143 13628 19451 13637
rect 19143 13626 19149 13628
rect 19205 13626 19229 13628
rect 19285 13626 19309 13628
rect 19365 13626 19389 13628
rect 19445 13626 19451 13628
rect 19205 13574 19207 13626
rect 19387 13574 19389 13626
rect 19143 13572 19149 13574
rect 19205 13572 19229 13574
rect 19285 13572 19309 13574
rect 19365 13572 19389 13574
rect 19445 13572 19451 13574
rect 19143 13563 19451 13572
rect 19064 13456 19116 13462
rect 19064 13398 19116 13404
rect 19616 13320 19668 13326
rect 19616 13262 19668 13268
rect 19064 13184 19116 13190
rect 19064 13126 19116 13132
rect 19076 12986 19104 13126
rect 19064 12980 19116 12986
rect 19064 12922 19116 12928
rect 19524 12844 19576 12850
rect 19524 12786 19576 12792
rect 19064 12640 19116 12646
rect 19064 12582 19116 12588
rect 19076 12434 19104 12582
rect 19143 12540 19451 12549
rect 19143 12538 19149 12540
rect 19205 12538 19229 12540
rect 19285 12538 19309 12540
rect 19365 12538 19389 12540
rect 19445 12538 19451 12540
rect 19205 12486 19207 12538
rect 19387 12486 19389 12538
rect 19143 12484 19149 12486
rect 19205 12484 19229 12486
rect 19285 12484 19309 12486
rect 19365 12484 19389 12486
rect 19445 12484 19451 12486
rect 19143 12475 19451 12484
rect 19076 12406 19196 12434
rect 18972 12368 19024 12374
rect 18972 12310 19024 12316
rect 19062 12336 19118 12345
rect 18878 9752 18934 9761
rect 18878 9687 18934 9696
rect 18788 9376 18840 9382
rect 18788 9318 18840 9324
rect 18984 9058 19012 12310
rect 19062 12271 19118 12280
rect 19076 12238 19104 12271
rect 19064 12232 19116 12238
rect 19064 12174 19116 12180
rect 19076 11898 19104 12174
rect 19064 11892 19116 11898
rect 19064 11834 19116 11840
rect 19168 11642 19196 12406
rect 19432 12232 19484 12238
rect 19536 12220 19564 12786
rect 19628 12646 19656 13262
rect 19616 12640 19668 12646
rect 19616 12582 19668 12588
rect 19720 12434 19748 17711
rect 19798 16552 19854 16561
rect 19798 16487 19854 16496
rect 19812 15502 19840 16487
rect 19800 15496 19852 15502
rect 19800 15438 19852 15444
rect 19812 15162 19840 15438
rect 19800 15156 19852 15162
rect 19800 15098 19852 15104
rect 19800 14000 19852 14006
rect 19800 13942 19852 13948
rect 19812 12850 19840 13942
rect 19800 12844 19852 12850
rect 19800 12786 19852 12792
rect 19904 12782 19932 22066
rect 20076 21956 20128 21962
rect 20076 21898 20128 21904
rect 20088 21622 20116 21898
rect 20076 21616 20128 21622
rect 20076 21558 20128 21564
rect 20076 21344 20128 21350
rect 20076 21286 20128 21292
rect 19984 20256 20036 20262
rect 19984 20198 20036 20204
rect 19996 20058 20024 20198
rect 19984 20052 20036 20058
rect 19984 19994 20036 20000
rect 20088 19689 20116 21286
rect 20180 20466 20208 22066
rect 20168 20460 20220 20466
rect 20168 20402 20220 20408
rect 20272 19802 20300 22607
rect 20352 22228 20404 22234
rect 20352 22170 20404 22176
rect 20364 21350 20392 22170
rect 20352 21344 20404 21350
rect 20352 21286 20404 21292
rect 20352 21004 20404 21010
rect 20352 20946 20404 20952
rect 20364 19922 20392 20946
rect 20352 19916 20404 19922
rect 20352 19858 20404 19864
rect 20168 19780 20220 19786
rect 20272 19774 20392 19802
rect 20456 19786 20484 23190
rect 20640 21622 20668 23287
rect 20628 21616 20680 21622
rect 20628 21558 20680 21564
rect 20536 21344 20588 21350
rect 20536 21286 20588 21292
rect 20548 21146 20576 21286
rect 20536 21140 20588 21146
rect 20536 21082 20588 21088
rect 20628 20868 20680 20874
rect 20628 20810 20680 20816
rect 20640 20754 20668 20810
rect 20732 20754 20760 23462
rect 20824 22642 20852 27390
rect 20916 26382 20944 27814
rect 21008 27470 21036 28358
rect 21088 27872 21140 27878
rect 21086 27840 21088 27849
rect 21140 27840 21142 27849
rect 21086 27775 21142 27784
rect 20996 27464 21048 27470
rect 20996 27406 21048 27412
rect 20996 27328 21048 27334
rect 20996 27270 21048 27276
rect 20904 26376 20956 26382
rect 20904 26318 20956 26324
rect 20904 25900 20956 25906
rect 20904 25842 20956 25848
rect 20916 24954 20944 25842
rect 20904 24948 20956 24954
rect 20904 24890 20956 24896
rect 21008 24290 21036 27270
rect 21088 25696 21140 25702
rect 21088 25638 21140 25644
rect 21100 24410 21128 25638
rect 21088 24404 21140 24410
rect 21088 24346 21140 24352
rect 20916 24262 21036 24290
rect 20916 24206 20944 24262
rect 20904 24200 20956 24206
rect 20904 24142 20956 24148
rect 21088 24132 21140 24138
rect 21088 24074 21140 24080
rect 20996 24064 21048 24070
rect 20996 24006 21048 24012
rect 21008 23118 21036 24006
rect 20996 23112 21048 23118
rect 20996 23054 21048 23060
rect 20812 22636 20864 22642
rect 20812 22578 20864 22584
rect 20996 21888 21048 21894
rect 20996 21830 21048 21836
rect 20904 21548 20956 21554
rect 20904 21490 20956 21496
rect 20810 21312 20866 21321
rect 20810 21247 20866 21256
rect 20824 21146 20852 21247
rect 20812 21140 20864 21146
rect 20812 21082 20864 21088
rect 20640 20726 20760 20754
rect 20812 20596 20864 20602
rect 20812 20538 20864 20544
rect 20536 20256 20588 20262
rect 20536 20198 20588 20204
rect 20168 19722 20220 19728
rect 20074 19680 20130 19689
rect 20074 19615 20130 19624
rect 19982 19272 20038 19281
rect 19982 19207 20038 19216
rect 19996 16522 20024 19207
rect 20076 18420 20128 18426
rect 20076 18362 20128 18368
rect 19984 16516 20036 16522
rect 19984 16458 20036 16464
rect 20088 14006 20116 18362
rect 20180 16998 20208 19722
rect 20364 19334 20392 19774
rect 20444 19780 20496 19786
rect 20444 19722 20496 19728
rect 20272 19306 20392 19334
rect 20168 16992 20220 16998
rect 20168 16934 20220 16940
rect 20168 16584 20220 16590
rect 20168 16526 20220 16532
rect 20076 14000 20128 14006
rect 20076 13942 20128 13948
rect 19984 13320 20036 13326
rect 19984 13262 20036 13268
rect 19996 13161 20024 13262
rect 19982 13152 20038 13161
rect 19982 13087 20038 13096
rect 19892 12776 19944 12782
rect 19892 12718 19944 12724
rect 19984 12776 20036 12782
rect 19984 12718 20036 12724
rect 19800 12640 19852 12646
rect 19800 12582 19852 12588
rect 19484 12192 19564 12220
rect 19628 12406 19748 12434
rect 19432 12174 19484 12180
rect 19524 11892 19576 11898
rect 19524 11834 19576 11840
rect 19076 11614 19196 11642
rect 19076 10180 19104 11614
rect 19143 11452 19451 11461
rect 19143 11450 19149 11452
rect 19205 11450 19229 11452
rect 19285 11450 19309 11452
rect 19365 11450 19389 11452
rect 19445 11450 19451 11452
rect 19205 11398 19207 11450
rect 19387 11398 19389 11450
rect 19143 11396 19149 11398
rect 19205 11396 19229 11398
rect 19285 11396 19309 11398
rect 19365 11396 19389 11398
rect 19445 11396 19451 11398
rect 19143 11387 19451 11396
rect 19340 11280 19392 11286
rect 19340 11222 19392 11228
rect 19352 10810 19380 11222
rect 19340 10804 19392 10810
rect 19340 10746 19392 10752
rect 19432 10668 19484 10674
rect 19432 10610 19484 10616
rect 19444 10452 19472 10610
rect 19536 10606 19564 11834
rect 19628 10713 19656 12406
rect 19812 11898 19840 12582
rect 19996 12442 20024 12718
rect 20076 12640 20128 12646
rect 20076 12582 20128 12588
rect 20088 12442 20116 12582
rect 19984 12436 20036 12442
rect 19984 12378 20036 12384
rect 20076 12436 20128 12442
rect 20076 12378 20128 12384
rect 19892 12232 19944 12238
rect 19892 12174 19944 12180
rect 19984 12232 20036 12238
rect 20180 12220 20208 16526
rect 19984 12174 20036 12180
rect 20088 12192 20208 12220
rect 19800 11892 19852 11898
rect 19800 11834 19852 11840
rect 19800 11756 19852 11762
rect 19800 11698 19852 11704
rect 19812 11354 19840 11698
rect 19800 11348 19852 11354
rect 19800 11290 19852 11296
rect 19708 11280 19760 11286
rect 19708 11222 19760 11228
rect 19720 11150 19748 11222
rect 19708 11144 19760 11150
rect 19708 11086 19760 11092
rect 19708 11008 19760 11014
rect 19708 10950 19760 10956
rect 19614 10704 19670 10713
rect 19614 10639 19670 10648
rect 19524 10600 19576 10606
rect 19576 10560 19656 10588
rect 19524 10542 19576 10548
rect 19444 10424 19564 10452
rect 19143 10364 19451 10373
rect 19143 10362 19149 10364
rect 19205 10362 19229 10364
rect 19285 10362 19309 10364
rect 19365 10362 19389 10364
rect 19445 10362 19451 10364
rect 19205 10310 19207 10362
rect 19387 10310 19389 10362
rect 19143 10308 19149 10310
rect 19205 10308 19229 10310
rect 19285 10308 19309 10310
rect 19365 10308 19389 10310
rect 19445 10308 19451 10310
rect 19143 10299 19451 10308
rect 19076 10152 19196 10180
rect 19064 10056 19116 10062
rect 19064 9998 19116 10004
rect 19076 9081 19104 9998
rect 19168 9586 19196 10152
rect 19248 10056 19300 10062
rect 19248 9998 19300 10004
rect 19260 9625 19288 9998
rect 19536 9722 19564 10424
rect 19524 9716 19576 9722
rect 19524 9658 19576 9664
rect 19628 9654 19656 10560
rect 19616 9648 19668 9654
rect 19246 9616 19302 9625
rect 19156 9580 19208 9586
rect 19616 9590 19668 9596
rect 19246 9551 19302 9560
rect 19156 9522 19208 9528
rect 19143 9276 19451 9285
rect 19143 9274 19149 9276
rect 19205 9274 19229 9276
rect 19285 9274 19309 9276
rect 19365 9274 19389 9276
rect 19445 9274 19451 9276
rect 19205 9222 19207 9274
rect 19387 9222 19389 9274
rect 19143 9220 19149 9222
rect 19205 9220 19229 9222
rect 19285 9220 19309 9222
rect 19365 9220 19389 9222
rect 19445 9220 19451 9222
rect 19143 9211 19451 9220
rect 19340 9172 19392 9178
rect 19720 9160 19748 10950
rect 19904 10810 19932 12174
rect 19996 11694 20024 12174
rect 20088 12084 20116 12192
rect 20088 12056 20208 12084
rect 19984 11688 20036 11694
rect 19984 11630 20036 11636
rect 20074 11656 20130 11665
rect 20074 11591 20130 11600
rect 19800 10804 19852 10810
rect 19800 10746 19852 10752
rect 19892 10804 19944 10810
rect 19892 10746 19944 10752
rect 19812 9994 19840 10746
rect 19800 9988 19852 9994
rect 19800 9930 19852 9936
rect 19812 9586 19840 9930
rect 19984 9648 20036 9654
rect 19984 9590 20036 9596
rect 19800 9580 19852 9586
rect 19800 9522 19852 9528
rect 19892 9580 19944 9586
rect 19892 9522 19944 9528
rect 19340 9114 19392 9120
rect 19628 9132 19748 9160
rect 18892 9030 19012 9058
rect 19062 9072 19118 9081
rect 18892 8242 18920 9030
rect 19062 9007 19118 9016
rect 18972 8968 19024 8974
rect 19352 8945 19380 9114
rect 19628 9024 19656 9132
rect 19628 8996 19748 9024
rect 19432 8968 19484 8974
rect 18972 8910 19024 8916
rect 19338 8936 19394 8945
rect 18984 8634 19012 8910
rect 19432 8910 19484 8916
rect 19524 8968 19576 8974
rect 19524 8910 19576 8916
rect 19338 8871 19394 8880
rect 19444 8838 19472 8910
rect 19432 8832 19484 8838
rect 19432 8774 19484 8780
rect 18972 8628 19024 8634
rect 18972 8570 19024 8576
rect 18970 8256 19026 8265
rect 18892 8214 18970 8242
rect 18970 8191 19026 8200
rect 19143 8188 19451 8197
rect 19143 8186 19149 8188
rect 19205 8186 19229 8188
rect 19285 8186 19309 8188
rect 19365 8186 19389 8188
rect 19445 8186 19451 8188
rect 19205 8134 19207 8186
rect 19387 8134 19389 8186
rect 19143 8132 19149 8134
rect 19205 8132 19229 8134
rect 19285 8132 19309 8134
rect 19365 8132 19389 8134
rect 19445 8132 19451 8134
rect 18878 8120 18934 8129
rect 19143 8123 19451 8132
rect 18878 8055 18934 8064
rect 18786 7712 18842 7721
rect 18786 7647 18842 7656
rect 18696 6656 18748 6662
rect 18696 6598 18748 6604
rect 18696 6452 18748 6458
rect 18696 6394 18748 6400
rect 18708 6361 18736 6394
rect 18694 6352 18750 6361
rect 18420 6316 18472 6322
rect 18800 6322 18828 7647
rect 18892 7410 18920 8055
rect 19432 7948 19484 7954
rect 19432 7890 19484 7896
rect 19076 7818 19380 7834
rect 19076 7812 19392 7818
rect 19076 7806 19340 7812
rect 18880 7404 18932 7410
rect 18880 7346 18932 7352
rect 18970 7304 19026 7313
rect 18970 7239 19026 7248
rect 18878 7032 18934 7041
rect 18878 6967 18934 6976
rect 18694 6287 18750 6296
rect 18788 6316 18840 6322
rect 18420 6258 18472 6264
rect 18788 6258 18840 6264
rect 18512 6248 18564 6254
rect 18512 6190 18564 6196
rect 18248 5902 18368 5930
rect 18144 5364 18196 5370
rect 18144 5306 18196 5312
rect 18248 5030 18276 5902
rect 18328 5840 18380 5846
rect 18328 5782 18380 5788
rect 18340 5681 18368 5782
rect 18524 5778 18552 6190
rect 18602 6080 18658 6089
rect 18602 6015 18658 6024
rect 18512 5772 18564 5778
rect 18512 5714 18564 5720
rect 18326 5672 18382 5681
rect 18326 5607 18382 5616
rect 18418 5536 18474 5545
rect 18418 5471 18474 5480
rect 18432 5302 18460 5471
rect 18512 5364 18564 5370
rect 18512 5306 18564 5312
rect 18420 5296 18472 5302
rect 18420 5238 18472 5244
rect 18236 5024 18288 5030
rect 18288 4984 18368 5012
rect 18236 4966 18288 4972
rect 18236 4752 18288 4758
rect 18236 4694 18288 4700
rect 18248 4457 18276 4694
rect 18234 4448 18290 4457
rect 18234 4383 18290 4392
rect 18234 4312 18290 4321
rect 18052 4276 18104 4282
rect 18234 4247 18290 4256
rect 18052 4218 18104 4224
rect 18064 4049 18092 4218
rect 18248 4146 18276 4247
rect 18236 4140 18288 4146
rect 18236 4082 18288 4088
rect 18050 4040 18106 4049
rect 18234 4040 18290 4049
rect 18050 3975 18106 3984
rect 18144 4004 18196 4010
rect 18234 3975 18290 3984
rect 18144 3946 18196 3952
rect 18052 3392 18104 3398
rect 18050 3360 18052 3369
rect 18104 3360 18106 3369
rect 18050 3295 18106 3304
rect 18156 3194 18184 3946
rect 18144 3188 18196 3194
rect 18144 3130 18196 3136
rect 18248 3058 18276 3975
rect 18340 3618 18368 4984
rect 18418 4992 18474 5001
rect 18418 4927 18474 4936
rect 18432 4010 18460 4927
rect 18420 4004 18472 4010
rect 18420 3946 18472 3952
rect 18418 3768 18474 3777
rect 18524 3738 18552 5306
rect 18616 4865 18644 6015
rect 18694 5944 18750 5953
rect 18694 5879 18750 5888
rect 18708 5642 18736 5879
rect 18892 5710 18920 6967
rect 18984 6866 19012 7239
rect 18972 6860 19024 6866
rect 18972 6802 19024 6808
rect 19076 6746 19104 7806
rect 19340 7754 19392 7760
rect 19444 7410 19472 7890
rect 19536 7546 19564 8910
rect 19616 8356 19668 8362
rect 19616 8298 19668 8304
rect 19524 7540 19576 7546
rect 19524 7482 19576 7488
rect 19432 7404 19484 7410
rect 19432 7346 19484 7352
rect 19143 7100 19451 7109
rect 19143 7098 19149 7100
rect 19205 7098 19229 7100
rect 19285 7098 19309 7100
rect 19365 7098 19389 7100
rect 19445 7098 19451 7100
rect 19205 7046 19207 7098
rect 19387 7046 19389 7098
rect 19143 7044 19149 7046
rect 19205 7044 19229 7046
rect 19285 7044 19309 7046
rect 19365 7044 19389 7046
rect 19445 7044 19451 7046
rect 19143 7035 19451 7044
rect 19248 6928 19300 6934
rect 19248 6870 19300 6876
rect 18984 6718 19104 6746
rect 19260 6730 19288 6870
rect 19628 6798 19656 8298
rect 19340 6792 19392 6798
rect 19340 6734 19392 6740
rect 19616 6792 19668 6798
rect 19616 6734 19668 6740
rect 19248 6724 19300 6730
rect 18788 5704 18840 5710
rect 18786 5672 18788 5681
rect 18880 5704 18932 5710
rect 18840 5672 18842 5681
rect 18696 5636 18748 5642
rect 18880 5646 18932 5652
rect 18786 5607 18842 5616
rect 18696 5578 18748 5584
rect 18696 5364 18748 5370
rect 18696 5306 18748 5312
rect 18602 4856 18658 4865
rect 18602 4791 18658 4800
rect 18604 4480 18656 4486
rect 18604 4422 18656 4428
rect 18616 4214 18644 4422
rect 18604 4208 18656 4214
rect 18604 4150 18656 4156
rect 18708 4146 18736 5306
rect 18984 4570 19012 6718
rect 19248 6666 19300 6672
rect 19064 6656 19116 6662
rect 19064 6598 19116 6604
rect 19156 6656 19208 6662
rect 19156 6598 19208 6604
rect 19076 5642 19104 6598
rect 19168 6497 19196 6598
rect 19154 6488 19210 6497
rect 19154 6423 19210 6432
rect 19248 6452 19300 6458
rect 19248 6394 19300 6400
rect 19260 6361 19288 6394
rect 19246 6352 19302 6361
rect 19246 6287 19302 6296
rect 19352 6186 19380 6734
rect 19340 6180 19392 6186
rect 19340 6122 19392 6128
rect 19143 6012 19451 6021
rect 19143 6010 19149 6012
rect 19205 6010 19229 6012
rect 19285 6010 19309 6012
rect 19365 6010 19389 6012
rect 19445 6010 19451 6012
rect 19205 5958 19207 6010
rect 19387 5958 19389 6010
rect 19143 5956 19149 5958
rect 19205 5956 19229 5958
rect 19285 5956 19309 5958
rect 19365 5956 19389 5958
rect 19445 5956 19451 5958
rect 19143 5947 19451 5956
rect 19156 5840 19208 5846
rect 19720 5794 19748 8996
rect 19904 8566 19932 9522
rect 19996 8906 20024 9590
rect 19984 8900 20036 8906
rect 19984 8842 20036 8848
rect 19892 8560 19944 8566
rect 19892 8502 19944 8508
rect 19800 8492 19852 8498
rect 19800 8434 19852 8440
rect 19812 7993 19840 8434
rect 19996 8430 20024 8842
rect 20088 8514 20116 11591
rect 20180 9586 20208 12056
rect 20272 10266 20300 19306
rect 20444 19168 20496 19174
rect 20444 19110 20496 19116
rect 20352 18896 20404 18902
rect 20352 18838 20404 18844
rect 20364 18426 20392 18838
rect 20456 18426 20484 19110
rect 20548 18970 20576 20198
rect 20628 19372 20680 19378
rect 20628 19314 20680 19320
rect 20536 18964 20588 18970
rect 20536 18906 20588 18912
rect 20536 18692 20588 18698
rect 20536 18634 20588 18640
rect 20548 18426 20576 18634
rect 20640 18630 20668 19314
rect 20720 19168 20772 19174
rect 20720 19110 20772 19116
rect 20628 18624 20680 18630
rect 20628 18566 20680 18572
rect 20352 18420 20404 18426
rect 20352 18362 20404 18368
rect 20444 18420 20496 18426
rect 20444 18362 20496 18368
rect 20536 18420 20588 18426
rect 20536 18362 20588 18368
rect 20640 18306 20668 18566
rect 20732 18426 20760 19110
rect 20720 18420 20772 18426
rect 20720 18362 20772 18368
rect 20548 18278 20668 18306
rect 20548 17678 20576 18278
rect 20720 18080 20772 18086
rect 20720 18022 20772 18028
rect 20628 17740 20680 17746
rect 20628 17682 20680 17688
rect 20536 17672 20588 17678
rect 20536 17614 20588 17620
rect 20352 17536 20404 17542
rect 20352 17478 20404 17484
rect 20364 17066 20392 17478
rect 20352 17060 20404 17066
rect 20352 17002 20404 17008
rect 20364 16794 20392 17002
rect 20640 16998 20668 17682
rect 20732 17202 20760 18022
rect 20824 17898 20852 20538
rect 20916 19854 20944 21490
rect 21008 20466 21036 21830
rect 20996 20460 21048 20466
rect 20996 20402 21048 20408
rect 20904 19848 20956 19854
rect 20904 19790 20956 19796
rect 20996 19168 21048 19174
rect 20996 19110 21048 19116
rect 20824 17882 20944 17898
rect 21008 17882 21036 19110
rect 21100 18850 21128 24074
rect 21192 23254 21220 29446
rect 21284 29170 21312 30903
rect 21364 30864 21416 30870
rect 21364 30806 21416 30812
rect 21272 29164 21324 29170
rect 21272 29106 21324 29112
rect 21272 28076 21324 28082
rect 21272 28018 21324 28024
rect 21284 27130 21312 28018
rect 21272 27124 21324 27130
rect 21272 27066 21324 27072
rect 21272 26920 21324 26926
rect 21272 26862 21324 26868
rect 21284 26586 21312 26862
rect 21272 26580 21324 26586
rect 21376 26568 21404 30806
rect 21456 30048 21508 30054
rect 21454 30016 21456 30025
rect 21508 30016 21510 30025
rect 21454 29951 21510 29960
rect 21456 28960 21508 28966
rect 21454 28928 21456 28937
rect 21508 28928 21510 28937
rect 21454 28863 21510 28872
rect 21456 27872 21508 27878
rect 21456 27814 21508 27820
rect 21468 27033 21496 27814
rect 21454 27024 21510 27033
rect 21454 26959 21510 26968
rect 21376 26540 21496 26568
rect 21272 26522 21324 26528
rect 21468 26364 21496 26540
rect 21376 26336 21496 26364
rect 21272 26308 21324 26314
rect 21272 26250 21324 26256
rect 21284 25294 21312 26250
rect 21272 25288 21324 25294
rect 21272 25230 21324 25236
rect 21180 23248 21232 23254
rect 21180 23190 21232 23196
rect 21376 23100 21404 26336
rect 21456 25696 21508 25702
rect 21454 25664 21456 25673
rect 21508 25664 21510 25673
rect 21454 25599 21510 25608
rect 21456 24608 21508 24614
rect 21454 24576 21456 24585
rect 21508 24576 21510 24585
rect 21454 24511 21510 24520
rect 21560 24138 21588 31855
rect 21652 30258 21680 32982
rect 21742 32668 22050 32677
rect 21742 32666 21748 32668
rect 21804 32666 21828 32668
rect 21884 32666 21908 32668
rect 21964 32666 21988 32668
rect 22044 32666 22050 32668
rect 21804 32614 21806 32666
rect 21986 32614 21988 32666
rect 21742 32612 21748 32614
rect 21804 32612 21828 32614
rect 21884 32612 21908 32614
rect 21964 32612 21988 32614
rect 22044 32612 22050 32614
rect 21742 32603 22050 32612
rect 21742 31580 22050 31589
rect 21742 31578 21748 31580
rect 21804 31578 21828 31580
rect 21884 31578 21908 31580
rect 21964 31578 21988 31580
rect 22044 31578 22050 31580
rect 21804 31526 21806 31578
rect 21986 31526 21988 31578
rect 21742 31524 21748 31526
rect 21804 31524 21828 31526
rect 21884 31524 21908 31526
rect 21964 31524 21988 31526
rect 22044 31524 22050 31526
rect 21742 31515 22050 31524
rect 21742 30492 22050 30501
rect 21742 30490 21748 30492
rect 21804 30490 21828 30492
rect 21884 30490 21908 30492
rect 21964 30490 21988 30492
rect 22044 30490 22050 30492
rect 21804 30438 21806 30490
rect 21986 30438 21988 30490
rect 21742 30436 21748 30438
rect 21804 30436 21828 30438
rect 21884 30436 21908 30438
rect 21964 30436 21988 30438
rect 22044 30436 22050 30438
rect 21742 30427 22050 30436
rect 21640 30252 21692 30258
rect 21640 30194 21692 30200
rect 21742 29404 22050 29413
rect 21742 29402 21748 29404
rect 21804 29402 21828 29404
rect 21884 29402 21908 29404
rect 21964 29402 21988 29404
rect 22044 29402 22050 29404
rect 21804 29350 21806 29402
rect 21986 29350 21988 29402
rect 21742 29348 21748 29350
rect 21804 29348 21828 29350
rect 21884 29348 21908 29350
rect 21964 29348 21988 29350
rect 22044 29348 22050 29350
rect 21742 29339 22050 29348
rect 21742 28316 22050 28325
rect 21742 28314 21748 28316
rect 21804 28314 21828 28316
rect 21884 28314 21908 28316
rect 21964 28314 21988 28316
rect 22044 28314 22050 28316
rect 21804 28262 21806 28314
rect 21986 28262 21988 28314
rect 21742 28260 21748 28262
rect 21804 28260 21828 28262
rect 21884 28260 21908 28262
rect 21964 28260 21988 28262
rect 22044 28260 22050 28262
rect 21742 28251 22050 28260
rect 21640 27532 21692 27538
rect 21640 27474 21692 27480
rect 21548 24132 21600 24138
rect 21548 24074 21600 24080
rect 21546 23488 21602 23497
rect 21546 23423 21602 23432
rect 21560 23322 21588 23423
rect 21548 23316 21600 23322
rect 21548 23258 21600 23264
rect 21192 23072 21404 23100
rect 21192 21876 21220 23072
rect 21546 22808 21602 22817
rect 21546 22743 21602 22752
rect 21560 22574 21588 22743
rect 21652 22658 21680 27474
rect 21742 27228 22050 27237
rect 21742 27226 21748 27228
rect 21804 27226 21828 27228
rect 21884 27226 21908 27228
rect 21964 27226 21988 27228
rect 22044 27226 22050 27228
rect 21804 27174 21806 27226
rect 21986 27174 21988 27226
rect 21742 27172 21748 27174
rect 21804 27172 21828 27174
rect 21884 27172 21908 27174
rect 21964 27172 21988 27174
rect 22044 27172 22050 27174
rect 21742 27163 22050 27172
rect 21742 26140 22050 26149
rect 21742 26138 21748 26140
rect 21804 26138 21828 26140
rect 21884 26138 21908 26140
rect 21964 26138 21988 26140
rect 22044 26138 22050 26140
rect 21804 26086 21806 26138
rect 21986 26086 21988 26138
rect 21742 26084 21748 26086
rect 21804 26084 21828 26086
rect 21884 26084 21908 26086
rect 21964 26084 21988 26086
rect 22044 26084 22050 26086
rect 21742 26075 22050 26084
rect 21742 25052 22050 25061
rect 21742 25050 21748 25052
rect 21804 25050 21828 25052
rect 21884 25050 21908 25052
rect 21964 25050 21988 25052
rect 22044 25050 22050 25052
rect 21804 24998 21806 25050
rect 21986 24998 21988 25050
rect 21742 24996 21748 24998
rect 21804 24996 21828 24998
rect 21884 24996 21908 24998
rect 21964 24996 21988 24998
rect 22044 24996 22050 24998
rect 21742 24987 22050 24996
rect 22008 24948 22060 24954
rect 22008 24890 22060 24896
rect 22020 24154 22048 24890
rect 22112 24834 22140 33238
rect 22204 31754 22232 33374
rect 22296 32502 22324 34546
rect 22284 32496 22336 32502
rect 22284 32438 22336 32444
rect 22284 32360 22336 32366
rect 22284 32302 22336 32308
rect 22296 31872 22324 32302
rect 22296 31844 22416 31872
rect 22204 31726 22324 31754
rect 22192 31680 22244 31686
rect 22190 31648 22192 31657
rect 22244 31648 22246 31657
rect 22190 31583 22246 31592
rect 22296 30802 22324 31726
rect 22284 30796 22336 30802
rect 22284 30738 22336 30744
rect 22284 30660 22336 30666
rect 22284 30602 22336 30608
rect 22296 30569 22324 30602
rect 22282 30560 22338 30569
rect 22282 30495 22338 30504
rect 22192 29504 22244 29510
rect 22190 29472 22192 29481
rect 22244 29472 22246 29481
rect 22190 29407 22246 29416
rect 22192 29096 22244 29102
rect 22192 29038 22244 29044
rect 22204 28506 22232 29038
rect 22204 28478 22324 28506
rect 22192 28416 22244 28422
rect 22190 28384 22192 28393
rect 22244 28384 22246 28393
rect 22190 28319 22246 28328
rect 22192 27396 22244 27402
rect 22192 27338 22244 27344
rect 22204 27305 22232 27338
rect 22190 27296 22246 27305
rect 22190 27231 22246 27240
rect 22296 26466 22324 28478
rect 22204 26438 22324 26466
rect 22204 24954 22232 26438
rect 22284 26308 22336 26314
rect 22284 26250 22336 26256
rect 22296 26217 22324 26250
rect 22282 26208 22338 26217
rect 22282 26143 22338 26152
rect 22284 25220 22336 25226
rect 22284 25162 22336 25168
rect 22296 25129 22324 25162
rect 22282 25120 22338 25129
rect 22282 25055 22338 25064
rect 22192 24948 22244 24954
rect 22192 24890 22244 24896
rect 22112 24806 22324 24834
rect 22020 24126 22140 24154
rect 21742 23964 22050 23973
rect 21742 23962 21748 23964
rect 21804 23962 21828 23964
rect 21884 23962 21908 23964
rect 21964 23962 21988 23964
rect 22044 23962 22050 23964
rect 21804 23910 21806 23962
rect 21986 23910 21988 23962
rect 21742 23908 21748 23910
rect 21804 23908 21828 23910
rect 21884 23908 21908 23910
rect 21964 23908 21988 23910
rect 22044 23908 22050 23910
rect 21742 23899 22050 23908
rect 21742 22876 22050 22885
rect 21742 22874 21748 22876
rect 21804 22874 21828 22876
rect 21884 22874 21908 22876
rect 21964 22874 21988 22876
rect 22044 22874 22050 22876
rect 21804 22822 21806 22874
rect 21986 22822 21988 22874
rect 21742 22820 21748 22822
rect 21804 22820 21828 22822
rect 21884 22820 21908 22822
rect 21964 22820 21988 22822
rect 22044 22820 22050 22822
rect 21742 22811 22050 22820
rect 21916 22704 21968 22710
rect 21652 22642 21772 22658
rect 22112 22658 22140 24126
rect 22192 24064 22244 24070
rect 22190 24032 22192 24041
rect 22244 24032 22246 24041
rect 22190 23967 22246 23976
rect 22190 22944 22246 22953
rect 22190 22879 22246 22888
rect 22204 22778 22232 22879
rect 22192 22772 22244 22778
rect 22192 22714 22244 22720
rect 21916 22646 21968 22652
rect 21652 22636 21784 22642
rect 21652 22630 21732 22636
rect 21732 22578 21784 22584
rect 21548 22568 21600 22574
rect 21548 22510 21600 22516
rect 21272 22500 21324 22506
rect 21272 22442 21324 22448
rect 21284 22030 21312 22442
rect 21364 22432 21416 22438
rect 21364 22374 21416 22380
rect 21454 22400 21510 22409
rect 21376 22030 21404 22374
rect 21454 22335 21510 22344
rect 21468 22234 21496 22335
rect 21456 22228 21508 22234
rect 21456 22170 21508 22176
rect 21546 22128 21602 22137
rect 21456 22094 21508 22098
rect 21456 22092 21546 22094
rect 21508 22072 21546 22092
rect 21928 22094 21956 22646
rect 22020 22630 22140 22658
rect 22190 22672 22246 22681
rect 22020 22137 22048 22630
rect 22190 22607 22246 22616
rect 22098 22536 22154 22545
rect 22098 22471 22154 22480
rect 21508 22066 21602 22072
rect 21546 22063 21602 22066
rect 21652 22066 21956 22094
rect 22006 22128 22062 22137
rect 21456 22034 21508 22040
rect 21272 22024 21324 22030
rect 21272 21966 21324 21972
rect 21364 22024 21416 22030
rect 21468 22003 21496 22034
rect 21548 22024 21600 22030
rect 21364 21966 21416 21972
rect 21548 21966 21600 21972
rect 21192 21848 21496 21876
rect 21364 21480 21416 21486
rect 21364 21422 21416 21428
rect 21180 21344 21232 21350
rect 21180 21286 21232 21292
rect 21272 21344 21324 21350
rect 21272 21286 21324 21292
rect 21192 20602 21220 21286
rect 21284 20942 21312 21286
rect 21272 20936 21324 20942
rect 21272 20878 21324 20884
rect 21270 20768 21326 20777
rect 21270 20703 21326 20712
rect 21180 20596 21232 20602
rect 21180 20538 21232 20544
rect 21180 20256 21232 20262
rect 21180 20198 21232 20204
rect 21192 19854 21220 20198
rect 21180 19848 21232 19854
rect 21180 19790 21232 19796
rect 21180 19372 21232 19378
rect 21180 19314 21232 19320
rect 21192 18970 21220 19314
rect 21180 18964 21232 18970
rect 21180 18906 21232 18912
rect 21100 18822 21220 18850
rect 20824 17876 20956 17882
rect 20824 17870 20904 17876
rect 20904 17818 20956 17824
rect 20996 17876 21048 17882
rect 20996 17818 21048 17824
rect 20812 17808 20864 17814
rect 20812 17750 20864 17756
rect 20720 17196 20772 17202
rect 20720 17138 20772 17144
rect 20536 16992 20588 16998
rect 20536 16934 20588 16940
rect 20628 16992 20680 16998
rect 20628 16934 20680 16940
rect 20352 16788 20404 16794
rect 20352 16730 20404 16736
rect 20352 14816 20404 14822
rect 20352 14758 20404 14764
rect 20364 14618 20392 14758
rect 20352 14612 20404 14618
rect 20352 14554 20404 14560
rect 20548 12238 20576 16934
rect 20720 16584 20772 16590
rect 20720 16526 20772 16532
rect 20732 16250 20760 16526
rect 20824 16250 20852 17750
rect 20904 17536 20956 17542
rect 20904 17478 20956 17484
rect 20916 17338 20944 17478
rect 20904 17332 20956 17338
rect 20904 17274 20956 17280
rect 20904 16652 20956 16658
rect 20904 16594 20956 16600
rect 20720 16244 20772 16250
rect 20720 16186 20772 16192
rect 20812 16244 20864 16250
rect 20812 16186 20864 16192
rect 20732 15502 20760 16186
rect 20916 15706 20944 16594
rect 21088 16584 21140 16590
rect 21088 16526 21140 16532
rect 20996 16448 21048 16454
rect 20996 16390 21048 16396
rect 21008 16250 21036 16390
rect 21100 16250 21128 16526
rect 20996 16244 21048 16250
rect 20996 16186 21048 16192
rect 21088 16244 21140 16250
rect 21088 16186 21140 16192
rect 20904 15700 20956 15706
rect 20904 15642 20956 15648
rect 21192 15502 21220 18822
rect 21284 17678 21312 20703
rect 21376 19854 21404 21422
rect 21468 20806 21496 21848
rect 21456 20800 21508 20806
rect 21456 20742 21508 20748
rect 21456 20256 21508 20262
rect 21454 20224 21456 20233
rect 21508 20224 21510 20233
rect 21454 20159 21510 20168
rect 21364 19848 21416 19854
rect 21364 19790 21416 19796
rect 21362 19408 21418 19417
rect 21362 19343 21418 19352
rect 21272 17672 21324 17678
rect 21272 17614 21324 17620
rect 21270 17232 21326 17241
rect 21270 17167 21326 17176
rect 20720 15496 20772 15502
rect 20720 15438 20772 15444
rect 21180 15496 21232 15502
rect 21180 15438 21232 15444
rect 21088 15428 21140 15434
rect 21088 15370 21140 15376
rect 20720 15360 20772 15366
rect 20720 15302 20772 15308
rect 20810 15328 20866 15337
rect 20732 15162 20760 15302
rect 20810 15263 20866 15272
rect 20720 15156 20772 15162
rect 20720 15098 20772 15104
rect 20720 13932 20772 13938
rect 20720 13874 20772 13880
rect 20732 13326 20760 13874
rect 20824 13530 20852 15263
rect 20904 15020 20956 15026
rect 20904 14962 20956 14968
rect 20916 14618 20944 14962
rect 20996 14816 21048 14822
rect 20996 14758 21048 14764
rect 21008 14618 21036 14758
rect 20904 14612 20956 14618
rect 20904 14554 20956 14560
rect 20996 14612 21048 14618
rect 20996 14554 21048 14560
rect 21100 14414 21128 15370
rect 21088 14408 21140 14414
rect 21088 14350 21140 14356
rect 21180 14272 21232 14278
rect 21180 14214 21232 14220
rect 21192 14074 21220 14214
rect 21088 14068 21140 14074
rect 21088 14010 21140 14016
rect 21180 14068 21232 14074
rect 21180 14010 21232 14016
rect 20812 13524 20864 13530
rect 20812 13466 20864 13472
rect 20720 13320 20772 13326
rect 20720 13262 20772 13268
rect 20628 13184 20680 13190
rect 20628 13126 20680 13132
rect 21100 13138 21128 14010
rect 21178 13968 21234 13977
rect 21178 13903 21234 13912
rect 21192 13546 21220 13903
rect 21284 13734 21312 17167
rect 21272 13728 21324 13734
rect 21272 13670 21324 13676
rect 21192 13518 21312 13546
rect 20640 12918 20668 13126
rect 21100 13110 21220 13138
rect 20628 12912 20680 12918
rect 20628 12854 20680 12860
rect 20640 12306 20668 12854
rect 20904 12776 20956 12782
rect 20904 12718 20956 12724
rect 20720 12640 20772 12646
rect 20720 12582 20772 12588
rect 20628 12300 20680 12306
rect 20628 12242 20680 12248
rect 20732 12238 20760 12582
rect 20916 12442 20944 12718
rect 21088 12640 21140 12646
rect 21086 12608 21088 12617
rect 21140 12608 21142 12617
rect 21086 12543 21142 12552
rect 20904 12436 20956 12442
rect 20904 12378 20956 12384
rect 20996 12368 21048 12374
rect 20810 12336 20866 12345
rect 20996 12310 21048 12316
rect 20810 12271 20866 12280
rect 20444 12232 20496 12238
rect 20444 12174 20496 12180
rect 20536 12232 20588 12238
rect 20536 12174 20588 12180
rect 20720 12232 20772 12238
rect 20720 12174 20772 12180
rect 20352 12096 20404 12102
rect 20352 12038 20404 12044
rect 20364 11898 20392 12038
rect 20456 11898 20484 12174
rect 20628 12164 20680 12170
rect 20628 12106 20680 12112
rect 20640 12050 20668 12106
rect 20640 12022 20760 12050
rect 20352 11892 20404 11898
rect 20352 11834 20404 11840
rect 20444 11892 20496 11898
rect 20444 11834 20496 11840
rect 20732 10742 20760 12022
rect 20720 10736 20772 10742
rect 20720 10678 20772 10684
rect 20352 10464 20404 10470
rect 20352 10406 20404 10412
rect 20364 10266 20392 10406
rect 20260 10260 20312 10266
rect 20260 10202 20312 10208
rect 20352 10260 20404 10266
rect 20352 10202 20404 10208
rect 20260 9920 20312 9926
rect 20260 9862 20312 9868
rect 20536 9920 20588 9926
rect 20536 9862 20588 9868
rect 20272 9586 20300 9862
rect 20168 9580 20220 9586
rect 20168 9522 20220 9528
rect 20260 9580 20312 9586
rect 20260 9522 20312 9528
rect 20272 9024 20300 9522
rect 20352 9444 20404 9450
rect 20352 9386 20404 9392
rect 20180 8996 20300 9024
rect 20180 8906 20208 8996
rect 20258 8936 20314 8945
rect 20168 8900 20220 8906
rect 20258 8871 20314 8880
rect 20168 8842 20220 8848
rect 20272 8838 20300 8871
rect 20260 8832 20312 8838
rect 20260 8774 20312 8780
rect 20088 8486 20208 8514
rect 19984 8424 20036 8430
rect 19984 8366 20036 8372
rect 19798 7984 19854 7993
rect 19798 7919 19854 7928
rect 19984 7744 20036 7750
rect 19984 7686 20036 7692
rect 19892 7404 19944 7410
rect 19892 7346 19944 7352
rect 19800 7336 19852 7342
rect 19800 7278 19852 7284
rect 19208 5788 19748 5794
rect 19156 5782 19748 5788
rect 19168 5766 19748 5782
rect 19154 5672 19210 5681
rect 19064 5636 19116 5642
rect 19210 5630 19380 5658
rect 19154 5607 19210 5616
rect 19064 5578 19116 5584
rect 19352 5522 19380 5630
rect 19352 5494 19564 5522
rect 19536 5166 19564 5494
rect 19524 5160 19576 5166
rect 19524 5102 19576 5108
rect 19064 5024 19116 5030
rect 19064 4966 19116 4972
rect 19076 4758 19104 4966
rect 19143 4924 19451 4933
rect 19143 4922 19149 4924
rect 19205 4922 19229 4924
rect 19285 4922 19309 4924
rect 19365 4922 19389 4924
rect 19445 4922 19451 4924
rect 19205 4870 19207 4922
rect 19387 4870 19389 4922
rect 19143 4868 19149 4870
rect 19205 4868 19229 4870
rect 19285 4868 19309 4870
rect 19365 4868 19389 4870
rect 19445 4868 19451 4870
rect 19143 4859 19451 4868
rect 19536 4826 19564 5102
rect 19524 4820 19576 4826
rect 19524 4762 19576 4768
rect 19064 4752 19116 4758
rect 19064 4694 19116 4700
rect 19340 4684 19392 4690
rect 19340 4626 19392 4632
rect 19248 4616 19300 4622
rect 18984 4542 19196 4570
rect 19248 4558 19300 4564
rect 19064 4480 19116 4486
rect 19064 4422 19116 4428
rect 18696 4140 18748 4146
rect 18696 4082 18748 4088
rect 18972 4140 19024 4146
rect 18972 4082 19024 4088
rect 18788 3936 18840 3942
rect 18788 3878 18840 3884
rect 18878 3904 18934 3913
rect 18800 3738 18828 3878
rect 18878 3839 18934 3848
rect 18418 3703 18420 3712
rect 18472 3703 18474 3712
rect 18512 3732 18564 3738
rect 18420 3674 18472 3680
rect 18512 3674 18564 3680
rect 18788 3732 18840 3738
rect 18788 3674 18840 3680
rect 18340 3590 18552 3618
rect 18328 3528 18380 3534
rect 18328 3470 18380 3476
rect 18340 3369 18368 3470
rect 18420 3392 18472 3398
rect 18326 3360 18382 3369
rect 18420 3334 18472 3340
rect 18326 3295 18382 3304
rect 18432 3176 18460 3334
rect 18524 3194 18552 3590
rect 18604 3528 18656 3534
rect 18604 3470 18656 3476
rect 18696 3528 18748 3534
rect 18696 3470 18748 3476
rect 18616 3233 18644 3470
rect 18602 3224 18658 3233
rect 18340 3148 18460 3176
rect 18512 3188 18564 3194
rect 17960 3052 18012 3058
rect 17960 2994 18012 3000
rect 18236 3052 18288 3058
rect 18236 2994 18288 3000
rect 18052 2984 18104 2990
rect 17958 2952 18014 2961
rect 18340 2938 18368 3148
rect 18602 3159 18658 3168
rect 18512 3130 18564 3136
rect 18420 3052 18472 3058
rect 18420 2994 18472 3000
rect 18104 2932 18368 2938
rect 18052 2926 18368 2932
rect 18064 2910 18368 2926
rect 17958 2887 18014 2896
rect 17776 2848 17828 2854
rect 17776 2790 17828 2796
rect 17590 2544 17646 2553
rect 17590 2479 17592 2488
rect 17644 2479 17646 2488
rect 17684 2508 17736 2514
rect 17592 2450 17644 2456
rect 17684 2450 17736 2456
rect 17696 2394 17724 2450
rect 17788 2446 17816 2790
rect 17604 2366 17724 2394
rect 17776 2440 17828 2446
rect 17776 2382 17828 2388
rect 17500 1012 17552 1018
rect 17500 954 17552 960
rect 17130 54 17264 82
rect 17130 -300 17186 54
rect 17314 -300 17370 160
rect 17498 82 17554 160
rect 17604 82 17632 2366
rect 17868 1964 17920 1970
rect 17868 1906 17920 1912
rect 17684 1284 17736 1290
rect 17684 1226 17736 1232
rect 17696 160 17724 1226
rect 17880 160 17908 1906
rect 17972 1426 18000 2887
rect 18052 2576 18104 2582
rect 18052 2518 18104 2524
rect 17960 1420 18012 1426
rect 17960 1362 18012 1368
rect 18064 160 18092 2518
rect 18328 2304 18380 2310
rect 18328 2246 18380 2252
rect 18340 1902 18368 2246
rect 18328 1896 18380 1902
rect 18328 1838 18380 1844
rect 18142 1592 18198 1601
rect 18142 1527 18198 1536
rect 18156 1222 18184 1527
rect 18144 1216 18196 1222
rect 18144 1158 18196 1164
rect 18432 218 18460 2994
rect 18602 2816 18658 2825
rect 18602 2751 18658 2760
rect 18510 2680 18566 2689
rect 18510 2615 18566 2624
rect 18524 2446 18552 2615
rect 18512 2440 18564 2446
rect 18512 2382 18564 2388
rect 18512 1420 18564 1426
rect 18512 1362 18564 1368
rect 18340 190 18460 218
rect 17498 54 17632 82
rect 17498 -300 17554 54
rect 17682 -300 17738 160
rect 17866 -300 17922 160
rect 18050 -300 18106 160
rect 18234 82 18290 160
rect 18340 82 18368 190
rect 18234 54 18368 82
rect 18418 82 18474 160
rect 18524 82 18552 1362
rect 18616 1340 18644 2751
rect 18708 2553 18736 3470
rect 18892 2854 18920 3839
rect 18880 2848 18932 2854
rect 18880 2790 18932 2796
rect 18694 2544 18750 2553
rect 18694 2479 18750 2488
rect 18696 2440 18748 2446
rect 18694 2408 18696 2417
rect 18748 2408 18750 2417
rect 18694 2343 18750 2352
rect 18880 2100 18932 2106
rect 18880 2042 18932 2048
rect 18788 2032 18840 2038
rect 18788 1974 18840 1980
rect 18696 1352 18748 1358
rect 18616 1312 18696 1340
rect 18696 1294 18748 1300
rect 18604 1216 18656 1222
rect 18604 1158 18656 1164
rect 18616 160 18644 1158
rect 18800 160 18828 1974
rect 18892 1884 18920 2042
rect 18984 2009 19012 4082
rect 19076 3058 19104 4422
rect 19168 4282 19196 4542
rect 19156 4276 19208 4282
rect 19156 4218 19208 4224
rect 19260 4049 19288 4558
rect 19352 4282 19380 4626
rect 19524 4616 19576 4622
rect 19522 4584 19524 4593
rect 19576 4584 19578 4593
rect 19522 4519 19578 4528
rect 19524 4480 19576 4486
rect 19524 4422 19576 4428
rect 19616 4480 19668 4486
rect 19616 4422 19668 4428
rect 19340 4276 19392 4282
rect 19340 4218 19392 4224
rect 19246 4040 19302 4049
rect 19246 3975 19302 3984
rect 19143 3836 19451 3845
rect 19143 3834 19149 3836
rect 19205 3834 19229 3836
rect 19285 3834 19309 3836
rect 19365 3834 19389 3836
rect 19445 3834 19451 3836
rect 19205 3782 19207 3834
rect 19387 3782 19389 3834
rect 19143 3780 19149 3782
rect 19205 3780 19229 3782
rect 19285 3780 19309 3782
rect 19365 3780 19389 3782
rect 19445 3780 19451 3782
rect 19143 3771 19451 3780
rect 19536 3058 19564 4422
rect 19628 3194 19656 4422
rect 19708 4208 19760 4214
rect 19708 4150 19760 4156
rect 19616 3188 19668 3194
rect 19616 3130 19668 3136
rect 19064 3052 19116 3058
rect 19064 2994 19116 3000
rect 19524 3052 19576 3058
rect 19524 2994 19576 3000
rect 19352 2922 19564 2938
rect 19340 2916 19564 2922
rect 19392 2910 19564 2916
rect 19340 2858 19392 2864
rect 19064 2848 19116 2854
rect 19064 2790 19116 2796
rect 18970 2000 19026 2009
rect 18970 1935 19026 1944
rect 18892 1856 19012 1884
rect 18984 160 19012 1856
rect 18418 54 18552 82
rect 18234 -300 18290 54
rect 18418 -300 18474 54
rect 18602 -300 18658 160
rect 18786 -300 18842 160
rect 18970 -300 19026 160
rect 19076 82 19104 2790
rect 19143 2748 19451 2757
rect 19143 2746 19149 2748
rect 19205 2746 19229 2748
rect 19285 2746 19309 2748
rect 19365 2746 19389 2748
rect 19445 2746 19451 2748
rect 19205 2694 19207 2746
rect 19387 2694 19389 2746
rect 19143 2692 19149 2694
rect 19205 2692 19229 2694
rect 19285 2692 19309 2694
rect 19365 2692 19389 2694
rect 19445 2692 19451 2694
rect 19143 2683 19451 2692
rect 19143 1660 19451 1669
rect 19143 1658 19149 1660
rect 19205 1658 19229 1660
rect 19285 1658 19309 1660
rect 19365 1658 19389 1660
rect 19445 1658 19451 1660
rect 19205 1606 19207 1658
rect 19387 1606 19389 1658
rect 19143 1604 19149 1606
rect 19205 1604 19229 1606
rect 19285 1604 19309 1606
rect 19365 1604 19389 1606
rect 19445 1604 19451 1606
rect 19143 1595 19451 1604
rect 19536 218 19564 2910
rect 19720 2774 19748 4150
rect 19812 3380 19840 7278
rect 19904 6322 19932 7346
rect 19996 7206 20024 7686
rect 20076 7404 20128 7410
rect 20076 7346 20128 7352
rect 19984 7200 20036 7206
rect 19984 7142 20036 7148
rect 19892 6316 19944 6322
rect 19892 6258 19944 6264
rect 19904 4690 19932 6258
rect 19996 5710 20024 7142
rect 20088 6934 20116 7346
rect 20076 6928 20128 6934
rect 20076 6870 20128 6876
rect 20180 6746 20208 8486
rect 20088 6718 20208 6746
rect 19984 5704 20036 5710
rect 19984 5646 20036 5652
rect 19892 4684 19944 4690
rect 19892 4626 19944 4632
rect 19904 3942 19932 4626
rect 20088 4321 20116 6718
rect 20168 6384 20220 6390
rect 20168 6326 20220 6332
rect 20180 5817 20208 6326
rect 20166 5808 20222 5817
rect 20166 5743 20222 5752
rect 20272 5234 20300 8774
rect 20364 8566 20392 9386
rect 20352 8560 20404 8566
rect 20352 8502 20404 8508
rect 20352 8288 20404 8294
rect 20352 8230 20404 8236
rect 20260 5228 20312 5234
rect 20260 5170 20312 5176
rect 20074 4312 20130 4321
rect 20074 4247 20130 4256
rect 19984 4208 20036 4214
rect 19984 4150 20036 4156
rect 19892 3936 19944 3942
rect 19892 3878 19944 3884
rect 19904 3534 19932 3878
rect 19892 3528 19944 3534
rect 19892 3470 19944 3476
rect 19996 3398 20024 4150
rect 20074 4040 20130 4049
rect 20074 3975 20130 3984
rect 19984 3392 20036 3398
rect 19812 3352 19932 3380
rect 19800 2984 19852 2990
rect 19800 2926 19852 2932
rect 19444 190 19564 218
rect 19628 2746 19748 2774
rect 19154 82 19210 160
rect 19076 54 19210 82
rect 19154 -300 19210 54
rect 19338 82 19394 160
rect 19444 82 19472 190
rect 19338 54 19472 82
rect 19522 82 19578 160
rect 19628 82 19656 2746
rect 19522 54 19656 82
rect 19706 82 19762 160
rect 19812 82 19840 2926
rect 19904 2774 19932 3352
rect 19984 3334 20036 3340
rect 20088 3194 20116 3975
rect 20260 3936 20312 3942
rect 20166 3904 20222 3913
rect 20260 3878 20312 3884
rect 20166 3839 20222 3848
rect 20076 3188 20128 3194
rect 20076 3130 20128 3136
rect 19904 2746 20116 2774
rect 20088 2514 20116 2746
rect 20076 2508 20128 2514
rect 20076 2450 20128 2456
rect 20180 2378 20208 3839
rect 20168 2372 20220 2378
rect 20168 2314 20220 2320
rect 19706 54 19840 82
rect 19890 82 19946 160
rect 20272 82 20300 3878
rect 20364 2038 20392 8230
rect 20444 3732 20496 3738
rect 20444 3674 20496 3680
rect 20456 3058 20484 3674
rect 20444 3052 20496 3058
rect 20444 2994 20496 3000
rect 20548 2922 20576 9862
rect 20628 8832 20680 8838
rect 20628 8774 20680 8780
rect 20640 8634 20668 8774
rect 20628 8628 20680 8634
rect 20628 8570 20680 8576
rect 20824 8378 20852 12271
rect 21008 11778 21036 12310
rect 21088 12096 21140 12102
rect 21088 12038 21140 12044
rect 20916 11750 21036 11778
rect 20916 10554 20944 11750
rect 20996 11620 21048 11626
rect 20996 11562 21048 11568
rect 21008 11257 21036 11562
rect 21100 11529 21128 12038
rect 21192 11762 21220 13110
rect 21180 11756 21232 11762
rect 21180 11698 21232 11704
rect 21086 11520 21142 11529
rect 21086 11455 21142 11464
rect 20994 11248 21050 11257
rect 20994 11183 21050 11192
rect 21284 10713 21312 13518
rect 21376 13274 21404 19343
rect 21456 19168 21508 19174
rect 21454 19136 21456 19145
rect 21508 19136 21510 19145
rect 21454 19071 21510 19080
rect 21456 18080 21508 18086
rect 21454 18048 21456 18057
rect 21508 18048 21510 18057
rect 21454 17983 21510 17992
rect 21456 16992 21508 16998
rect 21454 16960 21456 16969
rect 21508 16960 21510 16969
rect 21454 16895 21510 16904
rect 21456 16652 21508 16658
rect 21456 16594 21508 16600
rect 21468 16561 21496 16594
rect 21454 16552 21510 16561
rect 21454 16487 21510 16496
rect 21456 15904 21508 15910
rect 21454 15872 21456 15881
rect 21508 15872 21510 15881
rect 21454 15807 21510 15816
rect 21560 14929 21588 21966
rect 21546 14920 21602 14929
rect 21546 14855 21602 14864
rect 21456 14816 21508 14822
rect 21454 14784 21456 14793
rect 21508 14784 21510 14793
rect 21454 14719 21510 14728
rect 21456 13728 21508 13734
rect 21454 13696 21456 13705
rect 21508 13696 21510 13705
rect 21454 13631 21510 13640
rect 21652 13512 21680 22066
rect 22006 22063 22062 22072
rect 21742 21788 22050 21797
rect 21742 21786 21748 21788
rect 21804 21786 21828 21788
rect 21884 21786 21908 21788
rect 21964 21786 21988 21788
rect 22044 21786 22050 21788
rect 21804 21734 21806 21786
rect 21986 21734 21988 21786
rect 21742 21732 21748 21734
rect 21804 21732 21828 21734
rect 21884 21732 21908 21734
rect 21964 21732 21988 21734
rect 22044 21732 22050 21734
rect 21742 21723 22050 21732
rect 22112 20913 22140 22471
rect 22204 22030 22232 22607
rect 22192 22024 22244 22030
rect 22192 21966 22244 21972
rect 22192 21888 22244 21894
rect 22190 21856 22192 21865
rect 22244 21856 22246 21865
rect 22190 21791 22246 21800
rect 22098 20904 22154 20913
rect 22098 20839 22154 20848
rect 22192 20868 22244 20874
rect 22192 20810 22244 20816
rect 22204 20777 22232 20810
rect 22190 20768 22246 20777
rect 21742 20700 22050 20709
rect 22190 20703 22246 20712
rect 21742 20698 21748 20700
rect 21804 20698 21828 20700
rect 21884 20698 21908 20700
rect 21964 20698 21988 20700
rect 22044 20698 22050 20700
rect 21804 20646 21806 20698
rect 21986 20646 21988 20698
rect 21742 20644 21748 20646
rect 21804 20644 21828 20646
rect 21884 20644 21908 20646
rect 21964 20644 21988 20646
rect 22044 20644 22050 20646
rect 21742 20635 22050 20644
rect 22098 19816 22154 19825
rect 22098 19751 22154 19760
rect 21742 19612 22050 19621
rect 21742 19610 21748 19612
rect 21804 19610 21828 19612
rect 21884 19610 21908 19612
rect 21964 19610 21988 19612
rect 22044 19610 22050 19612
rect 21804 19558 21806 19610
rect 21986 19558 21988 19610
rect 21742 19556 21748 19558
rect 21804 19556 21828 19558
rect 21884 19556 21908 19558
rect 21964 19556 21988 19558
rect 22044 19556 22050 19558
rect 21742 19547 22050 19556
rect 21742 18524 22050 18533
rect 21742 18522 21748 18524
rect 21804 18522 21828 18524
rect 21884 18522 21908 18524
rect 21964 18522 21988 18524
rect 22044 18522 22050 18524
rect 21804 18470 21806 18522
rect 21986 18470 21988 18522
rect 21742 18468 21748 18470
rect 21804 18468 21828 18470
rect 21884 18468 21908 18470
rect 21964 18468 21988 18470
rect 22044 18468 22050 18470
rect 21742 18459 22050 18468
rect 21742 17436 22050 17445
rect 21742 17434 21748 17436
rect 21804 17434 21828 17436
rect 21884 17434 21908 17436
rect 21964 17434 21988 17436
rect 22044 17434 22050 17436
rect 21804 17382 21806 17434
rect 21986 17382 21988 17434
rect 21742 17380 21748 17382
rect 21804 17380 21828 17382
rect 21884 17380 21908 17382
rect 21964 17380 21988 17382
rect 22044 17380 22050 17382
rect 21742 17371 22050 17380
rect 22112 17354 22140 19751
rect 22192 19712 22244 19718
rect 22190 19680 22192 19689
rect 22244 19680 22246 19689
rect 22190 19615 22246 19624
rect 22192 18624 22244 18630
rect 22190 18592 22192 18601
rect 22244 18592 22246 18601
rect 22190 18527 22246 18536
rect 22192 17536 22244 17542
rect 22190 17504 22192 17513
rect 22244 17504 22246 17513
rect 22190 17439 22246 17448
rect 22112 17326 22232 17354
rect 21742 16348 22050 16357
rect 21742 16346 21748 16348
rect 21804 16346 21828 16348
rect 21884 16346 21908 16348
rect 21964 16346 21988 16348
rect 22044 16346 22050 16348
rect 21804 16294 21806 16346
rect 21986 16294 21988 16346
rect 21742 16292 21748 16294
rect 21804 16292 21828 16294
rect 21884 16292 21908 16294
rect 21964 16292 21988 16294
rect 22044 16292 22050 16294
rect 21742 16283 22050 16292
rect 21742 15260 22050 15269
rect 21742 15258 21748 15260
rect 21804 15258 21828 15260
rect 21884 15258 21908 15260
rect 21964 15258 21988 15260
rect 22044 15258 22050 15260
rect 21804 15206 21806 15258
rect 21986 15206 21988 15258
rect 22204 15230 22232 17326
rect 21742 15204 21748 15206
rect 21804 15204 21828 15206
rect 21884 15204 21908 15206
rect 21964 15204 21988 15206
rect 22044 15204 22050 15206
rect 21742 15195 22050 15204
rect 22192 15224 22244 15230
rect 22192 15166 22244 15172
rect 22192 14272 22244 14278
rect 22190 14240 22192 14249
rect 22244 14240 22246 14249
rect 21742 14172 22050 14181
rect 22190 14175 22246 14184
rect 21742 14170 21748 14172
rect 21804 14170 21828 14172
rect 21884 14170 21908 14172
rect 21964 14170 21988 14172
rect 22044 14170 22050 14172
rect 21804 14118 21806 14170
rect 21986 14118 21988 14170
rect 21742 14116 21748 14118
rect 21804 14116 21828 14118
rect 21884 14116 21908 14118
rect 21964 14116 21988 14118
rect 22044 14116 22050 14118
rect 21742 14107 22050 14116
rect 21560 13484 21680 13512
rect 21376 13246 21496 13274
rect 21364 13184 21416 13190
rect 21364 13126 21416 13132
rect 21376 12986 21404 13126
rect 21364 12980 21416 12986
rect 21364 12922 21416 12928
rect 21468 11506 21496 13246
rect 21376 11478 21496 11506
rect 21376 11393 21404 11478
rect 21362 11384 21418 11393
rect 21560 11336 21588 13484
rect 22190 13152 22246 13161
rect 21742 13084 22050 13093
rect 22190 13087 22246 13096
rect 21742 13082 21748 13084
rect 21804 13082 21828 13084
rect 21884 13082 21908 13084
rect 21964 13082 21988 13084
rect 22044 13082 22050 13084
rect 21804 13030 21806 13082
rect 21986 13030 21988 13082
rect 21742 13028 21748 13030
rect 21804 13028 21828 13030
rect 21884 13028 21908 13030
rect 21964 13028 21988 13030
rect 22044 13028 22050 13030
rect 21742 13019 22050 13028
rect 22204 12510 22232 13087
rect 22192 12504 22244 12510
rect 22192 12446 22244 12452
rect 22192 12164 22244 12170
rect 22192 12106 22244 12112
rect 22204 12073 22232 12106
rect 22190 12064 22246 12073
rect 21742 11996 22050 12005
rect 22190 11999 22246 12008
rect 21742 11994 21748 11996
rect 21804 11994 21828 11996
rect 21884 11994 21908 11996
rect 21964 11994 21988 11996
rect 22044 11994 22050 11996
rect 21804 11942 21806 11994
rect 21986 11942 21988 11994
rect 21742 11940 21748 11942
rect 21804 11940 21828 11942
rect 21884 11940 21908 11942
rect 21964 11940 21988 11942
rect 22044 11940 22050 11942
rect 21742 11931 22050 11940
rect 21362 11319 21418 11328
rect 21468 11308 21588 11336
rect 21364 11008 21416 11014
rect 21364 10950 21416 10956
rect 21270 10704 21326 10713
rect 21270 10639 21326 10648
rect 20916 10526 21036 10554
rect 20902 10432 20958 10441
rect 20902 10367 20958 10376
rect 20916 10266 20944 10367
rect 20904 10260 20956 10266
rect 20904 10202 20956 10208
rect 21008 9110 21036 10526
rect 21180 9988 21232 9994
rect 21180 9930 21232 9936
rect 21088 9580 21140 9586
rect 21088 9522 21140 9528
rect 20996 9104 21048 9110
rect 20996 9046 21048 9052
rect 20640 8350 20852 8378
rect 20640 3194 20668 8350
rect 21100 8090 21128 9522
rect 21192 8634 21220 9930
rect 21272 9580 21324 9586
rect 21272 9522 21324 9528
rect 21284 9178 21312 9522
rect 21376 9178 21404 10950
rect 21468 9432 21496 11308
rect 22190 10976 22246 10985
rect 21742 10908 22050 10917
rect 22190 10911 22246 10920
rect 21742 10906 21748 10908
rect 21804 10906 21828 10908
rect 21884 10906 21908 10908
rect 21964 10906 21988 10908
rect 22044 10906 22050 10908
rect 21804 10854 21806 10906
rect 21986 10854 21988 10906
rect 21742 10852 21748 10854
rect 21804 10852 21828 10854
rect 21884 10852 21908 10854
rect 21964 10852 21988 10854
rect 22044 10852 22050 10854
rect 21742 10843 22050 10852
rect 22204 10810 22232 10911
rect 22192 10804 22244 10810
rect 22192 10746 22244 10752
rect 21638 10704 21694 10713
rect 21638 10639 21694 10648
rect 21468 9404 21588 9432
rect 21454 9344 21510 9353
rect 21454 9279 21510 9288
rect 21468 9178 21496 9279
rect 21272 9172 21324 9178
rect 21272 9114 21324 9120
rect 21364 9172 21416 9178
rect 21364 9114 21416 9120
rect 21456 9172 21508 9178
rect 21456 9114 21508 9120
rect 21272 8968 21324 8974
rect 21272 8910 21324 8916
rect 21180 8628 21232 8634
rect 21180 8570 21232 8576
rect 21180 8356 21232 8362
rect 21180 8298 21232 8304
rect 21088 8084 21140 8090
rect 21088 8026 21140 8032
rect 20720 7880 20772 7886
rect 20772 7828 21036 7834
rect 20720 7822 21036 7828
rect 20732 7806 21036 7822
rect 20812 7744 20864 7750
rect 20812 7686 20864 7692
rect 20824 6458 20852 7686
rect 20904 6656 20956 6662
rect 20904 6598 20956 6604
rect 20916 6458 20944 6598
rect 20720 6452 20772 6458
rect 20720 6394 20772 6400
rect 20812 6452 20864 6458
rect 20812 6394 20864 6400
rect 20904 6452 20956 6458
rect 20904 6394 20956 6400
rect 20732 5302 20760 6394
rect 21008 6338 21036 7806
rect 21192 6866 21220 8298
rect 21180 6860 21232 6866
rect 21180 6802 21232 6808
rect 21088 6792 21140 6798
rect 21088 6734 21140 6740
rect 21178 6760 21234 6769
rect 20824 6310 21036 6338
rect 20824 5574 20852 6310
rect 20904 6112 20956 6118
rect 20904 6054 20956 6060
rect 20812 5568 20864 5574
rect 20812 5510 20864 5516
rect 20720 5296 20772 5302
rect 20720 5238 20772 5244
rect 20916 5234 20944 6054
rect 21100 5914 21128 6734
rect 21178 6695 21234 6704
rect 21088 5908 21140 5914
rect 21088 5850 21140 5856
rect 20994 5808 21050 5817
rect 20994 5743 20996 5752
rect 21048 5743 21050 5752
rect 20996 5714 21048 5720
rect 21192 5234 21220 6695
rect 21284 6662 21312 8910
rect 21456 7540 21508 7546
rect 21456 7482 21508 7488
rect 21364 7200 21416 7206
rect 21364 7142 21416 7148
rect 21272 6656 21324 6662
rect 21272 6598 21324 6604
rect 21376 5710 21404 7142
rect 21468 6458 21496 7482
rect 21560 7449 21588 9404
rect 21546 7440 21602 7449
rect 21546 7375 21602 7384
rect 21456 6452 21508 6458
rect 21456 6394 21508 6400
rect 21364 5704 21416 5710
rect 21364 5646 21416 5652
rect 20904 5228 20956 5234
rect 20904 5170 20956 5176
rect 21088 5228 21140 5234
rect 21088 5170 21140 5176
rect 21180 5228 21232 5234
rect 21180 5170 21232 5176
rect 21100 4729 21128 5170
rect 21180 4820 21232 4826
rect 21180 4762 21232 4768
rect 21086 4720 21142 4729
rect 21086 4655 21142 4664
rect 21088 4140 21140 4146
rect 21088 4082 21140 4088
rect 20996 3936 21048 3942
rect 20996 3878 21048 3884
rect 20718 3632 20774 3641
rect 20718 3567 20774 3576
rect 20732 3534 20760 3567
rect 20720 3528 20772 3534
rect 20720 3470 20772 3476
rect 20810 3496 20866 3505
rect 20810 3431 20866 3440
rect 20628 3188 20680 3194
rect 20628 3130 20680 3136
rect 20824 3058 20852 3431
rect 20904 3392 20956 3398
rect 20904 3334 20956 3340
rect 20916 3194 20944 3334
rect 20904 3188 20956 3194
rect 20904 3130 20956 3136
rect 21008 3097 21036 3878
rect 20994 3088 21050 3097
rect 20812 3052 20864 3058
rect 20994 3023 21050 3032
rect 20812 2994 20864 3000
rect 20536 2916 20588 2922
rect 20536 2858 20588 2864
rect 21100 2825 21128 4082
rect 21086 2816 21142 2825
rect 21086 2751 21142 2760
rect 21192 2514 21220 4762
rect 21364 4480 21416 4486
rect 21364 4422 21416 4428
rect 21376 4185 21404 4422
rect 21362 4176 21418 4185
rect 21272 4140 21324 4146
rect 21362 4111 21418 4120
rect 21272 4082 21324 4088
rect 21284 3738 21312 4082
rect 21364 3936 21416 3942
rect 21364 3878 21416 3884
rect 21272 3732 21324 3738
rect 21272 3674 21324 3680
rect 21376 3194 21404 3878
rect 21548 3460 21600 3466
rect 21548 3402 21600 3408
rect 21364 3188 21416 3194
rect 21364 3130 21416 3136
rect 21364 2848 21416 2854
rect 21364 2790 21416 2796
rect 21180 2508 21232 2514
rect 21180 2450 21232 2456
rect 21376 2394 21404 2790
rect 21376 2366 21496 2394
rect 20718 2272 20774 2281
rect 20718 2207 20774 2216
rect 20994 2272 21050 2281
rect 20994 2207 21050 2216
rect 21362 2272 21418 2281
rect 21362 2207 21418 2216
rect 20352 2032 20404 2038
rect 20352 1974 20404 1980
rect 20732 1970 20760 2207
rect 21008 2106 21036 2207
rect 21376 2106 21404 2207
rect 20996 2100 21048 2106
rect 20996 2042 21048 2048
rect 21364 2100 21416 2106
rect 21364 2042 21416 2048
rect 21468 2038 21496 2366
rect 21560 2145 21588 3402
rect 21652 2650 21680 10639
rect 22296 10112 22324 24806
rect 22388 22817 22416 31844
rect 22374 22808 22430 22817
rect 22374 22743 22430 22752
rect 22376 22636 22428 22642
rect 22376 22578 22428 22584
rect 22204 10084 22324 10112
rect 21742 9820 22050 9829
rect 21742 9818 21748 9820
rect 21804 9818 21828 9820
rect 21884 9818 21908 9820
rect 21964 9818 21988 9820
rect 22044 9818 22050 9820
rect 21804 9766 21806 9818
rect 21986 9766 21988 9818
rect 21742 9764 21748 9766
rect 21804 9764 21828 9766
rect 21884 9764 21908 9766
rect 21964 9764 21988 9766
rect 22044 9764 22050 9766
rect 21742 9755 22050 9764
rect 21742 8732 22050 8741
rect 21742 8730 21748 8732
rect 21804 8730 21828 8732
rect 21884 8730 21908 8732
rect 21964 8730 21988 8732
rect 22044 8730 22050 8732
rect 21804 8678 21806 8730
rect 21986 8678 21988 8730
rect 21742 8676 21748 8678
rect 21804 8676 21828 8678
rect 21884 8676 21908 8678
rect 21964 8676 21988 8678
rect 22044 8676 22050 8678
rect 21742 8667 22050 8676
rect 22100 8016 22152 8022
rect 22100 7958 22152 7964
rect 21742 7644 22050 7653
rect 21742 7642 21748 7644
rect 21804 7642 21828 7644
rect 21884 7642 21908 7644
rect 21964 7642 21988 7644
rect 22044 7642 22050 7644
rect 21804 7590 21806 7642
rect 21986 7590 21988 7642
rect 21742 7588 21748 7590
rect 21804 7588 21828 7590
rect 21884 7588 21908 7590
rect 21964 7588 21988 7590
rect 22044 7588 22050 7590
rect 21742 7579 22050 7588
rect 21742 6556 22050 6565
rect 21742 6554 21748 6556
rect 21804 6554 21828 6556
rect 21884 6554 21908 6556
rect 21964 6554 21988 6556
rect 22044 6554 22050 6556
rect 21804 6502 21806 6554
rect 21986 6502 21988 6554
rect 21742 6500 21748 6502
rect 21804 6500 21828 6502
rect 21884 6500 21908 6502
rect 21964 6500 21988 6502
rect 22044 6500 22050 6502
rect 21742 6491 22050 6500
rect 21742 5468 22050 5477
rect 21742 5466 21748 5468
rect 21804 5466 21828 5468
rect 21884 5466 21908 5468
rect 21964 5466 21988 5468
rect 22044 5466 22050 5468
rect 21804 5414 21806 5466
rect 21986 5414 21988 5466
rect 21742 5412 21748 5414
rect 21804 5412 21828 5414
rect 21884 5412 21908 5414
rect 21964 5412 21988 5414
rect 22044 5412 22050 5414
rect 21742 5403 22050 5412
rect 21742 4380 22050 4389
rect 21742 4378 21748 4380
rect 21804 4378 21828 4380
rect 21884 4378 21908 4380
rect 21964 4378 21988 4380
rect 22044 4378 22050 4380
rect 21804 4326 21806 4378
rect 21986 4326 21988 4378
rect 21742 4324 21748 4326
rect 21804 4324 21828 4326
rect 21884 4324 21908 4326
rect 21964 4324 21988 4326
rect 22044 4324 22050 4326
rect 21742 4315 22050 4324
rect 21742 3292 22050 3301
rect 21742 3290 21748 3292
rect 21804 3290 21828 3292
rect 21884 3290 21908 3292
rect 21964 3290 21988 3292
rect 22044 3290 22050 3292
rect 21804 3238 21806 3290
rect 21986 3238 21988 3290
rect 21742 3236 21748 3238
rect 21804 3236 21828 3238
rect 21884 3236 21908 3238
rect 21964 3236 21988 3238
rect 22044 3236 22050 3238
rect 21742 3227 22050 3236
rect 21640 2644 21692 2650
rect 21640 2586 21692 2592
rect 21742 2204 22050 2213
rect 21742 2202 21748 2204
rect 21804 2202 21828 2204
rect 21884 2202 21908 2204
rect 21964 2202 21988 2204
rect 22044 2202 22050 2204
rect 21804 2150 21806 2202
rect 21986 2150 21988 2202
rect 21742 2148 21748 2150
rect 21804 2148 21828 2150
rect 21884 2148 21908 2150
rect 21964 2148 21988 2150
rect 22044 2148 22050 2150
rect 21546 2136 21602 2145
rect 21742 2139 22050 2148
rect 21546 2071 21602 2080
rect 21456 2032 21508 2038
rect 21456 1974 21508 1980
rect 20720 1964 20772 1970
rect 20720 1906 20772 1912
rect 22112 1562 22140 7958
rect 22204 2990 22232 10084
rect 22284 9988 22336 9994
rect 22284 9930 22336 9936
rect 22296 9897 22324 9930
rect 22282 9888 22338 9897
rect 22282 9823 22338 9832
rect 22284 9376 22336 9382
rect 22284 9318 22336 9324
rect 22192 2984 22244 2990
rect 22192 2926 22244 2932
rect 22296 2774 22324 9318
rect 22388 5681 22416 22578
rect 22374 5672 22430 5681
rect 22374 5607 22430 5616
rect 22480 3602 22508 39850
rect 22572 31772 22600 41414
rect 22560 31766 22612 31772
rect 22560 31708 22612 31714
rect 22560 30796 22612 30802
rect 22560 30738 22612 30744
rect 22572 18578 22600 30738
rect 22664 30394 22692 41618
rect 22836 35624 22888 35630
rect 22836 35566 22888 35572
rect 22928 35624 22980 35630
rect 22928 35566 22980 35572
rect 22742 34096 22798 34105
rect 22742 34031 22798 34040
rect 22756 32366 22784 34031
rect 22848 32978 22876 35566
rect 22836 32972 22888 32978
rect 22836 32914 22888 32920
rect 22836 32836 22888 32842
rect 22836 32778 22888 32784
rect 22744 32360 22796 32366
rect 22744 32302 22796 32308
rect 22848 32298 22876 32778
rect 22836 32292 22888 32298
rect 22836 32234 22888 32240
rect 22940 32178 22968 35566
rect 22756 32150 22968 32178
rect 22652 30388 22704 30394
rect 22652 30330 22704 30336
rect 22652 26784 22704 26790
rect 22652 26726 22704 26732
rect 22664 22094 22692 26726
rect 22756 22710 22784 32150
rect 22836 32088 22888 32094
rect 22836 32030 22888 32036
rect 22744 22704 22796 22710
rect 22744 22646 22796 22652
rect 22664 22066 22784 22094
rect 22650 21992 22706 22001
rect 22650 21927 22706 21936
rect 22664 21010 22692 21927
rect 22652 21004 22704 21010
rect 22652 20946 22704 20952
rect 22650 20904 22706 20913
rect 22650 20839 22706 20848
rect 22664 18698 22692 20839
rect 22756 18766 22784 22066
rect 22744 18760 22796 18766
rect 22744 18702 22796 18708
rect 22652 18692 22704 18698
rect 22652 18634 22704 18640
rect 22572 18550 22784 18578
rect 22652 18488 22704 18494
rect 22652 18430 22704 18436
rect 22560 15428 22612 15434
rect 22560 15370 22612 15376
rect 22572 15337 22600 15370
rect 22558 15328 22614 15337
rect 22558 15263 22614 15272
rect 22560 15224 22612 15230
rect 22560 15166 22612 15172
rect 22468 3596 22520 3602
rect 22468 3538 22520 3544
rect 22572 3398 22600 15166
rect 22664 3738 22692 18430
rect 22756 15026 22784 18550
rect 22744 15020 22796 15026
rect 22744 14962 22796 14968
rect 22744 14884 22796 14890
rect 22744 14826 22796 14832
rect 22652 3732 22704 3738
rect 22652 3674 22704 3680
rect 22560 3392 22612 3398
rect 22560 3334 22612 3340
rect 22204 2746 22324 2774
rect 22100 1556 22152 1562
rect 22100 1498 22152 1504
rect 22204 1290 22232 2746
rect 22756 1358 22784 14826
rect 22848 12238 22876 32030
rect 22928 31816 22980 31822
rect 22928 31758 22980 31764
rect 22940 22234 22968 31758
rect 22928 22228 22980 22234
rect 22928 22170 22980 22176
rect 22928 20664 22980 20670
rect 22928 20606 22980 20612
rect 22836 12232 22888 12238
rect 22836 12174 22888 12180
rect 22834 11792 22890 11801
rect 22834 11727 22890 11736
rect 22848 1902 22876 11727
rect 22836 1896 22888 1902
rect 22836 1838 22888 1844
rect 22744 1352 22796 1358
rect 22744 1294 22796 1300
rect 22192 1284 22244 1290
rect 22192 1226 22244 1232
rect 21742 1116 22050 1125
rect 21742 1114 21748 1116
rect 21804 1114 21828 1116
rect 21884 1114 21908 1116
rect 21964 1114 21988 1116
rect 22044 1114 22050 1116
rect 21804 1062 21806 1114
rect 21986 1062 21988 1114
rect 21742 1060 21748 1062
rect 21804 1060 21828 1062
rect 21884 1060 21908 1062
rect 21964 1060 21988 1062
rect 22044 1060 22050 1062
rect 21742 1051 22050 1060
rect 22940 1018 22968 20606
rect 22928 1012 22980 1018
rect 22928 954 22980 960
rect 19890 54 20300 82
rect 19338 -300 19394 54
rect 19522 -300 19578 54
rect 19706 -300 19762 54
rect 19890 -300 19946 54
<< via2 >>
rect 2226 43832 2282 43888
rect 18 41384 74 41440
rect 294 35672 350 35728
rect 938 42200 994 42256
rect 478 35536 534 35592
rect 294 29552 350 29608
rect 294 29008 350 29064
rect 478 17584 534 17640
rect 846 42064 902 42120
rect 754 37848 810 37904
rect 754 31864 810 31920
rect 754 29960 810 30016
rect 754 28872 810 28928
rect 754 27784 810 27840
rect 662 27376 718 27432
rect 846 26152 902 26208
rect 846 24812 902 24848
rect 846 24792 848 24812
rect 848 24792 900 24812
rect 900 24792 902 24812
rect 754 23704 810 23760
rect 662 21936 718 21992
rect 754 21528 810 21584
rect 754 21004 810 21040
rect 754 20984 756 21004
rect 756 20984 808 21004
rect 808 20984 810 21004
rect 754 19896 810 19952
rect 662 14592 718 14648
rect 754 1400 810 1456
rect 1122 38664 1178 38720
rect 1398 39752 1454 39808
rect 1306 38936 1362 38992
rect 1306 37576 1362 37632
rect 1214 36896 1270 36952
rect 2226 41540 2282 41576
rect 2226 41520 2228 41540
rect 2228 41520 2280 41540
rect 2280 41520 2282 41540
rect 2134 40976 2190 41032
rect 1674 40024 1730 40080
rect 1214 34992 1270 35048
rect 1490 34992 1546 35048
rect 1490 33224 1546 33280
rect 2042 38528 2098 38584
rect 1950 37168 2006 37224
rect 1766 36080 1822 36136
rect 1674 35264 1730 35320
rect 1674 33904 1730 33960
rect 3882 43832 3938 43888
rect 3555 43002 3611 43004
rect 3635 43002 3691 43004
rect 3715 43002 3771 43004
rect 3795 43002 3851 43004
rect 3555 42950 3601 43002
rect 3601 42950 3611 43002
rect 3635 42950 3665 43002
rect 3665 42950 3677 43002
rect 3677 42950 3691 43002
rect 3715 42950 3729 43002
rect 3729 42950 3741 43002
rect 3741 42950 3771 43002
rect 3795 42950 3805 43002
rect 3805 42950 3851 43002
rect 3555 42948 3611 42950
rect 3635 42948 3691 42950
rect 3715 42948 3771 42950
rect 3795 42948 3851 42950
rect 2410 39752 2466 39808
rect 2502 39616 2558 39672
rect 2410 37848 2466 37904
rect 2778 39480 2834 39536
rect 2410 37732 2466 37768
rect 2410 37712 2412 37732
rect 2412 37712 2464 37732
rect 2464 37712 2466 37732
rect 2410 36896 2466 36952
rect 2686 38664 2742 38720
rect 2962 39208 3018 39264
rect 2962 38392 3018 38448
rect 2870 38256 2926 38312
rect 2778 37304 2834 37360
rect 3555 41914 3611 41916
rect 3635 41914 3691 41916
rect 3715 41914 3771 41916
rect 3795 41914 3851 41916
rect 3555 41862 3601 41914
rect 3601 41862 3611 41914
rect 3635 41862 3665 41914
rect 3665 41862 3677 41914
rect 3677 41862 3691 41914
rect 3715 41862 3729 41914
rect 3729 41862 3741 41914
rect 3741 41862 3771 41914
rect 3795 41862 3805 41914
rect 3805 41862 3851 41914
rect 3555 41860 3611 41862
rect 3635 41860 3691 41862
rect 3715 41860 3771 41862
rect 3795 41860 3851 41862
rect 4342 42880 4398 42936
rect 4250 41656 4306 41712
rect 3606 41384 3662 41440
rect 3555 40826 3611 40828
rect 3635 40826 3691 40828
rect 3715 40826 3771 40828
rect 3795 40826 3851 40828
rect 3555 40774 3601 40826
rect 3601 40774 3611 40826
rect 3635 40774 3665 40826
rect 3665 40774 3677 40826
rect 3677 40774 3691 40826
rect 3715 40774 3729 40826
rect 3729 40774 3741 40826
rect 3741 40774 3771 40826
rect 3795 40774 3805 40826
rect 3805 40774 3851 40826
rect 3555 40772 3611 40774
rect 3635 40772 3691 40774
rect 3715 40772 3771 40774
rect 3795 40772 3851 40774
rect 4526 41556 4528 41576
rect 4528 41556 4580 41576
rect 4580 41556 4582 41576
rect 4526 41520 4582 41556
rect 3974 40432 4030 40488
rect 2870 36216 2926 36272
rect 1858 33632 1914 33688
rect 1490 31592 1546 31648
rect 1490 31184 1546 31240
rect 1398 30368 1454 30424
rect 1490 29824 1546 29880
rect 1490 29144 1546 29200
rect 1858 32408 1914 32464
rect 1766 32272 1822 32328
rect 1858 32136 1914 32192
rect 1950 31864 2006 31920
rect 1858 31764 1860 31784
rect 1860 31764 1912 31784
rect 1912 31764 1914 31784
rect 1674 30504 1730 30560
rect 1858 31728 1914 31764
rect 2226 32408 2282 32464
rect 2134 31728 2190 31784
rect 1674 29144 1730 29200
rect 1950 29280 2006 29336
rect 1398 28328 1454 28384
rect 1214 27648 1270 27704
rect 1306 27240 1362 27296
rect 1306 27004 1308 27024
rect 1308 27004 1360 27024
rect 1360 27004 1362 27024
rect 1306 26968 1362 27004
rect 1490 27512 1546 27568
rect 1674 27940 1730 27976
rect 1674 27920 1676 27940
rect 1676 27920 1728 27940
rect 1728 27920 1730 27940
rect 1398 26832 1454 26888
rect 1214 26696 1270 26752
rect 1490 25064 1546 25120
rect 1490 24928 1546 24984
rect 1398 24384 1454 24440
rect 1858 27104 1914 27160
rect 1858 26560 1914 26616
rect 1766 26424 1822 26480
rect 1766 26288 1822 26344
rect 3054 35128 3110 35184
rect 3054 34992 3110 35048
rect 2594 31864 2650 31920
rect 2962 32680 3018 32736
rect 2962 32272 3018 32328
rect 2410 31184 2466 31240
rect 2594 31184 2650 31240
rect 2686 31048 2742 31104
rect 2594 30640 2650 30696
rect 2502 30096 2558 30152
rect 2870 30676 2872 30696
rect 2872 30676 2924 30696
rect 2924 30676 2926 30696
rect 2870 30640 2926 30676
rect 2778 29688 2834 29744
rect 2226 29280 2282 29336
rect 2410 28328 2466 28384
rect 3555 39738 3611 39740
rect 3635 39738 3691 39740
rect 3715 39738 3771 39740
rect 3795 39738 3851 39740
rect 3555 39686 3601 39738
rect 3601 39686 3611 39738
rect 3635 39686 3665 39738
rect 3665 39686 3677 39738
rect 3677 39686 3691 39738
rect 3715 39686 3729 39738
rect 3729 39686 3741 39738
rect 3741 39686 3771 39738
rect 3795 39686 3805 39738
rect 3805 39686 3851 39738
rect 3555 39684 3611 39686
rect 3635 39684 3691 39686
rect 3715 39684 3771 39686
rect 3795 39684 3851 39686
rect 3555 38650 3611 38652
rect 3635 38650 3691 38652
rect 3715 38650 3771 38652
rect 3795 38650 3851 38652
rect 3555 38598 3601 38650
rect 3601 38598 3611 38650
rect 3635 38598 3665 38650
rect 3665 38598 3677 38650
rect 3677 38598 3691 38650
rect 3715 38598 3729 38650
rect 3729 38598 3741 38650
rect 3741 38598 3771 38650
rect 3795 38598 3805 38650
rect 3805 38598 3851 38650
rect 3555 38596 3611 38598
rect 3635 38596 3691 38598
rect 3715 38596 3771 38598
rect 3795 38596 3851 38598
rect 4250 38528 4306 38584
rect 3422 37848 3478 37904
rect 3555 37562 3611 37564
rect 3635 37562 3691 37564
rect 3715 37562 3771 37564
rect 3795 37562 3851 37564
rect 3555 37510 3601 37562
rect 3601 37510 3611 37562
rect 3635 37510 3665 37562
rect 3665 37510 3677 37562
rect 3677 37510 3691 37562
rect 3715 37510 3729 37562
rect 3729 37510 3741 37562
rect 3741 37510 3771 37562
rect 3795 37510 3805 37562
rect 3805 37510 3851 37562
rect 3555 37508 3611 37510
rect 3635 37508 3691 37510
rect 3715 37508 3771 37510
rect 3795 37508 3851 37510
rect 3974 37712 4030 37768
rect 3238 34856 3294 34912
rect 3555 36474 3611 36476
rect 3635 36474 3691 36476
rect 3715 36474 3771 36476
rect 3795 36474 3851 36476
rect 3555 36422 3601 36474
rect 3601 36422 3611 36474
rect 3635 36422 3665 36474
rect 3665 36422 3677 36474
rect 3677 36422 3691 36474
rect 3715 36422 3729 36474
rect 3729 36422 3741 36474
rect 3741 36422 3771 36474
rect 3795 36422 3805 36474
rect 3805 36422 3851 36474
rect 3555 36420 3611 36422
rect 3635 36420 3691 36422
rect 3715 36420 3771 36422
rect 3795 36420 3851 36422
rect 3514 35536 3570 35592
rect 3555 35386 3611 35388
rect 3635 35386 3691 35388
rect 3715 35386 3771 35388
rect 3795 35386 3851 35388
rect 3555 35334 3601 35386
rect 3601 35334 3611 35386
rect 3635 35334 3665 35386
rect 3665 35334 3677 35386
rect 3677 35334 3691 35386
rect 3715 35334 3729 35386
rect 3729 35334 3741 35386
rect 3741 35334 3771 35386
rect 3795 35334 3805 35386
rect 3805 35334 3851 35386
rect 3555 35332 3611 35334
rect 3635 35332 3691 35334
rect 3715 35332 3771 35334
rect 3795 35332 3851 35334
rect 3422 35264 3478 35320
rect 3514 35128 3570 35184
rect 3514 34992 3570 35048
rect 3146 33768 3202 33824
rect 3330 32952 3386 33008
rect 3238 32816 3294 32872
rect 3238 31456 3294 31512
rect 3790 34584 3846 34640
rect 3555 34298 3611 34300
rect 3635 34298 3691 34300
rect 3715 34298 3771 34300
rect 3795 34298 3851 34300
rect 3555 34246 3601 34298
rect 3601 34246 3611 34298
rect 3635 34246 3665 34298
rect 3665 34246 3677 34298
rect 3677 34246 3691 34298
rect 3715 34246 3729 34298
rect 3729 34246 3741 34298
rect 3741 34246 3771 34298
rect 3795 34246 3805 34298
rect 3805 34246 3851 34298
rect 3555 34244 3611 34246
rect 3635 34244 3691 34246
rect 3715 34244 3771 34246
rect 3795 34244 3851 34246
rect 4250 35808 4306 35864
rect 4066 35128 4122 35184
rect 4250 34584 4306 34640
rect 4066 34040 4122 34096
rect 3882 33632 3938 33688
rect 3555 33210 3611 33212
rect 3635 33210 3691 33212
rect 3715 33210 3771 33212
rect 3795 33210 3851 33212
rect 3555 33158 3601 33210
rect 3601 33158 3611 33210
rect 3635 33158 3665 33210
rect 3665 33158 3677 33210
rect 3677 33158 3691 33210
rect 3715 33158 3729 33210
rect 3729 33158 3741 33210
rect 3741 33158 3771 33210
rect 3795 33158 3805 33210
rect 3805 33158 3851 33210
rect 3555 33156 3611 33158
rect 3635 33156 3691 33158
rect 3715 33156 3771 33158
rect 3795 33156 3851 33158
rect 3790 32952 3846 33008
rect 3555 32122 3611 32124
rect 3635 32122 3691 32124
rect 3715 32122 3771 32124
rect 3795 32122 3851 32124
rect 3555 32070 3601 32122
rect 3601 32070 3611 32122
rect 3635 32070 3665 32122
rect 3665 32070 3677 32122
rect 3677 32070 3691 32122
rect 3715 32070 3729 32122
rect 3729 32070 3741 32122
rect 3741 32070 3771 32122
rect 3795 32070 3805 32122
rect 3805 32070 3851 32122
rect 3555 32068 3611 32070
rect 3635 32068 3691 32070
rect 3715 32068 3771 32070
rect 3795 32068 3851 32070
rect 3698 31456 3754 31512
rect 3790 31320 3846 31376
rect 3555 31034 3611 31036
rect 3635 31034 3691 31036
rect 3715 31034 3771 31036
rect 3795 31034 3851 31036
rect 3555 30982 3601 31034
rect 3601 30982 3611 31034
rect 3635 30982 3665 31034
rect 3665 30982 3677 31034
rect 3677 30982 3691 31034
rect 3715 30982 3729 31034
rect 3729 30982 3741 31034
rect 3741 30982 3771 31034
rect 3795 30982 3805 31034
rect 3805 30982 3851 31034
rect 3555 30980 3611 30982
rect 3635 30980 3691 30982
rect 3715 30980 3771 30982
rect 3795 30980 3851 30982
rect 4066 32408 4122 32464
rect 4066 31764 4068 31784
rect 4068 31764 4120 31784
rect 4120 31764 4122 31784
rect 4066 31728 4122 31764
rect 4250 32000 4306 32056
rect 4066 30776 4122 30832
rect 4250 31456 4306 31512
rect 3238 29824 3294 29880
rect 3054 29144 3110 29200
rect 2594 28192 2650 28248
rect 2042 26424 2098 26480
rect 1950 26152 2006 26208
rect 2134 26016 2190 26072
rect 1858 24656 1914 24712
rect 1582 23976 1638 24032
rect 1398 23432 1454 23488
rect 1582 23024 1638 23080
rect 1306 22888 1362 22944
rect 1674 22772 1730 22808
rect 1674 22752 1676 22772
rect 1676 22752 1728 22772
rect 1728 22752 1730 22772
rect 1122 22616 1178 22672
rect 1122 22480 1178 22536
rect 938 18536 994 18592
rect 938 14728 994 14784
rect 938 13776 994 13832
rect 938 12960 994 13016
rect 1030 11464 1086 11520
rect 1030 10240 1086 10296
rect 1030 7248 1086 7304
rect 938 3576 994 3632
rect 1398 22092 1454 22128
rect 1398 22072 1400 22092
rect 1400 22072 1452 22092
rect 1452 22072 1454 22092
rect 1214 21800 1270 21856
rect 1674 21664 1730 21720
rect 1490 21256 1546 21312
rect 1306 20712 1362 20768
rect 1306 17312 1362 17368
rect 1582 20324 1638 20360
rect 1582 20304 1584 20324
rect 1584 20304 1636 20324
rect 1636 20304 1638 20324
rect 1490 20168 1546 20224
rect 1766 21392 1822 21448
rect 2686 27124 2742 27160
rect 2686 27104 2688 27124
rect 2688 27104 2740 27124
rect 2740 27104 2742 27124
rect 2502 26852 2558 26888
rect 2962 28056 3018 28112
rect 2502 26832 2504 26852
rect 2504 26832 2556 26852
rect 2556 26832 2558 26852
rect 2502 26460 2504 26480
rect 2504 26460 2556 26480
rect 2556 26460 2558 26480
rect 2502 26424 2558 26460
rect 2226 25472 2282 25528
rect 2134 25064 2190 25120
rect 2042 21800 2098 21856
rect 1950 21256 2006 21312
rect 1674 18828 1730 18864
rect 1674 18808 1676 18828
rect 1676 18808 1728 18828
rect 1728 18808 1730 18828
rect 1674 18536 1730 18592
rect 1490 17992 1546 18048
rect 1582 17856 1638 17912
rect 2502 24928 2558 24984
rect 2226 22616 2282 22672
rect 2410 22752 2466 22808
rect 2318 22344 2374 22400
rect 2778 25336 2834 25392
rect 2962 26988 3018 27024
rect 2962 26968 2964 26988
rect 2964 26968 3016 26988
rect 3016 26968 3018 26988
rect 2962 26696 3018 26752
rect 3146 28056 3202 28112
rect 3146 27276 3148 27296
rect 3148 27276 3200 27296
rect 3200 27276 3202 27296
rect 3146 27240 3202 27276
rect 3330 26560 3386 26616
rect 3606 30252 3662 30288
rect 3606 30232 3608 30252
rect 3608 30232 3660 30252
rect 3660 30232 3662 30252
rect 3882 30268 3884 30288
rect 3884 30268 3936 30288
rect 3936 30268 3938 30288
rect 3882 30232 3938 30268
rect 3555 29946 3611 29948
rect 3635 29946 3691 29948
rect 3715 29946 3771 29948
rect 3795 29946 3851 29948
rect 3555 29894 3601 29946
rect 3601 29894 3611 29946
rect 3635 29894 3665 29946
rect 3665 29894 3677 29946
rect 3677 29894 3691 29946
rect 3715 29894 3729 29946
rect 3729 29894 3741 29946
rect 3741 29894 3771 29946
rect 3795 29894 3805 29946
rect 3805 29894 3851 29946
rect 3555 29892 3611 29894
rect 3635 29892 3691 29894
rect 3715 29892 3771 29894
rect 3795 29892 3851 29894
rect 3514 29416 3570 29472
rect 3555 28858 3611 28860
rect 3635 28858 3691 28860
rect 3715 28858 3771 28860
rect 3795 28858 3851 28860
rect 3555 28806 3601 28858
rect 3601 28806 3611 28858
rect 3635 28806 3665 28858
rect 3665 28806 3677 28858
rect 3677 28806 3691 28858
rect 3715 28806 3729 28858
rect 3729 28806 3741 28858
rect 3741 28806 3771 28858
rect 3795 28806 3805 28858
rect 3805 28806 3851 28858
rect 3555 28804 3611 28806
rect 3635 28804 3691 28806
rect 3715 28804 3771 28806
rect 3795 28804 3851 28806
rect 3790 28600 3846 28656
rect 3606 28328 3662 28384
rect 4250 29960 4306 30016
rect 3555 27770 3611 27772
rect 3635 27770 3691 27772
rect 3715 27770 3771 27772
rect 3795 27770 3851 27772
rect 3555 27718 3601 27770
rect 3601 27718 3611 27770
rect 3635 27718 3665 27770
rect 3665 27718 3677 27770
rect 3677 27718 3691 27770
rect 3715 27718 3729 27770
rect 3729 27718 3741 27770
rect 3741 27718 3771 27770
rect 3795 27718 3805 27770
rect 3805 27718 3851 27770
rect 3555 27716 3611 27718
rect 3635 27716 3691 27718
rect 3715 27716 3771 27718
rect 3795 27716 3851 27718
rect 4158 28600 4214 28656
rect 4250 27920 4306 27976
rect 4066 27240 4122 27296
rect 4066 27104 4122 27160
rect 3555 26682 3611 26684
rect 3635 26682 3691 26684
rect 3715 26682 3771 26684
rect 3795 26682 3851 26684
rect 3555 26630 3601 26682
rect 3601 26630 3611 26682
rect 3635 26630 3665 26682
rect 3665 26630 3677 26682
rect 3677 26630 3691 26682
rect 3715 26630 3729 26682
rect 3729 26630 3741 26682
rect 3741 26630 3771 26682
rect 3795 26630 3805 26682
rect 3805 26630 3851 26682
rect 3555 26628 3611 26630
rect 3635 26628 3691 26630
rect 3715 26628 3771 26630
rect 3795 26628 3851 26630
rect 3330 26460 3332 26480
rect 3332 26460 3384 26480
rect 3384 26460 3386 26480
rect 3054 25608 3110 25664
rect 2778 23160 2834 23216
rect 2962 23432 3018 23488
rect 2594 22072 2650 22128
rect 2410 21120 2466 21176
rect 1950 19624 2006 19680
rect 2318 20596 2374 20632
rect 2318 20576 2320 20596
rect 2320 20576 2372 20596
rect 2372 20576 2374 20596
rect 2318 19916 2374 19952
rect 2318 19896 2320 19916
rect 2320 19896 2372 19916
rect 2372 19896 2374 19916
rect 2318 19780 2374 19816
rect 2318 19760 2320 19780
rect 2320 19760 2372 19780
rect 2372 19760 2374 19780
rect 2686 21120 2742 21176
rect 2594 20576 2650 20632
rect 2594 19760 2650 19816
rect 3054 21256 3110 21312
rect 3330 26424 3386 26460
rect 3514 26288 3570 26344
rect 3330 26152 3386 26208
rect 4618 34584 4674 34640
rect 4618 33496 4674 33552
rect 4342 27104 4398 27160
rect 3555 25594 3611 25596
rect 3635 25594 3691 25596
rect 3715 25594 3771 25596
rect 3795 25594 3851 25596
rect 3555 25542 3601 25594
rect 3601 25542 3611 25594
rect 3635 25542 3665 25594
rect 3665 25542 3677 25594
rect 3677 25542 3691 25594
rect 3715 25542 3729 25594
rect 3729 25542 3741 25594
rect 3741 25542 3771 25594
rect 3795 25542 3805 25594
rect 3805 25542 3851 25594
rect 3555 25540 3611 25542
rect 3635 25540 3691 25542
rect 3715 25540 3771 25542
rect 3795 25540 3851 25542
rect 3606 25336 3662 25392
rect 3238 24520 3294 24576
rect 3555 24506 3611 24508
rect 3635 24506 3691 24508
rect 3715 24506 3771 24508
rect 3795 24506 3851 24508
rect 3555 24454 3601 24506
rect 3601 24454 3611 24506
rect 3635 24454 3665 24506
rect 3665 24454 3677 24506
rect 3677 24454 3691 24506
rect 3715 24454 3729 24506
rect 3729 24454 3741 24506
rect 3741 24454 3771 24506
rect 3795 24454 3805 24506
rect 3805 24454 3851 24506
rect 3555 24452 3611 24454
rect 3635 24452 3691 24454
rect 3715 24452 3771 24454
rect 3795 24452 3851 24454
rect 3974 23704 4030 23760
rect 3555 23418 3611 23420
rect 3635 23418 3691 23420
rect 3715 23418 3771 23420
rect 3795 23418 3851 23420
rect 3555 23366 3601 23418
rect 3601 23366 3611 23418
rect 3635 23366 3665 23418
rect 3665 23366 3677 23418
rect 3677 23366 3691 23418
rect 3715 23366 3729 23418
rect 3729 23366 3741 23418
rect 3741 23366 3771 23418
rect 3795 23366 3805 23418
rect 3805 23366 3851 23418
rect 3555 23364 3611 23366
rect 3635 23364 3691 23366
rect 3715 23364 3771 23366
rect 3795 23364 3851 23366
rect 3606 23160 3662 23216
rect 3974 23604 3976 23624
rect 3976 23604 4028 23624
rect 4028 23604 4030 23624
rect 3974 23568 4030 23604
rect 3974 23432 4030 23488
rect 5354 42064 5410 42120
rect 6154 43546 6210 43548
rect 6234 43546 6290 43548
rect 6314 43546 6370 43548
rect 6394 43546 6450 43548
rect 6154 43494 6200 43546
rect 6200 43494 6210 43546
rect 6234 43494 6264 43546
rect 6264 43494 6276 43546
rect 6276 43494 6290 43546
rect 6314 43494 6328 43546
rect 6328 43494 6340 43546
rect 6340 43494 6370 43546
rect 6394 43494 6404 43546
rect 6404 43494 6450 43546
rect 6154 43492 6210 43494
rect 6234 43492 6290 43494
rect 6314 43492 6370 43494
rect 6394 43492 6450 43494
rect 5262 40160 5318 40216
rect 4894 37576 4950 37632
rect 4894 35572 4896 35592
rect 4896 35572 4948 35592
rect 4948 35572 4950 35592
rect 4894 35536 4950 35572
rect 4802 33224 4858 33280
rect 5354 37712 5410 37768
rect 5446 37576 5502 37632
rect 5262 36488 5318 36544
rect 5262 35264 5318 35320
rect 5446 36080 5502 36136
rect 6154 42458 6210 42460
rect 6234 42458 6290 42460
rect 6314 42458 6370 42460
rect 6394 42458 6450 42460
rect 6154 42406 6200 42458
rect 6200 42406 6210 42458
rect 6234 42406 6264 42458
rect 6264 42406 6276 42458
rect 6276 42406 6290 42458
rect 6314 42406 6328 42458
rect 6328 42406 6340 42458
rect 6340 42406 6370 42458
rect 6394 42406 6404 42458
rect 6404 42406 6450 42458
rect 6154 42404 6210 42406
rect 6234 42404 6290 42406
rect 6314 42404 6370 42406
rect 6394 42404 6450 42406
rect 6458 42200 6514 42256
rect 6154 41370 6210 41372
rect 6234 41370 6290 41372
rect 6314 41370 6370 41372
rect 6394 41370 6450 41372
rect 6154 41318 6200 41370
rect 6200 41318 6210 41370
rect 6234 41318 6264 41370
rect 6264 41318 6276 41370
rect 6276 41318 6290 41370
rect 6314 41318 6328 41370
rect 6328 41318 6340 41370
rect 6340 41318 6370 41370
rect 6394 41318 6404 41370
rect 6404 41318 6450 41370
rect 6154 41316 6210 41318
rect 6234 41316 6290 41318
rect 6314 41316 6370 41318
rect 6394 41316 6450 41318
rect 7378 41556 7380 41576
rect 7380 41556 7432 41576
rect 7432 41556 7434 41576
rect 7378 41520 7434 41556
rect 7286 41248 7342 41304
rect 7286 41132 7342 41168
rect 7562 41384 7618 41440
rect 7286 41112 7288 41132
rect 7288 41112 7340 41132
rect 7340 41112 7342 41132
rect 6550 40568 6606 40624
rect 7010 40432 7066 40488
rect 6154 40282 6210 40284
rect 6234 40282 6290 40284
rect 6314 40282 6370 40284
rect 6394 40282 6450 40284
rect 6154 40230 6200 40282
rect 6200 40230 6210 40282
rect 6234 40230 6264 40282
rect 6264 40230 6276 40282
rect 6276 40230 6290 40282
rect 6314 40230 6328 40282
rect 6328 40230 6340 40282
rect 6340 40230 6370 40282
rect 6394 40230 6404 40282
rect 6404 40230 6450 40282
rect 6154 40228 6210 40230
rect 6234 40228 6290 40230
rect 6314 40228 6370 40230
rect 6394 40228 6450 40230
rect 5998 39888 6054 39944
rect 6154 39194 6210 39196
rect 6234 39194 6290 39196
rect 6314 39194 6370 39196
rect 6394 39194 6450 39196
rect 6154 39142 6200 39194
rect 6200 39142 6210 39194
rect 6234 39142 6264 39194
rect 6264 39142 6276 39194
rect 6276 39142 6290 39194
rect 6314 39142 6328 39194
rect 6328 39142 6340 39194
rect 6340 39142 6370 39194
rect 6394 39142 6404 39194
rect 6404 39142 6450 39194
rect 6154 39140 6210 39142
rect 6234 39140 6290 39142
rect 6314 39140 6370 39142
rect 6394 39140 6450 39142
rect 5538 34040 5594 34096
rect 5814 35536 5870 35592
rect 4710 32136 4766 32192
rect 4618 29280 4674 29336
rect 4618 28872 4674 28928
rect 4250 24520 4306 24576
rect 4250 24404 4306 24440
rect 4250 24384 4252 24404
rect 4252 24384 4304 24404
rect 4304 24384 4306 24404
rect 2870 20848 2926 20904
rect 2778 19488 2834 19544
rect 2410 19216 2466 19272
rect 1858 18264 1914 18320
rect 1858 17856 1914 17912
rect 1582 15816 1638 15872
rect 1490 15680 1546 15736
rect 1398 15136 1454 15192
rect 1398 13796 1454 13832
rect 1398 13776 1400 13796
rect 1400 13776 1452 13796
rect 1452 13776 1454 13796
rect 1950 17176 2006 17232
rect 1766 16904 1822 16960
rect 2134 17620 2136 17640
rect 2136 17620 2188 17640
rect 2188 17620 2190 17640
rect 2134 17584 2190 17620
rect 1858 14456 1914 14512
rect 1674 14184 1730 14240
rect 1490 12164 1546 12200
rect 1490 12144 1492 12164
rect 1492 12144 1544 12164
rect 1544 12144 1546 12164
rect 1582 11892 1638 11928
rect 1582 11872 1584 11892
rect 1584 11872 1636 11892
rect 1636 11872 1638 11892
rect 1582 11736 1638 11792
rect 1490 11600 1546 11656
rect 1766 13932 1822 13968
rect 1766 13912 1768 13932
rect 1768 13912 1820 13932
rect 1820 13912 1822 13932
rect 1766 13504 1822 13560
rect 2502 18128 2558 18184
rect 2318 16768 2374 16824
rect 2870 19080 2926 19136
rect 3146 20712 3202 20768
rect 3555 22330 3611 22332
rect 3635 22330 3691 22332
rect 3715 22330 3771 22332
rect 3795 22330 3851 22332
rect 3555 22278 3601 22330
rect 3601 22278 3611 22330
rect 3635 22278 3665 22330
rect 3665 22278 3677 22330
rect 3677 22278 3691 22330
rect 3715 22278 3729 22330
rect 3729 22278 3741 22330
rect 3741 22278 3771 22330
rect 3795 22278 3805 22330
rect 3805 22278 3851 22330
rect 3555 22276 3611 22278
rect 3635 22276 3691 22278
rect 3715 22276 3771 22278
rect 3795 22276 3851 22278
rect 3555 21242 3611 21244
rect 3635 21242 3691 21244
rect 3715 21242 3771 21244
rect 3795 21242 3851 21244
rect 3555 21190 3601 21242
rect 3601 21190 3611 21242
rect 3635 21190 3665 21242
rect 3665 21190 3677 21242
rect 3677 21190 3691 21242
rect 3715 21190 3729 21242
rect 3729 21190 3741 21242
rect 3741 21190 3771 21242
rect 3795 21190 3805 21242
rect 3805 21190 3851 21242
rect 3555 21188 3611 21190
rect 3635 21188 3691 21190
rect 3715 21188 3771 21190
rect 3795 21188 3851 21190
rect 3238 20440 3294 20496
rect 3238 19916 3294 19952
rect 3238 19896 3240 19916
rect 3240 19896 3292 19916
rect 3292 19896 3294 19916
rect 3330 19488 3386 19544
rect 3238 19352 3294 19408
rect 2778 17992 2834 18048
rect 2686 17856 2742 17912
rect 2778 17720 2834 17776
rect 3555 20154 3611 20156
rect 3635 20154 3691 20156
rect 3715 20154 3771 20156
rect 3795 20154 3851 20156
rect 3555 20102 3601 20154
rect 3601 20102 3611 20154
rect 3635 20102 3665 20154
rect 3665 20102 3677 20154
rect 3677 20102 3691 20154
rect 3715 20102 3729 20154
rect 3729 20102 3741 20154
rect 3741 20102 3771 20154
rect 3795 20102 3805 20154
rect 3805 20102 3851 20154
rect 3555 20100 3611 20102
rect 3635 20100 3691 20102
rect 3715 20100 3771 20102
rect 3795 20100 3851 20102
rect 3555 19066 3611 19068
rect 3635 19066 3691 19068
rect 3715 19066 3771 19068
rect 3795 19066 3851 19068
rect 3555 19014 3601 19066
rect 3601 19014 3611 19066
rect 3635 19014 3665 19066
rect 3665 19014 3677 19066
rect 3677 19014 3691 19066
rect 3715 19014 3729 19066
rect 3729 19014 3741 19066
rect 3741 19014 3771 19066
rect 3795 19014 3805 19066
rect 3805 19014 3851 19066
rect 3555 19012 3611 19014
rect 3635 19012 3691 19014
rect 3715 19012 3771 19014
rect 3795 19012 3851 19014
rect 4342 24132 4398 24168
rect 4342 24112 4344 24132
rect 4344 24112 4396 24132
rect 4396 24112 4398 24132
rect 4526 25764 4582 25800
rect 4526 25744 4528 25764
rect 4528 25744 4580 25764
rect 4580 25744 4582 25764
rect 4526 25608 4582 25664
rect 4250 23160 4306 23216
rect 4342 22208 4398 22264
rect 4250 21664 4306 21720
rect 5078 32952 5134 33008
rect 4894 27920 4950 27976
rect 4894 27240 4950 27296
rect 5170 32020 5226 32056
rect 5170 32000 5172 32020
rect 5172 32000 5224 32020
rect 5224 32000 5226 32020
rect 5262 31456 5318 31512
rect 5170 31048 5226 31104
rect 5354 30932 5410 30968
rect 5354 30912 5356 30932
rect 5356 30912 5408 30932
rect 5408 30912 5410 30932
rect 5170 30776 5226 30832
rect 5170 30096 5226 30152
rect 5170 29008 5226 29064
rect 5354 30096 5410 30152
rect 5262 28600 5318 28656
rect 5078 27648 5134 27704
rect 5078 27376 5134 27432
rect 5354 27376 5410 27432
rect 5262 26560 5318 26616
rect 5078 25200 5134 25256
rect 4986 24384 5042 24440
rect 4802 23976 4858 24032
rect 5170 24792 5226 24848
rect 6154 38106 6210 38108
rect 6234 38106 6290 38108
rect 6314 38106 6370 38108
rect 6394 38106 6450 38108
rect 6154 38054 6200 38106
rect 6200 38054 6210 38106
rect 6234 38054 6264 38106
rect 6264 38054 6276 38106
rect 6276 38054 6290 38106
rect 6314 38054 6328 38106
rect 6328 38054 6340 38106
rect 6340 38054 6370 38106
rect 6394 38054 6404 38106
rect 6404 38054 6450 38106
rect 6154 38052 6210 38054
rect 6234 38052 6290 38054
rect 6314 38052 6370 38054
rect 6394 38052 6450 38054
rect 6550 37032 6606 37088
rect 6154 37018 6210 37020
rect 6234 37018 6290 37020
rect 6314 37018 6370 37020
rect 6394 37018 6450 37020
rect 6154 36966 6200 37018
rect 6200 36966 6210 37018
rect 6234 36966 6264 37018
rect 6264 36966 6276 37018
rect 6276 36966 6290 37018
rect 6314 36966 6328 37018
rect 6328 36966 6340 37018
rect 6340 36966 6370 37018
rect 6394 36966 6404 37018
rect 6404 36966 6450 37018
rect 6154 36964 6210 36966
rect 6234 36964 6290 36966
rect 6314 36964 6370 36966
rect 6394 36964 6450 36966
rect 5998 36896 6054 36952
rect 6090 36760 6146 36816
rect 6366 36488 6422 36544
rect 6154 35930 6210 35932
rect 6234 35930 6290 35932
rect 6314 35930 6370 35932
rect 6394 35930 6450 35932
rect 6154 35878 6200 35930
rect 6200 35878 6210 35930
rect 6234 35878 6264 35930
rect 6264 35878 6276 35930
rect 6276 35878 6290 35930
rect 6314 35878 6328 35930
rect 6328 35878 6340 35930
rect 6340 35878 6370 35930
rect 6394 35878 6404 35930
rect 6404 35878 6450 35930
rect 6154 35876 6210 35878
rect 6234 35876 6290 35878
rect 6314 35876 6370 35878
rect 6394 35876 6450 35878
rect 5998 35536 6054 35592
rect 6918 36760 6974 36816
rect 6918 36080 6974 36136
rect 7102 38120 7158 38176
rect 5998 34892 6000 34912
rect 6000 34892 6052 34912
rect 6052 34892 6054 34912
rect 5998 34856 6054 34892
rect 6154 34842 6210 34844
rect 6234 34842 6290 34844
rect 6314 34842 6370 34844
rect 6394 34842 6450 34844
rect 6154 34790 6200 34842
rect 6200 34790 6210 34842
rect 6234 34790 6264 34842
rect 6264 34790 6276 34842
rect 6276 34790 6290 34842
rect 6314 34790 6328 34842
rect 6328 34790 6340 34842
rect 6340 34790 6370 34842
rect 6394 34790 6404 34842
rect 6404 34790 6450 34842
rect 6154 34788 6210 34790
rect 6234 34788 6290 34790
rect 6314 34788 6370 34790
rect 6394 34788 6450 34790
rect 5722 31728 5778 31784
rect 6458 34176 6514 34232
rect 6826 34584 6882 34640
rect 6154 33754 6210 33756
rect 6234 33754 6290 33756
rect 6314 33754 6370 33756
rect 6394 33754 6450 33756
rect 6154 33702 6200 33754
rect 6200 33702 6210 33754
rect 6234 33702 6264 33754
rect 6264 33702 6276 33754
rect 6276 33702 6290 33754
rect 6314 33702 6328 33754
rect 6328 33702 6340 33754
rect 6340 33702 6370 33754
rect 6394 33702 6404 33754
rect 6404 33702 6450 33754
rect 6154 33700 6210 33702
rect 6234 33700 6290 33702
rect 6314 33700 6370 33702
rect 6394 33700 6450 33702
rect 6154 32666 6210 32668
rect 6234 32666 6290 32668
rect 6314 32666 6370 32668
rect 6394 32666 6450 32668
rect 6154 32614 6200 32666
rect 6200 32614 6210 32666
rect 6234 32614 6264 32666
rect 6264 32614 6276 32666
rect 6276 32614 6290 32666
rect 6314 32614 6328 32666
rect 6328 32614 6340 32666
rect 6340 32614 6370 32666
rect 6394 32614 6404 32666
rect 6404 32614 6450 32666
rect 6154 32612 6210 32614
rect 6234 32612 6290 32614
rect 6314 32612 6370 32614
rect 6394 32612 6450 32614
rect 5998 32272 6054 32328
rect 5906 30504 5962 30560
rect 5538 28056 5594 28112
rect 5538 26968 5594 27024
rect 5722 27920 5778 27976
rect 5262 23432 5318 23488
rect 5078 23296 5134 23352
rect 4618 22500 4674 22536
rect 4618 22480 4620 22500
rect 4620 22480 4672 22500
rect 4672 22480 4674 22500
rect 4618 21800 4674 21856
rect 4434 21256 4490 21312
rect 4066 20440 4122 20496
rect 4066 20168 4122 20224
rect 2686 17332 2742 17368
rect 2686 17312 2688 17332
rect 2688 17312 2740 17332
rect 2740 17312 2742 17332
rect 2134 15272 2190 15328
rect 2410 15136 2466 15192
rect 2594 15000 2650 15056
rect 1766 11772 1768 11792
rect 1768 11772 1820 11792
rect 1820 11772 1822 11792
rect 1766 11736 1822 11772
rect 1674 11328 1730 11384
rect 1674 9832 1730 9888
rect 1490 9424 1546 9480
rect 1582 9288 1638 9344
rect 1398 8744 1454 8800
rect 1398 8336 1454 8392
rect 1490 7928 1546 7984
rect 1214 6296 1270 6352
rect 1306 4664 1362 4720
rect 1490 7520 1546 7576
rect 1490 5344 1546 5400
rect 2318 11600 2374 11656
rect 2226 11056 2282 11112
rect 2594 13504 2650 13560
rect 2594 12688 2650 12744
rect 3054 15952 3110 16008
rect 4066 18264 4122 18320
rect 4342 20848 4398 20904
rect 4618 21120 4674 21176
rect 4618 19488 4674 19544
rect 3555 17978 3611 17980
rect 3635 17978 3691 17980
rect 3715 17978 3771 17980
rect 3795 17978 3851 17980
rect 3555 17926 3601 17978
rect 3601 17926 3611 17978
rect 3635 17926 3665 17978
rect 3665 17926 3677 17978
rect 3677 17926 3691 17978
rect 3715 17926 3729 17978
rect 3729 17926 3741 17978
rect 3741 17926 3771 17978
rect 3795 17926 3805 17978
rect 3805 17926 3851 17978
rect 3555 17924 3611 17926
rect 3635 17924 3691 17926
rect 3715 17924 3771 17926
rect 3795 17924 3851 17926
rect 3514 17584 3570 17640
rect 4066 17856 4122 17912
rect 4342 17720 4398 17776
rect 4158 17312 4214 17368
rect 3882 17040 3938 17096
rect 4066 17040 4122 17096
rect 3555 16890 3611 16892
rect 3635 16890 3691 16892
rect 3715 16890 3771 16892
rect 3795 16890 3851 16892
rect 3555 16838 3601 16890
rect 3601 16838 3611 16890
rect 3635 16838 3665 16890
rect 3665 16838 3677 16890
rect 3677 16838 3691 16890
rect 3715 16838 3729 16890
rect 3729 16838 3741 16890
rect 3741 16838 3771 16890
rect 3795 16838 3805 16890
rect 3805 16838 3851 16890
rect 3555 16836 3611 16838
rect 3635 16836 3691 16838
rect 3715 16836 3771 16838
rect 3795 16836 3851 16838
rect 3422 16768 3478 16824
rect 3606 16632 3662 16688
rect 2870 13676 2872 13696
rect 2872 13676 2924 13696
rect 2924 13676 2926 13696
rect 2870 13640 2926 13676
rect 3054 14048 3110 14104
rect 3974 16396 3976 16416
rect 3976 16396 4028 16416
rect 4028 16396 4030 16416
rect 3974 16360 4030 16396
rect 3555 15802 3611 15804
rect 3635 15802 3691 15804
rect 3715 15802 3771 15804
rect 3795 15802 3851 15804
rect 3555 15750 3601 15802
rect 3601 15750 3611 15802
rect 3635 15750 3665 15802
rect 3665 15750 3677 15802
rect 3677 15750 3691 15802
rect 3715 15750 3729 15802
rect 3729 15750 3741 15802
rect 3741 15750 3771 15802
rect 3795 15750 3805 15802
rect 3805 15750 3851 15802
rect 3555 15748 3611 15750
rect 3635 15748 3691 15750
rect 3715 15748 3771 15750
rect 3795 15748 3851 15750
rect 3555 14714 3611 14716
rect 3635 14714 3691 14716
rect 3715 14714 3771 14716
rect 3795 14714 3851 14716
rect 3555 14662 3601 14714
rect 3601 14662 3611 14714
rect 3635 14662 3665 14714
rect 3665 14662 3677 14714
rect 3677 14662 3691 14714
rect 3715 14662 3729 14714
rect 3729 14662 3741 14714
rect 3741 14662 3771 14714
rect 3795 14662 3805 14714
rect 3805 14662 3851 14714
rect 3555 14660 3611 14662
rect 3635 14660 3691 14662
rect 3715 14660 3771 14662
rect 3795 14660 3851 14662
rect 3882 14456 3938 14512
rect 3238 14320 3294 14376
rect 3882 14184 3938 14240
rect 2870 13096 2926 13152
rect 2778 12824 2834 12880
rect 2686 11600 2742 11656
rect 2594 11328 2650 11384
rect 2686 11056 2742 11112
rect 1766 8608 1822 8664
rect 1766 6976 1822 7032
rect 2226 9696 2282 9752
rect 2134 7792 2190 7848
rect 1490 3304 1546 3360
rect 1858 5072 1914 5128
rect 2686 10784 2742 10840
rect 2502 9288 2558 9344
rect 2410 8064 2466 8120
rect 2226 7112 2282 7168
rect 3054 12824 3110 12880
rect 3555 13626 3611 13628
rect 3635 13626 3691 13628
rect 3715 13626 3771 13628
rect 3795 13626 3851 13628
rect 3555 13574 3601 13626
rect 3601 13574 3611 13626
rect 3635 13574 3665 13626
rect 3665 13574 3677 13626
rect 3677 13574 3691 13626
rect 3715 13574 3729 13626
rect 3729 13574 3741 13626
rect 3741 13574 3771 13626
rect 3795 13574 3805 13626
rect 3805 13574 3851 13626
rect 3555 13572 3611 13574
rect 3635 13572 3691 13574
rect 3715 13572 3771 13574
rect 3795 13572 3851 13574
rect 3054 12552 3110 12608
rect 2778 10104 2834 10160
rect 3054 10240 3110 10296
rect 2870 7248 2926 7304
rect 2502 6704 2558 6760
rect 2502 6296 2558 6352
rect 2410 6160 2466 6216
rect 2042 3168 2098 3224
rect 2502 5616 2558 5672
rect 2778 6160 2834 6216
rect 2686 4528 2742 4584
rect 2870 3304 2926 3360
rect 3790 13268 3792 13288
rect 3792 13268 3844 13288
rect 3844 13268 3846 13288
rect 3790 13232 3846 13268
rect 3555 12538 3611 12540
rect 3635 12538 3691 12540
rect 3715 12538 3771 12540
rect 3795 12538 3851 12540
rect 3555 12486 3601 12538
rect 3601 12486 3611 12538
rect 3635 12486 3665 12538
rect 3665 12486 3677 12538
rect 3677 12486 3691 12538
rect 3715 12486 3729 12538
rect 3729 12486 3741 12538
rect 3741 12486 3771 12538
rect 3795 12486 3805 12538
rect 3805 12486 3851 12538
rect 3555 12484 3611 12486
rect 3635 12484 3691 12486
rect 3715 12484 3771 12486
rect 3795 12484 3851 12486
rect 3974 12552 4030 12608
rect 4250 14592 4306 14648
rect 5078 22888 5134 22944
rect 4526 16768 4582 16824
rect 4526 15580 4528 15600
rect 4528 15580 4580 15600
rect 4580 15580 4582 15600
rect 4526 15544 4582 15580
rect 4710 16088 4766 16144
rect 4434 14728 4490 14784
rect 3974 12280 4030 12336
rect 3555 11450 3611 11452
rect 3635 11450 3691 11452
rect 3715 11450 3771 11452
rect 3795 11450 3851 11452
rect 3555 11398 3601 11450
rect 3601 11398 3611 11450
rect 3635 11398 3665 11450
rect 3665 11398 3677 11450
rect 3677 11398 3691 11450
rect 3715 11398 3729 11450
rect 3729 11398 3741 11450
rect 3741 11398 3771 11450
rect 3795 11398 3805 11450
rect 3805 11398 3851 11450
rect 3555 11396 3611 11398
rect 3635 11396 3691 11398
rect 3715 11396 3771 11398
rect 3795 11396 3851 11398
rect 3330 9560 3386 9616
rect 4066 12008 4122 12064
rect 4158 11872 4214 11928
rect 3882 11192 3938 11248
rect 4066 10920 4122 10976
rect 3974 10648 4030 10704
rect 3555 10362 3611 10364
rect 3635 10362 3691 10364
rect 3715 10362 3771 10364
rect 3795 10362 3851 10364
rect 3555 10310 3601 10362
rect 3601 10310 3611 10362
rect 3635 10310 3665 10362
rect 3665 10310 3677 10362
rect 3677 10310 3691 10362
rect 3715 10310 3729 10362
rect 3729 10310 3741 10362
rect 3741 10310 3771 10362
rect 3795 10310 3805 10362
rect 3805 10310 3851 10362
rect 3555 10308 3611 10310
rect 3635 10308 3691 10310
rect 3715 10308 3771 10310
rect 3795 10308 3851 10310
rect 3974 10104 4030 10160
rect 4158 10648 4214 10704
rect 3882 9696 3938 9752
rect 3555 9274 3611 9276
rect 3635 9274 3691 9276
rect 3715 9274 3771 9276
rect 3795 9274 3851 9276
rect 3555 9222 3601 9274
rect 3601 9222 3611 9274
rect 3635 9222 3665 9274
rect 3665 9222 3677 9274
rect 3677 9222 3691 9274
rect 3715 9222 3729 9274
rect 3729 9222 3741 9274
rect 3741 9222 3771 9274
rect 3795 9222 3805 9274
rect 3805 9222 3851 9274
rect 3555 9220 3611 9222
rect 3635 9220 3691 9222
rect 3715 9220 3771 9222
rect 3795 9220 3851 9222
rect 3974 9152 4030 9208
rect 4618 15272 4674 15328
rect 4526 13640 4582 13696
rect 4434 13368 4490 13424
rect 4894 17856 4950 17912
rect 4986 17484 4988 17504
rect 4988 17484 5040 17504
rect 5040 17484 5042 17504
rect 4986 17448 5042 17484
rect 4894 16360 4950 16416
rect 4894 15816 4950 15872
rect 4894 15680 4950 15736
rect 5446 22752 5502 22808
rect 6154 31578 6210 31580
rect 6234 31578 6290 31580
rect 6314 31578 6370 31580
rect 6394 31578 6450 31580
rect 6154 31526 6200 31578
rect 6200 31526 6210 31578
rect 6234 31526 6264 31578
rect 6264 31526 6276 31578
rect 6276 31526 6290 31578
rect 6314 31526 6328 31578
rect 6328 31526 6340 31578
rect 6340 31526 6370 31578
rect 6394 31526 6404 31578
rect 6404 31526 6450 31578
rect 6154 31524 6210 31526
rect 6234 31524 6290 31526
rect 6314 31524 6370 31526
rect 6394 31524 6450 31526
rect 6366 31184 6422 31240
rect 6090 30776 6146 30832
rect 6826 32272 6882 32328
rect 6154 30490 6210 30492
rect 6234 30490 6290 30492
rect 6314 30490 6370 30492
rect 6394 30490 6450 30492
rect 6154 30438 6200 30490
rect 6200 30438 6210 30490
rect 6234 30438 6264 30490
rect 6264 30438 6276 30490
rect 6276 30438 6290 30490
rect 6314 30438 6328 30490
rect 6328 30438 6340 30490
rect 6340 30438 6370 30490
rect 6394 30438 6404 30490
rect 6404 30438 6450 30490
rect 6154 30436 6210 30438
rect 6234 30436 6290 30438
rect 6314 30436 6370 30438
rect 6394 30436 6450 30438
rect 6090 30232 6146 30288
rect 6366 29824 6422 29880
rect 5998 29416 6054 29472
rect 6154 29402 6210 29404
rect 6234 29402 6290 29404
rect 6314 29402 6370 29404
rect 6394 29402 6450 29404
rect 6154 29350 6200 29402
rect 6200 29350 6210 29402
rect 6234 29350 6264 29402
rect 6264 29350 6276 29402
rect 6276 29350 6290 29402
rect 6314 29350 6328 29402
rect 6328 29350 6340 29402
rect 6340 29350 6370 29402
rect 6394 29350 6404 29402
rect 6404 29350 6450 29402
rect 6154 29348 6210 29350
rect 6234 29348 6290 29350
rect 6314 29348 6370 29350
rect 6394 29348 6450 29350
rect 5998 29008 6054 29064
rect 6154 28314 6210 28316
rect 6234 28314 6290 28316
rect 6314 28314 6370 28316
rect 6394 28314 6450 28316
rect 6154 28262 6200 28314
rect 6200 28262 6210 28314
rect 6234 28262 6264 28314
rect 6264 28262 6276 28314
rect 6276 28262 6290 28314
rect 6314 28262 6328 28314
rect 6328 28262 6340 28314
rect 6340 28262 6370 28314
rect 6394 28262 6404 28314
rect 6404 28262 6450 28314
rect 6154 28260 6210 28262
rect 6234 28260 6290 28262
rect 6314 28260 6370 28262
rect 6394 28260 6450 28262
rect 6154 27226 6210 27228
rect 6234 27226 6290 27228
rect 6314 27226 6370 27228
rect 6394 27226 6450 27228
rect 6154 27174 6200 27226
rect 6200 27174 6210 27226
rect 6234 27174 6264 27226
rect 6264 27174 6276 27226
rect 6276 27174 6290 27226
rect 6314 27174 6328 27226
rect 6328 27174 6340 27226
rect 6340 27174 6370 27226
rect 6394 27174 6404 27226
rect 6404 27174 6450 27226
rect 6154 27172 6210 27174
rect 6234 27172 6290 27174
rect 6314 27172 6370 27174
rect 6394 27172 6450 27174
rect 6734 30096 6790 30152
rect 6642 28736 6698 28792
rect 5906 26152 5962 26208
rect 6366 26288 6422 26344
rect 6154 26138 6210 26140
rect 6234 26138 6290 26140
rect 6314 26138 6370 26140
rect 6394 26138 6450 26140
rect 6154 26086 6200 26138
rect 6200 26086 6210 26138
rect 6234 26086 6264 26138
rect 6264 26086 6276 26138
rect 6276 26086 6290 26138
rect 6314 26086 6328 26138
rect 6328 26086 6340 26138
rect 6340 26086 6370 26138
rect 6394 26086 6404 26138
rect 6404 26086 6450 26138
rect 6154 26084 6210 26086
rect 6234 26084 6290 26086
rect 6314 26084 6370 26086
rect 6394 26084 6450 26086
rect 7102 31728 7158 31784
rect 7102 30912 7158 30968
rect 7194 30232 7250 30288
rect 7010 29824 7066 29880
rect 6918 28464 6974 28520
rect 6826 26696 6882 26752
rect 7654 41148 7656 41168
rect 7656 41148 7708 41168
rect 7708 41148 7710 41168
rect 7654 41112 7710 41148
rect 8390 41656 8446 41712
rect 8942 43152 8998 43208
rect 8753 43002 8809 43004
rect 8833 43002 8889 43004
rect 8913 43002 8969 43004
rect 8993 43002 9049 43004
rect 8753 42950 8799 43002
rect 8799 42950 8809 43002
rect 8833 42950 8863 43002
rect 8863 42950 8875 43002
rect 8875 42950 8889 43002
rect 8913 42950 8927 43002
rect 8927 42950 8939 43002
rect 8939 42950 8969 43002
rect 8993 42950 9003 43002
rect 9003 42950 9049 43002
rect 8753 42948 8809 42950
rect 8833 42948 8889 42950
rect 8913 42948 8969 42950
rect 8993 42948 9049 42950
rect 8574 42608 8630 42664
rect 8390 41268 8446 41304
rect 8390 41248 8392 41268
rect 8392 41248 8444 41268
rect 8444 41248 8446 41268
rect 9402 42608 9458 42664
rect 9126 42336 9182 42392
rect 8942 42084 8998 42120
rect 8942 42064 8944 42084
rect 8944 42064 8996 42084
rect 8996 42064 8998 42084
rect 8753 41914 8809 41916
rect 8833 41914 8889 41916
rect 8913 41914 8969 41916
rect 8993 41914 9049 41916
rect 8753 41862 8799 41914
rect 8799 41862 8809 41914
rect 8833 41862 8863 41914
rect 8863 41862 8875 41914
rect 8875 41862 8889 41914
rect 8913 41862 8927 41914
rect 8927 41862 8939 41914
rect 8939 41862 8969 41914
rect 8993 41862 9003 41914
rect 9003 41862 9049 41914
rect 8753 41860 8809 41862
rect 8833 41860 8889 41862
rect 8913 41860 8969 41862
rect 8993 41860 9049 41862
rect 7562 38528 7618 38584
rect 7562 37848 7618 37904
rect 8022 40024 8078 40080
rect 7838 38120 7894 38176
rect 7838 37304 7894 37360
rect 7746 37068 7748 37088
rect 7748 37068 7800 37088
rect 7800 37068 7802 37088
rect 7746 37032 7802 37068
rect 7562 36780 7618 36816
rect 7562 36760 7564 36780
rect 7564 36760 7616 36780
rect 7616 36760 7618 36780
rect 7746 35944 7802 36000
rect 7654 35128 7710 35184
rect 7654 32816 7710 32872
rect 7654 32000 7710 32056
rect 7562 31048 7618 31104
rect 7562 29960 7618 30016
rect 7378 29008 7434 29064
rect 7102 27784 7158 27840
rect 7010 26560 7066 26616
rect 6826 26288 6882 26344
rect 6734 25608 6790 25664
rect 6642 25472 6698 25528
rect 6550 25200 6606 25256
rect 5998 25064 6054 25120
rect 6154 25050 6210 25052
rect 6234 25050 6290 25052
rect 6314 25050 6370 25052
rect 6394 25050 6450 25052
rect 6154 24998 6200 25050
rect 6200 24998 6210 25050
rect 6234 24998 6264 25050
rect 6264 24998 6276 25050
rect 6276 24998 6290 25050
rect 6314 24998 6328 25050
rect 6328 24998 6340 25050
rect 6340 24998 6370 25050
rect 6394 24998 6404 25050
rect 6404 24998 6450 25050
rect 6154 24996 6210 24998
rect 6234 24996 6290 24998
rect 6314 24996 6370 24998
rect 6394 24996 6450 24998
rect 5814 24384 5870 24440
rect 5814 24248 5870 24304
rect 5722 22480 5778 22536
rect 5538 21392 5594 21448
rect 5078 15136 5134 15192
rect 5354 19896 5410 19952
rect 5262 19488 5318 19544
rect 5262 18692 5318 18728
rect 5262 18672 5264 18692
rect 5264 18672 5316 18692
rect 5316 18672 5318 18692
rect 5538 19624 5594 19680
rect 5446 18128 5502 18184
rect 5446 17856 5502 17912
rect 5722 18128 5778 18184
rect 5538 16396 5540 16416
rect 5540 16396 5592 16416
rect 5592 16396 5594 16416
rect 5538 16360 5594 16396
rect 5078 14048 5134 14104
rect 5262 14184 5318 14240
rect 4894 13504 4950 13560
rect 4618 13232 4674 13288
rect 4986 13232 5042 13288
rect 4342 10920 4398 10976
rect 4618 10920 4674 10976
rect 4342 10784 4398 10840
rect 4066 8744 4122 8800
rect 3330 8200 3386 8256
rect 3238 7792 3294 7848
rect 3054 5072 3110 5128
rect 3330 6740 3332 6760
rect 3332 6740 3384 6760
rect 3384 6740 3386 6760
rect 3330 6704 3386 6740
rect 3555 8186 3611 8188
rect 3635 8186 3691 8188
rect 3715 8186 3771 8188
rect 3795 8186 3851 8188
rect 3555 8134 3601 8186
rect 3601 8134 3611 8186
rect 3635 8134 3665 8186
rect 3665 8134 3677 8186
rect 3677 8134 3691 8186
rect 3715 8134 3729 8186
rect 3729 8134 3741 8186
rect 3741 8134 3771 8186
rect 3795 8134 3805 8186
rect 3805 8134 3851 8186
rect 3555 8132 3611 8134
rect 3635 8132 3691 8134
rect 3715 8132 3771 8134
rect 3795 8132 3851 8134
rect 3790 7828 3792 7848
rect 3792 7828 3844 7848
rect 3844 7828 3846 7848
rect 3790 7792 3846 7828
rect 4158 7656 4214 7712
rect 4802 10512 4858 10568
rect 4802 9968 4858 10024
rect 4710 9288 4766 9344
rect 4710 9016 4766 9072
rect 4526 8336 4582 8392
rect 4526 8064 4582 8120
rect 4158 7384 4214 7440
rect 3555 7098 3611 7100
rect 3635 7098 3691 7100
rect 3715 7098 3771 7100
rect 3795 7098 3851 7100
rect 3555 7046 3601 7098
rect 3601 7046 3611 7098
rect 3635 7046 3665 7098
rect 3665 7046 3677 7098
rect 3677 7046 3691 7098
rect 3715 7046 3729 7098
rect 3729 7046 3741 7098
rect 3741 7046 3771 7098
rect 3795 7046 3805 7098
rect 3805 7046 3851 7098
rect 3555 7044 3611 7046
rect 3635 7044 3691 7046
rect 3715 7044 3771 7046
rect 3795 7044 3851 7046
rect 3330 5616 3386 5672
rect 3514 6160 3570 6216
rect 3790 6704 3846 6760
rect 3882 6432 3938 6488
rect 3555 6010 3611 6012
rect 3635 6010 3691 6012
rect 3715 6010 3771 6012
rect 3795 6010 3851 6012
rect 3555 5958 3601 6010
rect 3601 5958 3611 6010
rect 3635 5958 3665 6010
rect 3665 5958 3677 6010
rect 3677 5958 3691 6010
rect 3715 5958 3729 6010
rect 3729 5958 3741 6010
rect 3741 5958 3771 6010
rect 3795 5958 3805 6010
rect 3805 5958 3851 6010
rect 3555 5956 3611 5958
rect 3635 5956 3691 5958
rect 3715 5956 3771 5958
rect 3795 5956 3851 5958
rect 4066 6840 4122 6896
rect 4250 6876 4252 6896
rect 4252 6876 4304 6896
rect 4304 6876 4306 6896
rect 4250 6840 4306 6876
rect 4250 6740 4252 6760
rect 4252 6740 4304 6760
rect 4304 6740 4306 6760
rect 4250 6704 4306 6740
rect 4158 6296 4214 6352
rect 4434 7384 4490 7440
rect 4526 7112 4582 7168
rect 4710 7404 4766 7440
rect 4710 7384 4712 7404
rect 4712 7384 4764 7404
rect 4764 7384 4766 7404
rect 5078 12280 5134 12336
rect 4986 11464 5042 11520
rect 4986 10784 5042 10840
rect 4618 6704 4674 6760
rect 4618 6568 4674 6624
rect 4434 6160 4490 6216
rect 4066 5752 4122 5808
rect 4158 5652 4160 5672
rect 4160 5652 4212 5672
rect 4212 5652 4214 5672
rect 4158 5616 4214 5652
rect 3555 4922 3611 4924
rect 3635 4922 3691 4924
rect 3715 4922 3771 4924
rect 3795 4922 3851 4924
rect 3555 4870 3601 4922
rect 3601 4870 3611 4922
rect 3635 4870 3665 4922
rect 3665 4870 3677 4922
rect 3677 4870 3691 4922
rect 3715 4870 3729 4922
rect 3729 4870 3741 4922
rect 3741 4870 3771 4922
rect 3795 4870 3805 4922
rect 3805 4870 3851 4922
rect 3555 4868 3611 4870
rect 3635 4868 3691 4870
rect 3715 4868 3771 4870
rect 3795 4868 3851 4870
rect 3606 4528 3662 4584
rect 3698 4392 3754 4448
rect 4066 5480 4122 5536
rect 4066 5208 4122 5264
rect 3555 3834 3611 3836
rect 3635 3834 3691 3836
rect 3715 3834 3771 3836
rect 3795 3834 3851 3836
rect 3555 3782 3601 3834
rect 3601 3782 3611 3834
rect 3635 3782 3665 3834
rect 3665 3782 3677 3834
rect 3677 3782 3691 3834
rect 3715 3782 3729 3834
rect 3729 3782 3741 3834
rect 3741 3782 3771 3834
rect 3795 3782 3805 3834
rect 3805 3782 3851 3834
rect 3555 3780 3611 3782
rect 3635 3780 3691 3782
rect 3715 3780 3771 3782
rect 3795 3780 3851 3782
rect 4158 3576 4214 3632
rect 4066 2896 4122 2952
rect 3555 2746 3611 2748
rect 3635 2746 3691 2748
rect 3715 2746 3771 2748
rect 3795 2746 3851 2748
rect 2870 2488 2926 2544
rect 1490 720 1546 776
rect 3555 2694 3601 2746
rect 3601 2694 3611 2746
rect 3635 2694 3665 2746
rect 3665 2694 3677 2746
rect 3677 2694 3691 2746
rect 3715 2694 3729 2746
rect 3729 2694 3741 2746
rect 3741 2694 3771 2746
rect 3795 2694 3805 2746
rect 3805 2694 3851 2746
rect 3555 2692 3611 2694
rect 3635 2692 3691 2694
rect 3715 2692 3771 2694
rect 3795 2692 3851 2694
rect 5354 13232 5410 13288
rect 5354 12008 5410 12064
rect 5354 11464 5410 11520
rect 6090 24520 6146 24576
rect 6154 23962 6210 23964
rect 6234 23962 6290 23964
rect 6314 23962 6370 23964
rect 6394 23962 6450 23964
rect 6154 23910 6200 23962
rect 6200 23910 6210 23962
rect 6234 23910 6264 23962
rect 6264 23910 6276 23962
rect 6276 23910 6290 23962
rect 6314 23910 6328 23962
rect 6328 23910 6340 23962
rect 6340 23910 6370 23962
rect 6394 23910 6404 23962
rect 6404 23910 6450 23962
rect 6154 23908 6210 23910
rect 6234 23908 6290 23910
rect 6314 23908 6370 23910
rect 6394 23908 6450 23910
rect 6550 23160 6606 23216
rect 6154 22874 6210 22876
rect 6234 22874 6290 22876
rect 6314 22874 6370 22876
rect 6394 22874 6450 22876
rect 6154 22822 6200 22874
rect 6200 22822 6210 22874
rect 6234 22822 6264 22874
rect 6264 22822 6276 22874
rect 6276 22822 6290 22874
rect 6314 22822 6328 22874
rect 6328 22822 6340 22874
rect 6340 22822 6370 22874
rect 6394 22822 6404 22874
rect 6404 22822 6450 22874
rect 6154 22820 6210 22822
rect 6234 22820 6290 22822
rect 6314 22820 6370 22822
rect 6394 22820 6450 22822
rect 6458 22208 6514 22264
rect 6274 21936 6330 21992
rect 6154 21786 6210 21788
rect 6234 21786 6290 21788
rect 6314 21786 6370 21788
rect 6394 21786 6450 21788
rect 6154 21734 6200 21786
rect 6200 21734 6210 21786
rect 6234 21734 6264 21786
rect 6264 21734 6276 21786
rect 6276 21734 6290 21786
rect 6314 21734 6328 21786
rect 6328 21734 6340 21786
rect 6340 21734 6370 21786
rect 6394 21734 6404 21786
rect 6404 21734 6450 21786
rect 6154 21732 6210 21734
rect 6234 21732 6290 21734
rect 6314 21732 6370 21734
rect 6394 21732 6450 21734
rect 6182 20848 6238 20904
rect 6154 20698 6210 20700
rect 6234 20698 6290 20700
rect 6314 20698 6370 20700
rect 6394 20698 6450 20700
rect 6154 20646 6200 20698
rect 6200 20646 6210 20698
rect 6234 20646 6264 20698
rect 6264 20646 6276 20698
rect 6276 20646 6290 20698
rect 6314 20646 6328 20698
rect 6328 20646 6340 20698
rect 6340 20646 6370 20698
rect 6394 20646 6404 20698
rect 6404 20646 6450 20698
rect 6154 20644 6210 20646
rect 6234 20644 6290 20646
rect 6314 20644 6370 20646
rect 6394 20644 6450 20646
rect 6458 20476 6460 20496
rect 6460 20476 6512 20496
rect 6512 20476 6514 20496
rect 6458 20440 6514 20476
rect 7286 27648 7342 27704
rect 7562 29008 7618 29064
rect 7930 35128 7986 35184
rect 8298 38392 8354 38448
rect 8298 35672 8354 35728
rect 8206 34720 8262 34776
rect 8022 33924 8078 33960
rect 8022 33904 8024 33924
rect 8024 33904 8076 33924
rect 8076 33904 8078 33924
rect 8206 33904 8262 33960
rect 7930 32136 7986 32192
rect 8114 31728 8170 31784
rect 7838 28636 7840 28656
rect 7840 28636 7892 28656
rect 7892 28636 7894 28656
rect 7838 28600 7894 28636
rect 7746 27920 7802 27976
rect 7654 27648 7710 27704
rect 7378 26988 7434 27024
rect 7378 26968 7380 26988
rect 7380 26968 7432 26988
rect 7432 26968 7434 26988
rect 7010 25472 7066 25528
rect 7194 24112 7250 24168
rect 7838 26324 7840 26344
rect 7840 26324 7892 26344
rect 7892 26324 7894 26344
rect 7838 26288 7894 26324
rect 7746 25608 7802 25664
rect 7286 23160 7342 23216
rect 7286 21256 7342 21312
rect 6918 20712 6974 20768
rect 6154 19610 6210 19612
rect 6234 19610 6290 19612
rect 6314 19610 6370 19612
rect 6394 19610 6450 19612
rect 6154 19558 6200 19610
rect 6200 19558 6210 19610
rect 6234 19558 6264 19610
rect 6264 19558 6276 19610
rect 6276 19558 6290 19610
rect 6314 19558 6328 19610
rect 6328 19558 6340 19610
rect 6340 19558 6370 19610
rect 6394 19558 6404 19610
rect 6404 19558 6450 19610
rect 6154 19556 6210 19558
rect 6234 19556 6290 19558
rect 6314 19556 6370 19558
rect 6394 19556 6450 19558
rect 6154 18522 6210 18524
rect 6234 18522 6290 18524
rect 6314 18522 6370 18524
rect 6394 18522 6450 18524
rect 6154 18470 6200 18522
rect 6200 18470 6210 18522
rect 6234 18470 6264 18522
rect 6264 18470 6276 18522
rect 6276 18470 6290 18522
rect 6314 18470 6328 18522
rect 6328 18470 6340 18522
rect 6340 18470 6370 18522
rect 6394 18470 6404 18522
rect 6404 18470 6450 18522
rect 6154 18468 6210 18470
rect 6234 18468 6290 18470
rect 6314 18468 6370 18470
rect 6394 18468 6450 18470
rect 6642 18536 6698 18592
rect 6182 17876 6238 17912
rect 6182 17856 6184 17876
rect 6184 17856 6236 17876
rect 6236 17856 6238 17876
rect 6154 17434 6210 17436
rect 6234 17434 6290 17436
rect 6314 17434 6370 17436
rect 6394 17434 6450 17436
rect 6154 17382 6200 17434
rect 6200 17382 6210 17434
rect 6234 17382 6264 17434
rect 6264 17382 6276 17434
rect 6276 17382 6290 17434
rect 6314 17382 6328 17434
rect 6328 17382 6340 17434
rect 6340 17382 6370 17434
rect 6394 17382 6404 17434
rect 6404 17382 6450 17434
rect 6154 17380 6210 17382
rect 6234 17380 6290 17382
rect 6314 17380 6370 17382
rect 6394 17380 6450 17382
rect 5722 14864 5778 14920
rect 5906 16652 5962 16688
rect 5906 16632 5908 16652
rect 5908 16632 5960 16652
rect 5960 16632 5962 16652
rect 6154 16346 6210 16348
rect 6234 16346 6290 16348
rect 6314 16346 6370 16348
rect 6394 16346 6450 16348
rect 6154 16294 6200 16346
rect 6200 16294 6210 16346
rect 6234 16294 6264 16346
rect 6264 16294 6276 16346
rect 6276 16294 6290 16346
rect 6314 16294 6328 16346
rect 6328 16294 6340 16346
rect 6340 16294 6370 16346
rect 6394 16294 6404 16346
rect 6404 16294 6450 16346
rect 6154 16292 6210 16294
rect 6234 16292 6290 16294
rect 6314 16292 6370 16294
rect 6394 16292 6450 16294
rect 5998 15308 6000 15328
rect 6000 15308 6052 15328
rect 6052 15308 6054 15328
rect 5998 15272 6054 15308
rect 6154 15258 6210 15260
rect 6234 15258 6290 15260
rect 6314 15258 6370 15260
rect 6394 15258 6450 15260
rect 6154 15206 6200 15258
rect 6200 15206 6210 15258
rect 6234 15206 6264 15258
rect 6264 15206 6276 15258
rect 6276 15206 6290 15258
rect 6314 15206 6328 15258
rect 6328 15206 6340 15258
rect 6340 15206 6370 15258
rect 6394 15206 6404 15258
rect 6404 15206 6450 15258
rect 6154 15204 6210 15206
rect 6234 15204 6290 15206
rect 6314 15204 6370 15206
rect 6394 15204 6450 15206
rect 6458 14728 6514 14784
rect 6154 14170 6210 14172
rect 6234 14170 6290 14172
rect 6314 14170 6370 14172
rect 6394 14170 6450 14172
rect 6154 14118 6200 14170
rect 6200 14118 6210 14170
rect 6234 14118 6264 14170
rect 6264 14118 6276 14170
rect 6276 14118 6290 14170
rect 6314 14118 6328 14170
rect 6328 14118 6340 14170
rect 6340 14118 6370 14170
rect 6394 14118 6404 14170
rect 6404 14118 6450 14170
rect 6154 14116 6210 14118
rect 6234 14116 6290 14118
rect 6314 14116 6370 14118
rect 6394 14116 6450 14118
rect 5906 13504 5962 13560
rect 5722 13268 5724 13288
rect 5724 13268 5776 13288
rect 5776 13268 5778 13288
rect 5722 13232 5778 13268
rect 6274 13368 6330 13424
rect 6154 13082 6210 13084
rect 6234 13082 6290 13084
rect 6314 13082 6370 13084
rect 6394 13082 6450 13084
rect 6154 13030 6200 13082
rect 6200 13030 6210 13082
rect 6234 13030 6264 13082
rect 6264 13030 6276 13082
rect 6276 13030 6290 13082
rect 6314 13030 6328 13082
rect 6328 13030 6340 13082
rect 6340 13030 6370 13082
rect 6394 13030 6404 13082
rect 6404 13030 6450 13082
rect 6154 13028 6210 13030
rect 6234 13028 6290 13030
rect 6314 13028 6370 13030
rect 6394 13028 6450 13030
rect 5722 12416 5778 12472
rect 5630 11736 5686 11792
rect 6274 12280 6330 12336
rect 5998 12008 6054 12064
rect 6154 11994 6210 11996
rect 6234 11994 6290 11996
rect 6314 11994 6370 11996
rect 6394 11994 6450 11996
rect 6154 11942 6200 11994
rect 6200 11942 6210 11994
rect 6234 11942 6264 11994
rect 6264 11942 6276 11994
rect 6276 11942 6290 11994
rect 6314 11942 6328 11994
rect 6328 11942 6340 11994
rect 6340 11942 6370 11994
rect 6394 11942 6404 11994
rect 6404 11942 6450 11994
rect 6154 11940 6210 11942
rect 6234 11940 6290 11942
rect 6314 11940 6370 11942
rect 6394 11940 6450 11942
rect 7102 18400 7158 18456
rect 7286 20576 7342 20632
rect 7378 19760 7434 19816
rect 7194 18264 7250 18320
rect 7102 18128 7158 18184
rect 7010 17856 7066 17912
rect 7010 17604 7066 17640
rect 7010 17584 7012 17604
rect 7012 17584 7064 17604
rect 7064 17584 7066 17604
rect 6734 14320 6790 14376
rect 7562 22208 7618 22264
rect 7378 17448 7434 17504
rect 7194 15544 7250 15600
rect 6918 12416 6974 12472
rect 7286 14728 7342 14784
rect 7286 12960 7342 13016
rect 7378 12860 7380 12880
rect 7380 12860 7432 12880
rect 7432 12860 7434 12880
rect 7378 12824 7434 12860
rect 5078 9968 5134 10024
rect 5078 9832 5134 9888
rect 6366 11464 6422 11520
rect 5630 10648 5686 10704
rect 5630 9696 5686 9752
rect 4986 6976 5042 7032
rect 5354 8608 5410 8664
rect 4894 4936 4950 4992
rect 4342 4548 4398 4584
rect 4342 4528 4344 4548
rect 4344 4528 4396 4548
rect 4396 4528 4398 4548
rect 3330 1128 3386 1184
rect 4986 4528 5042 4584
rect 4158 2488 4214 2544
rect 3555 1658 3611 1660
rect 3635 1658 3691 1660
rect 3715 1658 3771 1660
rect 3795 1658 3851 1660
rect 3555 1606 3601 1658
rect 3601 1606 3611 1658
rect 3635 1606 3665 1658
rect 3665 1606 3677 1658
rect 3677 1606 3691 1658
rect 3715 1606 3729 1658
rect 3729 1606 3741 1658
rect 3741 1606 3771 1658
rect 3795 1606 3805 1658
rect 3805 1606 3851 1658
rect 3555 1604 3611 1606
rect 3635 1604 3691 1606
rect 3715 1604 3771 1606
rect 3795 1604 3851 1606
rect 3514 1264 3570 1320
rect 4802 2216 4858 2272
rect 4802 720 4858 776
rect 5262 8064 5318 8120
rect 5722 9560 5778 9616
rect 5722 9288 5778 9344
rect 5446 7112 5502 7168
rect 5446 6840 5502 6896
rect 5262 6296 5318 6352
rect 5446 6568 5502 6624
rect 5170 3984 5226 4040
rect 5262 3576 5318 3632
rect 5446 3168 5502 3224
rect 5446 3052 5502 3088
rect 5446 3032 5448 3052
rect 5448 3032 5500 3052
rect 5500 3032 5502 3052
rect 5446 2216 5502 2272
rect 6154 10906 6210 10908
rect 6234 10906 6290 10908
rect 6314 10906 6370 10908
rect 6394 10906 6450 10908
rect 6154 10854 6200 10906
rect 6200 10854 6210 10906
rect 6234 10854 6264 10906
rect 6264 10854 6276 10906
rect 6276 10854 6290 10906
rect 6314 10854 6328 10906
rect 6328 10854 6340 10906
rect 6340 10854 6370 10906
rect 6394 10854 6404 10906
rect 6404 10854 6450 10906
rect 6154 10852 6210 10854
rect 6234 10852 6290 10854
rect 6314 10852 6370 10854
rect 6394 10852 6450 10854
rect 6090 10648 6146 10704
rect 6550 10240 6606 10296
rect 6154 9818 6210 9820
rect 6234 9818 6290 9820
rect 6314 9818 6370 9820
rect 6394 9818 6450 9820
rect 6154 9766 6200 9818
rect 6200 9766 6210 9818
rect 6234 9766 6264 9818
rect 6264 9766 6276 9818
rect 6276 9766 6290 9818
rect 6314 9766 6328 9818
rect 6328 9766 6340 9818
rect 6340 9766 6370 9818
rect 6394 9766 6404 9818
rect 6404 9766 6450 9818
rect 6154 9764 6210 9766
rect 6234 9764 6290 9766
rect 6314 9764 6370 9766
rect 6394 9764 6450 9766
rect 6458 9016 6514 9072
rect 6154 8730 6210 8732
rect 6234 8730 6290 8732
rect 6314 8730 6370 8732
rect 6394 8730 6450 8732
rect 6154 8678 6200 8730
rect 6200 8678 6210 8730
rect 6234 8678 6264 8730
rect 6264 8678 6276 8730
rect 6276 8678 6290 8730
rect 6314 8678 6328 8730
rect 6328 8678 6340 8730
rect 6340 8678 6370 8730
rect 6394 8678 6404 8730
rect 6404 8678 6450 8730
rect 6154 8676 6210 8678
rect 6234 8676 6290 8678
rect 6314 8676 6370 8678
rect 6394 8676 6450 8678
rect 6274 8492 6330 8528
rect 6274 8472 6276 8492
rect 6276 8472 6328 8492
rect 6328 8472 6330 8492
rect 6154 7642 6210 7644
rect 6234 7642 6290 7644
rect 6314 7642 6370 7644
rect 6394 7642 6450 7644
rect 6154 7590 6200 7642
rect 6200 7590 6210 7642
rect 6234 7590 6264 7642
rect 6264 7590 6276 7642
rect 6276 7590 6290 7642
rect 6314 7590 6328 7642
rect 6328 7590 6340 7642
rect 6340 7590 6370 7642
rect 6394 7590 6404 7642
rect 6404 7590 6450 7642
rect 6154 7588 6210 7590
rect 6234 7588 6290 7590
rect 6314 7588 6370 7590
rect 6394 7588 6450 7590
rect 6090 7112 6146 7168
rect 5906 6860 5962 6896
rect 5906 6840 5908 6860
rect 5908 6840 5960 6860
rect 5960 6840 5962 6860
rect 6154 6554 6210 6556
rect 6234 6554 6290 6556
rect 6314 6554 6370 6556
rect 6394 6554 6450 6556
rect 6154 6502 6200 6554
rect 6200 6502 6210 6554
rect 6234 6502 6264 6554
rect 6264 6502 6276 6554
rect 6276 6502 6290 6554
rect 6314 6502 6328 6554
rect 6328 6502 6340 6554
rect 6340 6502 6370 6554
rect 6394 6502 6404 6554
rect 6404 6502 6450 6554
rect 6154 6500 6210 6502
rect 6234 6500 6290 6502
rect 6314 6500 6370 6502
rect 6394 6500 6450 6502
rect 6182 6160 6238 6216
rect 5998 6060 6000 6080
rect 6000 6060 6052 6080
rect 6052 6060 6054 6080
rect 5998 6024 6054 6060
rect 6274 6024 6330 6080
rect 6826 10668 6882 10704
rect 6826 10648 6828 10668
rect 6828 10648 6880 10668
rect 6880 10648 6882 10668
rect 7378 12280 7434 12336
rect 7194 12008 7250 12064
rect 6918 10412 6920 10432
rect 6920 10412 6972 10432
rect 6972 10412 6974 10432
rect 6918 10376 6974 10412
rect 7010 9696 7066 9752
rect 6918 9424 6974 9480
rect 7010 8608 7066 8664
rect 6826 7792 6882 7848
rect 6734 7656 6790 7712
rect 7102 7828 7104 7848
rect 7104 7828 7156 7848
rect 7156 7828 7158 7848
rect 7102 7792 7158 7828
rect 6918 7112 6974 7168
rect 6642 6160 6698 6216
rect 6154 5466 6210 5468
rect 6234 5466 6290 5468
rect 6314 5466 6370 5468
rect 6394 5466 6450 5468
rect 6154 5414 6200 5466
rect 6200 5414 6210 5466
rect 6234 5414 6264 5466
rect 6264 5414 6276 5466
rect 6276 5414 6290 5466
rect 6314 5414 6328 5466
rect 6328 5414 6340 5466
rect 6340 5414 6370 5466
rect 6394 5414 6404 5466
rect 6404 5414 6450 5466
rect 6154 5412 6210 5414
rect 6234 5412 6290 5414
rect 6314 5412 6370 5414
rect 6394 5412 6450 5414
rect 5998 5228 6054 5264
rect 5998 5208 6000 5228
rect 6000 5208 6052 5228
rect 6052 5208 6054 5228
rect 5722 3304 5778 3360
rect 5630 2488 5686 2544
rect 5722 2100 5778 2136
rect 5722 2080 5724 2100
rect 5724 2080 5776 2100
rect 5776 2080 5778 2100
rect 6154 4378 6210 4380
rect 6234 4378 6290 4380
rect 6314 4378 6370 4380
rect 6394 4378 6450 4380
rect 6154 4326 6200 4378
rect 6200 4326 6210 4378
rect 6234 4326 6264 4378
rect 6264 4326 6276 4378
rect 6276 4326 6290 4378
rect 6314 4326 6328 4378
rect 6328 4326 6340 4378
rect 6340 4326 6370 4378
rect 6394 4326 6404 4378
rect 6404 4326 6450 4378
rect 6154 4324 6210 4326
rect 6234 4324 6290 4326
rect 6314 4324 6370 4326
rect 6394 4324 6450 4326
rect 6154 3290 6210 3292
rect 6234 3290 6290 3292
rect 6314 3290 6370 3292
rect 6394 3290 6450 3292
rect 6154 3238 6200 3290
rect 6200 3238 6210 3290
rect 6234 3238 6264 3290
rect 6264 3238 6276 3290
rect 6276 3238 6290 3290
rect 6314 3238 6328 3290
rect 6328 3238 6340 3290
rect 6340 3238 6370 3290
rect 6394 3238 6404 3290
rect 6404 3238 6450 3290
rect 6154 3236 6210 3238
rect 6234 3236 6290 3238
rect 6314 3236 6370 3238
rect 6394 3236 6450 3238
rect 6550 2488 6606 2544
rect 6274 2372 6330 2408
rect 6274 2352 6276 2372
rect 6276 2352 6328 2372
rect 6328 2352 6330 2372
rect 6154 2202 6210 2204
rect 6234 2202 6290 2204
rect 6314 2202 6370 2204
rect 6394 2202 6450 2204
rect 6154 2150 6200 2202
rect 6200 2150 6210 2202
rect 6234 2150 6264 2202
rect 6264 2150 6276 2202
rect 6276 2150 6290 2202
rect 6314 2150 6328 2202
rect 6328 2150 6340 2202
rect 6340 2150 6370 2202
rect 6394 2150 6404 2202
rect 6404 2150 6450 2202
rect 6154 2148 6210 2150
rect 6234 2148 6290 2150
rect 6314 2148 6370 2150
rect 6394 2148 6450 2150
rect 6154 1114 6210 1116
rect 6234 1114 6290 1116
rect 6314 1114 6370 1116
rect 6394 1114 6450 1116
rect 6154 1062 6200 1114
rect 6200 1062 6210 1114
rect 6234 1062 6264 1114
rect 6264 1062 6276 1114
rect 6276 1062 6290 1114
rect 6314 1062 6328 1114
rect 6328 1062 6340 1114
rect 6340 1062 6370 1114
rect 6394 1062 6404 1114
rect 6404 1062 6450 1114
rect 6154 1060 6210 1062
rect 6234 1060 6290 1062
rect 6314 1060 6370 1062
rect 6394 1060 6450 1062
rect 7378 10920 7434 10976
rect 7378 8064 7434 8120
rect 7378 6160 7434 6216
rect 7378 4936 7434 4992
rect 8574 38256 8630 38312
rect 8482 37612 8484 37632
rect 8484 37612 8536 37632
rect 8536 37612 8538 37632
rect 8482 37576 8538 37612
rect 8753 40826 8809 40828
rect 8833 40826 8889 40828
rect 8913 40826 8969 40828
rect 8993 40826 9049 40828
rect 8753 40774 8799 40826
rect 8799 40774 8809 40826
rect 8833 40774 8863 40826
rect 8863 40774 8875 40826
rect 8875 40774 8889 40826
rect 8913 40774 8927 40826
rect 8927 40774 8939 40826
rect 8939 40774 8969 40826
rect 8993 40774 9003 40826
rect 9003 40774 9049 40826
rect 8753 40772 8809 40774
rect 8833 40772 8889 40774
rect 8913 40772 8969 40774
rect 8993 40772 9049 40774
rect 9402 42064 9458 42120
rect 8753 39738 8809 39740
rect 8833 39738 8889 39740
rect 8913 39738 8969 39740
rect 8993 39738 9049 39740
rect 8753 39686 8799 39738
rect 8799 39686 8809 39738
rect 8833 39686 8863 39738
rect 8863 39686 8875 39738
rect 8875 39686 8889 39738
rect 8913 39686 8927 39738
rect 8927 39686 8939 39738
rect 8939 39686 8969 39738
rect 8993 39686 9003 39738
rect 9003 39686 9049 39738
rect 8753 39684 8809 39686
rect 8833 39684 8889 39686
rect 8913 39684 8969 39686
rect 8993 39684 9049 39686
rect 9586 41792 9642 41848
rect 8753 38650 8809 38652
rect 8833 38650 8889 38652
rect 8913 38650 8969 38652
rect 8993 38650 9049 38652
rect 8753 38598 8799 38650
rect 8799 38598 8809 38650
rect 8833 38598 8863 38650
rect 8863 38598 8875 38650
rect 8875 38598 8889 38650
rect 8913 38598 8927 38650
rect 8927 38598 8939 38650
rect 8939 38598 8969 38650
rect 8993 38598 9003 38650
rect 9003 38598 9049 38650
rect 8753 38596 8809 38598
rect 8833 38596 8889 38598
rect 8913 38596 8969 38598
rect 8993 38596 9049 38598
rect 8753 37562 8809 37564
rect 8833 37562 8889 37564
rect 8913 37562 8969 37564
rect 8993 37562 9049 37564
rect 8753 37510 8799 37562
rect 8799 37510 8809 37562
rect 8833 37510 8863 37562
rect 8863 37510 8875 37562
rect 8875 37510 8889 37562
rect 8913 37510 8927 37562
rect 8927 37510 8939 37562
rect 8939 37510 8969 37562
rect 8993 37510 9003 37562
rect 9003 37510 9049 37562
rect 8753 37508 8809 37510
rect 8833 37508 8889 37510
rect 8913 37508 8969 37510
rect 8993 37508 9049 37510
rect 8753 36474 8809 36476
rect 8833 36474 8889 36476
rect 8913 36474 8969 36476
rect 8993 36474 9049 36476
rect 8753 36422 8799 36474
rect 8799 36422 8809 36474
rect 8833 36422 8863 36474
rect 8863 36422 8875 36474
rect 8875 36422 8889 36474
rect 8913 36422 8927 36474
rect 8927 36422 8939 36474
rect 8939 36422 8969 36474
rect 8993 36422 9003 36474
rect 9003 36422 9049 36474
rect 8753 36420 8809 36422
rect 8833 36420 8889 36422
rect 8913 36420 8969 36422
rect 8993 36420 9049 36422
rect 8666 36080 8722 36136
rect 8666 35808 8722 35864
rect 8574 35708 8576 35728
rect 8576 35708 8628 35728
rect 8628 35708 8630 35728
rect 8574 35672 8630 35708
rect 8482 35400 8538 35456
rect 8753 35386 8809 35388
rect 8833 35386 8889 35388
rect 8913 35386 8969 35388
rect 8993 35386 9049 35388
rect 8753 35334 8799 35386
rect 8799 35334 8809 35386
rect 8833 35334 8863 35386
rect 8863 35334 8875 35386
rect 8875 35334 8889 35386
rect 8913 35334 8927 35386
rect 8927 35334 8939 35386
rect 8939 35334 8969 35386
rect 8993 35334 9003 35386
rect 9003 35334 9049 35386
rect 8753 35332 8809 35334
rect 8833 35332 8889 35334
rect 8913 35332 8969 35334
rect 8993 35332 9049 35334
rect 8574 34720 8630 34776
rect 8022 28736 8078 28792
rect 8022 28056 8078 28112
rect 7930 24248 7986 24304
rect 8114 26560 8170 26616
rect 8753 34298 8809 34300
rect 8833 34298 8889 34300
rect 8913 34298 8969 34300
rect 8993 34298 9049 34300
rect 8753 34246 8799 34298
rect 8799 34246 8809 34298
rect 8833 34246 8863 34298
rect 8863 34246 8875 34298
rect 8875 34246 8889 34298
rect 8913 34246 8927 34298
rect 8927 34246 8939 34298
rect 8939 34246 8969 34298
rect 8993 34246 9003 34298
rect 9003 34246 9049 34298
rect 8753 34244 8809 34246
rect 8833 34244 8889 34246
rect 8913 34244 8969 34246
rect 8993 34244 9049 34246
rect 8574 32272 8630 32328
rect 8482 32000 8538 32056
rect 8482 31764 8484 31784
rect 8484 31764 8536 31784
rect 8536 31764 8538 31784
rect 8482 31728 8538 31764
rect 8482 31184 8538 31240
rect 8298 28056 8354 28112
rect 8206 26288 8262 26344
rect 8574 28872 8630 28928
rect 8482 28464 8538 28520
rect 8753 33210 8809 33212
rect 8833 33210 8889 33212
rect 8913 33210 8969 33212
rect 8993 33210 9049 33212
rect 8753 33158 8799 33210
rect 8799 33158 8809 33210
rect 8833 33158 8863 33210
rect 8863 33158 8875 33210
rect 8875 33158 8889 33210
rect 8913 33158 8927 33210
rect 8927 33158 8939 33210
rect 8939 33158 8969 33210
rect 8993 33158 9003 33210
rect 9003 33158 9049 33210
rect 8753 33156 8809 33158
rect 8833 33156 8889 33158
rect 8913 33156 8969 33158
rect 8993 33156 9049 33158
rect 8942 32680 8998 32736
rect 9770 41384 9826 41440
rect 10046 41928 10102 41984
rect 9954 41112 10010 41168
rect 10506 42508 10508 42528
rect 10508 42508 10560 42528
rect 10560 42508 10562 42528
rect 10506 42472 10562 42508
rect 11352 43546 11408 43548
rect 11432 43546 11488 43548
rect 11512 43546 11568 43548
rect 11592 43546 11648 43548
rect 11352 43494 11398 43546
rect 11398 43494 11408 43546
rect 11432 43494 11462 43546
rect 11462 43494 11474 43546
rect 11474 43494 11488 43546
rect 11512 43494 11526 43546
rect 11526 43494 11538 43546
rect 11538 43494 11568 43546
rect 11592 43494 11602 43546
rect 11602 43494 11648 43546
rect 11352 43492 11408 43494
rect 11432 43492 11488 43494
rect 11512 43492 11568 43494
rect 11592 43492 11648 43494
rect 11150 43052 11152 43072
rect 11152 43052 11204 43072
rect 11204 43052 11206 43072
rect 11150 43016 11206 43052
rect 10690 42336 10746 42392
rect 10230 41384 10286 41440
rect 9586 38256 9642 38312
rect 9402 35944 9458 36000
rect 9402 35808 9458 35864
rect 9954 37324 10010 37360
rect 9954 37304 9956 37324
rect 9956 37304 10008 37324
rect 10008 37304 10010 37324
rect 9862 36524 9864 36544
rect 9864 36524 9916 36544
rect 9916 36524 9918 36544
rect 9862 36488 9918 36524
rect 9218 34040 9274 34096
rect 8753 32122 8809 32124
rect 8833 32122 8889 32124
rect 8913 32122 8969 32124
rect 8993 32122 9049 32124
rect 8753 32070 8799 32122
rect 8799 32070 8809 32122
rect 8833 32070 8863 32122
rect 8863 32070 8875 32122
rect 8875 32070 8889 32122
rect 8913 32070 8927 32122
rect 8927 32070 8939 32122
rect 8939 32070 8969 32122
rect 8993 32070 9003 32122
rect 9003 32070 9049 32122
rect 8753 32068 8809 32070
rect 8833 32068 8889 32070
rect 8913 32068 8969 32070
rect 8993 32068 9049 32070
rect 9402 35400 9458 35456
rect 9494 35264 9550 35320
rect 9770 35264 9826 35320
rect 9954 35808 10010 35864
rect 9678 34620 9680 34640
rect 9680 34620 9732 34640
rect 9732 34620 9734 34640
rect 9678 34584 9734 34620
rect 8753 31034 8809 31036
rect 8833 31034 8889 31036
rect 8913 31034 8969 31036
rect 8993 31034 9049 31036
rect 8753 30982 8799 31034
rect 8799 30982 8809 31034
rect 8833 30982 8863 31034
rect 8863 30982 8875 31034
rect 8875 30982 8889 31034
rect 8913 30982 8927 31034
rect 8927 30982 8939 31034
rect 8939 30982 8969 31034
rect 8993 30982 9003 31034
rect 9003 30982 9049 31034
rect 8753 30980 8809 30982
rect 8833 30980 8889 30982
rect 8913 30980 8969 30982
rect 8993 30980 9049 30982
rect 9034 30504 9090 30560
rect 8753 29946 8809 29948
rect 8833 29946 8889 29948
rect 8913 29946 8969 29948
rect 8993 29946 9049 29948
rect 8753 29894 8799 29946
rect 8799 29894 8809 29946
rect 8833 29894 8863 29946
rect 8863 29894 8875 29946
rect 8875 29894 8889 29946
rect 8913 29894 8927 29946
rect 8927 29894 8939 29946
rect 8939 29894 8969 29946
rect 8993 29894 9003 29946
rect 9003 29894 9049 29946
rect 8753 29892 8809 29894
rect 8833 29892 8889 29894
rect 8913 29892 8969 29894
rect 8993 29892 9049 29894
rect 8753 28858 8809 28860
rect 8833 28858 8889 28860
rect 8913 28858 8969 28860
rect 8993 28858 9049 28860
rect 8753 28806 8799 28858
rect 8799 28806 8809 28858
rect 8833 28806 8863 28858
rect 8863 28806 8875 28858
rect 8875 28806 8889 28858
rect 8913 28806 8927 28858
rect 8927 28806 8939 28858
rect 8939 28806 8969 28858
rect 8993 28806 9003 28858
rect 9003 28806 9049 28858
rect 8753 28804 8809 28806
rect 8833 28804 8889 28806
rect 8913 28804 8969 28806
rect 8993 28804 9049 28806
rect 8850 28192 8906 28248
rect 8942 27920 8998 27976
rect 8753 27770 8809 27772
rect 8833 27770 8889 27772
rect 8913 27770 8969 27772
rect 8993 27770 9049 27772
rect 8753 27718 8799 27770
rect 8799 27718 8809 27770
rect 8833 27718 8863 27770
rect 8863 27718 8875 27770
rect 8875 27718 8889 27770
rect 8913 27718 8927 27770
rect 8927 27718 8939 27770
rect 8939 27718 8969 27770
rect 8993 27718 9003 27770
rect 9003 27718 9049 27770
rect 8753 27716 8809 27718
rect 8833 27716 8889 27718
rect 8913 27716 8969 27718
rect 8993 27716 9049 27718
rect 9770 32272 9826 32328
rect 9586 31048 9642 31104
rect 9310 28736 9366 28792
rect 8574 27104 8630 27160
rect 8298 25336 8354 25392
rect 8206 24384 8262 24440
rect 8114 22072 8170 22128
rect 8022 21256 8078 21312
rect 8666 26988 8722 27024
rect 8666 26968 8668 26988
rect 8668 26968 8720 26988
rect 8720 26968 8722 26988
rect 8666 26832 8722 26888
rect 9126 27512 9182 27568
rect 8753 26682 8809 26684
rect 8833 26682 8889 26684
rect 8913 26682 8969 26684
rect 8993 26682 9049 26684
rect 8753 26630 8799 26682
rect 8799 26630 8809 26682
rect 8833 26630 8863 26682
rect 8863 26630 8875 26682
rect 8875 26630 8889 26682
rect 8913 26630 8927 26682
rect 8927 26630 8939 26682
rect 8939 26630 8969 26682
rect 8993 26630 9003 26682
rect 9003 26630 9049 26682
rect 8753 26628 8809 26630
rect 8833 26628 8889 26630
rect 8913 26628 8969 26630
rect 8993 26628 9049 26630
rect 9586 28328 9642 28384
rect 9494 27920 9550 27976
rect 8753 25594 8809 25596
rect 8833 25594 8889 25596
rect 8913 25594 8969 25596
rect 8993 25594 9049 25596
rect 8753 25542 8799 25594
rect 8799 25542 8809 25594
rect 8833 25542 8863 25594
rect 8863 25542 8875 25594
rect 8875 25542 8889 25594
rect 8913 25542 8927 25594
rect 8927 25542 8939 25594
rect 8939 25542 8969 25594
rect 8993 25542 9003 25594
rect 9003 25542 9049 25594
rect 8753 25540 8809 25542
rect 8833 25540 8889 25542
rect 8913 25540 8969 25542
rect 8993 25540 9049 25542
rect 8753 24506 8809 24508
rect 8833 24506 8889 24508
rect 8913 24506 8969 24508
rect 8993 24506 9049 24508
rect 8753 24454 8799 24506
rect 8799 24454 8809 24506
rect 8833 24454 8863 24506
rect 8863 24454 8875 24506
rect 8875 24454 8889 24506
rect 8913 24454 8927 24506
rect 8927 24454 8939 24506
rect 8939 24454 8969 24506
rect 8993 24454 9003 24506
rect 9003 24454 9049 24506
rect 8753 24452 8809 24454
rect 8833 24452 8889 24454
rect 8913 24452 8969 24454
rect 8993 24452 9049 24454
rect 9770 31184 9826 31240
rect 9954 34604 10010 34640
rect 10230 36624 10286 36680
rect 10322 35808 10378 35864
rect 10598 36488 10654 36544
rect 10230 35536 10286 35592
rect 10322 35128 10378 35184
rect 9954 34584 9956 34604
rect 9956 34584 10008 34604
rect 10008 34584 10010 34604
rect 9954 31764 9956 31784
rect 9956 31764 10008 31784
rect 10008 31764 10010 31784
rect 9954 31728 10010 31764
rect 9862 30232 9918 30288
rect 10414 32136 10470 32192
rect 9954 28872 10010 28928
rect 10414 30912 10470 30968
rect 10414 28872 10470 28928
rect 10046 27376 10102 27432
rect 10138 27104 10194 27160
rect 8753 23418 8809 23420
rect 8833 23418 8889 23420
rect 8913 23418 8969 23420
rect 8993 23418 9049 23420
rect 8753 23366 8799 23418
rect 8799 23366 8809 23418
rect 8833 23366 8863 23418
rect 8863 23366 8875 23418
rect 8875 23366 8889 23418
rect 8913 23366 8927 23418
rect 8927 23366 8939 23418
rect 8939 23366 8969 23418
rect 8993 23366 9003 23418
rect 9003 23366 9049 23418
rect 8753 23364 8809 23366
rect 8833 23364 8889 23366
rect 8913 23364 8969 23366
rect 8993 23364 9049 23366
rect 8390 22072 8446 22128
rect 8206 21936 8262 21992
rect 8298 21120 8354 21176
rect 8298 20168 8354 20224
rect 7838 18944 7894 19000
rect 7838 18400 7894 18456
rect 8114 16088 8170 16144
rect 7838 13640 7894 13696
rect 7746 13232 7802 13288
rect 7930 13096 7986 13152
rect 7654 12552 7710 12608
rect 7654 12416 7710 12472
rect 7654 12008 7710 12064
rect 8390 17720 8446 17776
rect 8390 15136 8446 15192
rect 8206 14592 8262 14648
rect 8298 14456 8354 14512
rect 8206 13776 8262 13832
rect 7930 11872 7986 11928
rect 8298 11636 8300 11656
rect 8300 11636 8352 11656
rect 8352 11636 8354 11656
rect 8298 11600 8354 11636
rect 7654 9580 7710 9616
rect 7654 9560 7656 9580
rect 7656 9560 7708 9580
rect 7708 9560 7710 9580
rect 7562 9424 7618 9480
rect 7654 8916 7656 8936
rect 7656 8916 7708 8936
rect 7708 8916 7710 8936
rect 7654 8880 7710 8916
rect 8022 8336 8078 8392
rect 7838 7384 7894 7440
rect 8753 22330 8809 22332
rect 8833 22330 8889 22332
rect 8913 22330 8969 22332
rect 8993 22330 9049 22332
rect 8753 22278 8799 22330
rect 8799 22278 8809 22330
rect 8833 22278 8863 22330
rect 8863 22278 8875 22330
rect 8875 22278 8889 22330
rect 8913 22278 8927 22330
rect 8927 22278 8939 22330
rect 8939 22278 8969 22330
rect 8993 22278 9003 22330
rect 9003 22278 9049 22330
rect 8753 22276 8809 22278
rect 8833 22276 8889 22278
rect 8913 22276 8969 22278
rect 8993 22276 9049 22278
rect 9310 24112 9366 24168
rect 9586 23296 9642 23352
rect 9586 22888 9642 22944
rect 9862 25900 9918 25936
rect 9862 25880 9864 25900
rect 9864 25880 9916 25900
rect 9916 25880 9918 25900
rect 9862 22924 9864 22944
rect 9864 22924 9916 22944
rect 9916 22924 9918 22944
rect 9862 22888 9918 22924
rect 9402 21936 9458 21992
rect 8753 21242 8809 21244
rect 8833 21242 8889 21244
rect 8913 21242 8969 21244
rect 8993 21242 9049 21244
rect 8753 21190 8799 21242
rect 8799 21190 8809 21242
rect 8833 21190 8863 21242
rect 8863 21190 8875 21242
rect 8875 21190 8889 21242
rect 8913 21190 8927 21242
rect 8927 21190 8939 21242
rect 8939 21190 8969 21242
rect 8993 21190 9003 21242
rect 9003 21190 9049 21242
rect 8753 21188 8809 21190
rect 8833 21188 8889 21190
rect 8913 21188 8969 21190
rect 8993 21188 9049 21190
rect 9402 21256 9458 21312
rect 9126 20984 9182 21040
rect 8753 20154 8809 20156
rect 8833 20154 8889 20156
rect 8913 20154 8969 20156
rect 8993 20154 9049 20156
rect 8753 20102 8799 20154
rect 8799 20102 8809 20154
rect 8833 20102 8863 20154
rect 8863 20102 8875 20154
rect 8875 20102 8889 20154
rect 8913 20102 8927 20154
rect 8927 20102 8939 20154
rect 8939 20102 8969 20154
rect 8993 20102 9003 20154
rect 9003 20102 9049 20154
rect 8753 20100 8809 20102
rect 8833 20100 8889 20102
rect 8913 20100 8969 20102
rect 8993 20100 9049 20102
rect 8574 17992 8630 18048
rect 8753 19066 8809 19068
rect 8833 19066 8889 19068
rect 8913 19066 8969 19068
rect 8993 19066 9049 19068
rect 8753 19014 8799 19066
rect 8799 19014 8809 19066
rect 8833 19014 8863 19066
rect 8863 19014 8875 19066
rect 8875 19014 8889 19066
rect 8913 19014 8927 19066
rect 8927 19014 8939 19066
rect 8939 19014 8969 19066
rect 8993 19014 9003 19066
rect 9003 19014 9049 19066
rect 8753 19012 8809 19014
rect 8833 19012 8889 19014
rect 8913 19012 8969 19014
rect 8993 19012 9049 19014
rect 9402 19896 9458 19952
rect 9310 19760 9366 19816
rect 8753 17978 8809 17980
rect 8833 17978 8889 17980
rect 8913 17978 8969 17980
rect 8993 17978 9049 17980
rect 8753 17926 8799 17978
rect 8799 17926 8809 17978
rect 8833 17926 8863 17978
rect 8863 17926 8875 17978
rect 8875 17926 8889 17978
rect 8913 17926 8927 17978
rect 8927 17926 8939 17978
rect 8939 17926 8969 17978
rect 8993 17926 9003 17978
rect 9003 17926 9049 17978
rect 8753 17924 8809 17926
rect 8833 17924 8889 17926
rect 8913 17924 8969 17926
rect 8993 17924 9049 17926
rect 8574 17584 8630 17640
rect 8758 17484 8760 17504
rect 8760 17484 8812 17504
rect 8812 17484 8814 17504
rect 8758 17448 8814 17484
rect 8753 16890 8809 16892
rect 8833 16890 8889 16892
rect 8913 16890 8969 16892
rect 8993 16890 9049 16892
rect 8753 16838 8799 16890
rect 8799 16838 8809 16890
rect 8833 16838 8863 16890
rect 8863 16838 8875 16890
rect 8875 16838 8889 16890
rect 8913 16838 8927 16890
rect 8927 16838 8939 16890
rect 8939 16838 8969 16890
rect 8993 16838 9003 16890
rect 9003 16838 9049 16890
rect 8753 16836 8809 16838
rect 8833 16836 8889 16838
rect 8913 16836 8969 16838
rect 8993 16836 9049 16838
rect 9218 17856 9274 17912
rect 9494 19624 9550 19680
rect 10046 23976 10102 24032
rect 10046 22888 10102 22944
rect 9954 21684 10010 21720
rect 9954 21664 9956 21684
rect 9956 21664 10008 21684
rect 10008 21664 10010 21684
rect 9770 19488 9826 19544
rect 9770 19080 9826 19136
rect 9586 17720 9642 17776
rect 9126 16088 9182 16144
rect 8753 15802 8809 15804
rect 8833 15802 8889 15804
rect 8913 15802 8969 15804
rect 8993 15802 9049 15804
rect 8753 15750 8799 15802
rect 8799 15750 8809 15802
rect 8833 15750 8863 15802
rect 8863 15750 8875 15802
rect 8875 15750 8889 15802
rect 8913 15750 8927 15802
rect 8927 15750 8939 15802
rect 8939 15750 8969 15802
rect 8993 15750 9003 15802
rect 9003 15750 9049 15802
rect 8753 15748 8809 15750
rect 8833 15748 8889 15750
rect 8913 15748 8969 15750
rect 8993 15748 9049 15750
rect 9126 15000 9182 15056
rect 8753 14714 8809 14716
rect 8833 14714 8889 14716
rect 8913 14714 8969 14716
rect 8993 14714 9049 14716
rect 8753 14662 8799 14714
rect 8799 14662 8809 14714
rect 8833 14662 8863 14714
rect 8863 14662 8875 14714
rect 8875 14662 8889 14714
rect 8913 14662 8927 14714
rect 8927 14662 8939 14714
rect 8939 14662 8969 14714
rect 8993 14662 9003 14714
rect 9003 14662 9049 14714
rect 8753 14660 8809 14662
rect 8833 14660 8889 14662
rect 8913 14660 8969 14662
rect 8993 14660 9049 14662
rect 8574 8628 8630 8664
rect 8574 8608 8576 8628
rect 8576 8608 8628 8628
rect 8628 8608 8630 8628
rect 8390 7964 8392 7984
rect 8392 7964 8444 7984
rect 8444 7964 8446 7984
rect 8390 7928 8446 7964
rect 7746 6976 7802 7032
rect 7838 6568 7894 6624
rect 8753 13626 8809 13628
rect 8833 13626 8889 13628
rect 8913 13626 8969 13628
rect 8993 13626 9049 13628
rect 8753 13574 8799 13626
rect 8799 13574 8809 13626
rect 8833 13574 8863 13626
rect 8863 13574 8875 13626
rect 8875 13574 8889 13626
rect 8913 13574 8927 13626
rect 8927 13574 8939 13626
rect 8939 13574 8969 13626
rect 8993 13574 9003 13626
rect 9003 13574 9049 13626
rect 8753 13572 8809 13574
rect 8833 13572 8889 13574
rect 8913 13572 8969 13574
rect 8993 13572 9049 13574
rect 9034 12688 9090 12744
rect 8753 12538 8809 12540
rect 8833 12538 8889 12540
rect 8913 12538 8969 12540
rect 8993 12538 9049 12540
rect 8753 12486 8799 12538
rect 8799 12486 8809 12538
rect 8833 12486 8863 12538
rect 8863 12486 8875 12538
rect 8875 12486 8889 12538
rect 8913 12486 8927 12538
rect 8927 12486 8939 12538
rect 8939 12486 8969 12538
rect 8993 12486 9003 12538
rect 9003 12486 9049 12538
rect 8753 12484 8809 12486
rect 8833 12484 8889 12486
rect 8913 12484 8969 12486
rect 8993 12484 9049 12486
rect 8753 11450 8809 11452
rect 8833 11450 8889 11452
rect 8913 11450 8969 11452
rect 8993 11450 9049 11452
rect 8753 11398 8799 11450
rect 8799 11398 8809 11450
rect 8833 11398 8863 11450
rect 8863 11398 8875 11450
rect 8875 11398 8889 11450
rect 8913 11398 8927 11450
rect 8927 11398 8939 11450
rect 8939 11398 8969 11450
rect 8993 11398 9003 11450
rect 9003 11398 9049 11450
rect 8753 11396 8809 11398
rect 8833 11396 8889 11398
rect 8913 11396 8969 11398
rect 8993 11396 9049 11398
rect 8753 10362 8809 10364
rect 8833 10362 8889 10364
rect 8913 10362 8969 10364
rect 8993 10362 9049 10364
rect 8753 10310 8799 10362
rect 8799 10310 8809 10362
rect 8833 10310 8863 10362
rect 8863 10310 8875 10362
rect 8875 10310 8889 10362
rect 8913 10310 8927 10362
rect 8927 10310 8939 10362
rect 8939 10310 8969 10362
rect 8993 10310 9003 10362
rect 9003 10310 9049 10362
rect 8753 10308 8809 10310
rect 8833 10308 8889 10310
rect 8913 10308 8969 10310
rect 8993 10308 9049 10310
rect 8758 9696 8814 9752
rect 8753 9274 8809 9276
rect 8833 9274 8889 9276
rect 8913 9274 8969 9276
rect 8993 9274 9049 9276
rect 8753 9222 8799 9274
rect 8799 9222 8809 9274
rect 8833 9222 8863 9274
rect 8863 9222 8875 9274
rect 8875 9222 8889 9274
rect 8913 9222 8927 9274
rect 8927 9222 8939 9274
rect 8939 9222 8969 9274
rect 8993 9222 9003 9274
rect 9003 9222 9049 9274
rect 8753 9220 8809 9222
rect 8833 9220 8889 9222
rect 8913 9220 8969 9222
rect 8993 9220 9049 9222
rect 8753 8186 8809 8188
rect 8833 8186 8889 8188
rect 8913 8186 8969 8188
rect 8993 8186 9049 8188
rect 8753 8134 8799 8186
rect 8799 8134 8809 8186
rect 8833 8134 8863 8186
rect 8863 8134 8875 8186
rect 8875 8134 8889 8186
rect 8913 8134 8927 8186
rect 8927 8134 8939 8186
rect 8939 8134 8969 8186
rect 8993 8134 9003 8186
rect 9003 8134 9049 8186
rect 8753 8132 8809 8134
rect 8833 8132 8889 8134
rect 8913 8132 8969 8134
rect 8993 8132 9049 8134
rect 8850 7792 8906 7848
rect 8758 7656 8814 7712
rect 8390 6024 8446 6080
rect 7470 3984 7526 4040
rect 7286 3848 7342 3904
rect 7010 1808 7066 1864
rect 7194 2644 7250 2680
rect 7194 2624 7196 2644
rect 7196 2624 7248 2644
rect 7248 2624 7250 2644
rect 7194 1400 7250 1456
rect 7378 1300 7380 1320
rect 7380 1300 7432 1320
rect 7432 1300 7434 1320
rect 7378 1264 7434 1300
rect 7930 2644 7986 2680
rect 7930 2624 7932 2644
rect 7932 2624 7984 2644
rect 7984 2624 7986 2644
rect 7654 1808 7710 1864
rect 8753 7098 8809 7100
rect 8833 7098 8889 7100
rect 8913 7098 8969 7100
rect 8993 7098 9049 7100
rect 8753 7046 8799 7098
rect 8799 7046 8809 7098
rect 8833 7046 8863 7098
rect 8863 7046 8875 7098
rect 8875 7046 8889 7098
rect 8913 7046 8927 7098
rect 8927 7046 8939 7098
rect 8939 7046 8969 7098
rect 8993 7046 9003 7098
rect 9003 7046 9049 7098
rect 8753 7044 8809 7046
rect 8833 7044 8889 7046
rect 8913 7044 8969 7046
rect 8993 7044 9049 7046
rect 8753 6010 8809 6012
rect 8833 6010 8889 6012
rect 8913 6010 8969 6012
rect 8993 6010 9049 6012
rect 8753 5958 8799 6010
rect 8799 5958 8809 6010
rect 8833 5958 8863 6010
rect 8863 5958 8875 6010
rect 8875 5958 8889 6010
rect 8913 5958 8927 6010
rect 8927 5958 8939 6010
rect 8939 5958 8969 6010
rect 8993 5958 9003 6010
rect 9003 5958 9049 6010
rect 8753 5956 8809 5958
rect 8833 5956 8889 5958
rect 8913 5956 8969 5958
rect 8993 5956 9049 5958
rect 8942 5616 8998 5672
rect 8753 4922 8809 4924
rect 8833 4922 8889 4924
rect 8913 4922 8969 4924
rect 8993 4922 9049 4924
rect 8753 4870 8799 4922
rect 8799 4870 8809 4922
rect 8833 4870 8863 4922
rect 8863 4870 8875 4922
rect 8875 4870 8889 4922
rect 8913 4870 8927 4922
rect 8927 4870 8939 4922
rect 8939 4870 8969 4922
rect 8993 4870 9003 4922
rect 9003 4870 9049 4922
rect 8753 4868 8809 4870
rect 8833 4868 8889 4870
rect 8913 4868 8969 4870
rect 8993 4868 9049 4870
rect 9218 4664 9274 4720
rect 8753 3834 8809 3836
rect 8833 3834 8889 3836
rect 8913 3834 8969 3836
rect 8993 3834 9049 3836
rect 8753 3782 8799 3834
rect 8799 3782 8809 3834
rect 8833 3782 8863 3834
rect 8863 3782 8875 3834
rect 8875 3782 8889 3834
rect 8913 3782 8927 3834
rect 8927 3782 8939 3834
rect 8939 3782 8969 3834
rect 8993 3782 9003 3834
rect 9003 3782 9049 3834
rect 8753 3780 8809 3782
rect 8833 3780 8889 3782
rect 8913 3780 8969 3782
rect 8993 3780 9049 3782
rect 9678 16496 9734 16552
rect 9586 15816 9642 15872
rect 9586 13504 9642 13560
rect 10046 20168 10102 20224
rect 9954 18536 10010 18592
rect 10322 24248 10378 24304
rect 10322 23840 10378 23896
rect 10322 22344 10378 22400
rect 10322 21292 10324 21312
rect 10324 21292 10376 21312
rect 10376 21292 10378 21312
rect 10322 21256 10378 21292
rect 10874 42472 10930 42528
rect 11352 42458 11408 42460
rect 11432 42458 11488 42460
rect 11512 42458 11568 42460
rect 11592 42458 11648 42460
rect 11352 42406 11398 42458
rect 11398 42406 11408 42458
rect 11432 42406 11462 42458
rect 11462 42406 11474 42458
rect 11474 42406 11488 42458
rect 11512 42406 11526 42458
rect 11526 42406 11538 42458
rect 11538 42406 11568 42458
rect 11592 42406 11602 42458
rect 11602 42406 11648 42458
rect 11352 42404 11408 42406
rect 11432 42404 11488 42406
rect 11512 42404 11568 42406
rect 11592 42404 11648 42406
rect 11150 42200 11206 42256
rect 12070 43152 12126 43208
rect 11352 41370 11408 41372
rect 11432 41370 11488 41372
rect 11512 41370 11568 41372
rect 11592 41370 11648 41372
rect 11352 41318 11398 41370
rect 11398 41318 11408 41370
rect 11432 41318 11462 41370
rect 11462 41318 11474 41370
rect 11474 41318 11488 41370
rect 11512 41318 11526 41370
rect 11526 41318 11538 41370
rect 11538 41318 11568 41370
rect 11592 41318 11602 41370
rect 11602 41318 11648 41370
rect 11352 41316 11408 41318
rect 11432 41316 11488 41318
rect 11512 41316 11568 41318
rect 11592 41316 11648 41318
rect 11058 38392 11114 38448
rect 11352 40282 11408 40284
rect 11432 40282 11488 40284
rect 11512 40282 11568 40284
rect 11592 40282 11648 40284
rect 11352 40230 11398 40282
rect 11398 40230 11408 40282
rect 11432 40230 11462 40282
rect 11462 40230 11474 40282
rect 11474 40230 11488 40282
rect 11512 40230 11526 40282
rect 11526 40230 11538 40282
rect 11538 40230 11568 40282
rect 11592 40230 11602 40282
rect 11602 40230 11648 40282
rect 11352 40228 11408 40230
rect 11432 40228 11488 40230
rect 11512 40228 11568 40230
rect 11592 40228 11648 40230
rect 11352 39194 11408 39196
rect 11432 39194 11488 39196
rect 11512 39194 11568 39196
rect 11592 39194 11648 39196
rect 11352 39142 11398 39194
rect 11398 39142 11408 39194
rect 11432 39142 11462 39194
rect 11462 39142 11474 39194
rect 11474 39142 11488 39194
rect 11512 39142 11526 39194
rect 11526 39142 11538 39194
rect 11538 39142 11568 39194
rect 11592 39142 11602 39194
rect 11602 39142 11648 39194
rect 11352 39140 11408 39142
rect 11432 39140 11488 39142
rect 11512 39140 11568 39142
rect 11592 39140 11648 39142
rect 10966 35944 11022 36000
rect 10874 35128 10930 35184
rect 10874 34448 10930 34504
rect 11352 38106 11408 38108
rect 11432 38106 11488 38108
rect 11512 38106 11568 38108
rect 11592 38106 11648 38108
rect 11352 38054 11398 38106
rect 11398 38054 11408 38106
rect 11432 38054 11462 38106
rect 11462 38054 11474 38106
rect 11474 38054 11488 38106
rect 11512 38054 11526 38106
rect 11526 38054 11538 38106
rect 11538 38054 11568 38106
rect 11592 38054 11602 38106
rect 11602 38054 11648 38106
rect 11352 38052 11408 38054
rect 11432 38052 11488 38054
rect 11512 38052 11568 38054
rect 11592 38052 11648 38054
rect 11334 37168 11390 37224
rect 11352 37018 11408 37020
rect 11432 37018 11488 37020
rect 11512 37018 11568 37020
rect 11592 37018 11648 37020
rect 11352 36966 11398 37018
rect 11398 36966 11408 37018
rect 11432 36966 11462 37018
rect 11462 36966 11474 37018
rect 11474 36966 11488 37018
rect 11512 36966 11526 37018
rect 11526 36966 11538 37018
rect 11538 36966 11568 37018
rect 11592 36966 11602 37018
rect 11602 36966 11648 37018
rect 11352 36964 11408 36966
rect 11432 36964 11488 36966
rect 11512 36964 11568 36966
rect 11592 36964 11648 36966
rect 11352 35930 11408 35932
rect 11432 35930 11488 35932
rect 11512 35930 11568 35932
rect 11592 35930 11648 35932
rect 11352 35878 11398 35930
rect 11398 35878 11408 35930
rect 11432 35878 11462 35930
rect 11462 35878 11474 35930
rect 11474 35878 11488 35930
rect 11512 35878 11526 35930
rect 11526 35878 11538 35930
rect 11538 35878 11568 35930
rect 11592 35878 11602 35930
rect 11602 35878 11648 35930
rect 11352 35876 11408 35878
rect 11432 35876 11488 35878
rect 11512 35876 11568 35878
rect 11592 35876 11648 35878
rect 11610 35672 11666 35728
rect 10782 33360 10838 33416
rect 11352 34842 11408 34844
rect 11432 34842 11488 34844
rect 11512 34842 11568 34844
rect 11592 34842 11648 34844
rect 11352 34790 11398 34842
rect 11398 34790 11408 34842
rect 11432 34790 11462 34842
rect 11462 34790 11474 34842
rect 11474 34790 11488 34842
rect 11512 34790 11526 34842
rect 11526 34790 11538 34842
rect 11538 34790 11568 34842
rect 11592 34790 11602 34842
rect 11602 34790 11648 34842
rect 11352 34788 11408 34790
rect 11432 34788 11488 34790
rect 11512 34788 11568 34790
rect 11592 34788 11648 34790
rect 11242 33904 11298 33960
rect 11794 34584 11850 34640
rect 11702 34040 11758 34096
rect 11886 34040 11942 34096
rect 11352 33754 11408 33756
rect 11432 33754 11488 33756
rect 11512 33754 11568 33756
rect 11592 33754 11648 33756
rect 11352 33702 11398 33754
rect 11398 33702 11408 33754
rect 11432 33702 11462 33754
rect 11462 33702 11474 33754
rect 11474 33702 11488 33754
rect 11512 33702 11526 33754
rect 11526 33702 11538 33754
rect 11538 33702 11568 33754
rect 11592 33702 11602 33754
rect 11602 33702 11648 33754
rect 11352 33700 11408 33702
rect 11432 33700 11488 33702
rect 11512 33700 11568 33702
rect 11592 33700 11648 33702
rect 11794 33632 11850 33688
rect 11058 33360 11114 33416
rect 10690 32428 10746 32464
rect 10690 32408 10692 32428
rect 10692 32408 10744 32428
rect 10744 32408 10746 32428
rect 11058 32680 11114 32736
rect 10966 32272 11022 32328
rect 11794 33088 11850 33144
rect 11352 32666 11408 32668
rect 11432 32666 11488 32668
rect 11512 32666 11568 32668
rect 11592 32666 11648 32668
rect 11352 32614 11398 32666
rect 11398 32614 11408 32666
rect 11432 32614 11462 32666
rect 11462 32614 11474 32666
rect 11474 32614 11488 32666
rect 11512 32614 11526 32666
rect 11526 32614 11538 32666
rect 11538 32614 11568 32666
rect 11592 32614 11602 32666
rect 11602 32614 11648 32666
rect 11352 32612 11408 32614
rect 11432 32612 11488 32614
rect 11512 32612 11568 32614
rect 11592 32612 11648 32614
rect 10966 30368 11022 30424
rect 10782 29552 10838 29608
rect 10874 28192 10930 28248
rect 11058 28736 11114 28792
rect 10598 24656 10654 24712
rect 10506 23840 10562 23896
rect 10874 26324 10876 26344
rect 10876 26324 10928 26344
rect 10928 26324 10930 26344
rect 10874 26288 10930 26324
rect 10782 25880 10838 25936
rect 10230 18808 10286 18864
rect 9954 17448 10010 17504
rect 9770 13776 9826 13832
rect 10690 20304 10746 20360
rect 10690 17992 10746 18048
rect 10506 16632 10562 16688
rect 9862 12960 9918 13016
rect 9494 12044 9496 12064
rect 9496 12044 9548 12064
rect 9548 12044 9550 12064
rect 9494 12008 9550 12044
rect 9862 12688 9918 12744
rect 9862 11192 9918 11248
rect 9494 10512 9550 10568
rect 10230 12960 10286 13016
rect 10230 12824 10286 12880
rect 10690 16768 10746 16824
rect 11352 31578 11408 31580
rect 11432 31578 11488 31580
rect 11512 31578 11568 31580
rect 11592 31578 11648 31580
rect 11352 31526 11398 31578
rect 11398 31526 11408 31578
rect 11432 31526 11462 31578
rect 11462 31526 11474 31578
rect 11474 31526 11488 31578
rect 11512 31526 11526 31578
rect 11526 31526 11538 31578
rect 11538 31526 11568 31578
rect 11592 31526 11602 31578
rect 11602 31526 11648 31578
rect 11352 31524 11408 31526
rect 11432 31524 11488 31526
rect 11512 31524 11568 31526
rect 11592 31524 11648 31526
rect 11886 32680 11942 32736
rect 11886 32272 11942 32328
rect 11702 31320 11758 31376
rect 11352 30490 11408 30492
rect 11432 30490 11488 30492
rect 11512 30490 11568 30492
rect 11592 30490 11648 30492
rect 11352 30438 11398 30490
rect 11398 30438 11408 30490
rect 11432 30438 11462 30490
rect 11462 30438 11474 30490
rect 11474 30438 11488 30490
rect 11512 30438 11526 30490
rect 11526 30438 11538 30490
rect 11538 30438 11568 30490
rect 11592 30438 11602 30490
rect 11602 30438 11648 30490
rect 11352 30436 11408 30438
rect 11432 30436 11488 30438
rect 11512 30436 11568 30438
rect 11592 30436 11648 30438
rect 11610 30252 11666 30288
rect 11610 30232 11612 30252
rect 11612 30232 11664 30252
rect 11664 30232 11666 30252
rect 11794 31048 11850 31104
rect 11334 29824 11390 29880
rect 11794 29416 11850 29472
rect 11352 29402 11408 29404
rect 11432 29402 11488 29404
rect 11512 29402 11568 29404
rect 11592 29402 11648 29404
rect 11352 29350 11398 29402
rect 11398 29350 11408 29402
rect 11432 29350 11462 29402
rect 11462 29350 11474 29402
rect 11474 29350 11488 29402
rect 11512 29350 11526 29402
rect 11526 29350 11538 29402
rect 11538 29350 11568 29402
rect 11592 29350 11602 29402
rect 11602 29350 11648 29402
rect 11352 29348 11408 29350
rect 11432 29348 11488 29350
rect 11512 29348 11568 29350
rect 11592 29348 11648 29350
rect 11702 29144 11758 29200
rect 11352 28314 11408 28316
rect 11432 28314 11488 28316
rect 11512 28314 11568 28316
rect 11592 28314 11648 28316
rect 11352 28262 11398 28314
rect 11398 28262 11408 28314
rect 11432 28262 11462 28314
rect 11462 28262 11474 28314
rect 11474 28262 11488 28314
rect 11512 28262 11526 28314
rect 11526 28262 11538 28314
rect 11538 28262 11568 28314
rect 11592 28262 11602 28314
rect 11602 28262 11648 28314
rect 11352 28260 11408 28262
rect 11432 28260 11488 28262
rect 11512 28260 11568 28262
rect 11592 28260 11648 28262
rect 11610 27920 11666 27976
rect 11352 27226 11408 27228
rect 11432 27226 11488 27228
rect 11512 27226 11568 27228
rect 11592 27226 11648 27228
rect 11352 27174 11398 27226
rect 11398 27174 11408 27226
rect 11432 27174 11462 27226
rect 11462 27174 11474 27226
rect 11474 27174 11488 27226
rect 11512 27174 11526 27226
rect 11526 27174 11538 27226
rect 11538 27174 11568 27226
rect 11592 27174 11602 27226
rect 11602 27174 11648 27226
rect 11352 27172 11408 27174
rect 11432 27172 11488 27174
rect 11512 27172 11568 27174
rect 11592 27172 11648 27174
rect 11352 26138 11408 26140
rect 11432 26138 11488 26140
rect 11512 26138 11568 26140
rect 11592 26138 11648 26140
rect 11352 26086 11398 26138
rect 11398 26086 11408 26138
rect 11432 26086 11462 26138
rect 11462 26086 11474 26138
rect 11474 26086 11488 26138
rect 11512 26086 11526 26138
rect 11526 26086 11538 26138
rect 11538 26086 11568 26138
rect 11592 26086 11602 26138
rect 11602 26086 11648 26138
rect 11352 26084 11408 26086
rect 11432 26084 11488 26086
rect 11512 26084 11568 26086
rect 11592 26084 11648 26086
rect 11352 25050 11408 25052
rect 11432 25050 11488 25052
rect 11512 25050 11568 25052
rect 11592 25050 11648 25052
rect 11352 24998 11398 25050
rect 11398 24998 11408 25050
rect 11432 24998 11462 25050
rect 11462 24998 11474 25050
rect 11474 24998 11488 25050
rect 11512 24998 11526 25050
rect 11526 24998 11538 25050
rect 11538 24998 11568 25050
rect 11592 24998 11602 25050
rect 11602 24998 11648 25050
rect 11352 24996 11408 24998
rect 11432 24996 11488 24998
rect 11512 24996 11568 24998
rect 11592 24996 11648 24998
rect 13082 42880 13138 42936
rect 13450 43172 13506 43208
rect 13450 43152 13452 43172
rect 13452 43152 13504 43172
rect 13504 43152 13506 43172
rect 12254 41520 12310 41576
rect 12162 37168 12218 37224
rect 12070 32544 12126 32600
rect 12162 32408 12218 32464
rect 11702 24792 11758 24848
rect 11352 23962 11408 23964
rect 11432 23962 11488 23964
rect 11512 23962 11568 23964
rect 11592 23962 11648 23964
rect 11352 23910 11398 23962
rect 11398 23910 11408 23962
rect 11432 23910 11462 23962
rect 11462 23910 11474 23962
rect 11474 23910 11488 23962
rect 11512 23910 11526 23962
rect 11526 23910 11538 23962
rect 11538 23910 11568 23962
rect 11592 23910 11602 23962
rect 11602 23910 11648 23962
rect 11352 23908 11408 23910
rect 11432 23908 11488 23910
rect 11512 23908 11568 23910
rect 11592 23908 11648 23910
rect 10874 23432 10930 23488
rect 11426 23568 11482 23624
rect 10966 22652 10968 22672
rect 10968 22652 11020 22672
rect 11020 22652 11022 22672
rect 10966 22616 11022 22652
rect 11150 22888 11206 22944
rect 11150 22752 11206 22808
rect 11352 22874 11408 22876
rect 11432 22874 11488 22876
rect 11512 22874 11568 22876
rect 11592 22874 11648 22876
rect 11352 22822 11398 22874
rect 11398 22822 11408 22874
rect 11432 22822 11462 22874
rect 11462 22822 11474 22874
rect 11474 22822 11488 22874
rect 11512 22822 11526 22874
rect 11526 22822 11538 22874
rect 11538 22822 11568 22874
rect 11592 22822 11602 22874
rect 11602 22822 11648 22874
rect 11352 22820 11408 22822
rect 11432 22820 11488 22822
rect 11512 22820 11568 22822
rect 11592 22820 11648 22822
rect 10966 22344 11022 22400
rect 11150 22208 11206 22264
rect 11886 25336 11942 25392
rect 11352 21786 11408 21788
rect 11432 21786 11488 21788
rect 11512 21786 11568 21788
rect 11592 21786 11648 21788
rect 11352 21734 11398 21786
rect 11398 21734 11408 21786
rect 11432 21734 11462 21786
rect 11462 21734 11474 21786
rect 11474 21734 11488 21786
rect 11512 21734 11526 21786
rect 11526 21734 11538 21786
rect 11538 21734 11568 21786
rect 11592 21734 11602 21786
rect 11602 21734 11648 21786
rect 11352 21732 11408 21734
rect 11432 21732 11488 21734
rect 11512 21732 11568 21734
rect 11592 21732 11648 21734
rect 10966 20848 11022 20904
rect 11426 21392 11482 21448
rect 11058 20712 11114 20768
rect 11058 20576 11114 20632
rect 11794 21120 11850 21176
rect 11352 20698 11408 20700
rect 11432 20698 11488 20700
rect 11512 20698 11568 20700
rect 11592 20698 11648 20700
rect 11352 20646 11398 20698
rect 11398 20646 11408 20698
rect 11432 20646 11462 20698
rect 11462 20646 11474 20698
rect 11474 20646 11488 20698
rect 11512 20646 11526 20698
rect 11526 20646 11538 20698
rect 11538 20646 11568 20698
rect 11592 20646 11602 20698
rect 11602 20646 11648 20698
rect 11352 20644 11408 20646
rect 11432 20644 11488 20646
rect 11512 20644 11568 20646
rect 11592 20644 11648 20646
rect 11426 20304 11482 20360
rect 10874 18672 10930 18728
rect 11242 19760 11298 19816
rect 11058 19488 11114 19544
rect 11150 18128 11206 18184
rect 10966 16768 11022 16824
rect 11352 19610 11408 19612
rect 11432 19610 11488 19612
rect 11512 19610 11568 19612
rect 11592 19610 11648 19612
rect 11352 19558 11398 19610
rect 11398 19558 11408 19610
rect 11432 19558 11462 19610
rect 11462 19558 11474 19610
rect 11474 19558 11488 19610
rect 11512 19558 11526 19610
rect 11526 19558 11538 19610
rect 11538 19558 11568 19610
rect 11592 19558 11602 19610
rect 11602 19558 11648 19610
rect 11352 19556 11408 19558
rect 11432 19556 11488 19558
rect 11512 19556 11568 19558
rect 11592 19556 11648 19558
rect 11702 19352 11758 19408
rect 11610 18672 11666 18728
rect 11352 18522 11408 18524
rect 11432 18522 11488 18524
rect 11512 18522 11568 18524
rect 11592 18522 11648 18524
rect 11352 18470 11398 18522
rect 11398 18470 11408 18522
rect 11432 18470 11462 18522
rect 11462 18470 11474 18522
rect 11474 18470 11488 18522
rect 11512 18470 11526 18522
rect 11526 18470 11538 18522
rect 11538 18470 11568 18522
rect 11592 18470 11602 18522
rect 11602 18470 11648 18522
rect 11352 18468 11408 18470
rect 11432 18468 11488 18470
rect 11512 18468 11568 18470
rect 11592 18468 11648 18470
rect 11886 18808 11942 18864
rect 11886 18400 11942 18456
rect 11242 17584 11298 17640
rect 11352 17434 11408 17436
rect 11432 17434 11488 17436
rect 11512 17434 11568 17436
rect 11592 17434 11648 17436
rect 11352 17382 11398 17434
rect 11398 17382 11408 17434
rect 11432 17382 11462 17434
rect 11462 17382 11474 17434
rect 11474 17382 11488 17434
rect 11512 17382 11526 17434
rect 11526 17382 11538 17434
rect 11538 17382 11568 17434
rect 11592 17382 11602 17434
rect 11602 17382 11648 17434
rect 11352 17380 11408 17382
rect 11432 17380 11488 17382
rect 11512 17380 11568 17382
rect 11592 17380 11648 17382
rect 11150 17312 11206 17368
rect 11150 17040 11206 17096
rect 11058 16224 11114 16280
rect 12254 30504 12310 30560
rect 12254 29844 12310 29880
rect 12254 29824 12256 29844
rect 12256 29824 12308 29844
rect 12308 29824 12310 29844
rect 12438 42064 12494 42120
rect 12530 36216 12586 36272
rect 12530 32852 12532 32872
rect 12532 32852 12584 32872
rect 12584 32852 12586 32872
rect 12530 32816 12586 32852
rect 13082 37324 13138 37360
rect 13082 37304 13084 37324
rect 13084 37304 13136 37324
rect 13136 37304 13138 37324
rect 13082 35536 13138 35592
rect 14002 43832 14058 43888
rect 13910 43288 13966 43344
rect 13951 43002 14007 43004
rect 14031 43002 14087 43004
rect 14111 43002 14167 43004
rect 14191 43002 14247 43004
rect 13951 42950 13997 43002
rect 13997 42950 14007 43002
rect 14031 42950 14061 43002
rect 14061 42950 14073 43002
rect 14073 42950 14087 43002
rect 14111 42950 14125 43002
rect 14125 42950 14137 43002
rect 14137 42950 14167 43002
rect 14191 42950 14201 43002
rect 14201 42950 14247 43002
rect 13951 42948 14007 42950
rect 14031 42948 14087 42950
rect 14111 42948 14167 42950
rect 14191 42948 14247 42950
rect 14002 42064 14058 42120
rect 13951 41914 14007 41916
rect 14031 41914 14087 41916
rect 14111 41914 14167 41916
rect 14191 41914 14247 41916
rect 13951 41862 13997 41914
rect 13997 41862 14007 41914
rect 14031 41862 14061 41914
rect 14061 41862 14073 41914
rect 14073 41862 14087 41914
rect 14111 41862 14125 41914
rect 14125 41862 14137 41914
rect 14137 41862 14167 41914
rect 14191 41862 14201 41914
rect 14201 41862 14247 41914
rect 13951 41860 14007 41862
rect 14031 41860 14087 41862
rect 14111 41860 14167 41862
rect 14191 41860 14247 41862
rect 14186 41656 14242 41712
rect 12990 33496 13046 33552
rect 13174 32272 13230 32328
rect 13174 32000 13230 32056
rect 12438 30776 12494 30832
rect 12346 29416 12402 29472
rect 12162 27240 12218 27296
rect 12070 18672 12126 18728
rect 11352 16346 11408 16348
rect 11432 16346 11488 16348
rect 11512 16346 11568 16348
rect 11592 16346 11648 16348
rect 11352 16294 11398 16346
rect 11398 16294 11408 16346
rect 11432 16294 11462 16346
rect 11462 16294 11474 16346
rect 11474 16294 11488 16346
rect 11512 16294 11526 16346
rect 11526 16294 11538 16346
rect 11538 16294 11568 16346
rect 11592 16294 11602 16346
rect 11602 16294 11648 16346
rect 11352 16292 11408 16294
rect 11432 16292 11488 16294
rect 11512 16292 11568 16294
rect 11592 16292 11648 16294
rect 11352 15258 11408 15260
rect 11432 15258 11488 15260
rect 11512 15258 11568 15260
rect 11592 15258 11648 15260
rect 11352 15206 11398 15258
rect 11398 15206 11408 15258
rect 11432 15206 11462 15258
rect 11462 15206 11474 15258
rect 11474 15206 11488 15258
rect 11512 15206 11526 15258
rect 11526 15206 11538 15258
rect 11538 15206 11568 15258
rect 11592 15206 11602 15258
rect 11602 15206 11648 15258
rect 11352 15204 11408 15206
rect 11432 15204 11488 15206
rect 11512 15204 11568 15206
rect 11592 15204 11648 15206
rect 10782 14456 10838 14512
rect 11352 14170 11408 14172
rect 11432 14170 11488 14172
rect 11512 14170 11568 14172
rect 11592 14170 11648 14172
rect 11352 14118 11398 14170
rect 11398 14118 11408 14170
rect 11432 14118 11462 14170
rect 11462 14118 11474 14170
rect 11474 14118 11488 14170
rect 11512 14118 11526 14170
rect 11526 14118 11538 14170
rect 11538 14118 11568 14170
rect 11592 14118 11602 14170
rect 11602 14118 11648 14170
rect 11352 14116 11408 14118
rect 11432 14116 11488 14118
rect 11512 14116 11568 14118
rect 11592 14116 11648 14118
rect 10598 12960 10654 13016
rect 10322 12688 10378 12744
rect 10322 11872 10378 11928
rect 9586 8336 9642 8392
rect 9494 7792 9550 7848
rect 8206 2896 8262 2952
rect 8206 2216 8262 2272
rect 8206 1400 8262 1456
rect 8758 3168 8814 3224
rect 9218 3168 9274 3224
rect 8574 3032 8630 3088
rect 8753 2746 8809 2748
rect 8833 2746 8889 2748
rect 8913 2746 8969 2748
rect 8993 2746 9049 2748
rect 8753 2694 8799 2746
rect 8799 2694 8809 2746
rect 8833 2694 8863 2746
rect 8863 2694 8875 2746
rect 8875 2694 8889 2746
rect 8913 2694 8927 2746
rect 8927 2694 8939 2746
rect 8939 2694 8969 2746
rect 8993 2694 9003 2746
rect 9003 2694 9049 2746
rect 8753 2692 8809 2694
rect 8833 2692 8889 2694
rect 8913 2692 8969 2694
rect 8993 2692 9049 2694
rect 8758 2488 8814 2544
rect 8753 1658 8809 1660
rect 8833 1658 8889 1660
rect 8913 1658 8969 1660
rect 8993 1658 9049 1660
rect 8753 1606 8799 1658
rect 8799 1606 8809 1658
rect 8833 1606 8863 1658
rect 8863 1606 8875 1658
rect 8875 1606 8889 1658
rect 8913 1606 8927 1658
rect 8927 1606 8939 1658
rect 8939 1606 8969 1658
rect 8993 1606 9003 1658
rect 9003 1606 9049 1658
rect 8753 1604 8809 1606
rect 8833 1604 8889 1606
rect 8913 1604 8969 1606
rect 8993 1604 9049 1606
rect 9494 3052 9550 3088
rect 9494 3032 9496 3052
rect 9496 3032 9548 3052
rect 9548 3032 9550 3052
rect 9402 1400 9458 1456
rect 9770 6024 9826 6080
rect 10046 9016 10102 9072
rect 10046 8608 10102 8664
rect 10506 9716 10562 9752
rect 10506 9696 10508 9716
rect 10508 9696 10560 9716
rect 10560 9696 10562 9716
rect 11150 12960 11206 13016
rect 11058 12144 11114 12200
rect 11352 13082 11408 13084
rect 11432 13082 11488 13084
rect 11512 13082 11568 13084
rect 11592 13082 11648 13084
rect 11352 13030 11398 13082
rect 11398 13030 11408 13082
rect 11432 13030 11462 13082
rect 11462 13030 11474 13082
rect 11474 13030 11488 13082
rect 11512 13030 11526 13082
rect 11526 13030 11538 13082
rect 11538 13030 11568 13082
rect 11592 13030 11602 13082
rect 11602 13030 11648 13082
rect 11352 13028 11408 13030
rect 11432 13028 11488 13030
rect 11512 13028 11568 13030
rect 11592 13028 11648 13030
rect 11352 11994 11408 11996
rect 11432 11994 11488 11996
rect 11512 11994 11568 11996
rect 11592 11994 11648 11996
rect 11352 11942 11398 11994
rect 11398 11942 11408 11994
rect 11432 11942 11462 11994
rect 11462 11942 11474 11994
rect 11474 11942 11488 11994
rect 11512 11942 11526 11994
rect 11526 11942 11538 11994
rect 11538 11942 11568 11994
rect 11592 11942 11602 11994
rect 11602 11942 11648 11994
rect 11352 11940 11408 11942
rect 11432 11940 11488 11942
rect 11512 11940 11568 11942
rect 11592 11940 11648 11942
rect 11334 11212 11390 11248
rect 11334 11192 11336 11212
rect 11336 11192 11388 11212
rect 11388 11192 11390 11212
rect 10966 10956 10968 10976
rect 10968 10956 11020 10976
rect 11020 10956 11022 10976
rect 10966 10920 11022 10956
rect 10874 10784 10930 10840
rect 10782 10512 10838 10568
rect 10230 7384 10286 7440
rect 9770 1944 9826 2000
rect 10966 10240 11022 10296
rect 10782 8200 10838 8256
rect 10782 6160 10838 6216
rect 10506 3440 10562 3496
rect 10138 1944 10194 2000
rect 9862 1300 9864 1320
rect 9864 1300 9916 1320
rect 9916 1300 9918 1320
rect 9862 1264 9918 1300
rect 8942 40 8998 96
rect 10966 6976 11022 7032
rect 12898 31592 12954 31648
rect 13082 31456 13138 31512
rect 12806 28056 12862 28112
rect 12622 27240 12678 27296
rect 12990 26732 12992 26752
rect 12992 26732 13044 26752
rect 13044 26732 13046 26752
rect 12990 26696 13046 26732
rect 12530 24812 12586 24848
rect 12530 24792 12532 24812
rect 12532 24792 12584 24812
rect 12584 24792 12586 24812
rect 11978 12688 12034 12744
rect 11352 10906 11408 10908
rect 11432 10906 11488 10908
rect 11512 10906 11568 10908
rect 11592 10906 11648 10908
rect 11352 10854 11398 10906
rect 11398 10854 11408 10906
rect 11432 10854 11462 10906
rect 11462 10854 11474 10906
rect 11474 10854 11488 10906
rect 11512 10854 11526 10906
rect 11526 10854 11538 10906
rect 11538 10854 11568 10906
rect 11592 10854 11602 10906
rect 11602 10854 11648 10906
rect 11352 10852 11408 10854
rect 11432 10852 11488 10854
rect 11512 10852 11568 10854
rect 11592 10852 11648 10854
rect 11242 10376 11298 10432
rect 11794 10648 11850 10704
rect 11352 9818 11408 9820
rect 11432 9818 11488 9820
rect 11512 9818 11568 9820
rect 11592 9818 11648 9820
rect 11352 9766 11398 9818
rect 11398 9766 11408 9818
rect 11432 9766 11462 9818
rect 11462 9766 11474 9818
rect 11474 9766 11488 9818
rect 11512 9766 11526 9818
rect 11526 9766 11538 9818
rect 11538 9766 11568 9818
rect 11592 9766 11602 9818
rect 11602 9766 11648 9818
rect 11352 9764 11408 9766
rect 11432 9764 11488 9766
rect 11512 9764 11568 9766
rect 11592 9764 11648 9766
rect 11352 8730 11408 8732
rect 11432 8730 11488 8732
rect 11512 8730 11568 8732
rect 11592 8730 11648 8732
rect 11352 8678 11398 8730
rect 11398 8678 11408 8730
rect 11432 8678 11462 8730
rect 11462 8678 11474 8730
rect 11474 8678 11488 8730
rect 11512 8678 11526 8730
rect 11526 8678 11538 8730
rect 11538 8678 11568 8730
rect 11592 8678 11602 8730
rect 11602 8678 11648 8730
rect 11352 8676 11408 8678
rect 11432 8676 11488 8678
rect 11512 8676 11568 8678
rect 11592 8676 11648 8678
rect 12070 11348 12126 11384
rect 12070 11328 12072 11348
rect 12072 11328 12124 11348
rect 12124 11328 12126 11348
rect 11978 9560 12034 9616
rect 11794 9424 11850 9480
rect 11886 9288 11942 9344
rect 10966 5616 11022 5672
rect 12622 24656 12678 24712
rect 12898 25880 12954 25936
rect 12622 23296 12678 23352
rect 12438 22208 12494 22264
rect 12438 20304 12494 20360
rect 12622 21936 12678 21992
rect 12898 23024 12954 23080
rect 12622 20440 12678 20496
rect 13266 30504 13322 30560
rect 13266 30232 13322 30288
rect 13951 40826 14007 40828
rect 14031 40826 14087 40828
rect 14111 40826 14167 40828
rect 14191 40826 14247 40828
rect 13951 40774 13997 40826
rect 13997 40774 14007 40826
rect 14031 40774 14061 40826
rect 14061 40774 14073 40826
rect 14073 40774 14087 40826
rect 14111 40774 14125 40826
rect 14125 40774 14137 40826
rect 14137 40774 14167 40826
rect 14191 40774 14201 40826
rect 14201 40774 14247 40826
rect 13951 40772 14007 40774
rect 14031 40772 14087 40774
rect 14111 40772 14167 40774
rect 14191 40772 14247 40774
rect 13951 39738 14007 39740
rect 14031 39738 14087 39740
rect 14111 39738 14167 39740
rect 14191 39738 14247 39740
rect 13951 39686 13997 39738
rect 13997 39686 14007 39738
rect 14031 39686 14061 39738
rect 14061 39686 14073 39738
rect 14073 39686 14087 39738
rect 14111 39686 14125 39738
rect 14125 39686 14137 39738
rect 14137 39686 14167 39738
rect 14191 39686 14201 39738
rect 14201 39686 14247 39738
rect 13951 39684 14007 39686
rect 14031 39684 14087 39686
rect 14111 39684 14167 39686
rect 14191 39684 14247 39686
rect 14738 42200 14794 42256
rect 14646 41112 14702 41168
rect 15014 42880 15070 42936
rect 14462 39480 14518 39536
rect 14462 39344 14518 39400
rect 13951 38650 14007 38652
rect 14031 38650 14087 38652
rect 14111 38650 14167 38652
rect 14191 38650 14247 38652
rect 13951 38598 13997 38650
rect 13997 38598 14007 38650
rect 14031 38598 14061 38650
rect 14061 38598 14073 38650
rect 14073 38598 14087 38650
rect 14111 38598 14125 38650
rect 14125 38598 14137 38650
rect 14137 38598 14167 38650
rect 14191 38598 14201 38650
rect 14201 38598 14247 38650
rect 13951 38596 14007 38598
rect 14031 38596 14087 38598
rect 14111 38596 14167 38598
rect 14191 38596 14247 38598
rect 14186 37884 14188 37904
rect 14188 37884 14240 37904
rect 14240 37884 14242 37904
rect 14186 37848 14242 37884
rect 13951 37562 14007 37564
rect 14031 37562 14087 37564
rect 14111 37562 14167 37564
rect 14191 37562 14247 37564
rect 13951 37510 13997 37562
rect 13997 37510 14007 37562
rect 14031 37510 14061 37562
rect 14061 37510 14073 37562
rect 14073 37510 14087 37562
rect 14111 37510 14125 37562
rect 14125 37510 14137 37562
rect 14137 37510 14167 37562
rect 14191 37510 14201 37562
rect 14201 37510 14247 37562
rect 13951 37508 14007 37510
rect 14031 37508 14087 37510
rect 14111 37508 14167 37510
rect 14191 37508 14247 37510
rect 13910 36624 13966 36680
rect 13951 36474 14007 36476
rect 14031 36474 14087 36476
rect 14111 36474 14167 36476
rect 14191 36474 14247 36476
rect 13951 36422 13997 36474
rect 13997 36422 14007 36474
rect 14031 36422 14061 36474
rect 14061 36422 14073 36474
rect 14073 36422 14087 36474
rect 14111 36422 14125 36474
rect 14125 36422 14137 36474
rect 14137 36422 14167 36474
rect 14191 36422 14201 36474
rect 14201 36422 14247 36474
rect 13951 36420 14007 36422
rect 14031 36420 14087 36422
rect 14111 36420 14167 36422
rect 14191 36420 14247 36422
rect 13818 35672 13874 35728
rect 13951 35386 14007 35388
rect 14031 35386 14087 35388
rect 14111 35386 14167 35388
rect 14191 35386 14247 35388
rect 13951 35334 13997 35386
rect 13997 35334 14007 35386
rect 14031 35334 14061 35386
rect 14061 35334 14073 35386
rect 14073 35334 14087 35386
rect 14111 35334 14125 35386
rect 14125 35334 14137 35386
rect 14137 35334 14167 35386
rect 14191 35334 14201 35386
rect 14201 35334 14247 35386
rect 13951 35332 14007 35334
rect 14031 35332 14087 35334
rect 14111 35332 14167 35334
rect 14191 35332 14247 35334
rect 13726 34448 13782 34504
rect 13634 32952 13690 33008
rect 13634 31320 13690 31376
rect 13634 29552 13690 29608
rect 13266 28872 13322 28928
rect 13951 34298 14007 34300
rect 14031 34298 14087 34300
rect 14111 34298 14167 34300
rect 14191 34298 14247 34300
rect 13951 34246 13997 34298
rect 13997 34246 14007 34298
rect 14031 34246 14061 34298
rect 14061 34246 14073 34298
rect 14073 34246 14087 34298
rect 14111 34246 14125 34298
rect 14125 34246 14137 34298
rect 14137 34246 14167 34298
rect 14191 34246 14201 34298
rect 14201 34246 14247 34298
rect 13951 34244 14007 34246
rect 14031 34244 14087 34246
rect 14111 34244 14167 34246
rect 14191 34244 14247 34246
rect 13951 33210 14007 33212
rect 14031 33210 14087 33212
rect 14111 33210 14167 33212
rect 14191 33210 14247 33212
rect 13951 33158 13997 33210
rect 13997 33158 14007 33210
rect 14031 33158 14061 33210
rect 14061 33158 14073 33210
rect 14073 33158 14087 33210
rect 14111 33158 14125 33210
rect 14125 33158 14137 33210
rect 14137 33158 14167 33210
rect 14191 33158 14201 33210
rect 14201 33158 14247 33210
rect 13951 33156 14007 33158
rect 14031 33156 14087 33158
rect 14111 33156 14167 33158
rect 14191 33156 14247 33158
rect 14646 38664 14702 38720
rect 14554 33360 14610 33416
rect 14002 32272 14058 32328
rect 13951 32122 14007 32124
rect 14031 32122 14087 32124
rect 14111 32122 14167 32124
rect 14191 32122 14247 32124
rect 13951 32070 13997 32122
rect 13997 32070 14007 32122
rect 14031 32070 14061 32122
rect 14061 32070 14073 32122
rect 14073 32070 14087 32122
rect 14111 32070 14125 32122
rect 14125 32070 14137 32122
rect 14137 32070 14167 32122
rect 14191 32070 14201 32122
rect 14201 32070 14247 32122
rect 13951 32068 14007 32070
rect 14031 32068 14087 32070
rect 14111 32068 14167 32070
rect 14191 32068 14247 32070
rect 13910 31900 13912 31920
rect 13912 31900 13964 31920
rect 13964 31900 13966 31920
rect 13910 31864 13966 31900
rect 13951 31034 14007 31036
rect 14031 31034 14087 31036
rect 14111 31034 14167 31036
rect 14191 31034 14247 31036
rect 13951 30982 13997 31034
rect 13997 30982 14007 31034
rect 14031 30982 14061 31034
rect 14061 30982 14073 31034
rect 14073 30982 14087 31034
rect 14111 30982 14125 31034
rect 14125 30982 14137 31034
rect 14137 30982 14167 31034
rect 14191 30982 14201 31034
rect 14201 30982 14247 31034
rect 13951 30980 14007 30982
rect 14031 30980 14087 30982
rect 14111 30980 14167 30982
rect 14191 30980 14247 30982
rect 14186 30660 14242 30696
rect 14186 30640 14188 30660
rect 14188 30640 14240 30660
rect 14240 30640 14242 30660
rect 13951 29946 14007 29948
rect 14031 29946 14087 29948
rect 14111 29946 14167 29948
rect 14191 29946 14247 29948
rect 13951 29894 13997 29946
rect 13997 29894 14007 29946
rect 14031 29894 14061 29946
rect 14061 29894 14073 29946
rect 14073 29894 14087 29946
rect 14111 29894 14125 29946
rect 14125 29894 14137 29946
rect 14137 29894 14167 29946
rect 14191 29894 14201 29946
rect 14201 29894 14247 29946
rect 13951 29892 14007 29894
rect 14031 29892 14087 29894
rect 14111 29892 14167 29894
rect 14191 29892 14247 29894
rect 13910 29708 13966 29744
rect 13910 29688 13912 29708
rect 13912 29688 13964 29708
rect 13964 29688 13966 29708
rect 13726 29280 13782 29336
rect 13450 26288 13506 26344
rect 13951 28858 14007 28860
rect 14031 28858 14087 28860
rect 14111 28858 14167 28860
rect 14191 28858 14247 28860
rect 13951 28806 13997 28858
rect 13997 28806 14007 28858
rect 14031 28806 14061 28858
rect 14061 28806 14073 28858
rect 14073 28806 14087 28858
rect 14111 28806 14125 28858
rect 14125 28806 14137 28858
rect 14137 28806 14167 28858
rect 14191 28806 14201 28858
rect 14201 28806 14247 28858
rect 13951 28804 14007 28806
rect 14031 28804 14087 28806
rect 14111 28804 14167 28806
rect 14191 28804 14247 28806
rect 13726 28736 13782 28792
rect 13082 22752 13138 22808
rect 13082 22072 13138 22128
rect 13174 21664 13230 21720
rect 12990 20848 13046 20904
rect 13450 24520 13506 24576
rect 13634 25200 13690 25256
rect 14002 28500 14004 28520
rect 14004 28500 14056 28520
rect 14056 28500 14058 28520
rect 14002 28464 14058 28500
rect 14094 27920 14150 27976
rect 13951 27770 14007 27772
rect 14031 27770 14087 27772
rect 14111 27770 14167 27772
rect 14191 27770 14247 27772
rect 13951 27718 13997 27770
rect 13997 27718 14007 27770
rect 14031 27718 14061 27770
rect 14061 27718 14073 27770
rect 14073 27718 14087 27770
rect 14111 27718 14125 27770
rect 14125 27718 14137 27770
rect 14137 27718 14167 27770
rect 14191 27718 14201 27770
rect 14201 27718 14247 27770
rect 13951 27716 14007 27718
rect 14031 27716 14087 27718
rect 14111 27716 14167 27718
rect 14191 27716 14247 27718
rect 13951 26682 14007 26684
rect 14031 26682 14087 26684
rect 14111 26682 14167 26684
rect 14191 26682 14247 26684
rect 13951 26630 13997 26682
rect 13997 26630 14007 26682
rect 14031 26630 14061 26682
rect 14061 26630 14073 26682
rect 14073 26630 14087 26682
rect 14111 26630 14125 26682
rect 14125 26630 14137 26682
rect 14137 26630 14167 26682
rect 14191 26630 14201 26682
rect 14201 26630 14247 26682
rect 13951 26628 14007 26630
rect 14031 26628 14087 26630
rect 14111 26628 14167 26630
rect 14191 26628 14247 26630
rect 14554 33224 14610 33280
rect 14830 35264 14886 35320
rect 14830 34448 14886 34504
rect 15198 41656 15254 41712
rect 15658 43832 15714 43888
rect 15382 41520 15438 41576
rect 15474 41420 15476 41440
rect 15476 41420 15528 41440
rect 15528 41420 15530 41440
rect 15474 41384 15530 41420
rect 15934 41656 15990 41712
rect 16026 41520 16082 41576
rect 14922 32816 14978 32872
rect 14922 32544 14978 32600
rect 14830 31728 14886 31784
rect 14646 31048 14702 31104
rect 14646 30232 14702 30288
rect 14738 28736 14794 28792
rect 14462 27784 14518 27840
rect 13951 25594 14007 25596
rect 14031 25594 14087 25596
rect 14111 25594 14167 25596
rect 14191 25594 14247 25596
rect 13951 25542 13997 25594
rect 13997 25542 14007 25594
rect 14031 25542 14061 25594
rect 14061 25542 14073 25594
rect 14073 25542 14087 25594
rect 14111 25542 14125 25594
rect 14125 25542 14137 25594
rect 14137 25542 14167 25594
rect 14191 25542 14201 25594
rect 14201 25542 14247 25594
rect 13951 25540 14007 25542
rect 14031 25540 14087 25542
rect 14111 25540 14167 25542
rect 14191 25540 14247 25542
rect 13951 24506 14007 24508
rect 14031 24506 14087 24508
rect 14111 24506 14167 24508
rect 14191 24506 14247 24508
rect 13951 24454 13997 24506
rect 13997 24454 14007 24506
rect 14031 24454 14061 24506
rect 14061 24454 14073 24506
rect 14073 24454 14087 24506
rect 14111 24454 14125 24506
rect 14125 24454 14137 24506
rect 14137 24454 14167 24506
rect 14191 24454 14201 24506
rect 14201 24454 14247 24506
rect 13951 24452 14007 24454
rect 14031 24452 14087 24454
rect 14111 24452 14167 24454
rect 14191 24452 14247 24454
rect 15382 33088 15438 33144
rect 15382 31592 15438 31648
rect 15198 30912 15254 30968
rect 14922 27648 14978 27704
rect 15198 29552 15254 29608
rect 14922 26424 14978 26480
rect 14646 24656 14702 24712
rect 13726 23568 13782 23624
rect 13450 22072 13506 22128
rect 13450 21800 13506 21856
rect 12806 19080 12862 19136
rect 12530 18264 12586 18320
rect 12438 15408 12494 15464
rect 12346 13776 12402 13832
rect 12806 17720 12862 17776
rect 12622 16088 12678 16144
rect 12530 13640 12586 13696
rect 12254 11872 12310 11928
rect 13174 20596 13230 20632
rect 13174 20576 13176 20596
rect 13176 20576 13228 20596
rect 13228 20576 13230 20596
rect 12714 14476 12770 14512
rect 12714 14456 12716 14476
rect 12716 14456 12768 14476
rect 12768 14456 12770 14476
rect 12898 12708 12954 12744
rect 13358 18264 13414 18320
rect 13266 15408 13322 15464
rect 13951 23418 14007 23420
rect 14031 23418 14087 23420
rect 14111 23418 14167 23420
rect 14191 23418 14247 23420
rect 13951 23366 13997 23418
rect 13997 23366 14007 23418
rect 14031 23366 14061 23418
rect 14061 23366 14073 23418
rect 14073 23366 14087 23418
rect 14111 23366 14125 23418
rect 14125 23366 14137 23418
rect 14137 23366 14167 23418
rect 14191 23366 14201 23418
rect 14201 23366 14247 23418
rect 13951 23364 14007 23366
rect 14031 23364 14087 23366
rect 14111 23364 14167 23366
rect 14191 23364 14247 23366
rect 13951 22330 14007 22332
rect 14031 22330 14087 22332
rect 14111 22330 14167 22332
rect 14191 22330 14247 22332
rect 13951 22278 13997 22330
rect 13997 22278 14007 22330
rect 14031 22278 14061 22330
rect 14061 22278 14073 22330
rect 14073 22278 14087 22330
rect 14111 22278 14125 22330
rect 14125 22278 14137 22330
rect 14137 22278 14167 22330
rect 14191 22278 14201 22330
rect 14201 22278 14247 22330
rect 13951 22276 14007 22278
rect 14031 22276 14087 22278
rect 14111 22276 14167 22278
rect 14191 22276 14247 22278
rect 14462 23976 14518 24032
rect 14278 21392 14334 21448
rect 13951 21242 14007 21244
rect 14031 21242 14087 21244
rect 14111 21242 14167 21244
rect 14191 21242 14247 21244
rect 13951 21190 13997 21242
rect 13997 21190 14007 21242
rect 14031 21190 14061 21242
rect 14061 21190 14073 21242
rect 14073 21190 14087 21242
rect 14111 21190 14125 21242
rect 14125 21190 14137 21242
rect 14137 21190 14167 21242
rect 14191 21190 14201 21242
rect 14201 21190 14247 21242
rect 13951 21188 14007 21190
rect 14031 21188 14087 21190
rect 14111 21188 14167 21190
rect 14191 21188 14247 21190
rect 13726 18944 13782 19000
rect 13910 20848 13966 20904
rect 13951 20154 14007 20156
rect 14031 20154 14087 20156
rect 14111 20154 14167 20156
rect 14191 20154 14247 20156
rect 13951 20102 13997 20154
rect 13997 20102 14007 20154
rect 14031 20102 14061 20154
rect 14061 20102 14073 20154
rect 14073 20102 14087 20154
rect 14111 20102 14125 20154
rect 14125 20102 14137 20154
rect 14137 20102 14167 20154
rect 14191 20102 14201 20154
rect 14201 20102 14247 20154
rect 13951 20100 14007 20102
rect 14031 20100 14087 20102
rect 14111 20100 14167 20102
rect 14191 20100 14247 20102
rect 14094 19896 14150 19952
rect 14278 19896 14334 19952
rect 14094 19624 14150 19680
rect 13951 19066 14007 19068
rect 14031 19066 14087 19068
rect 14111 19066 14167 19068
rect 14191 19066 14247 19068
rect 13951 19014 13997 19066
rect 13997 19014 14007 19066
rect 14031 19014 14061 19066
rect 14061 19014 14073 19066
rect 14073 19014 14087 19066
rect 14111 19014 14125 19066
rect 14125 19014 14137 19066
rect 14137 19014 14167 19066
rect 14191 19014 14201 19066
rect 14201 19014 14247 19066
rect 13951 19012 14007 19014
rect 14031 19012 14087 19014
rect 14111 19012 14167 19014
rect 14191 19012 14247 19014
rect 13726 17992 13782 18048
rect 13951 17978 14007 17980
rect 14031 17978 14087 17980
rect 14111 17978 14167 17980
rect 14191 17978 14247 17980
rect 13951 17926 13997 17978
rect 13997 17926 14007 17978
rect 14031 17926 14061 17978
rect 14061 17926 14073 17978
rect 14073 17926 14087 17978
rect 14111 17926 14125 17978
rect 14125 17926 14137 17978
rect 14137 17926 14167 17978
rect 14191 17926 14201 17978
rect 14201 17926 14247 17978
rect 13951 17924 14007 17926
rect 14031 17924 14087 17926
rect 14111 17924 14167 17926
rect 14191 17924 14247 17926
rect 13951 16890 14007 16892
rect 14031 16890 14087 16892
rect 14111 16890 14167 16892
rect 14191 16890 14247 16892
rect 13951 16838 13997 16890
rect 13997 16838 14007 16890
rect 14031 16838 14061 16890
rect 14061 16838 14073 16890
rect 14073 16838 14087 16890
rect 14111 16838 14125 16890
rect 14125 16838 14137 16890
rect 14137 16838 14167 16890
rect 14191 16838 14201 16890
rect 14201 16838 14247 16890
rect 13951 16836 14007 16838
rect 14031 16836 14087 16838
rect 14111 16836 14167 16838
rect 14191 16836 14247 16838
rect 13951 15802 14007 15804
rect 14031 15802 14087 15804
rect 14111 15802 14167 15804
rect 14191 15802 14247 15804
rect 13951 15750 13997 15802
rect 13997 15750 14007 15802
rect 14031 15750 14061 15802
rect 14061 15750 14073 15802
rect 14073 15750 14087 15802
rect 14111 15750 14125 15802
rect 14125 15750 14137 15802
rect 14137 15750 14167 15802
rect 14191 15750 14201 15802
rect 14201 15750 14247 15802
rect 13951 15748 14007 15750
rect 14031 15748 14087 15750
rect 14111 15748 14167 15750
rect 14191 15748 14247 15750
rect 13174 12960 13230 13016
rect 12898 12688 12900 12708
rect 12900 12688 12952 12708
rect 12952 12688 12954 12708
rect 12806 12416 12862 12472
rect 12622 12008 12678 12064
rect 12346 9288 12402 9344
rect 12346 9016 12402 9072
rect 12530 9696 12586 9752
rect 12438 8336 12494 8392
rect 11352 7642 11408 7644
rect 11432 7642 11488 7644
rect 11512 7642 11568 7644
rect 11592 7642 11648 7644
rect 11352 7590 11398 7642
rect 11398 7590 11408 7642
rect 11432 7590 11462 7642
rect 11462 7590 11474 7642
rect 11474 7590 11488 7642
rect 11512 7590 11526 7642
rect 11526 7590 11538 7642
rect 11538 7590 11568 7642
rect 11592 7590 11602 7642
rect 11602 7590 11648 7642
rect 11352 7588 11408 7590
rect 11432 7588 11488 7590
rect 11512 7588 11568 7590
rect 11592 7588 11648 7590
rect 11352 6554 11408 6556
rect 11432 6554 11488 6556
rect 11512 6554 11568 6556
rect 11592 6554 11648 6556
rect 11352 6502 11398 6554
rect 11398 6502 11408 6554
rect 11432 6502 11462 6554
rect 11462 6502 11474 6554
rect 11474 6502 11488 6554
rect 11512 6502 11526 6554
rect 11526 6502 11538 6554
rect 11538 6502 11568 6554
rect 11592 6502 11602 6554
rect 11602 6502 11648 6554
rect 11352 6500 11408 6502
rect 11432 6500 11488 6502
rect 11512 6500 11568 6502
rect 11592 6500 11648 6502
rect 11352 5466 11408 5468
rect 11432 5466 11488 5468
rect 11512 5466 11568 5468
rect 11592 5466 11648 5468
rect 11352 5414 11398 5466
rect 11398 5414 11408 5466
rect 11432 5414 11462 5466
rect 11462 5414 11474 5466
rect 11474 5414 11488 5466
rect 11512 5414 11526 5466
rect 11526 5414 11538 5466
rect 11538 5414 11568 5466
rect 11592 5414 11602 5466
rect 11602 5414 11648 5466
rect 11352 5412 11408 5414
rect 11432 5412 11488 5414
rect 11512 5412 11568 5414
rect 11592 5412 11648 5414
rect 11352 4378 11408 4380
rect 11432 4378 11488 4380
rect 11512 4378 11568 4380
rect 11592 4378 11648 4380
rect 11352 4326 11398 4378
rect 11398 4326 11408 4378
rect 11432 4326 11462 4378
rect 11462 4326 11474 4378
rect 11474 4326 11488 4378
rect 11512 4326 11526 4378
rect 11526 4326 11538 4378
rect 11538 4326 11568 4378
rect 11592 4326 11602 4378
rect 11602 4326 11648 4378
rect 11352 4324 11408 4326
rect 11432 4324 11488 4326
rect 11512 4324 11568 4326
rect 11592 4324 11648 4326
rect 11352 3290 11408 3292
rect 11432 3290 11488 3292
rect 11512 3290 11568 3292
rect 11592 3290 11648 3292
rect 11352 3238 11398 3290
rect 11398 3238 11408 3290
rect 11432 3238 11462 3290
rect 11462 3238 11474 3290
rect 11474 3238 11488 3290
rect 11512 3238 11526 3290
rect 11526 3238 11538 3290
rect 11538 3238 11568 3290
rect 11592 3238 11602 3290
rect 11602 3238 11648 3290
rect 11352 3236 11408 3238
rect 11432 3236 11488 3238
rect 11512 3236 11568 3238
rect 11592 3236 11648 3238
rect 12070 7520 12126 7576
rect 12530 7248 12586 7304
rect 12346 7112 12402 7168
rect 12254 6976 12310 7032
rect 12162 5480 12218 5536
rect 12530 6840 12586 6896
rect 12254 5208 12310 5264
rect 12714 9016 12770 9072
rect 12990 9832 13046 9888
rect 12990 9560 13046 9616
rect 12898 7248 12954 7304
rect 12806 6024 12862 6080
rect 15290 25744 15346 25800
rect 16550 43546 16606 43548
rect 16630 43546 16686 43548
rect 16710 43546 16766 43548
rect 16790 43546 16846 43548
rect 16550 43494 16596 43546
rect 16596 43494 16606 43546
rect 16630 43494 16660 43546
rect 16660 43494 16672 43546
rect 16672 43494 16686 43546
rect 16710 43494 16724 43546
rect 16724 43494 16736 43546
rect 16736 43494 16766 43546
rect 16790 43494 16800 43546
rect 16800 43494 16846 43546
rect 16550 43492 16606 43494
rect 16630 43492 16686 43494
rect 16710 43492 16766 43494
rect 16790 43492 16846 43494
rect 16302 41792 16358 41848
rect 16550 42458 16606 42460
rect 16630 42458 16686 42460
rect 16710 42458 16766 42460
rect 16790 42458 16846 42460
rect 16550 42406 16596 42458
rect 16596 42406 16606 42458
rect 16630 42406 16660 42458
rect 16660 42406 16672 42458
rect 16672 42406 16686 42458
rect 16710 42406 16724 42458
rect 16724 42406 16736 42458
rect 16736 42406 16766 42458
rect 16790 42406 16800 42458
rect 16800 42406 16846 42458
rect 16550 42404 16606 42406
rect 16630 42404 16686 42406
rect 16710 42404 16766 42406
rect 16790 42404 16846 42406
rect 16854 41656 16910 41712
rect 16670 41556 16672 41576
rect 16672 41556 16724 41576
rect 16724 41556 16726 41576
rect 16670 41520 16726 41556
rect 16854 41520 16910 41576
rect 17498 42472 17554 42528
rect 16550 41370 16606 41372
rect 16630 41370 16686 41372
rect 16710 41370 16766 41372
rect 16790 41370 16846 41372
rect 16550 41318 16596 41370
rect 16596 41318 16606 41370
rect 16630 41318 16660 41370
rect 16660 41318 16672 41370
rect 16672 41318 16686 41370
rect 16710 41318 16724 41370
rect 16724 41318 16736 41370
rect 16736 41318 16766 41370
rect 16790 41318 16800 41370
rect 16800 41318 16846 41370
rect 16550 41316 16606 41318
rect 16630 41316 16686 41318
rect 16710 41316 16766 41318
rect 16790 41316 16846 41318
rect 16578 41012 16580 41032
rect 16580 41012 16632 41032
rect 16632 41012 16634 41032
rect 16578 40976 16634 41012
rect 17038 41112 17094 41168
rect 16550 40282 16606 40284
rect 16630 40282 16686 40284
rect 16710 40282 16766 40284
rect 16790 40282 16846 40284
rect 16550 40230 16596 40282
rect 16596 40230 16606 40282
rect 16630 40230 16660 40282
rect 16660 40230 16672 40282
rect 16672 40230 16686 40282
rect 16710 40230 16724 40282
rect 16724 40230 16736 40282
rect 16736 40230 16766 40282
rect 16790 40230 16800 40282
rect 16800 40230 16846 40282
rect 16550 40228 16606 40230
rect 16630 40228 16686 40230
rect 16710 40228 16766 40230
rect 16790 40228 16846 40230
rect 16550 39194 16606 39196
rect 16630 39194 16686 39196
rect 16710 39194 16766 39196
rect 16790 39194 16846 39196
rect 16550 39142 16596 39194
rect 16596 39142 16606 39194
rect 16630 39142 16660 39194
rect 16660 39142 16672 39194
rect 16672 39142 16686 39194
rect 16710 39142 16724 39194
rect 16724 39142 16736 39194
rect 16736 39142 16766 39194
rect 16790 39142 16800 39194
rect 16800 39142 16846 39194
rect 16550 39140 16606 39142
rect 16630 39140 16686 39142
rect 16710 39140 16766 39142
rect 16790 39140 16846 39142
rect 16486 38936 16542 38992
rect 16550 38106 16606 38108
rect 16630 38106 16686 38108
rect 16710 38106 16766 38108
rect 16790 38106 16846 38108
rect 16550 38054 16596 38106
rect 16596 38054 16606 38106
rect 16630 38054 16660 38106
rect 16660 38054 16672 38106
rect 16672 38054 16686 38106
rect 16710 38054 16724 38106
rect 16724 38054 16736 38106
rect 16736 38054 16766 38106
rect 16790 38054 16800 38106
rect 16800 38054 16846 38106
rect 16550 38052 16606 38054
rect 16630 38052 16686 38054
rect 16710 38052 16766 38054
rect 16790 38052 16846 38054
rect 17222 40160 17278 40216
rect 16550 37018 16606 37020
rect 16630 37018 16686 37020
rect 16710 37018 16766 37020
rect 16790 37018 16846 37020
rect 16550 36966 16596 37018
rect 16596 36966 16606 37018
rect 16630 36966 16660 37018
rect 16660 36966 16672 37018
rect 16672 36966 16686 37018
rect 16710 36966 16724 37018
rect 16724 36966 16736 37018
rect 16736 36966 16766 37018
rect 16790 36966 16800 37018
rect 16800 36966 16846 37018
rect 16550 36964 16606 36966
rect 16630 36964 16686 36966
rect 16710 36964 16766 36966
rect 16790 36964 16846 36966
rect 15842 33768 15898 33824
rect 15750 32952 15806 33008
rect 15474 27376 15530 27432
rect 14922 24656 14978 24712
rect 14830 22208 14886 22264
rect 14646 18844 14648 18864
rect 14648 18844 14700 18864
rect 14700 18844 14702 18864
rect 14646 18808 14702 18844
rect 15382 23296 15438 23352
rect 15474 23160 15530 23216
rect 15014 22480 15070 22536
rect 15382 23024 15438 23080
rect 14738 17584 14794 17640
rect 14738 17076 14740 17096
rect 14740 17076 14792 17096
rect 14792 17076 14794 17096
rect 14738 17040 14794 17076
rect 14738 16652 14794 16688
rect 14738 16632 14740 16652
rect 14740 16632 14792 16652
rect 14792 16632 14794 16652
rect 13951 14714 14007 14716
rect 14031 14714 14087 14716
rect 14111 14714 14167 14716
rect 14191 14714 14247 14716
rect 13951 14662 13997 14714
rect 13997 14662 14007 14714
rect 14031 14662 14061 14714
rect 14061 14662 14073 14714
rect 14073 14662 14087 14714
rect 14111 14662 14125 14714
rect 14125 14662 14137 14714
rect 14137 14662 14167 14714
rect 14191 14662 14201 14714
rect 14201 14662 14247 14714
rect 13951 14660 14007 14662
rect 14031 14660 14087 14662
rect 14111 14660 14167 14662
rect 14191 14660 14247 14662
rect 13951 13626 14007 13628
rect 14031 13626 14087 13628
rect 14111 13626 14167 13628
rect 14191 13626 14247 13628
rect 13951 13574 13997 13626
rect 13997 13574 14007 13626
rect 14031 13574 14061 13626
rect 14061 13574 14073 13626
rect 14073 13574 14087 13626
rect 14111 13574 14125 13626
rect 14125 13574 14137 13626
rect 14137 13574 14167 13626
rect 14191 13574 14201 13626
rect 14201 13574 14247 13626
rect 13951 13572 14007 13574
rect 14031 13572 14087 13574
rect 14111 13572 14167 13574
rect 14191 13572 14247 13574
rect 13818 12844 13874 12880
rect 13818 12824 13820 12844
rect 13820 12824 13872 12844
rect 13872 12824 13874 12844
rect 13542 11756 13598 11792
rect 13542 11736 13544 11756
rect 13544 11736 13596 11756
rect 13596 11736 13598 11756
rect 13951 12538 14007 12540
rect 14031 12538 14087 12540
rect 14111 12538 14167 12540
rect 14191 12538 14247 12540
rect 13951 12486 13997 12538
rect 13997 12486 14007 12538
rect 14031 12486 14061 12538
rect 14061 12486 14073 12538
rect 14073 12486 14087 12538
rect 14111 12486 14125 12538
rect 14125 12486 14137 12538
rect 14137 12486 14167 12538
rect 14191 12486 14201 12538
rect 14201 12486 14247 12538
rect 13951 12484 14007 12486
rect 14031 12484 14087 12486
rect 14111 12484 14167 12486
rect 14191 12484 14247 12486
rect 13910 12144 13966 12200
rect 13951 11450 14007 11452
rect 14031 11450 14087 11452
rect 14111 11450 14167 11452
rect 14191 11450 14247 11452
rect 13951 11398 13997 11450
rect 13997 11398 14007 11450
rect 14031 11398 14061 11450
rect 14061 11398 14073 11450
rect 14073 11398 14087 11450
rect 14111 11398 14125 11450
rect 14125 11398 14137 11450
rect 14137 11398 14167 11450
rect 14191 11398 14201 11450
rect 14201 11398 14247 11450
rect 13951 11396 14007 11398
rect 14031 11396 14087 11398
rect 14111 11396 14167 11398
rect 14191 11396 14247 11398
rect 13542 10124 13598 10160
rect 13542 10104 13544 10124
rect 13544 10104 13596 10124
rect 13596 10104 13598 10124
rect 13358 9696 13414 9752
rect 13266 8336 13322 8392
rect 13174 5208 13230 5264
rect 11352 2202 11408 2204
rect 11432 2202 11488 2204
rect 11512 2202 11568 2204
rect 11592 2202 11648 2204
rect 11352 2150 11398 2202
rect 11398 2150 11408 2202
rect 11432 2150 11462 2202
rect 11462 2150 11474 2202
rect 11474 2150 11488 2202
rect 11512 2150 11526 2202
rect 11526 2150 11538 2202
rect 11538 2150 11568 2202
rect 11592 2150 11602 2202
rect 11602 2150 11648 2202
rect 11352 2148 11408 2150
rect 11432 2148 11488 2150
rect 11512 2148 11568 2150
rect 11592 2148 11648 2150
rect 11352 1114 11408 1116
rect 11432 1114 11488 1116
rect 11512 1114 11568 1116
rect 11592 1114 11648 1116
rect 11352 1062 11398 1114
rect 11398 1062 11408 1114
rect 11432 1062 11462 1114
rect 11462 1062 11474 1114
rect 11474 1062 11488 1114
rect 11512 1062 11526 1114
rect 11526 1062 11538 1114
rect 11538 1062 11568 1114
rect 11592 1062 11602 1114
rect 11602 1062 11648 1114
rect 11352 1060 11408 1062
rect 11432 1060 11488 1062
rect 11512 1060 11568 1062
rect 11592 1060 11648 1062
rect 11978 1944 12034 2000
rect 12714 1964 12770 2000
rect 12714 1944 12716 1964
rect 12716 1944 12768 1964
rect 12768 1944 12770 1964
rect 13450 9324 13452 9344
rect 13452 9324 13504 9344
rect 13504 9324 13506 9344
rect 13450 9288 13506 9324
rect 13910 11056 13966 11112
rect 14278 10648 14334 10704
rect 13951 10362 14007 10364
rect 14031 10362 14087 10364
rect 14111 10362 14167 10364
rect 14191 10362 14247 10364
rect 13951 10310 13997 10362
rect 13997 10310 14007 10362
rect 14031 10310 14061 10362
rect 14061 10310 14073 10362
rect 14073 10310 14087 10362
rect 14111 10310 14125 10362
rect 14125 10310 14137 10362
rect 14137 10310 14167 10362
rect 14191 10310 14201 10362
rect 14201 10310 14247 10362
rect 13951 10308 14007 10310
rect 14031 10308 14087 10310
rect 14111 10308 14167 10310
rect 14191 10308 14247 10310
rect 15290 20848 15346 20904
rect 15106 19916 15162 19952
rect 15106 19896 15108 19916
rect 15108 19896 15160 19916
rect 15160 19896 15162 19916
rect 15198 19624 15254 19680
rect 15106 17312 15162 17368
rect 15014 17176 15070 17232
rect 14554 10104 14610 10160
rect 13951 9274 14007 9276
rect 14031 9274 14087 9276
rect 14111 9274 14167 9276
rect 14191 9274 14247 9276
rect 13951 9222 13997 9274
rect 13997 9222 14007 9274
rect 14031 9222 14061 9274
rect 14061 9222 14073 9274
rect 14073 9222 14087 9274
rect 14111 9222 14125 9274
rect 14125 9222 14137 9274
rect 14137 9222 14167 9274
rect 14191 9222 14201 9274
rect 14201 9222 14247 9274
rect 13951 9220 14007 9222
rect 14031 9220 14087 9222
rect 14111 9220 14167 9222
rect 14191 9220 14247 9222
rect 14186 8608 14242 8664
rect 14646 9968 14702 10024
rect 13951 8186 14007 8188
rect 14031 8186 14087 8188
rect 14111 8186 14167 8188
rect 14191 8186 14247 8188
rect 13951 8134 13997 8186
rect 13997 8134 14007 8186
rect 14031 8134 14061 8186
rect 14061 8134 14073 8186
rect 14073 8134 14087 8186
rect 14111 8134 14125 8186
rect 14125 8134 14137 8186
rect 14137 8134 14167 8186
rect 14191 8134 14201 8186
rect 14201 8134 14247 8186
rect 13951 8132 14007 8134
rect 14031 8132 14087 8134
rect 14111 8132 14167 8134
rect 14191 8132 14247 8134
rect 13634 4392 13690 4448
rect 14002 7828 14004 7848
rect 14004 7828 14056 7848
rect 14056 7828 14058 7848
rect 14002 7792 14058 7828
rect 13951 7098 14007 7100
rect 14031 7098 14087 7100
rect 14111 7098 14167 7100
rect 14191 7098 14247 7100
rect 13951 7046 13997 7098
rect 13997 7046 14007 7098
rect 14031 7046 14061 7098
rect 14061 7046 14073 7098
rect 14073 7046 14087 7098
rect 14111 7046 14125 7098
rect 14125 7046 14137 7098
rect 14137 7046 14167 7098
rect 14191 7046 14201 7098
rect 14201 7046 14247 7098
rect 13951 7044 14007 7046
rect 14031 7044 14087 7046
rect 14111 7044 14167 7046
rect 14191 7044 14247 7046
rect 14278 6568 14334 6624
rect 14554 7520 14610 7576
rect 15290 16768 15346 16824
rect 15290 12688 15346 12744
rect 15198 12280 15254 12336
rect 15014 9288 15070 9344
rect 14738 8608 14794 8664
rect 14738 8336 14794 8392
rect 15290 9596 15292 9616
rect 15292 9596 15344 9616
rect 15344 9596 15346 9616
rect 15290 9560 15346 9596
rect 13951 6010 14007 6012
rect 14031 6010 14087 6012
rect 14111 6010 14167 6012
rect 14191 6010 14247 6012
rect 13951 5958 13997 6010
rect 13997 5958 14007 6010
rect 14031 5958 14061 6010
rect 14061 5958 14073 6010
rect 14073 5958 14087 6010
rect 14111 5958 14125 6010
rect 14125 5958 14137 6010
rect 14137 5958 14167 6010
rect 14191 5958 14201 6010
rect 14201 5958 14247 6010
rect 13951 5956 14007 5958
rect 14031 5956 14087 5958
rect 14111 5956 14167 5958
rect 14191 5956 14247 5958
rect 13951 4922 14007 4924
rect 14031 4922 14087 4924
rect 14111 4922 14167 4924
rect 14191 4922 14247 4924
rect 13951 4870 13997 4922
rect 13997 4870 14007 4922
rect 14031 4870 14061 4922
rect 14061 4870 14073 4922
rect 14073 4870 14087 4922
rect 14111 4870 14125 4922
rect 14125 4870 14137 4922
rect 14137 4870 14167 4922
rect 14191 4870 14201 4922
rect 14201 4870 14247 4922
rect 13951 4868 14007 4870
rect 14031 4868 14087 4870
rect 14111 4868 14167 4870
rect 14191 4868 14247 4870
rect 14554 6160 14610 6216
rect 14830 8200 14886 8256
rect 14554 5208 14610 5264
rect 13951 3834 14007 3836
rect 14031 3834 14087 3836
rect 14111 3834 14167 3836
rect 14191 3834 14247 3836
rect 13951 3782 13997 3834
rect 13997 3782 14007 3834
rect 14031 3782 14061 3834
rect 14061 3782 14073 3834
rect 14073 3782 14087 3834
rect 14111 3782 14125 3834
rect 14125 3782 14137 3834
rect 14137 3782 14167 3834
rect 14191 3782 14201 3834
rect 14201 3782 14247 3834
rect 13951 3780 14007 3782
rect 14031 3780 14087 3782
rect 14111 3780 14167 3782
rect 14191 3780 14247 3782
rect 14922 4800 14978 4856
rect 14738 4120 14794 4176
rect 13450 1944 13506 2000
rect 14370 3712 14426 3768
rect 14094 3576 14150 3632
rect 14646 3848 14702 3904
rect 15106 6840 15162 6896
rect 15106 5752 15162 5808
rect 16550 35930 16606 35932
rect 16630 35930 16686 35932
rect 16710 35930 16766 35932
rect 16790 35930 16846 35932
rect 16550 35878 16596 35930
rect 16596 35878 16606 35930
rect 16630 35878 16660 35930
rect 16660 35878 16672 35930
rect 16672 35878 16686 35930
rect 16710 35878 16724 35930
rect 16724 35878 16736 35930
rect 16736 35878 16766 35930
rect 16790 35878 16800 35930
rect 16800 35878 16846 35930
rect 16550 35876 16606 35878
rect 16630 35876 16686 35878
rect 16710 35876 16766 35878
rect 16790 35876 16846 35878
rect 16550 34842 16606 34844
rect 16630 34842 16686 34844
rect 16710 34842 16766 34844
rect 16790 34842 16846 34844
rect 16550 34790 16596 34842
rect 16596 34790 16606 34842
rect 16630 34790 16660 34842
rect 16660 34790 16672 34842
rect 16672 34790 16686 34842
rect 16710 34790 16724 34842
rect 16724 34790 16736 34842
rect 16736 34790 16766 34842
rect 16790 34790 16800 34842
rect 16800 34790 16846 34842
rect 16550 34788 16606 34790
rect 16630 34788 16686 34790
rect 16710 34788 16766 34790
rect 16790 34788 16846 34790
rect 15934 29960 15990 30016
rect 15934 29280 15990 29336
rect 15934 26288 15990 26344
rect 15934 25336 15990 25392
rect 16302 30676 16304 30696
rect 16304 30676 16356 30696
rect 16356 30676 16358 30696
rect 16302 30640 16358 30676
rect 16550 33754 16606 33756
rect 16630 33754 16686 33756
rect 16710 33754 16766 33756
rect 16790 33754 16846 33756
rect 16550 33702 16596 33754
rect 16596 33702 16606 33754
rect 16630 33702 16660 33754
rect 16660 33702 16672 33754
rect 16672 33702 16686 33754
rect 16710 33702 16724 33754
rect 16724 33702 16736 33754
rect 16736 33702 16766 33754
rect 16790 33702 16800 33754
rect 16800 33702 16846 33754
rect 16550 33700 16606 33702
rect 16630 33700 16686 33702
rect 16710 33700 16766 33702
rect 16790 33700 16846 33702
rect 16550 32666 16606 32668
rect 16630 32666 16686 32668
rect 16710 32666 16766 32668
rect 16790 32666 16846 32668
rect 16550 32614 16596 32666
rect 16596 32614 16606 32666
rect 16630 32614 16660 32666
rect 16660 32614 16672 32666
rect 16672 32614 16686 32666
rect 16710 32614 16724 32666
rect 16724 32614 16736 32666
rect 16736 32614 16766 32666
rect 16790 32614 16800 32666
rect 16800 32614 16846 32666
rect 16550 32612 16606 32614
rect 16630 32612 16686 32614
rect 16710 32612 16766 32614
rect 16790 32612 16846 32614
rect 17222 38664 17278 38720
rect 17498 40840 17554 40896
rect 17866 41792 17922 41848
rect 17774 41556 17776 41576
rect 17776 41556 17828 41576
rect 17828 41556 17830 41576
rect 17774 41520 17830 41556
rect 18326 43152 18382 43208
rect 17958 40976 18014 41032
rect 17774 40568 17830 40624
rect 18050 40296 18106 40352
rect 18602 42880 18658 42936
rect 19149 43002 19205 43004
rect 19229 43002 19285 43004
rect 19309 43002 19365 43004
rect 19389 43002 19445 43004
rect 19149 42950 19195 43002
rect 19195 42950 19205 43002
rect 19229 42950 19259 43002
rect 19259 42950 19271 43002
rect 19271 42950 19285 43002
rect 19309 42950 19323 43002
rect 19323 42950 19335 43002
rect 19335 42950 19365 43002
rect 19389 42950 19399 43002
rect 19399 42950 19445 43002
rect 19149 42948 19205 42950
rect 19229 42948 19285 42950
rect 19309 42948 19365 42950
rect 19389 42948 19445 42950
rect 18970 42472 19026 42528
rect 22374 43560 22430 43616
rect 21748 43546 21804 43548
rect 21828 43546 21884 43548
rect 21908 43546 21964 43548
rect 21988 43546 22044 43548
rect 21748 43494 21794 43546
rect 21794 43494 21804 43546
rect 21828 43494 21858 43546
rect 21858 43494 21870 43546
rect 21870 43494 21884 43546
rect 21908 43494 21922 43546
rect 21922 43494 21934 43546
rect 21934 43494 21964 43546
rect 21988 43494 21998 43546
rect 21998 43494 22044 43546
rect 21748 43492 21804 43494
rect 21828 43492 21884 43494
rect 21908 43492 21964 43494
rect 21988 43492 22044 43494
rect 20534 43016 20590 43072
rect 19522 42064 19578 42120
rect 18970 41792 19026 41848
rect 18326 41248 18382 41304
rect 18234 41132 18290 41168
rect 18234 41112 18236 41132
rect 18236 41112 18288 41132
rect 18288 41112 18290 41132
rect 17314 35264 17370 35320
rect 17222 33360 17278 33416
rect 16550 31578 16606 31580
rect 16630 31578 16686 31580
rect 16710 31578 16766 31580
rect 16790 31578 16846 31580
rect 16550 31526 16596 31578
rect 16596 31526 16606 31578
rect 16630 31526 16660 31578
rect 16660 31526 16672 31578
rect 16672 31526 16686 31578
rect 16710 31526 16724 31578
rect 16724 31526 16736 31578
rect 16736 31526 16766 31578
rect 16790 31526 16800 31578
rect 16800 31526 16846 31578
rect 16550 31524 16606 31526
rect 16630 31524 16686 31526
rect 16710 31524 16766 31526
rect 16790 31524 16846 31526
rect 16550 30490 16606 30492
rect 16630 30490 16686 30492
rect 16710 30490 16766 30492
rect 16790 30490 16846 30492
rect 16550 30438 16596 30490
rect 16596 30438 16606 30490
rect 16630 30438 16660 30490
rect 16660 30438 16672 30490
rect 16672 30438 16686 30490
rect 16710 30438 16724 30490
rect 16724 30438 16736 30490
rect 16736 30438 16766 30490
rect 16790 30438 16800 30490
rect 16800 30438 16846 30490
rect 16550 30436 16606 30438
rect 16630 30436 16686 30438
rect 16710 30436 16766 30438
rect 16790 30436 16846 30438
rect 16210 28736 16266 28792
rect 16210 28500 16212 28520
rect 16212 28500 16264 28520
rect 16264 28500 16266 28520
rect 16210 28464 16266 28500
rect 16550 29402 16606 29404
rect 16630 29402 16686 29404
rect 16710 29402 16766 29404
rect 16790 29402 16846 29404
rect 16550 29350 16596 29402
rect 16596 29350 16606 29402
rect 16630 29350 16660 29402
rect 16660 29350 16672 29402
rect 16672 29350 16686 29402
rect 16710 29350 16724 29402
rect 16724 29350 16736 29402
rect 16736 29350 16766 29402
rect 16790 29350 16800 29402
rect 16800 29350 16846 29402
rect 16550 29348 16606 29350
rect 16630 29348 16686 29350
rect 16710 29348 16766 29350
rect 16790 29348 16846 29350
rect 17038 28872 17094 28928
rect 16550 28314 16606 28316
rect 16630 28314 16686 28316
rect 16710 28314 16766 28316
rect 16790 28314 16846 28316
rect 16550 28262 16596 28314
rect 16596 28262 16606 28314
rect 16630 28262 16660 28314
rect 16660 28262 16672 28314
rect 16672 28262 16686 28314
rect 16710 28262 16724 28314
rect 16724 28262 16736 28314
rect 16736 28262 16766 28314
rect 16790 28262 16800 28314
rect 16800 28262 16846 28314
rect 16550 28260 16606 28262
rect 16630 28260 16686 28262
rect 16710 28260 16766 28262
rect 16790 28260 16846 28262
rect 17130 27920 17186 27976
rect 16550 27226 16606 27228
rect 16630 27226 16686 27228
rect 16710 27226 16766 27228
rect 16790 27226 16846 27228
rect 16550 27174 16596 27226
rect 16596 27174 16606 27226
rect 16630 27174 16660 27226
rect 16660 27174 16672 27226
rect 16672 27174 16686 27226
rect 16710 27174 16724 27226
rect 16724 27174 16736 27226
rect 16736 27174 16766 27226
rect 16790 27174 16800 27226
rect 16800 27174 16846 27226
rect 16550 27172 16606 27174
rect 16630 27172 16686 27174
rect 16710 27172 16766 27174
rect 16790 27172 16846 27174
rect 16550 26138 16606 26140
rect 16630 26138 16686 26140
rect 16710 26138 16766 26140
rect 16790 26138 16846 26140
rect 16550 26086 16596 26138
rect 16596 26086 16606 26138
rect 16630 26086 16660 26138
rect 16660 26086 16672 26138
rect 16672 26086 16686 26138
rect 16710 26086 16724 26138
rect 16724 26086 16736 26138
rect 16736 26086 16766 26138
rect 16790 26086 16800 26138
rect 16800 26086 16846 26138
rect 16550 26084 16606 26086
rect 16630 26084 16686 26086
rect 16710 26084 16766 26086
rect 16790 26084 16846 26086
rect 15658 24928 15714 24984
rect 15566 23024 15622 23080
rect 15566 22888 15622 22944
rect 15658 21120 15714 21176
rect 16550 25050 16606 25052
rect 16630 25050 16686 25052
rect 16710 25050 16766 25052
rect 16790 25050 16846 25052
rect 16550 24998 16596 25050
rect 16596 24998 16606 25050
rect 16630 24998 16660 25050
rect 16660 24998 16672 25050
rect 16672 24998 16686 25050
rect 16710 24998 16724 25050
rect 16724 24998 16736 25050
rect 16736 24998 16766 25050
rect 16790 24998 16800 25050
rect 16800 24998 16846 25050
rect 16550 24996 16606 24998
rect 16630 24996 16686 24998
rect 16710 24996 16766 24998
rect 16790 24996 16846 24998
rect 16946 24792 17002 24848
rect 16394 24384 16450 24440
rect 16550 23962 16606 23964
rect 16630 23962 16686 23964
rect 16710 23962 16766 23964
rect 16790 23962 16846 23964
rect 16550 23910 16596 23962
rect 16596 23910 16606 23962
rect 16630 23910 16660 23962
rect 16660 23910 16672 23962
rect 16672 23910 16686 23962
rect 16710 23910 16724 23962
rect 16724 23910 16736 23962
rect 16736 23910 16766 23962
rect 16790 23910 16800 23962
rect 16800 23910 16846 23962
rect 16550 23908 16606 23910
rect 16630 23908 16686 23910
rect 16710 23908 16766 23910
rect 16790 23908 16846 23910
rect 16302 22752 16358 22808
rect 16550 22874 16606 22876
rect 16630 22874 16686 22876
rect 16710 22874 16766 22876
rect 16790 22874 16846 22876
rect 16550 22822 16596 22874
rect 16596 22822 16606 22874
rect 16630 22822 16660 22874
rect 16660 22822 16672 22874
rect 16672 22822 16686 22874
rect 16710 22822 16724 22874
rect 16724 22822 16736 22874
rect 16736 22822 16766 22874
rect 16790 22822 16800 22874
rect 16800 22822 16846 22874
rect 16550 22820 16606 22822
rect 16630 22820 16686 22822
rect 16710 22820 16766 22822
rect 16790 22820 16846 22822
rect 17774 39480 17830 39536
rect 18418 40432 18474 40488
rect 18878 41112 18934 41168
rect 18602 40568 18658 40624
rect 19149 41914 19205 41916
rect 19229 41914 19285 41916
rect 19309 41914 19365 41916
rect 19389 41914 19445 41916
rect 19149 41862 19195 41914
rect 19195 41862 19205 41914
rect 19229 41862 19259 41914
rect 19259 41862 19271 41914
rect 19271 41862 19285 41914
rect 19309 41862 19323 41914
rect 19323 41862 19335 41914
rect 19335 41862 19365 41914
rect 19389 41862 19399 41914
rect 19399 41862 19445 41914
rect 19149 41860 19205 41862
rect 19229 41860 19285 41862
rect 19309 41860 19365 41862
rect 19389 41860 19445 41862
rect 20442 42336 20498 42392
rect 19246 40976 19302 41032
rect 19149 40826 19205 40828
rect 19229 40826 19285 40828
rect 19309 40826 19365 40828
rect 19389 40826 19445 40828
rect 19149 40774 19195 40826
rect 19195 40774 19205 40826
rect 19229 40774 19259 40826
rect 19259 40774 19271 40826
rect 19271 40774 19285 40826
rect 19309 40774 19323 40826
rect 19323 40774 19335 40826
rect 19335 40774 19365 40826
rect 19389 40774 19399 40826
rect 19399 40774 19445 40826
rect 19149 40772 19205 40774
rect 19229 40772 19285 40774
rect 19309 40772 19365 40774
rect 19389 40772 19445 40774
rect 19798 40704 19854 40760
rect 19062 40024 19118 40080
rect 19522 39888 19578 39944
rect 19149 39738 19205 39740
rect 19229 39738 19285 39740
rect 19309 39738 19365 39740
rect 19389 39738 19445 39740
rect 19149 39686 19195 39738
rect 19195 39686 19205 39738
rect 19229 39686 19259 39738
rect 19259 39686 19271 39738
rect 19271 39686 19285 39738
rect 19309 39686 19323 39738
rect 19323 39686 19335 39738
rect 19335 39686 19365 39738
rect 19389 39686 19399 39738
rect 19399 39686 19445 39738
rect 19149 39684 19205 39686
rect 19229 39684 19285 39686
rect 19309 39684 19365 39686
rect 19389 39684 19445 39686
rect 17682 27784 17738 27840
rect 18050 35536 18106 35592
rect 18326 35692 18382 35728
rect 18326 35672 18328 35692
rect 18328 35672 18380 35692
rect 18380 35672 18382 35692
rect 18418 35128 18474 35184
rect 18234 34992 18290 35048
rect 18326 33224 18382 33280
rect 17866 32408 17922 32464
rect 17130 23432 17186 23488
rect 15934 20304 15990 20360
rect 15658 17584 15714 17640
rect 16118 18400 16174 18456
rect 16210 18128 16266 18184
rect 15934 13912 15990 13968
rect 15658 13368 15714 13424
rect 15566 12960 15622 13016
rect 15658 10920 15714 10976
rect 15290 7656 15346 7712
rect 17038 21836 17040 21856
rect 17040 21836 17092 21856
rect 17092 21836 17094 21856
rect 17038 21800 17094 21836
rect 16550 21786 16606 21788
rect 16630 21786 16686 21788
rect 16710 21786 16766 21788
rect 16790 21786 16846 21788
rect 16550 21734 16596 21786
rect 16596 21734 16606 21786
rect 16630 21734 16660 21786
rect 16660 21734 16672 21786
rect 16672 21734 16686 21786
rect 16710 21734 16724 21786
rect 16724 21734 16736 21786
rect 16736 21734 16766 21786
rect 16790 21734 16800 21786
rect 16800 21734 16846 21786
rect 16550 21732 16606 21734
rect 16630 21732 16686 21734
rect 16710 21732 16766 21734
rect 16790 21732 16846 21734
rect 16550 20698 16606 20700
rect 16630 20698 16686 20700
rect 16710 20698 16766 20700
rect 16790 20698 16846 20700
rect 16550 20646 16596 20698
rect 16596 20646 16606 20698
rect 16630 20646 16660 20698
rect 16660 20646 16672 20698
rect 16672 20646 16686 20698
rect 16710 20646 16724 20698
rect 16724 20646 16736 20698
rect 16736 20646 16766 20698
rect 16790 20646 16800 20698
rect 16800 20646 16846 20698
rect 16550 20644 16606 20646
rect 16630 20644 16686 20646
rect 16710 20644 16766 20646
rect 16790 20644 16846 20646
rect 16946 20032 17002 20088
rect 16762 19896 16818 19952
rect 16550 19610 16606 19612
rect 16630 19610 16686 19612
rect 16710 19610 16766 19612
rect 16790 19610 16846 19612
rect 16550 19558 16596 19610
rect 16596 19558 16606 19610
rect 16630 19558 16660 19610
rect 16660 19558 16672 19610
rect 16672 19558 16686 19610
rect 16710 19558 16724 19610
rect 16724 19558 16736 19610
rect 16736 19558 16766 19610
rect 16790 19558 16800 19610
rect 16800 19558 16846 19610
rect 16550 19556 16606 19558
rect 16630 19556 16686 19558
rect 16710 19556 16766 19558
rect 16790 19556 16846 19558
rect 17406 23296 17462 23352
rect 18050 26968 18106 27024
rect 17130 20304 17186 20360
rect 17130 20032 17186 20088
rect 17130 19216 17186 19272
rect 16550 18522 16606 18524
rect 16630 18522 16686 18524
rect 16710 18522 16766 18524
rect 16790 18522 16846 18524
rect 16550 18470 16596 18522
rect 16596 18470 16606 18522
rect 16630 18470 16660 18522
rect 16660 18470 16672 18522
rect 16672 18470 16686 18522
rect 16710 18470 16724 18522
rect 16724 18470 16736 18522
rect 16736 18470 16766 18522
rect 16790 18470 16800 18522
rect 16800 18470 16846 18522
rect 16550 18468 16606 18470
rect 16630 18468 16686 18470
rect 16710 18468 16766 18470
rect 16790 18468 16846 18470
rect 16302 15544 16358 15600
rect 16550 17434 16606 17436
rect 16630 17434 16686 17436
rect 16710 17434 16766 17436
rect 16790 17434 16846 17436
rect 16550 17382 16596 17434
rect 16596 17382 16606 17434
rect 16630 17382 16660 17434
rect 16660 17382 16672 17434
rect 16672 17382 16686 17434
rect 16710 17382 16724 17434
rect 16724 17382 16736 17434
rect 16736 17382 16766 17434
rect 16790 17382 16800 17434
rect 16800 17382 16846 17434
rect 16550 17380 16606 17382
rect 16630 17380 16686 17382
rect 16710 17380 16766 17382
rect 16790 17380 16846 17382
rect 16762 16904 16818 16960
rect 16550 16346 16606 16348
rect 16630 16346 16686 16348
rect 16710 16346 16766 16348
rect 16790 16346 16846 16348
rect 16550 16294 16596 16346
rect 16596 16294 16606 16346
rect 16630 16294 16660 16346
rect 16660 16294 16672 16346
rect 16672 16294 16686 16346
rect 16710 16294 16724 16346
rect 16724 16294 16736 16346
rect 16736 16294 16766 16346
rect 16790 16294 16800 16346
rect 16800 16294 16846 16346
rect 16550 16292 16606 16294
rect 16630 16292 16686 16294
rect 16710 16292 16766 16294
rect 16790 16292 16846 16294
rect 16550 15258 16606 15260
rect 16630 15258 16686 15260
rect 16710 15258 16766 15260
rect 16790 15258 16846 15260
rect 16550 15206 16596 15258
rect 16596 15206 16606 15258
rect 16630 15206 16660 15258
rect 16660 15206 16672 15258
rect 16672 15206 16686 15258
rect 16710 15206 16724 15258
rect 16724 15206 16736 15258
rect 16736 15206 16766 15258
rect 16790 15206 16800 15258
rect 16800 15206 16846 15258
rect 16550 15204 16606 15206
rect 16630 15204 16686 15206
rect 16710 15204 16766 15206
rect 16790 15204 16846 15206
rect 15842 11056 15898 11112
rect 15842 9016 15898 9072
rect 16026 9560 16082 9616
rect 16550 14170 16606 14172
rect 16630 14170 16686 14172
rect 16710 14170 16766 14172
rect 16790 14170 16846 14172
rect 16550 14118 16596 14170
rect 16596 14118 16606 14170
rect 16630 14118 16660 14170
rect 16660 14118 16672 14170
rect 16672 14118 16686 14170
rect 16710 14118 16724 14170
rect 16724 14118 16736 14170
rect 16736 14118 16766 14170
rect 16790 14118 16800 14170
rect 16800 14118 16846 14170
rect 16550 14116 16606 14118
rect 16630 14116 16686 14118
rect 16710 14116 16766 14118
rect 16790 14116 16846 14118
rect 17222 18264 17278 18320
rect 17682 20984 17738 21040
rect 16550 13082 16606 13084
rect 16630 13082 16686 13084
rect 16710 13082 16766 13084
rect 16790 13082 16846 13084
rect 16550 13030 16596 13082
rect 16596 13030 16606 13082
rect 16630 13030 16660 13082
rect 16660 13030 16672 13082
rect 16672 13030 16686 13082
rect 16710 13030 16724 13082
rect 16724 13030 16736 13082
rect 16736 13030 16766 13082
rect 16790 13030 16800 13082
rect 16800 13030 16846 13082
rect 16550 13028 16606 13030
rect 16630 13028 16686 13030
rect 16710 13028 16766 13030
rect 16790 13028 16846 13030
rect 16550 11994 16606 11996
rect 16630 11994 16686 11996
rect 16710 11994 16766 11996
rect 16790 11994 16846 11996
rect 16550 11942 16596 11994
rect 16596 11942 16606 11994
rect 16630 11942 16660 11994
rect 16660 11942 16672 11994
rect 16672 11942 16686 11994
rect 16710 11942 16724 11994
rect 16724 11942 16736 11994
rect 16736 11942 16766 11994
rect 16790 11942 16800 11994
rect 16800 11942 16846 11994
rect 16550 11940 16606 11942
rect 16630 11940 16686 11942
rect 16710 11940 16766 11942
rect 16790 11940 16846 11942
rect 16486 11736 16542 11792
rect 16302 11328 16358 11384
rect 16302 10240 16358 10296
rect 16550 10906 16606 10908
rect 16630 10906 16686 10908
rect 16710 10906 16766 10908
rect 16790 10906 16846 10908
rect 16550 10854 16596 10906
rect 16596 10854 16606 10906
rect 16630 10854 16660 10906
rect 16660 10854 16672 10906
rect 16672 10854 16686 10906
rect 16710 10854 16724 10906
rect 16724 10854 16736 10906
rect 16736 10854 16766 10906
rect 16790 10854 16800 10906
rect 16800 10854 16846 10906
rect 16550 10852 16606 10854
rect 16630 10852 16686 10854
rect 16710 10852 16766 10854
rect 16790 10852 16846 10854
rect 16762 10124 16818 10160
rect 16762 10104 16764 10124
rect 16764 10104 16816 10124
rect 16816 10104 16818 10124
rect 16550 9818 16606 9820
rect 16630 9818 16686 9820
rect 16710 9818 16766 9820
rect 16790 9818 16846 9820
rect 16550 9766 16596 9818
rect 16596 9766 16606 9818
rect 16630 9766 16660 9818
rect 16660 9766 16672 9818
rect 16672 9766 16686 9818
rect 16710 9766 16724 9818
rect 16724 9766 16736 9818
rect 16736 9766 16766 9818
rect 16790 9766 16800 9818
rect 16800 9766 16846 9818
rect 16550 9764 16606 9766
rect 16630 9764 16686 9766
rect 16710 9764 16766 9766
rect 16790 9764 16846 9766
rect 18234 26152 18290 26208
rect 18142 21800 18198 21856
rect 18142 19352 18198 19408
rect 17682 16904 17738 16960
rect 17958 16904 18014 16960
rect 18050 14864 18106 14920
rect 18050 14320 18106 14376
rect 17958 13640 18014 13696
rect 16394 8744 16450 8800
rect 16550 8730 16606 8732
rect 16630 8730 16686 8732
rect 16710 8730 16766 8732
rect 16790 8730 16846 8732
rect 16550 8678 16596 8730
rect 16596 8678 16606 8730
rect 16630 8678 16660 8730
rect 16660 8678 16672 8730
rect 16672 8678 16686 8730
rect 16710 8678 16724 8730
rect 16724 8678 16736 8730
rect 16736 8678 16766 8730
rect 16790 8678 16800 8730
rect 16800 8678 16846 8730
rect 16550 8676 16606 8678
rect 16630 8676 16686 8678
rect 16710 8676 16766 8678
rect 16790 8676 16846 8678
rect 16026 7792 16082 7848
rect 15382 5072 15438 5128
rect 14370 3052 14426 3088
rect 14370 3032 14372 3052
rect 14372 3032 14424 3052
rect 14424 3032 14426 3052
rect 13818 2896 13874 2952
rect 13951 2746 14007 2748
rect 14031 2746 14087 2748
rect 14111 2746 14167 2748
rect 14191 2746 14247 2748
rect 13951 2694 13997 2746
rect 13997 2694 14007 2746
rect 14031 2694 14061 2746
rect 14061 2694 14073 2746
rect 14073 2694 14087 2746
rect 14111 2694 14125 2746
rect 14125 2694 14137 2746
rect 14137 2694 14167 2746
rect 14191 2694 14201 2746
rect 14201 2694 14247 2746
rect 13951 2692 14007 2694
rect 14031 2692 14087 2694
rect 14111 2692 14167 2694
rect 14191 2692 14247 2694
rect 14370 2352 14426 2408
rect 14738 2896 14794 2952
rect 14554 2624 14610 2680
rect 13951 1658 14007 1660
rect 14031 1658 14087 1660
rect 14111 1658 14167 1660
rect 14191 1658 14247 1660
rect 13951 1606 13997 1658
rect 13997 1606 14007 1658
rect 14031 1606 14061 1658
rect 14061 1606 14073 1658
rect 14073 1606 14087 1658
rect 14111 1606 14125 1658
rect 14125 1606 14137 1658
rect 14137 1606 14167 1658
rect 14191 1606 14201 1658
rect 14201 1606 14247 1658
rect 13951 1604 14007 1606
rect 14031 1604 14087 1606
rect 14111 1604 14167 1606
rect 14191 1604 14247 1606
rect 14370 1400 14426 1456
rect 14554 1672 14610 1728
rect 16550 7642 16606 7644
rect 16630 7642 16686 7644
rect 16710 7642 16766 7644
rect 16790 7642 16846 7644
rect 16550 7590 16596 7642
rect 16596 7590 16606 7642
rect 16630 7590 16660 7642
rect 16660 7590 16672 7642
rect 16672 7590 16686 7642
rect 16710 7590 16724 7642
rect 16724 7590 16736 7642
rect 16736 7590 16766 7642
rect 16790 7590 16800 7642
rect 16800 7590 16846 7642
rect 16550 7588 16606 7590
rect 16630 7588 16686 7590
rect 16710 7588 16766 7590
rect 16790 7588 16846 7590
rect 16394 7520 16450 7576
rect 15750 5888 15806 5944
rect 15566 5480 15622 5536
rect 15934 4936 15990 4992
rect 17130 8916 17132 8936
rect 17132 8916 17184 8936
rect 17184 8916 17186 8936
rect 17130 8880 17186 8916
rect 17038 7384 17094 7440
rect 17498 12008 17554 12064
rect 16550 6554 16606 6556
rect 16630 6554 16686 6556
rect 16710 6554 16766 6556
rect 16790 6554 16846 6556
rect 16550 6502 16596 6554
rect 16596 6502 16606 6554
rect 16630 6502 16660 6554
rect 16660 6502 16672 6554
rect 16672 6502 16686 6554
rect 16710 6502 16724 6554
rect 16724 6502 16736 6554
rect 16736 6502 16766 6554
rect 16790 6502 16800 6554
rect 16800 6502 16846 6554
rect 16550 6500 16606 6502
rect 16630 6500 16686 6502
rect 16710 6500 16766 6502
rect 16790 6500 16846 6502
rect 16550 5466 16606 5468
rect 16630 5466 16686 5468
rect 16710 5466 16766 5468
rect 16790 5466 16846 5468
rect 16550 5414 16596 5466
rect 16596 5414 16606 5466
rect 16630 5414 16660 5466
rect 16660 5414 16672 5466
rect 16672 5414 16686 5466
rect 16710 5414 16724 5466
rect 16724 5414 16736 5466
rect 16736 5414 16766 5466
rect 16790 5414 16800 5466
rect 16800 5414 16846 5466
rect 16550 5412 16606 5414
rect 16630 5412 16686 5414
rect 16710 5412 16766 5414
rect 16790 5412 16846 5414
rect 15566 4664 15622 4720
rect 16118 4528 16174 4584
rect 15474 3576 15530 3632
rect 15106 3168 15162 3224
rect 14922 1536 14978 1592
rect 15658 3984 15714 4040
rect 16026 3848 16082 3904
rect 15750 3576 15806 3632
rect 15382 856 15438 912
rect 15842 3168 15898 3224
rect 15750 1536 15806 1592
rect 16118 2760 16174 2816
rect 16118 2624 16174 2680
rect 16302 4428 16304 4448
rect 16304 4428 16356 4448
rect 16356 4428 16358 4448
rect 16302 4392 16358 4428
rect 16550 4378 16606 4380
rect 16630 4378 16686 4380
rect 16710 4378 16766 4380
rect 16790 4378 16846 4380
rect 16550 4326 16596 4378
rect 16596 4326 16606 4378
rect 16630 4326 16660 4378
rect 16660 4326 16672 4378
rect 16672 4326 16686 4378
rect 16710 4326 16724 4378
rect 16724 4326 16736 4378
rect 16736 4326 16766 4378
rect 16790 4326 16800 4378
rect 16800 4326 16846 4378
rect 16550 4324 16606 4326
rect 16630 4324 16686 4326
rect 16710 4324 16766 4326
rect 16790 4324 16846 4326
rect 17222 4392 17278 4448
rect 16302 3440 16358 3496
rect 16302 3304 16358 3360
rect 16550 3290 16606 3292
rect 16630 3290 16686 3292
rect 16710 3290 16766 3292
rect 16790 3290 16846 3292
rect 16550 3238 16596 3290
rect 16596 3238 16606 3290
rect 16630 3238 16660 3290
rect 16660 3238 16672 3290
rect 16672 3238 16686 3290
rect 16710 3238 16724 3290
rect 16724 3238 16736 3290
rect 16736 3238 16766 3290
rect 16790 3238 16800 3290
rect 16800 3238 16846 3290
rect 16550 3236 16606 3238
rect 16630 3236 16686 3238
rect 16710 3236 16766 3238
rect 16790 3236 16846 3238
rect 16578 2624 16634 2680
rect 16550 2202 16606 2204
rect 16630 2202 16686 2204
rect 16710 2202 16766 2204
rect 16790 2202 16846 2204
rect 16550 2150 16596 2202
rect 16596 2150 16606 2202
rect 16630 2150 16660 2202
rect 16660 2150 16672 2202
rect 16672 2150 16686 2202
rect 16710 2150 16724 2202
rect 16724 2150 16736 2202
rect 16736 2150 16766 2202
rect 16790 2150 16800 2202
rect 16800 2150 16846 2202
rect 16550 2148 16606 2150
rect 16630 2148 16686 2150
rect 16710 2148 16766 2150
rect 16790 2148 16846 2150
rect 17590 11872 17646 11928
rect 17498 6568 17554 6624
rect 17682 9968 17738 10024
rect 17958 8492 18014 8528
rect 17958 8472 17960 8492
rect 17960 8472 18012 8492
rect 18012 8472 18014 8492
rect 18050 7792 18106 7848
rect 17774 7248 17830 7304
rect 17406 3304 17462 3360
rect 16854 1400 16910 1456
rect 16550 1114 16606 1116
rect 16630 1114 16686 1116
rect 16710 1114 16766 1116
rect 16790 1114 16846 1116
rect 16550 1062 16596 1114
rect 16596 1062 16606 1114
rect 16630 1062 16660 1114
rect 16660 1062 16672 1114
rect 16672 1062 16686 1114
rect 16710 1062 16724 1114
rect 16724 1062 16736 1114
rect 16736 1062 16766 1114
rect 16790 1062 16800 1114
rect 16800 1062 16846 1114
rect 16550 1060 16606 1062
rect 16630 1060 16686 1062
rect 16710 1060 16766 1062
rect 16790 1060 16846 1062
rect 17038 1672 17094 1728
rect 19890 40024 19946 40080
rect 18602 34448 18658 34504
rect 19338 39344 19394 39400
rect 19706 39208 19762 39264
rect 20626 41656 20682 41712
rect 20258 40568 20314 40624
rect 20442 41248 20498 41304
rect 20534 39208 20590 39264
rect 20258 38664 20314 38720
rect 19149 38650 19205 38652
rect 19229 38650 19285 38652
rect 19309 38650 19365 38652
rect 19389 38650 19445 38652
rect 19149 38598 19195 38650
rect 19195 38598 19205 38650
rect 19229 38598 19259 38650
rect 19259 38598 19271 38650
rect 19271 38598 19285 38650
rect 19309 38598 19323 38650
rect 19323 38598 19335 38650
rect 19335 38598 19365 38650
rect 19389 38598 19399 38650
rect 19399 38598 19445 38650
rect 19149 38596 19205 38598
rect 19229 38596 19285 38598
rect 19309 38596 19365 38598
rect 19389 38596 19445 38598
rect 19149 37562 19205 37564
rect 19229 37562 19285 37564
rect 19309 37562 19365 37564
rect 19389 37562 19445 37564
rect 19149 37510 19195 37562
rect 19195 37510 19205 37562
rect 19229 37510 19259 37562
rect 19259 37510 19271 37562
rect 19271 37510 19285 37562
rect 19309 37510 19323 37562
rect 19323 37510 19335 37562
rect 19335 37510 19365 37562
rect 19389 37510 19399 37562
rect 19399 37510 19445 37562
rect 19149 37508 19205 37510
rect 19229 37508 19285 37510
rect 19309 37508 19365 37510
rect 19389 37508 19445 37510
rect 19149 36474 19205 36476
rect 19229 36474 19285 36476
rect 19309 36474 19365 36476
rect 19389 36474 19445 36476
rect 19149 36422 19195 36474
rect 19195 36422 19205 36474
rect 19229 36422 19259 36474
rect 19259 36422 19271 36474
rect 19271 36422 19285 36474
rect 19309 36422 19323 36474
rect 19323 36422 19335 36474
rect 19335 36422 19365 36474
rect 19389 36422 19399 36474
rect 19399 36422 19445 36474
rect 19149 36420 19205 36422
rect 19229 36420 19285 36422
rect 19309 36420 19365 36422
rect 19389 36420 19445 36422
rect 19430 36216 19486 36272
rect 19149 35386 19205 35388
rect 19229 35386 19285 35388
rect 19309 35386 19365 35388
rect 19389 35386 19445 35388
rect 19149 35334 19195 35386
rect 19195 35334 19205 35386
rect 19229 35334 19259 35386
rect 19259 35334 19271 35386
rect 19271 35334 19285 35386
rect 19309 35334 19323 35386
rect 19323 35334 19335 35386
rect 19335 35334 19365 35386
rect 19389 35334 19399 35386
rect 19399 35334 19445 35386
rect 19149 35332 19205 35334
rect 19229 35332 19285 35334
rect 19309 35332 19365 35334
rect 19389 35332 19445 35334
rect 19982 38528 20038 38584
rect 20258 38256 20314 38312
rect 20074 37712 20130 37768
rect 20074 36760 20130 36816
rect 19982 36624 20038 36680
rect 19149 34298 19205 34300
rect 19229 34298 19285 34300
rect 19309 34298 19365 34300
rect 19389 34298 19445 34300
rect 19149 34246 19195 34298
rect 19195 34246 19205 34298
rect 19229 34246 19259 34298
rect 19259 34246 19271 34298
rect 19271 34246 19285 34298
rect 19309 34246 19323 34298
rect 19323 34246 19335 34298
rect 19335 34246 19365 34298
rect 19389 34246 19399 34298
rect 19399 34246 19445 34298
rect 19149 34244 19205 34246
rect 19229 34244 19285 34246
rect 19309 34244 19365 34246
rect 19389 34244 19445 34246
rect 19338 33516 19394 33552
rect 19338 33496 19340 33516
rect 19340 33496 19392 33516
rect 19392 33496 19394 33516
rect 19149 33210 19205 33212
rect 19229 33210 19285 33212
rect 19309 33210 19365 33212
rect 19389 33210 19445 33212
rect 19149 33158 19195 33210
rect 19195 33158 19205 33210
rect 19229 33158 19259 33210
rect 19259 33158 19271 33210
rect 19271 33158 19285 33210
rect 19309 33158 19323 33210
rect 19323 33158 19335 33210
rect 19335 33158 19365 33210
rect 19389 33158 19399 33210
rect 19399 33158 19445 33210
rect 19149 33156 19205 33158
rect 19229 33156 19285 33158
rect 19309 33156 19365 33158
rect 19389 33156 19445 33158
rect 18510 27376 18566 27432
rect 18970 32816 19026 32872
rect 18878 30776 18934 30832
rect 18418 24656 18474 24712
rect 18510 21936 18566 21992
rect 20166 35808 20222 35864
rect 20534 36760 20590 36816
rect 20534 36624 20590 36680
rect 20442 36216 20498 36272
rect 20442 35808 20498 35864
rect 20902 41112 20958 41168
rect 20902 40160 20958 40216
rect 22190 42472 22246 42528
rect 21748 42458 21804 42460
rect 21828 42458 21884 42460
rect 21908 42458 21964 42460
rect 21988 42458 22044 42460
rect 21748 42406 21794 42458
rect 21794 42406 21804 42458
rect 21828 42406 21858 42458
rect 21858 42406 21870 42458
rect 21870 42406 21884 42458
rect 21908 42406 21922 42458
rect 21922 42406 21934 42458
rect 21934 42406 21964 42458
rect 21988 42406 21998 42458
rect 21998 42406 22044 42458
rect 21748 42404 21804 42406
rect 21828 42404 21884 42406
rect 21908 42404 21964 42406
rect 21988 42404 22044 42406
rect 21914 41928 21970 41984
rect 22282 41384 22338 41440
rect 21748 41370 21804 41372
rect 21828 41370 21884 41372
rect 21908 41370 21964 41372
rect 21988 41370 22044 41372
rect 21748 41318 21794 41370
rect 21794 41318 21804 41370
rect 21828 41318 21858 41370
rect 21858 41318 21870 41370
rect 21870 41318 21884 41370
rect 21908 41318 21922 41370
rect 21922 41318 21934 41370
rect 21934 41318 21964 41370
rect 21988 41318 21998 41370
rect 21998 41318 22044 41370
rect 21748 41316 21804 41318
rect 21828 41316 21884 41318
rect 21908 41316 21964 41318
rect 21988 41316 22044 41318
rect 21546 40296 21602 40352
rect 21454 39788 21456 39808
rect 21456 39788 21508 39808
rect 21508 39788 21510 39808
rect 21454 39752 21510 39788
rect 21178 39344 21234 39400
rect 21454 38700 21456 38720
rect 21456 38700 21508 38720
rect 21508 38700 21510 38720
rect 21086 38528 21142 38584
rect 21454 38664 21510 38700
rect 21454 37612 21456 37632
rect 21456 37612 21508 37632
rect 21508 37612 21510 37632
rect 21454 37576 21510 37612
rect 21454 36524 21456 36544
rect 21456 36524 21508 36544
rect 21508 36524 21510 36544
rect 21454 36488 21510 36524
rect 19149 32122 19205 32124
rect 19229 32122 19285 32124
rect 19309 32122 19365 32124
rect 19389 32122 19445 32124
rect 19149 32070 19195 32122
rect 19195 32070 19205 32122
rect 19229 32070 19259 32122
rect 19259 32070 19271 32122
rect 19271 32070 19285 32122
rect 19309 32070 19323 32122
rect 19323 32070 19335 32122
rect 19335 32070 19365 32122
rect 19389 32070 19399 32122
rect 19399 32070 19445 32122
rect 19149 32068 19205 32070
rect 19229 32068 19285 32070
rect 19309 32068 19365 32070
rect 19389 32068 19445 32070
rect 19149 31034 19205 31036
rect 19229 31034 19285 31036
rect 19309 31034 19365 31036
rect 19389 31034 19445 31036
rect 19149 30982 19195 31034
rect 19195 30982 19205 31034
rect 19229 30982 19259 31034
rect 19259 30982 19271 31034
rect 19271 30982 19285 31034
rect 19309 30982 19323 31034
rect 19323 30982 19335 31034
rect 19335 30982 19365 31034
rect 19389 30982 19399 31034
rect 19399 30982 19445 31034
rect 19149 30980 19205 30982
rect 19229 30980 19285 30982
rect 19309 30980 19365 30982
rect 19389 30980 19445 30982
rect 19154 30676 19156 30696
rect 19156 30676 19208 30696
rect 19208 30676 19210 30696
rect 19154 30640 19210 30676
rect 19149 29946 19205 29948
rect 19229 29946 19285 29948
rect 19309 29946 19365 29948
rect 19389 29946 19445 29948
rect 19149 29894 19195 29946
rect 19195 29894 19205 29946
rect 19229 29894 19259 29946
rect 19259 29894 19271 29946
rect 19271 29894 19285 29946
rect 19309 29894 19323 29946
rect 19323 29894 19335 29946
rect 19335 29894 19365 29946
rect 19389 29894 19399 29946
rect 19399 29894 19445 29946
rect 19149 29892 19205 29894
rect 19229 29892 19285 29894
rect 19309 29892 19365 29894
rect 19389 29892 19445 29894
rect 18970 28872 19026 28928
rect 18878 26968 18934 27024
rect 19149 28858 19205 28860
rect 19229 28858 19285 28860
rect 19309 28858 19365 28860
rect 19389 28858 19445 28860
rect 19149 28806 19195 28858
rect 19195 28806 19205 28858
rect 19229 28806 19259 28858
rect 19259 28806 19271 28858
rect 19271 28806 19285 28858
rect 19309 28806 19323 28858
rect 19323 28806 19335 28858
rect 19335 28806 19365 28858
rect 19389 28806 19399 28858
rect 19399 28806 19445 28858
rect 19149 28804 19205 28806
rect 19229 28804 19285 28806
rect 19309 28804 19365 28806
rect 19389 28804 19445 28806
rect 19149 27770 19205 27772
rect 19229 27770 19285 27772
rect 19309 27770 19365 27772
rect 19389 27770 19445 27772
rect 19149 27718 19195 27770
rect 19195 27718 19205 27770
rect 19229 27718 19259 27770
rect 19259 27718 19271 27770
rect 19271 27718 19285 27770
rect 19309 27718 19323 27770
rect 19323 27718 19335 27770
rect 19335 27718 19365 27770
rect 19389 27718 19399 27770
rect 19399 27718 19445 27770
rect 19149 27716 19205 27718
rect 19229 27716 19285 27718
rect 19309 27716 19365 27718
rect 19389 27716 19445 27718
rect 19614 27920 19670 27976
rect 19149 26682 19205 26684
rect 19229 26682 19285 26684
rect 19309 26682 19365 26684
rect 19389 26682 19445 26684
rect 19149 26630 19195 26682
rect 19195 26630 19205 26682
rect 19229 26630 19259 26682
rect 19259 26630 19271 26682
rect 19271 26630 19285 26682
rect 19309 26630 19323 26682
rect 19323 26630 19335 26682
rect 19335 26630 19365 26682
rect 19389 26630 19399 26682
rect 19399 26630 19445 26682
rect 19149 26628 19205 26630
rect 19229 26628 19285 26630
rect 19309 26628 19365 26630
rect 19389 26628 19445 26630
rect 19149 25594 19205 25596
rect 19229 25594 19285 25596
rect 19309 25594 19365 25596
rect 19389 25594 19445 25596
rect 19149 25542 19195 25594
rect 19195 25542 19205 25594
rect 19229 25542 19259 25594
rect 19259 25542 19271 25594
rect 19271 25542 19285 25594
rect 19309 25542 19323 25594
rect 19323 25542 19335 25594
rect 19335 25542 19365 25594
rect 19389 25542 19399 25594
rect 19399 25542 19445 25594
rect 19149 25540 19205 25542
rect 19229 25540 19285 25542
rect 19309 25540 19365 25542
rect 19389 25540 19445 25542
rect 20074 31864 20130 31920
rect 19982 31320 20038 31376
rect 19890 26288 19946 26344
rect 19149 24506 19205 24508
rect 19229 24506 19285 24508
rect 19309 24506 19365 24508
rect 19389 24506 19445 24508
rect 19149 24454 19195 24506
rect 19195 24454 19205 24506
rect 19229 24454 19259 24506
rect 19259 24454 19271 24506
rect 19271 24454 19285 24506
rect 19309 24454 19323 24506
rect 19323 24454 19335 24506
rect 19335 24454 19365 24506
rect 19389 24454 19399 24506
rect 19399 24454 19445 24506
rect 19149 24452 19205 24454
rect 19229 24452 19285 24454
rect 19309 24452 19365 24454
rect 19389 24452 19445 24454
rect 18694 20712 18750 20768
rect 18326 19624 18382 19680
rect 18694 19352 18750 19408
rect 18326 13232 18382 13288
rect 19338 23724 19394 23760
rect 19338 23704 19340 23724
rect 19340 23704 19392 23724
rect 19392 23704 19394 23724
rect 19522 23432 19578 23488
rect 19149 23418 19205 23420
rect 19229 23418 19285 23420
rect 19309 23418 19365 23420
rect 19389 23418 19445 23420
rect 19149 23366 19195 23418
rect 19195 23366 19205 23418
rect 19229 23366 19259 23418
rect 19259 23366 19271 23418
rect 19271 23366 19285 23418
rect 19309 23366 19323 23418
rect 19323 23366 19335 23418
rect 19335 23366 19365 23418
rect 19389 23366 19399 23418
rect 19399 23366 19445 23418
rect 19149 23364 19205 23366
rect 19229 23364 19285 23366
rect 19309 23364 19365 23366
rect 19389 23364 19445 23366
rect 19522 23316 19578 23352
rect 19522 23296 19524 23316
rect 19524 23296 19576 23316
rect 19576 23296 19578 23316
rect 19338 23060 19340 23080
rect 19340 23060 19392 23080
rect 19392 23060 19394 23080
rect 19338 23024 19394 23060
rect 19338 22924 19346 22944
rect 19346 22924 19394 22944
rect 19338 22888 19394 22924
rect 19338 22752 19394 22808
rect 19149 22330 19205 22332
rect 19229 22330 19285 22332
rect 19309 22330 19365 22332
rect 19389 22330 19445 22332
rect 19149 22278 19195 22330
rect 19195 22278 19205 22330
rect 19229 22278 19259 22330
rect 19259 22278 19271 22330
rect 19271 22278 19285 22330
rect 19309 22278 19323 22330
rect 19323 22278 19335 22330
rect 19335 22278 19365 22330
rect 19389 22278 19399 22330
rect 19399 22278 19445 22330
rect 19149 22276 19205 22278
rect 19229 22276 19285 22278
rect 19309 22276 19365 22278
rect 19389 22276 19445 22278
rect 19890 23432 19946 23488
rect 19890 22888 19946 22944
rect 19798 22072 19854 22128
rect 20258 30232 20314 30288
rect 20442 31864 20498 31920
rect 20534 30368 20590 30424
rect 20074 29008 20130 29064
rect 20534 30232 20590 30288
rect 20258 24248 20314 24304
rect 21454 35436 21456 35456
rect 21456 35436 21508 35456
rect 21508 35436 21510 35456
rect 21454 35400 21510 35436
rect 21454 34348 21456 34368
rect 21456 34348 21508 34368
rect 21508 34348 21510 34368
rect 21454 34312 21510 34348
rect 21270 33260 21272 33280
rect 21272 33260 21324 33280
rect 21324 33260 21326 33280
rect 21270 33224 21326 33260
rect 21178 32952 21234 33008
rect 21546 33632 21602 33688
rect 22190 40876 22192 40896
rect 22192 40876 22244 40896
rect 22244 40876 22246 40896
rect 22190 40840 22246 40876
rect 22190 40332 22192 40352
rect 22192 40332 22244 40352
rect 22244 40332 22246 40352
rect 22190 40296 22246 40332
rect 21748 40282 21804 40284
rect 21828 40282 21884 40284
rect 21908 40282 21964 40284
rect 21988 40282 22044 40284
rect 21748 40230 21794 40282
rect 21794 40230 21804 40282
rect 21828 40230 21858 40282
rect 21858 40230 21870 40282
rect 21870 40230 21884 40282
rect 21908 40230 21922 40282
rect 21922 40230 21934 40282
rect 21934 40230 21964 40282
rect 21988 40230 21998 40282
rect 21998 40230 22044 40282
rect 21748 40228 21804 40230
rect 21828 40228 21884 40230
rect 21908 40228 21964 40230
rect 21988 40228 22044 40230
rect 22190 39244 22192 39264
rect 22192 39244 22244 39264
rect 22244 39244 22246 39264
rect 22190 39208 22246 39244
rect 21748 39194 21804 39196
rect 21828 39194 21884 39196
rect 21908 39194 21964 39196
rect 21988 39194 22044 39196
rect 21748 39142 21794 39194
rect 21794 39142 21804 39194
rect 21828 39142 21858 39194
rect 21858 39142 21870 39194
rect 21870 39142 21884 39194
rect 21908 39142 21922 39194
rect 21922 39142 21934 39194
rect 21934 39142 21964 39194
rect 21988 39142 21998 39194
rect 21998 39142 22044 39194
rect 21748 39140 21804 39142
rect 21828 39140 21884 39142
rect 21908 39140 21964 39142
rect 21988 39140 22044 39142
rect 22190 38156 22192 38176
rect 22192 38156 22244 38176
rect 22244 38156 22246 38176
rect 22190 38120 22246 38156
rect 21748 38106 21804 38108
rect 21828 38106 21884 38108
rect 21908 38106 21964 38108
rect 21988 38106 22044 38108
rect 21748 38054 21794 38106
rect 21794 38054 21804 38106
rect 21828 38054 21858 38106
rect 21858 38054 21870 38106
rect 21870 38054 21884 38106
rect 21908 38054 21922 38106
rect 21922 38054 21934 38106
rect 21934 38054 21964 38106
rect 21988 38054 21998 38106
rect 21998 38054 22044 38106
rect 21748 38052 21804 38054
rect 21828 38052 21884 38054
rect 21908 38052 21964 38054
rect 21988 38052 22044 38054
rect 22282 37032 22338 37088
rect 21748 37018 21804 37020
rect 21828 37018 21884 37020
rect 21908 37018 21964 37020
rect 21988 37018 22044 37020
rect 21748 36966 21794 37018
rect 21794 36966 21804 37018
rect 21828 36966 21858 37018
rect 21858 36966 21870 37018
rect 21870 36966 21884 37018
rect 21908 36966 21922 37018
rect 21922 36966 21934 37018
rect 21934 36966 21964 37018
rect 21988 36966 21998 37018
rect 21998 36966 22044 37018
rect 21748 36964 21804 36966
rect 21828 36964 21884 36966
rect 21908 36964 21964 36966
rect 21988 36964 22044 36966
rect 22282 35944 22338 36000
rect 21748 35930 21804 35932
rect 21828 35930 21884 35932
rect 21908 35930 21964 35932
rect 21988 35930 22044 35932
rect 21748 35878 21794 35930
rect 21794 35878 21804 35930
rect 21828 35878 21858 35930
rect 21858 35878 21870 35930
rect 21870 35878 21884 35930
rect 21908 35878 21922 35930
rect 21922 35878 21934 35930
rect 21934 35878 21964 35930
rect 21988 35878 21998 35930
rect 21998 35878 22044 35930
rect 21748 35876 21804 35878
rect 21828 35876 21884 35878
rect 21908 35876 21964 35878
rect 21988 35876 22044 35878
rect 21748 34842 21804 34844
rect 21828 34842 21884 34844
rect 21908 34842 21964 34844
rect 21988 34842 22044 34844
rect 21748 34790 21794 34842
rect 21794 34790 21804 34842
rect 21828 34790 21858 34842
rect 21858 34790 21870 34842
rect 21870 34790 21884 34842
rect 21908 34790 21922 34842
rect 21922 34790 21934 34842
rect 21934 34790 21964 34842
rect 21988 34790 21998 34842
rect 21998 34790 22044 34842
rect 21748 34788 21804 34790
rect 21828 34788 21884 34790
rect 21908 34788 21964 34790
rect 21988 34788 22044 34790
rect 21748 33754 21804 33756
rect 21828 33754 21884 33756
rect 21908 33754 21964 33756
rect 21988 33754 22044 33756
rect 21748 33702 21794 33754
rect 21794 33702 21804 33754
rect 21828 33702 21858 33754
rect 21858 33702 21870 33754
rect 21870 33702 21884 33754
rect 21908 33702 21922 33754
rect 21922 33702 21934 33754
rect 21934 33702 21964 33754
rect 21988 33702 21998 33754
rect 21998 33702 22044 33754
rect 21748 33700 21804 33702
rect 21828 33700 21884 33702
rect 21908 33700 21964 33702
rect 21988 33700 22044 33702
rect 22190 34892 22192 34912
rect 22192 34892 22244 34912
rect 22244 34892 22246 34912
rect 22190 34856 22246 34892
rect 22190 33804 22192 33824
rect 22192 33804 22244 33824
rect 22244 33804 22246 33824
rect 22190 33768 22246 33804
rect 21454 32172 21456 32192
rect 21456 32172 21508 32192
rect 21508 32172 21510 32192
rect 21454 32136 21510 32172
rect 21546 31864 21602 31920
rect 21454 31084 21456 31104
rect 21456 31084 21508 31104
rect 21508 31084 21510 31104
rect 21454 31048 21510 31084
rect 21270 30912 21326 30968
rect 20350 23432 20406 23488
rect 20626 23296 20682 23352
rect 20350 23024 20406 23080
rect 20258 22616 20314 22672
rect 19149 21242 19205 21244
rect 19229 21242 19285 21244
rect 19309 21242 19365 21244
rect 19389 21242 19445 21244
rect 19149 21190 19195 21242
rect 19195 21190 19205 21242
rect 19229 21190 19259 21242
rect 19259 21190 19271 21242
rect 19271 21190 19285 21242
rect 19309 21190 19323 21242
rect 19323 21190 19335 21242
rect 19335 21190 19365 21242
rect 19389 21190 19399 21242
rect 19399 21190 19445 21242
rect 19149 21188 19205 21190
rect 19229 21188 19285 21190
rect 19309 21188 19365 21190
rect 19389 21188 19445 21190
rect 19149 20154 19205 20156
rect 19229 20154 19285 20156
rect 19309 20154 19365 20156
rect 19389 20154 19445 20156
rect 19149 20102 19195 20154
rect 19195 20102 19205 20154
rect 19229 20102 19259 20154
rect 19259 20102 19271 20154
rect 19271 20102 19285 20154
rect 19309 20102 19323 20154
rect 19323 20102 19335 20154
rect 19335 20102 19365 20154
rect 19389 20102 19399 20154
rect 19399 20102 19445 20154
rect 19149 20100 19205 20102
rect 19229 20100 19285 20102
rect 19309 20100 19365 20102
rect 19389 20100 19445 20102
rect 19149 19066 19205 19068
rect 19229 19066 19285 19068
rect 19309 19066 19365 19068
rect 19389 19066 19445 19068
rect 19149 19014 19195 19066
rect 19195 19014 19205 19066
rect 19229 19014 19259 19066
rect 19259 19014 19271 19066
rect 19271 19014 19285 19066
rect 19309 19014 19323 19066
rect 19323 19014 19335 19066
rect 19335 19014 19365 19066
rect 19389 19014 19399 19066
rect 19399 19014 19445 19066
rect 19149 19012 19205 19014
rect 19229 19012 19285 19014
rect 19309 19012 19365 19014
rect 19389 19012 19445 19014
rect 19149 17978 19205 17980
rect 19229 17978 19285 17980
rect 19309 17978 19365 17980
rect 19389 17978 19445 17980
rect 19149 17926 19195 17978
rect 19195 17926 19205 17978
rect 19229 17926 19259 17978
rect 19259 17926 19271 17978
rect 19271 17926 19285 17978
rect 19309 17926 19323 17978
rect 19323 17926 19335 17978
rect 19335 17926 19365 17978
rect 19389 17926 19399 17978
rect 19399 17926 19445 17978
rect 19149 17924 19205 17926
rect 19229 17924 19285 17926
rect 19309 17924 19365 17926
rect 19389 17924 19445 17926
rect 18786 16496 18842 16552
rect 18694 15408 18750 15464
rect 19149 16890 19205 16892
rect 19229 16890 19285 16892
rect 19309 16890 19365 16892
rect 19389 16890 19445 16892
rect 19149 16838 19195 16890
rect 19195 16838 19205 16890
rect 19229 16838 19259 16890
rect 19259 16838 19271 16890
rect 19271 16838 19285 16890
rect 19309 16838 19323 16890
rect 19323 16838 19335 16890
rect 19335 16838 19365 16890
rect 19389 16838 19399 16890
rect 19399 16838 19445 16890
rect 19149 16836 19205 16838
rect 19229 16836 19285 16838
rect 19309 16836 19365 16838
rect 19389 16836 19445 16838
rect 19246 15972 19302 16008
rect 19246 15952 19248 15972
rect 19248 15952 19300 15972
rect 19300 15952 19302 15972
rect 19149 15802 19205 15804
rect 19229 15802 19285 15804
rect 19309 15802 19365 15804
rect 19389 15802 19445 15804
rect 19149 15750 19195 15802
rect 19195 15750 19205 15802
rect 19229 15750 19259 15802
rect 19259 15750 19271 15802
rect 19271 15750 19285 15802
rect 19309 15750 19323 15802
rect 19323 15750 19335 15802
rect 19335 15750 19365 15802
rect 19389 15750 19399 15802
rect 19399 15750 19445 15802
rect 19149 15748 19205 15750
rect 19229 15748 19285 15750
rect 19309 15748 19365 15750
rect 19389 15748 19445 15750
rect 19706 17720 19762 17776
rect 18326 12144 18382 12200
rect 18786 11736 18842 11792
rect 18418 9968 18474 10024
rect 18602 9016 18658 9072
rect 18418 7792 18474 7848
rect 18234 6432 18290 6488
rect 18234 6316 18290 6352
rect 18234 6296 18236 6316
rect 18236 6296 18288 6316
rect 18288 6296 18290 6316
rect 19149 14714 19205 14716
rect 19229 14714 19285 14716
rect 19309 14714 19365 14716
rect 19389 14714 19445 14716
rect 19149 14662 19195 14714
rect 19195 14662 19205 14714
rect 19229 14662 19259 14714
rect 19259 14662 19271 14714
rect 19271 14662 19285 14714
rect 19309 14662 19323 14714
rect 19323 14662 19335 14714
rect 19335 14662 19365 14714
rect 19389 14662 19399 14714
rect 19399 14662 19445 14714
rect 19149 14660 19205 14662
rect 19229 14660 19285 14662
rect 19309 14660 19365 14662
rect 19389 14660 19445 14662
rect 19149 13626 19205 13628
rect 19229 13626 19285 13628
rect 19309 13626 19365 13628
rect 19389 13626 19445 13628
rect 19149 13574 19195 13626
rect 19195 13574 19205 13626
rect 19229 13574 19259 13626
rect 19259 13574 19271 13626
rect 19271 13574 19285 13626
rect 19309 13574 19323 13626
rect 19323 13574 19335 13626
rect 19335 13574 19365 13626
rect 19389 13574 19399 13626
rect 19399 13574 19445 13626
rect 19149 13572 19205 13574
rect 19229 13572 19285 13574
rect 19309 13572 19365 13574
rect 19389 13572 19445 13574
rect 19149 12538 19205 12540
rect 19229 12538 19285 12540
rect 19309 12538 19365 12540
rect 19389 12538 19445 12540
rect 19149 12486 19195 12538
rect 19195 12486 19205 12538
rect 19229 12486 19259 12538
rect 19259 12486 19271 12538
rect 19271 12486 19285 12538
rect 19309 12486 19323 12538
rect 19323 12486 19335 12538
rect 19335 12486 19365 12538
rect 19389 12486 19399 12538
rect 19399 12486 19445 12538
rect 19149 12484 19205 12486
rect 19229 12484 19285 12486
rect 19309 12484 19365 12486
rect 19389 12484 19445 12486
rect 18878 9696 18934 9752
rect 19062 12280 19118 12336
rect 19798 16496 19854 16552
rect 21086 27820 21088 27840
rect 21088 27820 21140 27840
rect 21140 27820 21142 27840
rect 21086 27784 21142 27820
rect 20810 21256 20866 21312
rect 20074 19624 20130 19680
rect 19982 19216 20038 19272
rect 19982 13096 20038 13152
rect 19149 11450 19205 11452
rect 19229 11450 19285 11452
rect 19309 11450 19365 11452
rect 19389 11450 19445 11452
rect 19149 11398 19195 11450
rect 19195 11398 19205 11450
rect 19229 11398 19259 11450
rect 19259 11398 19271 11450
rect 19271 11398 19285 11450
rect 19309 11398 19323 11450
rect 19323 11398 19335 11450
rect 19335 11398 19365 11450
rect 19389 11398 19399 11450
rect 19399 11398 19445 11450
rect 19149 11396 19205 11398
rect 19229 11396 19285 11398
rect 19309 11396 19365 11398
rect 19389 11396 19445 11398
rect 19614 10648 19670 10704
rect 19149 10362 19205 10364
rect 19229 10362 19285 10364
rect 19309 10362 19365 10364
rect 19389 10362 19445 10364
rect 19149 10310 19195 10362
rect 19195 10310 19205 10362
rect 19229 10310 19259 10362
rect 19259 10310 19271 10362
rect 19271 10310 19285 10362
rect 19309 10310 19323 10362
rect 19323 10310 19335 10362
rect 19335 10310 19365 10362
rect 19389 10310 19399 10362
rect 19399 10310 19445 10362
rect 19149 10308 19205 10310
rect 19229 10308 19285 10310
rect 19309 10308 19365 10310
rect 19389 10308 19445 10310
rect 19246 9560 19302 9616
rect 19149 9274 19205 9276
rect 19229 9274 19285 9276
rect 19309 9274 19365 9276
rect 19389 9274 19445 9276
rect 19149 9222 19195 9274
rect 19195 9222 19205 9274
rect 19229 9222 19259 9274
rect 19259 9222 19271 9274
rect 19271 9222 19285 9274
rect 19309 9222 19323 9274
rect 19323 9222 19335 9274
rect 19335 9222 19365 9274
rect 19389 9222 19399 9274
rect 19399 9222 19445 9274
rect 19149 9220 19205 9222
rect 19229 9220 19285 9222
rect 19309 9220 19365 9222
rect 19389 9220 19445 9222
rect 20074 11600 20130 11656
rect 19062 9016 19118 9072
rect 19338 8880 19394 8936
rect 18970 8200 19026 8256
rect 19149 8186 19205 8188
rect 19229 8186 19285 8188
rect 19309 8186 19365 8188
rect 19389 8186 19445 8188
rect 19149 8134 19195 8186
rect 19195 8134 19205 8186
rect 19229 8134 19259 8186
rect 19259 8134 19271 8186
rect 19271 8134 19285 8186
rect 19309 8134 19323 8186
rect 19323 8134 19335 8186
rect 19335 8134 19365 8186
rect 19389 8134 19399 8186
rect 19399 8134 19445 8186
rect 19149 8132 19205 8134
rect 19229 8132 19285 8134
rect 19309 8132 19365 8134
rect 19389 8132 19445 8134
rect 18878 8064 18934 8120
rect 18786 7656 18842 7712
rect 18694 6296 18750 6352
rect 18970 7248 19026 7304
rect 18878 6976 18934 7032
rect 18602 6024 18658 6080
rect 18326 5616 18382 5672
rect 18418 5480 18474 5536
rect 18234 4392 18290 4448
rect 18234 4256 18290 4312
rect 18050 3984 18106 4040
rect 18234 3984 18290 4040
rect 18050 3340 18052 3360
rect 18052 3340 18104 3360
rect 18104 3340 18106 3360
rect 18050 3304 18106 3340
rect 18418 4936 18474 4992
rect 18418 3732 18474 3768
rect 18694 5888 18750 5944
rect 19149 7098 19205 7100
rect 19229 7098 19285 7100
rect 19309 7098 19365 7100
rect 19389 7098 19445 7100
rect 19149 7046 19195 7098
rect 19195 7046 19205 7098
rect 19229 7046 19259 7098
rect 19259 7046 19271 7098
rect 19271 7046 19285 7098
rect 19309 7046 19323 7098
rect 19323 7046 19335 7098
rect 19335 7046 19365 7098
rect 19389 7046 19399 7098
rect 19399 7046 19445 7098
rect 19149 7044 19205 7046
rect 19229 7044 19285 7046
rect 19309 7044 19365 7046
rect 19389 7044 19445 7046
rect 18786 5652 18788 5672
rect 18788 5652 18840 5672
rect 18840 5652 18842 5672
rect 18786 5616 18842 5652
rect 18602 4800 18658 4856
rect 19154 6432 19210 6488
rect 19246 6296 19302 6352
rect 19149 6010 19205 6012
rect 19229 6010 19285 6012
rect 19309 6010 19365 6012
rect 19389 6010 19445 6012
rect 19149 5958 19195 6010
rect 19195 5958 19205 6010
rect 19229 5958 19259 6010
rect 19259 5958 19271 6010
rect 19271 5958 19285 6010
rect 19309 5958 19323 6010
rect 19323 5958 19335 6010
rect 19335 5958 19365 6010
rect 19389 5958 19399 6010
rect 19399 5958 19445 6010
rect 19149 5956 19205 5958
rect 19229 5956 19285 5958
rect 19309 5956 19365 5958
rect 19389 5956 19445 5958
rect 21454 29996 21456 30016
rect 21456 29996 21508 30016
rect 21508 29996 21510 30016
rect 21454 29960 21510 29996
rect 21454 28908 21456 28928
rect 21456 28908 21508 28928
rect 21508 28908 21510 28928
rect 21454 28872 21510 28908
rect 21454 26968 21510 27024
rect 21454 25644 21456 25664
rect 21456 25644 21508 25664
rect 21508 25644 21510 25664
rect 21454 25608 21510 25644
rect 21454 24556 21456 24576
rect 21456 24556 21508 24576
rect 21508 24556 21510 24576
rect 21454 24520 21510 24556
rect 21748 32666 21804 32668
rect 21828 32666 21884 32668
rect 21908 32666 21964 32668
rect 21988 32666 22044 32668
rect 21748 32614 21794 32666
rect 21794 32614 21804 32666
rect 21828 32614 21858 32666
rect 21858 32614 21870 32666
rect 21870 32614 21884 32666
rect 21908 32614 21922 32666
rect 21922 32614 21934 32666
rect 21934 32614 21964 32666
rect 21988 32614 21998 32666
rect 21998 32614 22044 32666
rect 21748 32612 21804 32614
rect 21828 32612 21884 32614
rect 21908 32612 21964 32614
rect 21988 32612 22044 32614
rect 21748 31578 21804 31580
rect 21828 31578 21884 31580
rect 21908 31578 21964 31580
rect 21988 31578 22044 31580
rect 21748 31526 21794 31578
rect 21794 31526 21804 31578
rect 21828 31526 21858 31578
rect 21858 31526 21870 31578
rect 21870 31526 21884 31578
rect 21908 31526 21922 31578
rect 21922 31526 21934 31578
rect 21934 31526 21964 31578
rect 21988 31526 21998 31578
rect 21998 31526 22044 31578
rect 21748 31524 21804 31526
rect 21828 31524 21884 31526
rect 21908 31524 21964 31526
rect 21988 31524 22044 31526
rect 21748 30490 21804 30492
rect 21828 30490 21884 30492
rect 21908 30490 21964 30492
rect 21988 30490 22044 30492
rect 21748 30438 21794 30490
rect 21794 30438 21804 30490
rect 21828 30438 21858 30490
rect 21858 30438 21870 30490
rect 21870 30438 21884 30490
rect 21908 30438 21922 30490
rect 21922 30438 21934 30490
rect 21934 30438 21964 30490
rect 21988 30438 21998 30490
rect 21998 30438 22044 30490
rect 21748 30436 21804 30438
rect 21828 30436 21884 30438
rect 21908 30436 21964 30438
rect 21988 30436 22044 30438
rect 21748 29402 21804 29404
rect 21828 29402 21884 29404
rect 21908 29402 21964 29404
rect 21988 29402 22044 29404
rect 21748 29350 21794 29402
rect 21794 29350 21804 29402
rect 21828 29350 21858 29402
rect 21858 29350 21870 29402
rect 21870 29350 21884 29402
rect 21908 29350 21922 29402
rect 21922 29350 21934 29402
rect 21934 29350 21964 29402
rect 21988 29350 21998 29402
rect 21998 29350 22044 29402
rect 21748 29348 21804 29350
rect 21828 29348 21884 29350
rect 21908 29348 21964 29350
rect 21988 29348 22044 29350
rect 21748 28314 21804 28316
rect 21828 28314 21884 28316
rect 21908 28314 21964 28316
rect 21988 28314 22044 28316
rect 21748 28262 21794 28314
rect 21794 28262 21804 28314
rect 21828 28262 21858 28314
rect 21858 28262 21870 28314
rect 21870 28262 21884 28314
rect 21908 28262 21922 28314
rect 21922 28262 21934 28314
rect 21934 28262 21964 28314
rect 21988 28262 21998 28314
rect 21998 28262 22044 28314
rect 21748 28260 21804 28262
rect 21828 28260 21884 28262
rect 21908 28260 21964 28262
rect 21988 28260 22044 28262
rect 21546 23432 21602 23488
rect 21546 22752 21602 22808
rect 21748 27226 21804 27228
rect 21828 27226 21884 27228
rect 21908 27226 21964 27228
rect 21988 27226 22044 27228
rect 21748 27174 21794 27226
rect 21794 27174 21804 27226
rect 21828 27174 21858 27226
rect 21858 27174 21870 27226
rect 21870 27174 21884 27226
rect 21908 27174 21922 27226
rect 21922 27174 21934 27226
rect 21934 27174 21964 27226
rect 21988 27174 21998 27226
rect 21998 27174 22044 27226
rect 21748 27172 21804 27174
rect 21828 27172 21884 27174
rect 21908 27172 21964 27174
rect 21988 27172 22044 27174
rect 21748 26138 21804 26140
rect 21828 26138 21884 26140
rect 21908 26138 21964 26140
rect 21988 26138 22044 26140
rect 21748 26086 21794 26138
rect 21794 26086 21804 26138
rect 21828 26086 21858 26138
rect 21858 26086 21870 26138
rect 21870 26086 21884 26138
rect 21908 26086 21922 26138
rect 21922 26086 21934 26138
rect 21934 26086 21964 26138
rect 21988 26086 21998 26138
rect 21998 26086 22044 26138
rect 21748 26084 21804 26086
rect 21828 26084 21884 26086
rect 21908 26084 21964 26086
rect 21988 26084 22044 26086
rect 21748 25050 21804 25052
rect 21828 25050 21884 25052
rect 21908 25050 21964 25052
rect 21988 25050 22044 25052
rect 21748 24998 21794 25050
rect 21794 24998 21804 25050
rect 21828 24998 21858 25050
rect 21858 24998 21870 25050
rect 21870 24998 21884 25050
rect 21908 24998 21922 25050
rect 21922 24998 21934 25050
rect 21934 24998 21964 25050
rect 21988 24998 21998 25050
rect 21998 24998 22044 25050
rect 21748 24996 21804 24998
rect 21828 24996 21884 24998
rect 21908 24996 21964 24998
rect 21988 24996 22044 24998
rect 22190 31628 22192 31648
rect 22192 31628 22244 31648
rect 22244 31628 22246 31648
rect 22190 31592 22246 31628
rect 22282 30504 22338 30560
rect 22190 29452 22192 29472
rect 22192 29452 22244 29472
rect 22244 29452 22246 29472
rect 22190 29416 22246 29452
rect 22190 28364 22192 28384
rect 22192 28364 22244 28384
rect 22244 28364 22246 28384
rect 22190 28328 22246 28364
rect 22190 27240 22246 27296
rect 22282 26152 22338 26208
rect 22282 25064 22338 25120
rect 21748 23962 21804 23964
rect 21828 23962 21884 23964
rect 21908 23962 21964 23964
rect 21988 23962 22044 23964
rect 21748 23910 21794 23962
rect 21794 23910 21804 23962
rect 21828 23910 21858 23962
rect 21858 23910 21870 23962
rect 21870 23910 21884 23962
rect 21908 23910 21922 23962
rect 21922 23910 21934 23962
rect 21934 23910 21964 23962
rect 21988 23910 21998 23962
rect 21998 23910 22044 23962
rect 21748 23908 21804 23910
rect 21828 23908 21884 23910
rect 21908 23908 21964 23910
rect 21988 23908 22044 23910
rect 21748 22874 21804 22876
rect 21828 22874 21884 22876
rect 21908 22874 21964 22876
rect 21988 22874 22044 22876
rect 21748 22822 21794 22874
rect 21794 22822 21804 22874
rect 21828 22822 21858 22874
rect 21858 22822 21870 22874
rect 21870 22822 21884 22874
rect 21908 22822 21922 22874
rect 21922 22822 21934 22874
rect 21934 22822 21964 22874
rect 21988 22822 21998 22874
rect 21998 22822 22044 22874
rect 21748 22820 21804 22822
rect 21828 22820 21884 22822
rect 21908 22820 21964 22822
rect 21988 22820 22044 22822
rect 22190 24012 22192 24032
rect 22192 24012 22244 24032
rect 22244 24012 22246 24032
rect 22190 23976 22246 24012
rect 22190 22888 22246 22944
rect 21454 22344 21510 22400
rect 21546 22072 21602 22128
rect 22190 22616 22246 22672
rect 22098 22480 22154 22536
rect 22006 22072 22062 22128
rect 21270 20712 21326 20768
rect 21454 20204 21456 20224
rect 21456 20204 21508 20224
rect 21508 20204 21510 20224
rect 21454 20168 21510 20204
rect 21362 19352 21418 19408
rect 21270 17176 21326 17232
rect 20810 15272 20866 15328
rect 21178 13912 21234 13968
rect 21086 12588 21088 12608
rect 21088 12588 21140 12608
rect 21140 12588 21142 12608
rect 21086 12552 21142 12588
rect 20810 12280 20866 12336
rect 20258 8880 20314 8936
rect 19798 7928 19854 7984
rect 19154 5616 19210 5672
rect 19149 4922 19205 4924
rect 19229 4922 19285 4924
rect 19309 4922 19365 4924
rect 19389 4922 19445 4924
rect 19149 4870 19195 4922
rect 19195 4870 19205 4922
rect 19229 4870 19259 4922
rect 19259 4870 19271 4922
rect 19271 4870 19285 4922
rect 19309 4870 19323 4922
rect 19323 4870 19335 4922
rect 19335 4870 19365 4922
rect 19389 4870 19399 4922
rect 19399 4870 19445 4922
rect 19149 4868 19205 4870
rect 19229 4868 19285 4870
rect 19309 4868 19365 4870
rect 19389 4868 19445 4870
rect 18878 3848 18934 3904
rect 18418 3712 18420 3732
rect 18420 3712 18472 3732
rect 18472 3712 18474 3732
rect 18326 3304 18382 3360
rect 17958 2896 18014 2952
rect 18602 3168 18658 3224
rect 17590 2508 17646 2544
rect 17590 2488 17592 2508
rect 17592 2488 17644 2508
rect 17644 2488 17646 2508
rect 18142 1536 18198 1592
rect 18602 2760 18658 2816
rect 18510 2624 18566 2680
rect 18694 2488 18750 2544
rect 18694 2388 18696 2408
rect 18696 2388 18748 2408
rect 18748 2388 18750 2408
rect 18694 2352 18750 2388
rect 19522 4564 19524 4584
rect 19524 4564 19576 4584
rect 19576 4564 19578 4584
rect 19522 4528 19578 4564
rect 19246 3984 19302 4040
rect 19149 3834 19205 3836
rect 19229 3834 19285 3836
rect 19309 3834 19365 3836
rect 19389 3834 19445 3836
rect 19149 3782 19195 3834
rect 19195 3782 19205 3834
rect 19229 3782 19259 3834
rect 19259 3782 19271 3834
rect 19271 3782 19285 3834
rect 19309 3782 19323 3834
rect 19323 3782 19335 3834
rect 19335 3782 19365 3834
rect 19389 3782 19399 3834
rect 19399 3782 19445 3834
rect 19149 3780 19205 3782
rect 19229 3780 19285 3782
rect 19309 3780 19365 3782
rect 19389 3780 19445 3782
rect 18970 1944 19026 2000
rect 19149 2746 19205 2748
rect 19229 2746 19285 2748
rect 19309 2746 19365 2748
rect 19389 2746 19445 2748
rect 19149 2694 19195 2746
rect 19195 2694 19205 2746
rect 19229 2694 19259 2746
rect 19259 2694 19271 2746
rect 19271 2694 19285 2746
rect 19309 2694 19323 2746
rect 19323 2694 19335 2746
rect 19335 2694 19365 2746
rect 19389 2694 19399 2746
rect 19399 2694 19445 2746
rect 19149 2692 19205 2694
rect 19229 2692 19285 2694
rect 19309 2692 19365 2694
rect 19389 2692 19445 2694
rect 19149 1658 19205 1660
rect 19229 1658 19285 1660
rect 19309 1658 19365 1660
rect 19389 1658 19445 1660
rect 19149 1606 19195 1658
rect 19195 1606 19205 1658
rect 19229 1606 19259 1658
rect 19259 1606 19271 1658
rect 19271 1606 19285 1658
rect 19309 1606 19323 1658
rect 19323 1606 19335 1658
rect 19335 1606 19365 1658
rect 19389 1606 19399 1658
rect 19399 1606 19445 1658
rect 19149 1604 19205 1606
rect 19229 1604 19285 1606
rect 19309 1604 19365 1606
rect 19389 1604 19445 1606
rect 20166 5752 20222 5808
rect 20074 4256 20130 4312
rect 20074 3984 20130 4040
rect 20166 3848 20222 3904
rect 21086 11464 21142 11520
rect 20994 11192 21050 11248
rect 21454 19116 21456 19136
rect 21456 19116 21508 19136
rect 21508 19116 21510 19136
rect 21454 19080 21510 19116
rect 21454 18028 21456 18048
rect 21456 18028 21508 18048
rect 21508 18028 21510 18048
rect 21454 17992 21510 18028
rect 21454 16940 21456 16960
rect 21456 16940 21508 16960
rect 21508 16940 21510 16960
rect 21454 16904 21510 16940
rect 21454 16496 21510 16552
rect 21454 15852 21456 15872
rect 21456 15852 21508 15872
rect 21508 15852 21510 15872
rect 21454 15816 21510 15852
rect 21546 14864 21602 14920
rect 21454 14764 21456 14784
rect 21456 14764 21508 14784
rect 21508 14764 21510 14784
rect 21454 14728 21510 14764
rect 21454 13676 21456 13696
rect 21456 13676 21508 13696
rect 21508 13676 21510 13696
rect 21454 13640 21510 13676
rect 21748 21786 21804 21788
rect 21828 21786 21884 21788
rect 21908 21786 21964 21788
rect 21988 21786 22044 21788
rect 21748 21734 21794 21786
rect 21794 21734 21804 21786
rect 21828 21734 21858 21786
rect 21858 21734 21870 21786
rect 21870 21734 21884 21786
rect 21908 21734 21922 21786
rect 21922 21734 21934 21786
rect 21934 21734 21964 21786
rect 21988 21734 21998 21786
rect 21998 21734 22044 21786
rect 21748 21732 21804 21734
rect 21828 21732 21884 21734
rect 21908 21732 21964 21734
rect 21988 21732 22044 21734
rect 22190 21836 22192 21856
rect 22192 21836 22244 21856
rect 22244 21836 22246 21856
rect 22190 21800 22246 21836
rect 22098 20848 22154 20904
rect 22190 20712 22246 20768
rect 21748 20698 21804 20700
rect 21828 20698 21884 20700
rect 21908 20698 21964 20700
rect 21988 20698 22044 20700
rect 21748 20646 21794 20698
rect 21794 20646 21804 20698
rect 21828 20646 21858 20698
rect 21858 20646 21870 20698
rect 21870 20646 21884 20698
rect 21908 20646 21922 20698
rect 21922 20646 21934 20698
rect 21934 20646 21964 20698
rect 21988 20646 21998 20698
rect 21998 20646 22044 20698
rect 21748 20644 21804 20646
rect 21828 20644 21884 20646
rect 21908 20644 21964 20646
rect 21988 20644 22044 20646
rect 22098 19760 22154 19816
rect 21748 19610 21804 19612
rect 21828 19610 21884 19612
rect 21908 19610 21964 19612
rect 21988 19610 22044 19612
rect 21748 19558 21794 19610
rect 21794 19558 21804 19610
rect 21828 19558 21858 19610
rect 21858 19558 21870 19610
rect 21870 19558 21884 19610
rect 21908 19558 21922 19610
rect 21922 19558 21934 19610
rect 21934 19558 21964 19610
rect 21988 19558 21998 19610
rect 21998 19558 22044 19610
rect 21748 19556 21804 19558
rect 21828 19556 21884 19558
rect 21908 19556 21964 19558
rect 21988 19556 22044 19558
rect 21748 18522 21804 18524
rect 21828 18522 21884 18524
rect 21908 18522 21964 18524
rect 21988 18522 22044 18524
rect 21748 18470 21794 18522
rect 21794 18470 21804 18522
rect 21828 18470 21858 18522
rect 21858 18470 21870 18522
rect 21870 18470 21884 18522
rect 21908 18470 21922 18522
rect 21922 18470 21934 18522
rect 21934 18470 21964 18522
rect 21988 18470 21998 18522
rect 21998 18470 22044 18522
rect 21748 18468 21804 18470
rect 21828 18468 21884 18470
rect 21908 18468 21964 18470
rect 21988 18468 22044 18470
rect 21748 17434 21804 17436
rect 21828 17434 21884 17436
rect 21908 17434 21964 17436
rect 21988 17434 22044 17436
rect 21748 17382 21794 17434
rect 21794 17382 21804 17434
rect 21828 17382 21858 17434
rect 21858 17382 21870 17434
rect 21870 17382 21884 17434
rect 21908 17382 21922 17434
rect 21922 17382 21934 17434
rect 21934 17382 21964 17434
rect 21988 17382 21998 17434
rect 21998 17382 22044 17434
rect 21748 17380 21804 17382
rect 21828 17380 21884 17382
rect 21908 17380 21964 17382
rect 21988 17380 22044 17382
rect 22190 19660 22192 19680
rect 22192 19660 22244 19680
rect 22244 19660 22246 19680
rect 22190 19624 22246 19660
rect 22190 18572 22192 18592
rect 22192 18572 22244 18592
rect 22244 18572 22246 18592
rect 22190 18536 22246 18572
rect 22190 17484 22192 17504
rect 22192 17484 22244 17504
rect 22244 17484 22246 17504
rect 22190 17448 22246 17484
rect 21748 16346 21804 16348
rect 21828 16346 21884 16348
rect 21908 16346 21964 16348
rect 21988 16346 22044 16348
rect 21748 16294 21794 16346
rect 21794 16294 21804 16346
rect 21828 16294 21858 16346
rect 21858 16294 21870 16346
rect 21870 16294 21884 16346
rect 21908 16294 21922 16346
rect 21922 16294 21934 16346
rect 21934 16294 21964 16346
rect 21988 16294 21998 16346
rect 21998 16294 22044 16346
rect 21748 16292 21804 16294
rect 21828 16292 21884 16294
rect 21908 16292 21964 16294
rect 21988 16292 22044 16294
rect 21748 15258 21804 15260
rect 21828 15258 21884 15260
rect 21908 15258 21964 15260
rect 21988 15258 22044 15260
rect 21748 15206 21794 15258
rect 21794 15206 21804 15258
rect 21828 15206 21858 15258
rect 21858 15206 21870 15258
rect 21870 15206 21884 15258
rect 21908 15206 21922 15258
rect 21922 15206 21934 15258
rect 21934 15206 21964 15258
rect 21988 15206 21998 15258
rect 21998 15206 22044 15258
rect 21748 15204 21804 15206
rect 21828 15204 21884 15206
rect 21908 15204 21964 15206
rect 21988 15204 22044 15206
rect 22190 14220 22192 14240
rect 22192 14220 22244 14240
rect 22244 14220 22246 14240
rect 22190 14184 22246 14220
rect 21748 14170 21804 14172
rect 21828 14170 21884 14172
rect 21908 14170 21964 14172
rect 21988 14170 22044 14172
rect 21748 14118 21794 14170
rect 21794 14118 21804 14170
rect 21828 14118 21858 14170
rect 21858 14118 21870 14170
rect 21870 14118 21884 14170
rect 21908 14118 21922 14170
rect 21922 14118 21934 14170
rect 21934 14118 21964 14170
rect 21988 14118 21998 14170
rect 21998 14118 22044 14170
rect 21748 14116 21804 14118
rect 21828 14116 21884 14118
rect 21908 14116 21964 14118
rect 21988 14116 22044 14118
rect 21362 11328 21418 11384
rect 22190 13096 22246 13152
rect 21748 13082 21804 13084
rect 21828 13082 21884 13084
rect 21908 13082 21964 13084
rect 21988 13082 22044 13084
rect 21748 13030 21794 13082
rect 21794 13030 21804 13082
rect 21828 13030 21858 13082
rect 21858 13030 21870 13082
rect 21870 13030 21884 13082
rect 21908 13030 21922 13082
rect 21922 13030 21934 13082
rect 21934 13030 21964 13082
rect 21988 13030 21998 13082
rect 21998 13030 22044 13082
rect 21748 13028 21804 13030
rect 21828 13028 21884 13030
rect 21908 13028 21964 13030
rect 21988 13028 22044 13030
rect 22190 12008 22246 12064
rect 21748 11994 21804 11996
rect 21828 11994 21884 11996
rect 21908 11994 21964 11996
rect 21988 11994 22044 11996
rect 21748 11942 21794 11994
rect 21794 11942 21804 11994
rect 21828 11942 21858 11994
rect 21858 11942 21870 11994
rect 21870 11942 21884 11994
rect 21908 11942 21922 11994
rect 21922 11942 21934 11994
rect 21934 11942 21964 11994
rect 21988 11942 21998 11994
rect 21998 11942 22044 11994
rect 21748 11940 21804 11942
rect 21828 11940 21884 11942
rect 21908 11940 21964 11942
rect 21988 11940 22044 11942
rect 21270 10648 21326 10704
rect 20902 10376 20958 10432
rect 22190 10920 22246 10976
rect 21748 10906 21804 10908
rect 21828 10906 21884 10908
rect 21908 10906 21964 10908
rect 21988 10906 22044 10908
rect 21748 10854 21794 10906
rect 21794 10854 21804 10906
rect 21828 10854 21858 10906
rect 21858 10854 21870 10906
rect 21870 10854 21884 10906
rect 21908 10854 21922 10906
rect 21922 10854 21934 10906
rect 21934 10854 21964 10906
rect 21988 10854 21998 10906
rect 21998 10854 22044 10906
rect 21748 10852 21804 10854
rect 21828 10852 21884 10854
rect 21908 10852 21964 10854
rect 21988 10852 22044 10854
rect 21638 10648 21694 10704
rect 21454 9288 21510 9344
rect 21178 6704 21234 6760
rect 20994 5772 21050 5808
rect 20994 5752 20996 5772
rect 20996 5752 21048 5772
rect 21048 5752 21050 5772
rect 21546 7384 21602 7440
rect 21086 4664 21142 4720
rect 20718 3576 20774 3632
rect 20810 3440 20866 3496
rect 20994 3032 21050 3088
rect 21086 2760 21142 2816
rect 21362 4120 21418 4176
rect 20718 2216 20774 2272
rect 20994 2216 21050 2272
rect 21362 2216 21418 2272
rect 22374 22752 22430 22808
rect 21748 9818 21804 9820
rect 21828 9818 21884 9820
rect 21908 9818 21964 9820
rect 21988 9818 22044 9820
rect 21748 9766 21794 9818
rect 21794 9766 21804 9818
rect 21828 9766 21858 9818
rect 21858 9766 21870 9818
rect 21870 9766 21884 9818
rect 21908 9766 21922 9818
rect 21922 9766 21934 9818
rect 21934 9766 21964 9818
rect 21988 9766 21998 9818
rect 21998 9766 22044 9818
rect 21748 9764 21804 9766
rect 21828 9764 21884 9766
rect 21908 9764 21964 9766
rect 21988 9764 22044 9766
rect 21748 8730 21804 8732
rect 21828 8730 21884 8732
rect 21908 8730 21964 8732
rect 21988 8730 22044 8732
rect 21748 8678 21794 8730
rect 21794 8678 21804 8730
rect 21828 8678 21858 8730
rect 21858 8678 21870 8730
rect 21870 8678 21884 8730
rect 21908 8678 21922 8730
rect 21922 8678 21934 8730
rect 21934 8678 21964 8730
rect 21988 8678 21998 8730
rect 21998 8678 22044 8730
rect 21748 8676 21804 8678
rect 21828 8676 21884 8678
rect 21908 8676 21964 8678
rect 21988 8676 22044 8678
rect 21748 7642 21804 7644
rect 21828 7642 21884 7644
rect 21908 7642 21964 7644
rect 21988 7642 22044 7644
rect 21748 7590 21794 7642
rect 21794 7590 21804 7642
rect 21828 7590 21858 7642
rect 21858 7590 21870 7642
rect 21870 7590 21884 7642
rect 21908 7590 21922 7642
rect 21922 7590 21934 7642
rect 21934 7590 21964 7642
rect 21988 7590 21998 7642
rect 21998 7590 22044 7642
rect 21748 7588 21804 7590
rect 21828 7588 21884 7590
rect 21908 7588 21964 7590
rect 21988 7588 22044 7590
rect 21748 6554 21804 6556
rect 21828 6554 21884 6556
rect 21908 6554 21964 6556
rect 21988 6554 22044 6556
rect 21748 6502 21794 6554
rect 21794 6502 21804 6554
rect 21828 6502 21858 6554
rect 21858 6502 21870 6554
rect 21870 6502 21884 6554
rect 21908 6502 21922 6554
rect 21922 6502 21934 6554
rect 21934 6502 21964 6554
rect 21988 6502 21998 6554
rect 21998 6502 22044 6554
rect 21748 6500 21804 6502
rect 21828 6500 21884 6502
rect 21908 6500 21964 6502
rect 21988 6500 22044 6502
rect 21748 5466 21804 5468
rect 21828 5466 21884 5468
rect 21908 5466 21964 5468
rect 21988 5466 22044 5468
rect 21748 5414 21794 5466
rect 21794 5414 21804 5466
rect 21828 5414 21858 5466
rect 21858 5414 21870 5466
rect 21870 5414 21884 5466
rect 21908 5414 21922 5466
rect 21922 5414 21934 5466
rect 21934 5414 21964 5466
rect 21988 5414 21998 5466
rect 21998 5414 22044 5466
rect 21748 5412 21804 5414
rect 21828 5412 21884 5414
rect 21908 5412 21964 5414
rect 21988 5412 22044 5414
rect 21748 4378 21804 4380
rect 21828 4378 21884 4380
rect 21908 4378 21964 4380
rect 21988 4378 22044 4380
rect 21748 4326 21794 4378
rect 21794 4326 21804 4378
rect 21828 4326 21858 4378
rect 21858 4326 21870 4378
rect 21870 4326 21884 4378
rect 21908 4326 21922 4378
rect 21922 4326 21934 4378
rect 21934 4326 21964 4378
rect 21988 4326 21998 4378
rect 21998 4326 22044 4378
rect 21748 4324 21804 4326
rect 21828 4324 21884 4326
rect 21908 4324 21964 4326
rect 21988 4324 22044 4326
rect 21748 3290 21804 3292
rect 21828 3290 21884 3292
rect 21908 3290 21964 3292
rect 21988 3290 22044 3292
rect 21748 3238 21794 3290
rect 21794 3238 21804 3290
rect 21828 3238 21858 3290
rect 21858 3238 21870 3290
rect 21870 3238 21884 3290
rect 21908 3238 21922 3290
rect 21922 3238 21934 3290
rect 21934 3238 21964 3290
rect 21988 3238 21998 3290
rect 21998 3238 22044 3290
rect 21748 3236 21804 3238
rect 21828 3236 21884 3238
rect 21908 3236 21964 3238
rect 21988 3236 22044 3238
rect 21748 2202 21804 2204
rect 21828 2202 21884 2204
rect 21908 2202 21964 2204
rect 21988 2202 22044 2204
rect 21748 2150 21794 2202
rect 21794 2150 21804 2202
rect 21828 2150 21858 2202
rect 21858 2150 21870 2202
rect 21870 2150 21884 2202
rect 21908 2150 21922 2202
rect 21922 2150 21934 2202
rect 21934 2150 21964 2202
rect 21988 2150 21998 2202
rect 21998 2150 22044 2202
rect 21748 2148 21804 2150
rect 21828 2148 21884 2150
rect 21908 2148 21964 2150
rect 21988 2148 22044 2150
rect 21546 2080 21602 2136
rect 22282 9832 22338 9888
rect 22374 5616 22430 5672
rect 22742 34040 22798 34096
rect 22650 21936 22706 21992
rect 22650 20848 22706 20904
rect 22558 15272 22614 15328
rect 22834 11736 22890 11792
rect 21748 1114 21804 1116
rect 21828 1114 21884 1116
rect 21908 1114 21964 1116
rect 21988 1114 22044 1116
rect 21748 1062 21794 1114
rect 21794 1062 21804 1114
rect 21828 1062 21858 1114
rect 21858 1062 21870 1114
rect 21870 1062 21884 1114
rect 21908 1062 21922 1114
rect 21922 1062 21934 1114
rect 21934 1062 21964 1114
rect 21988 1062 21998 1114
rect 21998 1062 22044 1114
rect 21748 1060 21804 1062
rect 21828 1060 21884 1062
rect 21908 1060 21964 1062
rect 21988 1060 22044 1062
<< metal3 >>
rect 2221 43890 2287 43893
rect 3877 43890 3943 43893
rect 2221 43888 3943 43890
rect 2221 43832 2226 43888
rect 2282 43832 3882 43888
rect 3938 43832 3943 43888
rect 2221 43830 3943 43832
rect 2221 43827 2287 43830
rect 3877 43827 3943 43830
rect 13997 43890 14063 43893
rect 15653 43890 15719 43893
rect 13997 43888 15719 43890
rect 13997 43832 14002 43888
rect 14058 43832 15658 43888
rect 15714 43832 15719 43888
rect 13997 43830 15719 43832
rect 13997 43827 14063 43830
rect 15653 43827 15719 43830
rect 22369 43618 22435 43621
rect 22840 43618 23300 43648
rect 22369 43616 23300 43618
rect 22369 43560 22374 43616
rect 22430 43560 23300 43616
rect 22369 43558 23300 43560
rect 22369 43555 22435 43558
rect 6144 43552 6460 43553
rect 6144 43488 6150 43552
rect 6214 43488 6230 43552
rect 6294 43488 6310 43552
rect 6374 43488 6390 43552
rect 6454 43488 6460 43552
rect 6144 43487 6460 43488
rect 11342 43552 11658 43553
rect 11342 43488 11348 43552
rect 11412 43488 11428 43552
rect 11492 43488 11508 43552
rect 11572 43488 11588 43552
rect 11652 43488 11658 43552
rect 11342 43487 11658 43488
rect 16540 43552 16856 43553
rect 16540 43488 16546 43552
rect 16610 43488 16626 43552
rect 16690 43488 16706 43552
rect 16770 43488 16786 43552
rect 16850 43488 16856 43552
rect 16540 43487 16856 43488
rect 21738 43552 22054 43553
rect 21738 43488 21744 43552
rect 21808 43488 21824 43552
rect 21888 43488 21904 43552
rect 21968 43488 21984 43552
rect 22048 43488 22054 43552
rect 22840 43528 23300 43558
rect 21738 43487 22054 43488
rect 13905 43346 13971 43349
rect 12390 43344 13971 43346
rect 12390 43288 13910 43344
rect 13966 43288 13971 43344
rect 12390 43286 13971 43288
rect 8937 43210 9003 43213
rect 11830 43210 11836 43212
rect 8937 43208 11836 43210
rect 8937 43152 8942 43208
rect 8998 43152 11836 43208
rect 8937 43150 11836 43152
rect 8937 43147 9003 43150
rect 11830 43148 11836 43150
rect 11900 43148 11906 43212
rect 12065 43210 12131 43213
rect 12390 43210 12450 43286
rect 13905 43283 13971 43286
rect 12065 43208 12450 43210
rect 12065 43152 12070 43208
rect 12126 43152 12450 43208
rect 12065 43150 12450 43152
rect 13445 43210 13511 43213
rect 18321 43210 18387 43213
rect 13445 43208 18387 43210
rect 13445 43152 13450 43208
rect 13506 43152 18326 43208
rect 18382 43152 18387 43208
rect 13445 43150 18387 43152
rect 12065 43147 12131 43150
rect 13445 43147 13511 43150
rect 18321 43147 18387 43150
rect 11145 43074 11211 43077
rect 10918 43072 11211 43074
rect 10918 43016 11150 43072
rect 11206 43016 11211 43072
rect 10918 43014 11211 43016
rect 3545 43008 3861 43009
rect 3545 42944 3551 43008
rect 3615 42944 3631 43008
rect 3695 42944 3711 43008
rect 3775 42944 3791 43008
rect 3855 42944 3861 43008
rect 3545 42943 3861 42944
rect 8743 43008 9059 43009
rect 8743 42944 8749 43008
rect 8813 42944 8829 43008
rect 8893 42944 8909 43008
rect 8973 42944 8989 43008
rect 9053 42944 9059 43008
rect 8743 42943 9059 42944
rect 4337 42938 4403 42941
rect 5022 42938 5028 42940
rect 4337 42936 5028 42938
rect 4337 42880 4342 42936
rect 4398 42880 5028 42936
rect 4337 42878 5028 42880
rect 4337 42875 4403 42878
rect 5022 42876 5028 42878
rect 5092 42876 5098 42940
rect 8569 42666 8635 42669
rect 9397 42666 9463 42669
rect 8569 42664 9463 42666
rect 8569 42608 8574 42664
rect 8630 42608 9402 42664
rect 9458 42608 9463 42664
rect 8569 42606 9463 42608
rect 8569 42603 8635 42606
rect 9397 42603 9463 42606
rect 10918 42533 10978 43014
rect 11145 43011 11211 43014
rect 20529 43074 20595 43077
rect 22840 43074 23300 43104
rect 20529 43072 23300 43074
rect 20529 43016 20534 43072
rect 20590 43016 23300 43072
rect 20529 43014 23300 43016
rect 20529 43011 20595 43014
rect 13941 43008 14257 43009
rect 13941 42944 13947 43008
rect 14011 42944 14027 43008
rect 14091 42944 14107 43008
rect 14171 42944 14187 43008
rect 14251 42944 14257 43008
rect 13941 42943 14257 42944
rect 19139 43008 19455 43009
rect 19139 42944 19145 43008
rect 19209 42944 19225 43008
rect 19289 42944 19305 43008
rect 19369 42944 19385 43008
rect 19449 42944 19455 43008
rect 22840 42984 23300 43014
rect 19139 42943 19455 42944
rect 13077 42940 13143 42941
rect 13077 42936 13124 42940
rect 13188 42938 13194 42940
rect 15009 42938 15075 42941
rect 13077 42880 13082 42936
rect 13077 42876 13124 42880
rect 13188 42878 13234 42938
rect 14782 42936 15075 42938
rect 14782 42880 15014 42936
rect 15070 42880 15075 42936
rect 14782 42878 15075 42880
rect 13188 42876 13194 42878
rect 13077 42875 13143 42876
rect 6678 42468 6684 42532
rect 6748 42530 6754 42532
rect 10501 42530 10567 42533
rect 6748 42528 10567 42530
rect 6748 42472 10506 42528
rect 10562 42472 10567 42528
rect 6748 42470 10567 42472
rect 6748 42468 6754 42470
rect 10501 42467 10567 42470
rect 10869 42528 10978 42533
rect 10869 42472 10874 42528
rect 10930 42472 10978 42528
rect 10869 42470 10978 42472
rect 10869 42467 10935 42470
rect 6144 42464 6460 42465
rect 6144 42400 6150 42464
rect 6214 42400 6230 42464
rect 6294 42400 6310 42464
rect 6374 42400 6390 42464
rect 6454 42400 6460 42464
rect 6144 42399 6460 42400
rect 11342 42464 11658 42465
rect 11342 42400 11348 42464
rect 11412 42400 11428 42464
rect 11492 42400 11508 42464
rect 11572 42400 11588 42464
rect 11652 42400 11658 42464
rect 11342 42399 11658 42400
rect 9121 42394 9187 42397
rect 9254 42394 9260 42396
rect 9121 42392 9260 42394
rect 9121 42336 9126 42392
rect 9182 42336 9260 42392
rect 9121 42334 9260 42336
rect 9121 42331 9187 42334
rect 9254 42332 9260 42334
rect 9324 42332 9330 42396
rect 9438 42332 9444 42396
rect 9508 42394 9514 42396
rect 10685 42394 10751 42397
rect 9508 42392 10751 42394
rect 9508 42336 10690 42392
rect 10746 42336 10751 42392
rect 9508 42334 10751 42336
rect 9508 42332 9514 42334
rect 10685 42331 10751 42334
rect 14782 42261 14842 42878
rect 15009 42875 15075 42878
rect 17902 42876 17908 42940
rect 17972 42938 17978 42940
rect 18597 42938 18663 42941
rect 17972 42936 18663 42938
rect 17972 42880 18602 42936
rect 18658 42880 18663 42936
rect 17972 42878 18663 42880
rect 17972 42876 17978 42878
rect 18597 42875 18663 42878
rect 17493 42530 17559 42533
rect 18965 42530 19031 42533
rect 17493 42528 19031 42530
rect 17493 42472 17498 42528
rect 17554 42472 18970 42528
rect 19026 42472 19031 42528
rect 17493 42470 19031 42472
rect 17493 42467 17559 42470
rect 18965 42467 19031 42470
rect 22185 42530 22251 42533
rect 22840 42530 23300 42560
rect 22185 42528 23300 42530
rect 22185 42472 22190 42528
rect 22246 42472 23300 42528
rect 22185 42470 23300 42472
rect 22185 42467 22251 42470
rect 16540 42464 16856 42465
rect 16540 42400 16546 42464
rect 16610 42400 16626 42464
rect 16690 42400 16706 42464
rect 16770 42400 16786 42464
rect 16850 42400 16856 42464
rect 16540 42399 16856 42400
rect 21738 42464 22054 42465
rect 21738 42400 21744 42464
rect 21808 42400 21824 42464
rect 21888 42400 21904 42464
rect 21968 42400 21984 42464
rect 22048 42400 22054 42464
rect 22840 42440 23300 42470
rect 21738 42399 22054 42400
rect 19742 42332 19748 42396
rect 19812 42394 19818 42396
rect 20437 42394 20503 42397
rect 19812 42392 20503 42394
rect 19812 42336 20442 42392
rect 20498 42336 20503 42392
rect 19812 42334 20503 42336
rect 19812 42332 19818 42334
rect 20437 42331 20503 42334
rect 933 42258 999 42261
rect 6453 42258 6519 42261
rect 933 42256 6519 42258
rect 933 42200 938 42256
rect 994 42200 6458 42256
rect 6514 42200 6519 42256
rect 933 42198 6519 42200
rect 933 42195 999 42198
rect 6453 42195 6519 42198
rect 8334 42196 8340 42260
rect 8404 42258 8410 42260
rect 11145 42258 11211 42261
rect 8404 42256 11211 42258
rect 8404 42200 11150 42256
rect 11206 42200 11211 42256
rect 8404 42198 11211 42200
rect 8404 42196 8410 42198
rect 11145 42195 11211 42198
rect 14733 42256 14842 42261
rect 20478 42258 20484 42260
rect 14733 42200 14738 42256
rect 14794 42200 14842 42256
rect 14733 42198 14842 42200
rect 14966 42198 20484 42258
rect 14733 42195 14799 42198
rect 841 42122 907 42125
rect 5349 42122 5415 42125
rect 841 42120 5415 42122
rect 841 42064 846 42120
rect 902 42064 5354 42120
rect 5410 42064 5415 42120
rect 841 42062 5415 42064
rect 841 42059 907 42062
rect 5349 42059 5415 42062
rect 8937 42122 9003 42125
rect 9397 42122 9463 42125
rect 8937 42120 9463 42122
rect 8937 42064 8942 42120
rect 8998 42064 9402 42120
rect 9458 42064 9463 42120
rect 8937 42062 9463 42064
rect 8937 42059 9003 42062
rect 9397 42059 9463 42062
rect 12433 42122 12499 42125
rect 13997 42122 14063 42125
rect 12433 42120 14063 42122
rect 12433 42064 12438 42120
rect 12494 42064 14002 42120
rect 14058 42064 14063 42120
rect 12433 42062 14063 42064
rect 12433 42059 12499 42062
rect 13997 42059 14063 42062
rect 10041 41986 10107 41989
rect 10174 41986 10180 41988
rect 10041 41984 10180 41986
rect 10041 41928 10046 41984
rect 10102 41928 10180 41984
rect 10041 41926 10180 41928
rect 10041 41923 10107 41926
rect 10174 41924 10180 41926
rect 10244 41924 10250 41988
rect 3545 41920 3861 41921
rect 3545 41856 3551 41920
rect 3615 41856 3631 41920
rect 3695 41856 3711 41920
rect 3775 41856 3791 41920
rect 3855 41856 3861 41920
rect 3545 41855 3861 41856
rect 8743 41920 9059 41921
rect 8743 41856 8749 41920
rect 8813 41856 8829 41920
rect 8893 41856 8909 41920
rect 8973 41856 8989 41920
rect 9053 41856 9059 41920
rect 8743 41855 9059 41856
rect 13941 41920 14257 41921
rect 13941 41856 13947 41920
rect 14011 41856 14027 41920
rect 14091 41856 14107 41920
rect 14171 41856 14187 41920
rect 14251 41856 14257 41920
rect 13941 41855 14257 41856
rect 9581 41848 9647 41853
rect 9581 41792 9586 41848
rect 9642 41792 9647 41848
rect 9581 41787 9647 41792
rect 790 41652 796 41716
rect 860 41714 866 41716
rect 4245 41714 4311 41717
rect 860 41712 4311 41714
rect 860 41656 4250 41712
rect 4306 41656 4311 41712
rect 860 41654 4311 41656
rect 860 41652 866 41654
rect 4245 41651 4311 41654
rect 8385 41714 8451 41717
rect 9584 41714 9644 41787
rect 8385 41712 9644 41714
rect 8385 41656 8390 41712
rect 8446 41656 9644 41712
rect 8385 41654 9644 41656
rect 14181 41714 14247 41717
rect 14966 41714 15026 42198
rect 20478 42196 20484 42198
rect 20548 42196 20554 42260
rect 17718 42060 17724 42124
rect 17788 42122 17794 42124
rect 19517 42122 19583 42125
rect 17788 42120 19583 42122
rect 17788 42064 19522 42120
rect 19578 42064 19583 42120
rect 17788 42062 19583 42064
rect 17788 42060 17794 42062
rect 19517 42059 19583 42062
rect 21909 41986 21975 41989
rect 22840 41986 23300 42016
rect 21909 41984 23300 41986
rect 21909 41928 21914 41984
rect 21970 41928 23300 41984
rect 21909 41926 23300 41928
rect 21909 41923 21975 41926
rect 19139 41920 19455 41921
rect 19139 41856 19145 41920
rect 19209 41856 19225 41920
rect 19289 41856 19305 41920
rect 19369 41856 19385 41920
rect 19449 41856 19455 41920
rect 22840 41896 23300 41926
rect 19139 41855 19455 41856
rect 16297 41850 16363 41853
rect 17861 41850 17927 41853
rect 16297 41848 17927 41850
rect 16297 41792 16302 41848
rect 16358 41792 17866 41848
rect 17922 41792 17927 41848
rect 16297 41790 17927 41792
rect 16297 41787 16363 41790
rect 17861 41787 17927 41790
rect 18086 41788 18092 41852
rect 18156 41850 18162 41852
rect 18965 41850 19031 41853
rect 18156 41848 19031 41850
rect 18156 41792 18970 41848
rect 19026 41792 19031 41848
rect 18156 41790 19031 41792
rect 18156 41788 18162 41790
rect 18965 41787 19031 41790
rect 15193 41716 15259 41717
rect 15142 41714 15148 41716
rect 14181 41712 15026 41714
rect 14181 41656 14186 41712
rect 14242 41656 15026 41712
rect 14181 41654 15026 41656
rect 15102 41654 15148 41714
rect 15212 41712 15259 41716
rect 15254 41656 15259 41712
rect 8385 41651 8451 41654
rect 14181 41651 14247 41654
rect 15142 41652 15148 41654
rect 15212 41652 15259 41656
rect 15193 41651 15259 41652
rect 15929 41714 15995 41717
rect 16062 41714 16068 41716
rect 15929 41712 16068 41714
rect 15929 41656 15934 41712
rect 15990 41656 16068 41712
rect 15929 41654 16068 41656
rect 15929 41651 15995 41654
rect 16062 41652 16068 41654
rect 16132 41652 16138 41716
rect 16849 41714 16915 41717
rect 20621 41714 20687 41717
rect 16849 41712 20687 41714
rect 16849 41656 16854 41712
rect 16910 41656 20626 41712
rect 20682 41656 20687 41712
rect 16849 41654 20687 41656
rect 16849 41651 16915 41654
rect 20621 41651 20687 41654
rect 2221 41578 2287 41581
rect 4521 41578 4587 41581
rect 7373 41580 7439 41581
rect 4654 41578 4660 41580
rect 2221 41576 4354 41578
rect 2221 41520 2226 41576
rect 2282 41520 4354 41576
rect 2221 41518 4354 41520
rect 2221 41515 2287 41518
rect 13 41442 79 41445
rect 3601 41442 3667 41445
rect 13 41440 3667 41442
rect 13 41384 18 41440
rect 74 41384 3606 41440
rect 3662 41384 3667 41440
rect 13 41382 3667 41384
rect 4294 41442 4354 41518
rect 4521 41576 4660 41578
rect 4521 41520 4526 41576
rect 4582 41520 4660 41576
rect 4521 41518 4660 41520
rect 4521 41515 4587 41518
rect 4654 41516 4660 41518
rect 4724 41516 4730 41580
rect 4846 41518 6746 41578
rect 4846 41442 4906 41518
rect 4294 41382 4906 41442
rect 6686 41442 6746 41518
rect 7373 41576 7420 41580
rect 7484 41578 7490 41580
rect 12249 41578 12315 41581
rect 15377 41578 15443 41581
rect 7373 41520 7378 41576
rect 7373 41516 7420 41520
rect 7484 41518 7530 41578
rect 12249 41576 15443 41578
rect 12249 41520 12254 41576
rect 12310 41520 15382 41576
rect 15438 41520 15443 41576
rect 12249 41518 15443 41520
rect 7484 41516 7490 41518
rect 7373 41515 7439 41516
rect 12249 41515 12315 41518
rect 15377 41515 15443 41518
rect 16021 41578 16087 41581
rect 16665 41578 16731 41581
rect 16021 41576 16731 41578
rect 16021 41520 16026 41576
rect 16082 41520 16670 41576
rect 16726 41520 16731 41576
rect 16021 41518 16731 41520
rect 16021 41515 16087 41518
rect 16665 41515 16731 41518
rect 16849 41578 16915 41581
rect 16849 41576 17234 41578
rect 16849 41520 16854 41576
rect 16910 41520 17234 41576
rect 16849 41518 17234 41520
rect 16849 41515 16915 41518
rect 7557 41442 7623 41445
rect 6686 41440 7623 41442
rect 6686 41384 7562 41440
rect 7618 41384 7623 41440
rect 6686 41382 7623 41384
rect 13 41379 79 41382
rect 3601 41379 3667 41382
rect 7557 41379 7623 41382
rect 9765 41442 9831 41445
rect 10225 41442 10291 41445
rect 9765 41440 10291 41442
rect 9765 41384 9770 41440
rect 9826 41384 10230 41440
rect 10286 41384 10291 41440
rect 9765 41382 10291 41384
rect 9765 41379 9831 41382
rect 10225 41379 10291 41382
rect 15326 41380 15332 41444
rect 15396 41442 15402 41444
rect 15469 41442 15535 41445
rect 15396 41440 15535 41442
rect 15396 41384 15474 41440
rect 15530 41384 15535 41440
rect 15396 41382 15535 41384
rect 17174 41442 17234 41518
rect 17350 41516 17356 41580
rect 17420 41578 17426 41580
rect 17769 41578 17835 41581
rect 17420 41576 17835 41578
rect 17420 41520 17774 41576
rect 17830 41520 17835 41576
rect 17420 41518 17835 41520
rect 17420 41516 17426 41518
rect 17769 41515 17835 41518
rect 22277 41442 22343 41445
rect 22840 41442 23300 41472
rect 17174 41382 19442 41442
rect 15396 41380 15402 41382
rect 15469 41379 15535 41382
rect 6144 41376 6460 41377
rect 6144 41312 6150 41376
rect 6214 41312 6230 41376
rect 6294 41312 6310 41376
rect 6374 41312 6390 41376
rect 6454 41312 6460 41376
rect 6144 41311 6460 41312
rect 11342 41376 11658 41377
rect 11342 41312 11348 41376
rect 11412 41312 11428 41376
rect 11492 41312 11508 41376
rect 11572 41312 11588 41376
rect 11652 41312 11658 41376
rect 11342 41311 11658 41312
rect 16540 41376 16856 41377
rect 16540 41312 16546 41376
rect 16610 41312 16626 41376
rect 16690 41312 16706 41376
rect 16770 41312 16786 41376
rect 16850 41312 16856 41376
rect 16540 41311 16856 41312
rect 7281 41306 7347 41309
rect 8385 41306 8451 41309
rect 18321 41308 18387 41309
rect 18270 41306 18276 41308
rect 7281 41304 8451 41306
rect 7281 41248 7286 41304
rect 7342 41248 8390 41304
rect 8446 41248 8451 41304
rect 7281 41246 8451 41248
rect 18230 41246 18276 41306
rect 18340 41304 18387 41308
rect 18382 41248 18387 41304
rect 7281 41243 7347 41246
rect 8385 41243 8451 41246
rect 18270 41244 18276 41246
rect 18340 41244 18387 41248
rect 19382 41306 19442 41382
rect 22277 41440 23300 41442
rect 22277 41384 22282 41440
rect 22338 41384 23300 41440
rect 22277 41382 23300 41384
rect 22277 41379 22343 41382
rect 21738 41376 22054 41377
rect 21738 41312 21744 41376
rect 21808 41312 21824 41376
rect 21888 41312 21904 41376
rect 21968 41312 21984 41376
rect 22048 41312 22054 41376
rect 22840 41352 23300 41382
rect 21738 41311 22054 41312
rect 20437 41306 20503 41309
rect 19382 41304 20503 41306
rect 19382 41248 20442 41304
rect 20498 41248 20503 41304
rect 19382 41246 20503 41248
rect 18321 41243 18387 41244
rect 20437 41243 20503 41246
rect 7281 41170 7347 41173
rect 7649 41170 7715 41173
rect 7281 41168 7715 41170
rect 7281 41112 7286 41168
rect 7342 41112 7654 41168
rect 7710 41112 7715 41168
rect 7281 41110 7715 41112
rect 7281 41107 7347 41110
rect 7649 41107 7715 41110
rect 9949 41170 10015 41173
rect 14641 41170 14707 41173
rect 9949 41168 14707 41170
rect 9949 41112 9954 41168
rect 10010 41112 14646 41168
rect 14702 41112 14707 41168
rect 9949 41110 14707 41112
rect 9949 41107 10015 41110
rect 14641 41107 14707 41110
rect 17033 41170 17099 41173
rect 18229 41170 18295 41173
rect 17033 41168 18295 41170
rect 17033 41112 17038 41168
rect 17094 41112 18234 41168
rect 18290 41112 18295 41168
rect 17033 41110 18295 41112
rect 17033 41107 17099 41110
rect 18229 41107 18295 41110
rect 18873 41170 18939 41173
rect 20897 41170 20963 41173
rect 18873 41168 20963 41170
rect 18873 41112 18878 41168
rect 18934 41112 20902 41168
rect 20958 41112 20963 41168
rect 18873 41110 20963 41112
rect 18873 41107 18939 41110
rect 20897 41107 20963 41110
rect 2129 41034 2195 41037
rect 16573 41034 16639 41037
rect 2129 41032 16639 41034
rect 2129 40976 2134 41032
rect 2190 40976 16578 41032
rect 16634 40976 16639 41032
rect 2129 40974 16639 40976
rect 2129 40971 2195 40974
rect 16573 40971 16639 40974
rect 17953 41034 18019 41037
rect 19241 41034 19307 41037
rect 17953 41032 19307 41034
rect 17953 40976 17958 41032
rect 18014 40976 19246 41032
rect 19302 40976 19307 41032
rect 17953 40974 19307 40976
rect 17953 40971 18019 40974
rect 19241 40971 19307 40974
rect 17493 40898 17559 40901
rect 17718 40898 17724 40900
rect 17493 40896 17724 40898
rect 17493 40840 17498 40896
rect 17554 40840 17724 40896
rect 17493 40838 17724 40840
rect 17493 40835 17559 40838
rect 17718 40836 17724 40838
rect 17788 40836 17794 40900
rect 22185 40898 22251 40901
rect 22840 40898 23300 40928
rect 22185 40896 23300 40898
rect 22185 40840 22190 40896
rect 22246 40840 23300 40896
rect 22185 40838 23300 40840
rect 22185 40835 22251 40838
rect 3545 40832 3861 40833
rect 3545 40768 3551 40832
rect 3615 40768 3631 40832
rect 3695 40768 3711 40832
rect 3775 40768 3791 40832
rect 3855 40768 3861 40832
rect 3545 40767 3861 40768
rect 8743 40832 9059 40833
rect 8743 40768 8749 40832
rect 8813 40768 8829 40832
rect 8893 40768 8909 40832
rect 8973 40768 8989 40832
rect 9053 40768 9059 40832
rect 8743 40767 9059 40768
rect 13941 40832 14257 40833
rect 13941 40768 13947 40832
rect 14011 40768 14027 40832
rect 14091 40768 14107 40832
rect 14171 40768 14187 40832
rect 14251 40768 14257 40832
rect 13941 40767 14257 40768
rect 19139 40832 19455 40833
rect 19139 40768 19145 40832
rect 19209 40768 19225 40832
rect 19289 40768 19305 40832
rect 19369 40768 19385 40832
rect 19449 40768 19455 40832
rect 22840 40808 23300 40838
rect 19139 40767 19455 40768
rect 19793 40762 19859 40765
rect 19926 40762 19932 40764
rect 19793 40760 19932 40762
rect 19793 40704 19798 40760
rect 19854 40704 19932 40760
rect 19793 40702 19932 40704
rect 19793 40699 19859 40702
rect 19926 40700 19932 40702
rect 19996 40700 20002 40764
rect 606 40564 612 40628
rect 676 40626 682 40628
rect 6545 40626 6611 40629
rect 676 40624 6611 40626
rect 676 40568 6550 40624
rect 6606 40568 6611 40624
rect 676 40566 6611 40568
rect 676 40564 682 40566
rect 6545 40563 6611 40566
rect 17769 40626 17835 40629
rect 17902 40626 17908 40628
rect 17769 40624 17908 40626
rect 17769 40568 17774 40624
rect 17830 40568 17908 40624
rect 17769 40566 17908 40568
rect 17769 40563 17835 40566
rect 17902 40564 17908 40566
rect 17972 40564 17978 40628
rect 18597 40626 18663 40629
rect 20253 40626 20319 40629
rect 18597 40624 20319 40626
rect 18597 40568 18602 40624
rect 18658 40568 20258 40624
rect 20314 40568 20319 40624
rect 18597 40566 20319 40568
rect 18597 40563 18663 40566
rect 20253 40563 20319 40566
rect 3969 40490 4035 40493
rect 7005 40490 7071 40493
rect 3969 40488 7071 40490
rect 3969 40432 3974 40488
rect 4030 40432 7010 40488
rect 7066 40432 7071 40488
rect 3969 40430 7071 40432
rect 3969 40427 4035 40430
rect 7005 40427 7071 40430
rect 18413 40490 18479 40493
rect 19742 40490 19748 40492
rect 18413 40488 19748 40490
rect 18413 40432 18418 40488
rect 18474 40432 19748 40488
rect 18413 40430 19748 40432
rect 18413 40427 18479 40430
rect 19742 40428 19748 40430
rect 19812 40428 19818 40492
rect 18045 40354 18111 40357
rect 21541 40354 21607 40357
rect 18045 40352 21607 40354
rect 18045 40296 18050 40352
rect 18106 40296 21546 40352
rect 21602 40296 21607 40352
rect 18045 40294 21607 40296
rect 18045 40291 18111 40294
rect 21541 40291 21607 40294
rect 22185 40354 22251 40357
rect 22840 40354 23300 40384
rect 22185 40352 23300 40354
rect 22185 40296 22190 40352
rect 22246 40296 23300 40352
rect 22185 40294 23300 40296
rect 22185 40291 22251 40294
rect 6144 40288 6460 40289
rect 6144 40224 6150 40288
rect 6214 40224 6230 40288
rect 6294 40224 6310 40288
rect 6374 40224 6390 40288
rect 6454 40224 6460 40288
rect 6144 40223 6460 40224
rect 11342 40288 11658 40289
rect 11342 40224 11348 40288
rect 11412 40224 11428 40288
rect 11492 40224 11508 40288
rect 11572 40224 11588 40288
rect 11652 40224 11658 40288
rect 11342 40223 11658 40224
rect 16540 40288 16856 40289
rect 16540 40224 16546 40288
rect 16610 40224 16626 40288
rect 16690 40224 16706 40288
rect 16770 40224 16786 40288
rect 16850 40224 16856 40288
rect 16540 40223 16856 40224
rect 21738 40288 22054 40289
rect 21738 40224 21744 40288
rect 21808 40224 21824 40288
rect 21888 40224 21904 40288
rect 21968 40224 21984 40288
rect 22048 40224 22054 40288
rect 22840 40264 23300 40294
rect 21738 40223 22054 40224
rect 5257 40218 5323 40221
rect 5390 40218 5396 40220
rect 5257 40216 5396 40218
rect 5257 40160 5262 40216
rect 5318 40160 5396 40216
rect 5257 40158 5396 40160
rect 5257 40155 5323 40158
rect 5390 40156 5396 40158
rect 5460 40156 5466 40220
rect 17217 40218 17283 40221
rect 20897 40218 20963 40221
rect 17217 40216 20963 40218
rect 17217 40160 17222 40216
rect 17278 40160 20902 40216
rect 20958 40160 20963 40216
rect 17217 40158 20963 40160
rect 17217 40155 17283 40158
rect 20897 40155 20963 40158
rect 1669 40082 1735 40085
rect 8017 40082 8083 40085
rect 19057 40084 19123 40085
rect 19006 40082 19012 40084
rect 1669 40080 8083 40082
rect 1669 40024 1674 40080
rect 1730 40024 8022 40080
rect 8078 40024 8083 40080
rect 1669 40022 8083 40024
rect 18966 40022 19012 40082
rect 19076 40080 19123 40084
rect 19118 40024 19123 40080
rect 1669 40019 1735 40022
rect 8017 40019 8083 40022
rect 19006 40020 19012 40022
rect 19076 40020 19123 40024
rect 19558 40020 19564 40084
rect 19628 40082 19634 40084
rect 19885 40082 19951 40085
rect 19628 40080 19951 40082
rect 19628 40024 19890 40080
rect 19946 40024 19951 40080
rect 19628 40022 19951 40024
rect 19628 40020 19634 40022
rect 19057 40019 19123 40020
rect 19885 40019 19951 40022
rect 5022 39884 5028 39948
rect 5092 39946 5098 39948
rect 5993 39946 6059 39949
rect 5092 39944 6059 39946
rect 5092 39888 5998 39944
rect 6054 39888 6059 39944
rect 5092 39886 6059 39888
rect 5092 39884 5098 39886
rect 5993 39883 6059 39886
rect 19517 39946 19583 39949
rect 19926 39946 19932 39948
rect 19517 39944 19932 39946
rect 19517 39888 19522 39944
rect 19578 39888 19932 39944
rect 19517 39886 19932 39888
rect 19517 39883 19583 39886
rect 19926 39884 19932 39886
rect 19996 39884 20002 39948
rect 1393 39810 1459 39813
rect 2405 39810 2471 39813
rect 1393 39808 2471 39810
rect 1393 39752 1398 39808
rect 1454 39752 2410 39808
rect 2466 39752 2471 39808
rect 1393 39750 2471 39752
rect 1393 39747 1459 39750
rect 2405 39747 2471 39750
rect 21449 39810 21515 39813
rect 22840 39810 23300 39840
rect 21449 39808 23300 39810
rect 21449 39752 21454 39808
rect 21510 39752 23300 39808
rect 21449 39750 23300 39752
rect 21449 39747 21515 39750
rect 3545 39744 3861 39745
rect 3545 39680 3551 39744
rect 3615 39680 3631 39744
rect 3695 39680 3711 39744
rect 3775 39680 3791 39744
rect 3855 39680 3861 39744
rect 3545 39679 3861 39680
rect 8743 39744 9059 39745
rect 8743 39680 8749 39744
rect 8813 39680 8829 39744
rect 8893 39680 8909 39744
rect 8973 39680 8989 39744
rect 9053 39680 9059 39744
rect 8743 39679 9059 39680
rect 13941 39744 14257 39745
rect 13941 39680 13947 39744
rect 14011 39680 14027 39744
rect 14091 39680 14107 39744
rect 14171 39680 14187 39744
rect 14251 39680 14257 39744
rect 13941 39679 14257 39680
rect 19139 39744 19455 39745
rect 19139 39680 19145 39744
rect 19209 39680 19225 39744
rect 19289 39680 19305 39744
rect 19369 39680 19385 39744
rect 19449 39680 19455 39744
rect 22840 39720 23300 39750
rect 19139 39679 19455 39680
rect 2497 39674 2563 39677
rect 2497 39672 3434 39674
rect 2497 39616 2502 39672
rect 2558 39616 3434 39672
rect 2497 39614 3434 39616
rect 2497 39611 2563 39614
rect -300 39538 160 39568
rect 2773 39538 2839 39541
rect -300 39536 2839 39538
rect -300 39480 2778 39536
rect 2834 39480 2839 39536
rect -300 39478 2839 39480
rect 3374 39538 3434 39614
rect 14457 39538 14523 39541
rect 17769 39538 17835 39541
rect 3374 39478 12450 39538
rect -300 39448 160 39478
rect 2773 39475 2839 39478
rect 12390 39402 12450 39478
rect 14457 39536 17835 39538
rect 14457 39480 14462 39536
rect 14518 39480 17774 39536
rect 17830 39480 17835 39536
rect 14457 39478 17835 39480
rect 14457 39475 14523 39478
rect 17769 39475 17835 39478
rect 14457 39402 14523 39405
rect 12390 39400 14523 39402
rect 12390 39344 14462 39400
rect 14518 39344 14523 39400
rect 12390 39342 14523 39344
rect 14457 39339 14523 39342
rect 19333 39402 19399 39405
rect 21173 39402 21239 39405
rect 19333 39400 21239 39402
rect 19333 39344 19338 39400
rect 19394 39344 21178 39400
rect 21234 39344 21239 39400
rect 19333 39342 21239 39344
rect 19333 39339 19399 39342
rect 21173 39339 21239 39342
rect -300 39266 160 39296
rect 2957 39266 3023 39269
rect -300 39264 3023 39266
rect -300 39208 2962 39264
rect 3018 39208 3023 39264
rect -300 39206 3023 39208
rect -300 39176 160 39206
rect 2957 39203 3023 39206
rect 19701 39266 19767 39269
rect 20529 39266 20595 39269
rect 19701 39264 20595 39266
rect 19701 39208 19706 39264
rect 19762 39208 20534 39264
rect 20590 39208 20595 39264
rect 19701 39206 20595 39208
rect 19701 39203 19767 39206
rect 20529 39203 20595 39206
rect 22185 39266 22251 39269
rect 22840 39266 23300 39296
rect 22185 39264 23300 39266
rect 22185 39208 22190 39264
rect 22246 39208 23300 39264
rect 22185 39206 23300 39208
rect 22185 39203 22251 39206
rect 6144 39200 6460 39201
rect 6144 39136 6150 39200
rect 6214 39136 6230 39200
rect 6294 39136 6310 39200
rect 6374 39136 6390 39200
rect 6454 39136 6460 39200
rect 6144 39135 6460 39136
rect 11342 39200 11658 39201
rect 11342 39136 11348 39200
rect 11412 39136 11428 39200
rect 11492 39136 11508 39200
rect 11572 39136 11588 39200
rect 11652 39136 11658 39200
rect 11342 39135 11658 39136
rect 16540 39200 16856 39201
rect 16540 39136 16546 39200
rect 16610 39136 16626 39200
rect 16690 39136 16706 39200
rect 16770 39136 16786 39200
rect 16850 39136 16856 39200
rect 16540 39135 16856 39136
rect 21738 39200 22054 39201
rect 21738 39136 21744 39200
rect 21808 39136 21824 39200
rect 21888 39136 21904 39200
rect 21968 39136 21984 39200
rect 22048 39136 22054 39200
rect 22840 39176 23300 39206
rect 21738 39135 22054 39136
rect -300 38994 160 39024
rect 1301 38994 1367 38997
rect -300 38992 1367 38994
rect -300 38936 1306 38992
rect 1362 38936 1367 38992
rect -300 38934 1367 38936
rect -300 38904 160 38934
rect 1301 38931 1367 38934
rect 16481 38994 16547 38997
rect 18086 38994 18092 38996
rect 16481 38992 18092 38994
rect 16481 38936 16486 38992
rect 16542 38936 18092 38992
rect 16481 38934 18092 38936
rect 16481 38931 16547 38934
rect 18086 38932 18092 38934
rect 18156 38932 18162 38996
rect -300 38722 160 38752
rect 1117 38722 1183 38725
rect -300 38720 1183 38722
rect -300 38664 1122 38720
rect 1178 38664 1183 38720
rect -300 38662 1183 38664
rect -300 38632 160 38662
rect 1117 38659 1183 38662
rect 2262 38660 2268 38724
rect 2332 38722 2338 38724
rect 2681 38722 2747 38725
rect 2332 38720 2747 38722
rect 2332 38664 2686 38720
rect 2742 38664 2747 38720
rect 2332 38662 2747 38664
rect 2332 38660 2338 38662
rect 2681 38659 2747 38662
rect 14641 38722 14707 38725
rect 15326 38722 15332 38724
rect 14641 38720 15332 38722
rect 14641 38664 14646 38720
rect 14702 38664 15332 38720
rect 14641 38662 15332 38664
rect 14641 38659 14707 38662
rect 15326 38660 15332 38662
rect 15396 38660 15402 38724
rect 17217 38722 17283 38725
rect 18270 38722 18276 38724
rect 17217 38720 18276 38722
rect 17217 38664 17222 38720
rect 17278 38664 18276 38720
rect 17217 38662 18276 38664
rect 17217 38659 17283 38662
rect 18270 38660 18276 38662
rect 18340 38660 18346 38724
rect 20110 38660 20116 38724
rect 20180 38722 20186 38724
rect 20253 38722 20319 38725
rect 20180 38720 20319 38722
rect 20180 38664 20258 38720
rect 20314 38664 20319 38720
rect 20180 38662 20319 38664
rect 20180 38660 20186 38662
rect 20253 38659 20319 38662
rect 21449 38722 21515 38725
rect 22840 38722 23300 38752
rect 21449 38720 23300 38722
rect 21449 38664 21454 38720
rect 21510 38664 23300 38720
rect 21449 38662 23300 38664
rect 21449 38659 21515 38662
rect 3545 38656 3861 38657
rect 3545 38592 3551 38656
rect 3615 38592 3631 38656
rect 3695 38592 3711 38656
rect 3775 38592 3791 38656
rect 3855 38592 3861 38656
rect 3545 38591 3861 38592
rect 8743 38656 9059 38657
rect 8743 38592 8749 38656
rect 8813 38592 8829 38656
rect 8893 38592 8909 38656
rect 8973 38592 8989 38656
rect 9053 38592 9059 38656
rect 8743 38591 9059 38592
rect 13941 38656 14257 38657
rect 13941 38592 13947 38656
rect 14011 38592 14027 38656
rect 14091 38592 14107 38656
rect 14171 38592 14187 38656
rect 14251 38592 14257 38656
rect 13941 38591 14257 38592
rect 19139 38656 19455 38657
rect 19139 38592 19145 38656
rect 19209 38592 19225 38656
rect 19289 38592 19305 38656
rect 19369 38592 19385 38656
rect 19449 38592 19455 38656
rect 22840 38632 23300 38662
rect 19139 38591 19455 38592
rect 2037 38584 2103 38589
rect 2037 38528 2042 38584
rect 2098 38528 2103 38584
rect 2037 38523 2103 38528
rect 4245 38586 4311 38589
rect 7557 38586 7623 38589
rect 4245 38584 7623 38586
rect 4245 38528 4250 38584
rect 4306 38528 7562 38584
rect 7618 38528 7623 38584
rect 4245 38526 7623 38528
rect 4245 38523 4311 38526
rect 7557 38523 7623 38526
rect 19977 38586 20043 38589
rect 21081 38586 21147 38589
rect 19977 38584 21147 38586
rect 19977 38528 19982 38584
rect 20038 38528 21086 38584
rect 21142 38528 21147 38584
rect 19977 38526 21147 38528
rect 19977 38523 20043 38526
rect 21081 38523 21147 38526
rect -300 38450 160 38480
rect 2040 38450 2100 38523
rect -300 38390 2100 38450
rect 2957 38450 3023 38453
rect 8150 38450 8156 38452
rect 2957 38448 8156 38450
rect 2957 38392 2962 38448
rect 3018 38392 8156 38448
rect 2957 38390 8156 38392
rect -300 38360 160 38390
rect 2957 38387 3023 38390
rect 8150 38388 8156 38390
rect 8220 38450 8226 38452
rect 8293 38450 8359 38453
rect 8220 38448 8359 38450
rect 8220 38392 8298 38448
rect 8354 38392 8359 38448
rect 8220 38390 8359 38392
rect 8220 38388 8226 38390
rect 8293 38387 8359 38390
rect 11053 38450 11119 38453
rect 12566 38450 12572 38452
rect 11053 38448 12572 38450
rect 11053 38392 11058 38448
rect 11114 38392 12572 38448
rect 11053 38390 12572 38392
rect 11053 38387 11119 38390
rect 12566 38388 12572 38390
rect 12636 38388 12642 38452
rect 2865 38314 2931 38317
rect 8569 38314 8635 38317
rect 9581 38314 9647 38317
rect 20253 38314 20319 38317
rect 2730 38312 2931 38314
rect 2730 38256 2870 38312
rect 2926 38256 2931 38312
rect 2730 38254 2931 38256
rect -300 38178 160 38208
rect 2730 38178 2790 38254
rect 2865 38251 2931 38254
rect 5950 38312 9506 38314
rect 5950 38256 8574 38312
rect 8630 38256 9506 38312
rect 5950 38254 9506 38256
rect -300 38118 2790 38178
rect -300 38088 160 38118
rect 5950 38042 6010 38254
rect 8569 38251 8635 38254
rect 7097 38178 7163 38181
rect 7833 38178 7899 38181
rect 7097 38176 7899 38178
rect 7097 38120 7102 38176
rect 7158 38120 7838 38176
rect 7894 38120 7899 38176
rect 7097 38118 7899 38120
rect 7097 38115 7163 38118
rect 7833 38115 7899 38118
rect 6144 38112 6460 38113
rect 6144 38048 6150 38112
rect 6214 38048 6230 38112
rect 6294 38048 6310 38112
rect 6374 38048 6390 38112
rect 6454 38048 6460 38112
rect 6144 38047 6460 38048
rect 2730 37982 6010 38042
rect 9446 38042 9506 38254
rect 9581 38312 20319 38314
rect 9581 38256 9586 38312
rect 9642 38256 20258 38312
rect 20314 38256 20319 38312
rect 9581 38254 20319 38256
rect 9581 38251 9647 38254
rect 20253 38251 20319 38254
rect 22185 38178 22251 38181
rect 22840 38178 23300 38208
rect 22185 38176 23300 38178
rect 22185 38120 22190 38176
rect 22246 38120 23300 38176
rect 22185 38118 23300 38120
rect 22185 38115 22251 38118
rect 11342 38112 11658 38113
rect 11342 38048 11348 38112
rect 11412 38048 11428 38112
rect 11492 38048 11508 38112
rect 11572 38048 11588 38112
rect 11652 38048 11658 38112
rect 11342 38047 11658 38048
rect 16540 38112 16856 38113
rect 16540 38048 16546 38112
rect 16610 38048 16626 38112
rect 16690 38048 16706 38112
rect 16770 38048 16786 38112
rect 16850 38048 16856 38112
rect 16540 38047 16856 38048
rect 21738 38112 22054 38113
rect 21738 38048 21744 38112
rect 21808 38048 21824 38112
rect 21888 38048 21904 38112
rect 21968 38048 21984 38112
rect 22048 38048 22054 38112
rect 22840 38088 23300 38118
rect 21738 38047 22054 38048
rect 9446 37982 11208 38042
rect -300 37906 160 37936
rect 749 37906 815 37909
rect -300 37904 815 37906
rect -300 37848 754 37904
rect 810 37848 815 37904
rect -300 37846 815 37848
rect -300 37816 160 37846
rect 749 37843 815 37846
rect 2405 37906 2471 37909
rect 2730 37906 2790 37982
rect 2405 37904 2790 37906
rect 2405 37848 2410 37904
rect 2466 37848 2790 37904
rect 2405 37846 2790 37848
rect 3417 37906 3483 37909
rect 7557 37906 7623 37909
rect 11148 37906 11208 37982
rect 14181 37906 14247 37909
rect 3417 37904 10058 37906
rect 3417 37848 3422 37904
rect 3478 37848 7562 37904
rect 7618 37848 10058 37904
rect 3417 37846 10058 37848
rect 11148 37904 14247 37906
rect 11148 37848 14186 37904
rect 14242 37848 14247 37904
rect 11148 37846 14247 37848
rect 2405 37843 2471 37846
rect 3417 37843 3483 37846
rect 7557 37843 7623 37846
rect 2405 37770 2471 37773
rect 3969 37770 4035 37773
rect 2405 37768 4035 37770
rect 2405 37712 2410 37768
rect 2466 37712 3974 37768
rect 4030 37712 4035 37768
rect 2405 37710 4035 37712
rect 2405 37707 2471 37710
rect 3969 37707 4035 37710
rect 5349 37770 5415 37773
rect 9806 37770 9812 37772
rect 5349 37768 9812 37770
rect 5349 37712 5354 37768
rect 5410 37712 9812 37768
rect 5349 37710 9812 37712
rect 5349 37707 5415 37710
rect 9806 37708 9812 37710
rect 9876 37708 9882 37772
rect 9998 37770 10058 37846
rect 14181 37843 14247 37846
rect 20069 37770 20135 37773
rect 9998 37768 20135 37770
rect 9998 37712 20074 37768
rect 20130 37712 20135 37768
rect 9998 37710 20135 37712
rect 20069 37707 20135 37710
rect -300 37634 160 37664
rect 1301 37634 1367 37637
rect 4889 37636 4955 37637
rect -300 37632 1367 37634
rect -300 37576 1306 37632
rect 1362 37576 1367 37632
rect -300 37574 1367 37576
rect -300 37544 160 37574
rect 1301 37571 1367 37574
rect 4838 37572 4844 37636
rect 4908 37634 4955 37636
rect 5441 37634 5507 37637
rect 8477 37634 8543 37637
rect 4908 37632 5000 37634
rect 4950 37576 5000 37632
rect 4908 37574 5000 37576
rect 5441 37632 8543 37634
rect 5441 37576 5446 37632
rect 5502 37576 8482 37632
rect 8538 37576 8543 37632
rect 5441 37574 8543 37576
rect 4908 37572 4955 37574
rect 4889 37571 4955 37572
rect 5441 37571 5507 37574
rect 8477 37571 8543 37574
rect 21449 37634 21515 37637
rect 22840 37634 23300 37664
rect 21449 37632 23300 37634
rect 21449 37576 21454 37632
rect 21510 37576 23300 37632
rect 21449 37574 23300 37576
rect 21449 37571 21515 37574
rect 3545 37568 3861 37569
rect 3545 37504 3551 37568
rect 3615 37504 3631 37568
rect 3695 37504 3711 37568
rect 3775 37504 3791 37568
rect 3855 37504 3861 37568
rect 3545 37503 3861 37504
rect 8743 37568 9059 37569
rect 8743 37504 8749 37568
rect 8813 37504 8829 37568
rect 8893 37504 8909 37568
rect 8973 37504 8989 37568
rect 9053 37504 9059 37568
rect 8743 37503 9059 37504
rect 13941 37568 14257 37569
rect 13941 37504 13947 37568
rect 14011 37504 14027 37568
rect 14091 37504 14107 37568
rect 14171 37504 14187 37568
rect 14251 37504 14257 37568
rect 13941 37503 14257 37504
rect 19139 37568 19455 37569
rect 19139 37504 19145 37568
rect 19209 37504 19225 37568
rect 19289 37504 19305 37568
rect 19369 37504 19385 37568
rect 19449 37504 19455 37568
rect 22840 37544 23300 37574
rect 19139 37503 19455 37504
rect -300 37362 160 37392
rect 2773 37362 2839 37365
rect -300 37360 2839 37362
rect -300 37304 2778 37360
rect 2834 37304 2839 37360
rect -300 37302 2839 37304
rect -300 37272 160 37302
rect 2773 37299 2839 37302
rect 7833 37362 7899 37365
rect 7966 37362 7972 37364
rect 7833 37360 7972 37362
rect 7833 37304 7838 37360
rect 7894 37304 7972 37360
rect 7833 37302 7972 37304
rect 7833 37299 7899 37302
rect 7966 37300 7972 37302
rect 8036 37300 8042 37364
rect 9949 37362 10015 37365
rect 13077 37362 13143 37365
rect 9949 37360 13143 37362
rect 9949 37304 9954 37360
rect 10010 37304 13082 37360
rect 13138 37304 13143 37360
rect 9949 37302 13143 37304
rect 9949 37299 10015 37302
rect 13077 37299 13143 37302
rect 1945 37226 2011 37229
rect 8518 37226 8524 37228
rect 1350 37224 2011 37226
rect 1350 37168 1950 37224
rect 2006 37168 2011 37224
rect 1350 37166 2011 37168
rect -300 37090 160 37120
rect 1350 37090 1410 37166
rect 1945 37163 2011 37166
rect 7054 37166 8524 37226
rect -300 37030 1410 37090
rect 6545 37090 6611 37093
rect 7054 37090 7114 37166
rect 8518 37164 8524 37166
rect 8588 37226 8594 37228
rect 11329 37226 11395 37229
rect 8588 37224 11395 37226
rect 8588 37168 11334 37224
rect 11390 37168 11395 37224
rect 8588 37166 11395 37168
rect 8588 37164 8594 37166
rect 11329 37163 11395 37166
rect 12157 37226 12223 37229
rect 14406 37226 14412 37228
rect 12157 37224 14412 37226
rect 12157 37168 12162 37224
rect 12218 37168 14412 37224
rect 12157 37166 14412 37168
rect 12157 37163 12223 37166
rect 14406 37164 14412 37166
rect 14476 37164 14482 37228
rect 6545 37088 7114 37090
rect 6545 37032 6550 37088
rect 6606 37032 7114 37088
rect 6545 37030 7114 37032
rect 7741 37092 7807 37093
rect 7741 37088 7788 37092
rect 7852 37090 7858 37092
rect 22277 37090 22343 37093
rect 22840 37090 23300 37120
rect 7741 37032 7746 37088
rect -300 37000 160 37030
rect 6545 37027 6611 37030
rect 7741 37028 7788 37032
rect 7852 37030 7898 37090
rect 22277 37088 23300 37090
rect 22277 37032 22282 37088
rect 22338 37032 23300 37088
rect 22277 37030 23300 37032
rect 7852 37028 7858 37030
rect 7741 37027 7807 37028
rect 22277 37027 22343 37030
rect 6144 37024 6460 37025
rect 6144 36960 6150 37024
rect 6214 36960 6230 37024
rect 6294 36960 6310 37024
rect 6374 36960 6390 37024
rect 6454 36960 6460 37024
rect 6144 36959 6460 36960
rect 11342 37024 11658 37025
rect 11342 36960 11348 37024
rect 11412 36960 11428 37024
rect 11492 36960 11508 37024
rect 11572 36960 11588 37024
rect 11652 36960 11658 37024
rect 11342 36959 11658 36960
rect 16540 37024 16856 37025
rect 16540 36960 16546 37024
rect 16610 36960 16626 37024
rect 16690 36960 16706 37024
rect 16770 36960 16786 37024
rect 16850 36960 16856 37024
rect 16540 36959 16856 36960
rect 21738 37024 22054 37025
rect 21738 36960 21744 37024
rect 21808 36960 21824 37024
rect 21888 36960 21904 37024
rect 21968 36960 21984 37024
rect 22048 36960 22054 37024
rect 22840 37000 23300 37030
rect 21738 36959 22054 36960
rect 1209 36954 1275 36957
rect 798 36952 1275 36954
rect 798 36896 1214 36952
rect 1270 36896 1275 36952
rect 798 36894 1275 36896
rect -300 36818 160 36848
rect 798 36818 858 36894
rect 1209 36891 1275 36894
rect 2405 36954 2471 36957
rect 5993 36954 6059 36957
rect 2405 36952 6059 36954
rect 2405 36896 2410 36952
rect 2466 36896 5998 36952
rect 6054 36896 6059 36952
rect 2405 36894 6059 36896
rect 2405 36891 2471 36894
rect 5993 36891 6059 36894
rect -300 36758 858 36818
rect 6085 36818 6151 36821
rect 6913 36820 6979 36821
rect 6678 36818 6684 36820
rect 6085 36816 6684 36818
rect 6085 36760 6090 36816
rect 6146 36760 6684 36816
rect 6085 36758 6684 36760
rect -300 36728 160 36758
rect 6085 36755 6151 36758
rect 6678 36756 6684 36758
rect 6748 36756 6754 36820
rect 6862 36756 6868 36820
rect 6932 36818 6979 36820
rect 7557 36818 7623 36821
rect 20069 36818 20135 36821
rect 20529 36818 20595 36821
rect 6932 36816 7024 36818
rect 6974 36760 7024 36816
rect 6932 36758 7024 36760
rect 7557 36816 20595 36818
rect 7557 36760 7562 36816
rect 7618 36760 20074 36816
rect 20130 36760 20534 36816
rect 20590 36760 20595 36816
rect 7557 36758 20595 36760
rect 6932 36756 6979 36758
rect 6913 36755 6979 36756
rect 7557 36755 7623 36758
rect 20069 36755 20135 36758
rect 20529 36755 20595 36758
rect 2262 36620 2268 36684
rect 2332 36682 2338 36684
rect 7230 36682 7236 36684
rect 2332 36622 7236 36682
rect 2332 36620 2338 36622
rect 7230 36620 7236 36622
rect 7300 36682 7306 36684
rect 10225 36682 10291 36685
rect 7300 36680 10291 36682
rect 7300 36624 10230 36680
rect 10286 36624 10291 36680
rect 7300 36622 10291 36624
rect 7300 36620 7306 36622
rect 10225 36619 10291 36622
rect 13905 36682 13971 36685
rect 14774 36682 14780 36684
rect 13905 36680 14780 36682
rect 13905 36624 13910 36680
rect 13966 36624 14780 36680
rect 13905 36622 14780 36624
rect 13905 36619 13971 36622
rect 14774 36620 14780 36622
rect 14844 36682 14850 36684
rect 19977 36682 20043 36685
rect 20529 36682 20595 36685
rect 14844 36680 20595 36682
rect 14844 36624 19982 36680
rect 20038 36624 20534 36680
rect 20590 36624 20595 36680
rect 14844 36622 20595 36624
rect 14844 36620 14850 36622
rect 19977 36619 20043 36622
rect 20529 36619 20595 36622
rect -300 36546 160 36576
rect -300 36486 3250 36546
rect -300 36456 160 36486
rect -300 36274 160 36304
rect 2865 36274 2931 36277
rect -300 36272 2931 36274
rect -300 36216 2870 36272
rect 2926 36216 2931 36272
rect -300 36214 2931 36216
rect 3190 36274 3250 36486
rect 5022 36484 5028 36548
rect 5092 36546 5098 36548
rect 5257 36546 5323 36549
rect 5092 36544 5323 36546
rect 5092 36488 5262 36544
rect 5318 36488 5323 36544
rect 5092 36486 5323 36488
rect 5092 36484 5098 36486
rect 5257 36483 5323 36486
rect 6361 36544 6427 36549
rect 6361 36488 6366 36544
rect 6422 36488 6427 36544
rect 6361 36483 6427 36488
rect 9857 36546 9923 36549
rect 10593 36546 10659 36549
rect 9857 36544 10659 36546
rect 9857 36488 9862 36544
rect 9918 36488 10598 36544
rect 10654 36488 10659 36544
rect 9857 36486 10659 36488
rect 9857 36483 9923 36486
rect 10593 36483 10659 36486
rect 21449 36546 21515 36549
rect 22840 36546 23300 36576
rect 21449 36544 23300 36546
rect 21449 36488 21454 36544
rect 21510 36488 23300 36544
rect 21449 36486 23300 36488
rect 21449 36483 21515 36486
rect 3545 36480 3861 36481
rect 3545 36416 3551 36480
rect 3615 36416 3631 36480
rect 3695 36416 3711 36480
rect 3775 36416 3791 36480
rect 3855 36416 3861 36480
rect 3545 36415 3861 36416
rect 6364 36410 6424 36483
rect 8743 36480 9059 36481
rect 8743 36416 8749 36480
rect 8813 36416 8829 36480
rect 8893 36416 8909 36480
rect 8973 36416 8989 36480
rect 9053 36416 9059 36480
rect 8743 36415 9059 36416
rect 13941 36480 14257 36481
rect 13941 36416 13947 36480
rect 14011 36416 14027 36480
rect 14091 36416 14107 36480
rect 14171 36416 14187 36480
rect 14251 36416 14257 36480
rect 13941 36415 14257 36416
rect 19139 36480 19455 36481
rect 19139 36416 19145 36480
rect 19209 36416 19225 36480
rect 19289 36416 19305 36480
rect 19369 36416 19385 36480
rect 19449 36416 19455 36480
rect 22840 36456 23300 36486
rect 19139 36415 19455 36416
rect 3926 36350 6424 36410
rect 3926 36274 3986 36350
rect 3190 36214 3986 36274
rect 12525 36274 12591 36277
rect 15510 36274 15516 36276
rect 12525 36272 15516 36274
rect 12525 36216 12530 36272
rect 12586 36216 15516 36272
rect 12525 36214 15516 36216
rect -300 36184 160 36214
rect 2865 36211 2931 36214
rect 12525 36211 12591 36214
rect 15510 36212 15516 36214
rect 15580 36212 15586 36276
rect 17718 36212 17724 36276
rect 17788 36212 17794 36276
rect 19425 36274 19491 36277
rect 20437 36274 20503 36277
rect 19425 36272 20503 36274
rect 19425 36216 19430 36272
rect 19486 36216 20442 36272
rect 20498 36216 20503 36272
rect 19425 36214 20503 36216
rect 1761 36138 1827 36141
rect 982 36136 1827 36138
rect 982 36080 1766 36136
rect 1822 36080 1827 36136
rect 982 36078 1827 36080
rect -300 36002 160 36032
rect 982 36002 1042 36078
rect 1761 36075 1827 36078
rect 5441 36138 5507 36141
rect 6913 36138 6979 36141
rect 5441 36136 6979 36138
rect 5441 36080 5446 36136
rect 5502 36080 6918 36136
rect 6974 36080 6979 36136
rect 5441 36078 6979 36080
rect 5441 36075 5507 36078
rect 6913 36075 6979 36078
rect 8661 36138 8727 36141
rect 17726 36138 17786 36212
rect 19425 36211 19491 36214
rect 20437 36211 20503 36214
rect 8661 36136 17786 36138
rect 8661 36080 8666 36136
rect 8722 36080 17786 36136
rect 8661 36078 17786 36080
rect 8661 36075 8727 36078
rect -300 35942 1042 36002
rect -300 35912 160 35942
rect 7598 35940 7604 36004
rect 7668 36002 7674 36004
rect 7741 36002 7807 36005
rect 7668 36000 7807 36002
rect 7668 35944 7746 36000
rect 7802 35944 7807 36000
rect 7668 35942 7807 35944
rect 7668 35940 7674 35942
rect 7741 35939 7807 35942
rect 9397 36002 9463 36005
rect 9990 36002 9996 36004
rect 9397 36000 9996 36002
rect 9397 35944 9402 36000
rect 9458 35944 9996 36000
rect 9397 35942 9996 35944
rect 9397 35939 9463 35942
rect 9990 35940 9996 35942
rect 10060 35940 10066 36004
rect 10726 35940 10732 36004
rect 10796 36002 10802 36004
rect 10961 36002 11027 36005
rect 10796 36000 11027 36002
rect 10796 35944 10966 36000
rect 11022 35944 11027 36000
rect 10796 35942 11027 35944
rect 10796 35940 10802 35942
rect 10961 35939 11027 35942
rect 22277 36002 22343 36005
rect 22840 36002 23300 36032
rect 22277 36000 23300 36002
rect 22277 35944 22282 36000
rect 22338 35944 23300 36000
rect 22277 35942 23300 35944
rect 22277 35939 22343 35942
rect 6144 35936 6460 35937
rect 6144 35872 6150 35936
rect 6214 35872 6230 35936
rect 6294 35872 6310 35936
rect 6374 35872 6390 35936
rect 6454 35872 6460 35936
rect 6144 35871 6460 35872
rect 11342 35936 11658 35937
rect 11342 35872 11348 35936
rect 11412 35872 11428 35936
rect 11492 35872 11508 35936
rect 11572 35872 11588 35936
rect 11652 35872 11658 35936
rect 11342 35871 11658 35872
rect 16540 35936 16856 35937
rect 16540 35872 16546 35936
rect 16610 35872 16626 35936
rect 16690 35872 16706 35936
rect 16770 35872 16786 35936
rect 16850 35872 16856 35936
rect 16540 35871 16856 35872
rect 21738 35936 22054 35937
rect 21738 35872 21744 35936
rect 21808 35872 21824 35936
rect 21888 35872 21904 35936
rect 21968 35872 21984 35936
rect 22048 35872 22054 35936
rect 22840 35912 23300 35942
rect 21738 35871 22054 35872
rect 4245 35866 4311 35869
rect 5758 35866 5764 35868
rect 4245 35864 5764 35866
rect 4245 35808 4250 35864
rect 4306 35808 5764 35864
rect 4245 35806 5764 35808
rect 4245 35803 4311 35806
rect 5758 35804 5764 35806
rect 5828 35804 5834 35868
rect 8334 35804 8340 35868
rect 8404 35866 8410 35868
rect 8661 35866 8727 35869
rect 8404 35864 8727 35866
rect 8404 35808 8666 35864
rect 8722 35808 8727 35864
rect 8404 35806 8727 35808
rect 8404 35804 8410 35806
rect 8661 35803 8727 35806
rect 9397 35866 9463 35869
rect 9949 35866 10015 35869
rect 9397 35864 10015 35866
rect 9397 35808 9402 35864
rect 9458 35808 9954 35864
rect 10010 35808 10015 35864
rect 9397 35806 10015 35808
rect 9397 35803 9463 35806
rect 9949 35803 10015 35806
rect 10317 35866 10383 35869
rect 11094 35866 11100 35868
rect 10317 35864 11100 35866
rect 10317 35808 10322 35864
rect 10378 35808 11100 35864
rect 10317 35806 11100 35808
rect 10317 35803 10383 35806
rect 11094 35804 11100 35806
rect 11164 35804 11170 35868
rect 20161 35866 20227 35869
rect 20437 35866 20503 35869
rect 20161 35864 20503 35866
rect 20161 35808 20166 35864
rect 20222 35808 20442 35864
rect 20498 35808 20503 35864
rect 20161 35806 20503 35808
rect 20161 35803 20227 35806
rect 20437 35803 20503 35806
rect -300 35730 160 35760
rect 289 35730 355 35733
rect 8293 35730 8359 35733
rect -300 35728 355 35730
rect -300 35672 294 35728
rect 350 35672 355 35728
rect -300 35670 355 35672
rect -300 35640 160 35670
rect 289 35667 355 35670
rect 2730 35728 8359 35730
rect 2730 35672 8298 35728
rect 8354 35672 8359 35728
rect 2730 35670 8359 35672
rect 473 35594 539 35597
rect 2730 35594 2790 35670
rect 8293 35667 8359 35670
rect 8569 35730 8635 35733
rect 11605 35730 11671 35733
rect 8569 35728 11671 35730
rect 8569 35672 8574 35728
rect 8630 35672 11610 35728
rect 11666 35672 11671 35728
rect 8569 35670 11671 35672
rect 8569 35667 8635 35670
rect 11605 35667 11671 35670
rect 13813 35730 13879 35733
rect 18321 35730 18387 35733
rect 13813 35728 18387 35730
rect 13813 35672 13818 35728
rect 13874 35672 18326 35728
rect 18382 35672 18387 35728
rect 13813 35670 18387 35672
rect 13813 35667 13879 35670
rect 18321 35667 18387 35670
rect 3509 35594 3575 35597
rect 473 35592 2790 35594
rect 473 35536 478 35592
rect 534 35536 2790 35592
rect 473 35534 2790 35536
rect 3190 35592 3575 35594
rect 3190 35536 3514 35592
rect 3570 35536 3575 35592
rect 3190 35534 3575 35536
rect 473 35531 539 35534
rect -300 35458 160 35488
rect 3190 35458 3250 35534
rect 3509 35531 3575 35534
rect 4889 35594 4955 35597
rect 5809 35594 5875 35597
rect 4889 35592 5875 35594
rect 4889 35536 4894 35592
rect 4950 35536 5814 35592
rect 5870 35536 5875 35592
rect 4889 35534 5875 35536
rect 4889 35531 4955 35534
rect 5809 35531 5875 35534
rect 5993 35594 6059 35597
rect 10225 35594 10291 35597
rect 5993 35592 10291 35594
rect 5993 35536 5998 35592
rect 6054 35536 10230 35592
rect 10286 35536 10291 35592
rect 5993 35534 10291 35536
rect 5993 35531 6059 35534
rect 10225 35531 10291 35534
rect 13077 35594 13143 35597
rect 15326 35594 15332 35596
rect 13077 35592 15332 35594
rect 13077 35536 13082 35592
rect 13138 35536 15332 35592
rect 13077 35534 15332 35536
rect 13077 35531 13143 35534
rect 15326 35532 15332 35534
rect 15396 35594 15402 35596
rect 18045 35594 18111 35597
rect 15396 35592 18111 35594
rect 15396 35536 18050 35592
rect 18106 35536 18111 35592
rect 15396 35534 18111 35536
rect 15396 35532 15402 35534
rect 18045 35531 18111 35534
rect -300 35398 3250 35458
rect -300 35368 160 35398
rect 5390 35396 5396 35460
rect 5460 35458 5466 35460
rect 8477 35458 8543 35461
rect 9397 35460 9463 35461
rect 9397 35458 9444 35460
rect 5460 35456 8543 35458
rect 5460 35400 8482 35456
rect 8538 35400 8543 35456
rect 5460 35398 8543 35400
rect 9352 35456 9444 35458
rect 9352 35400 9402 35456
rect 9352 35398 9444 35400
rect 5460 35396 5466 35398
rect 8477 35395 8543 35398
rect 9397 35396 9444 35398
rect 9508 35396 9514 35460
rect 21449 35458 21515 35461
rect 22840 35458 23300 35488
rect 21449 35456 23300 35458
rect 21449 35400 21454 35456
rect 21510 35400 23300 35456
rect 21449 35398 23300 35400
rect 9397 35395 9463 35396
rect 21449 35395 21515 35398
rect 3545 35392 3861 35393
rect 3545 35328 3551 35392
rect 3615 35328 3631 35392
rect 3695 35328 3711 35392
rect 3775 35328 3791 35392
rect 3855 35328 3861 35392
rect 3545 35327 3861 35328
rect 8743 35392 9059 35393
rect 8743 35328 8749 35392
rect 8813 35328 8829 35392
rect 8893 35328 8909 35392
rect 8973 35328 8989 35392
rect 9053 35328 9059 35392
rect 8743 35327 9059 35328
rect 13941 35392 14257 35393
rect 13941 35328 13947 35392
rect 14011 35328 14027 35392
rect 14091 35328 14107 35392
rect 14171 35328 14187 35392
rect 14251 35328 14257 35392
rect 13941 35327 14257 35328
rect 19139 35392 19455 35393
rect 19139 35328 19145 35392
rect 19209 35328 19225 35392
rect 19289 35328 19305 35392
rect 19369 35328 19385 35392
rect 19449 35328 19455 35392
rect 22840 35368 23300 35398
rect 19139 35327 19455 35328
rect 1669 35324 1735 35325
rect 1669 35322 1716 35324
rect 1624 35320 1716 35322
rect 1624 35264 1674 35320
rect 1624 35262 1716 35264
rect 1669 35260 1716 35262
rect 1780 35260 1786 35324
rect 2446 35260 2452 35324
rect 2516 35322 2522 35324
rect 3417 35322 3483 35325
rect 2516 35320 3483 35322
rect 2516 35264 3422 35320
rect 3478 35264 3483 35320
rect 2516 35262 3483 35264
rect 2516 35260 2522 35262
rect 1669 35259 1735 35260
rect 3417 35259 3483 35262
rect 5257 35322 5323 35325
rect 9489 35322 9555 35325
rect 9765 35322 9831 35325
rect 5257 35320 7988 35322
rect 5257 35264 5262 35320
rect 5318 35264 7988 35320
rect 5257 35262 7988 35264
rect 5257 35259 5323 35262
rect -300 35186 160 35216
rect 7928 35189 7988 35262
rect 9489 35320 9831 35322
rect 9489 35264 9494 35320
rect 9550 35264 9770 35320
rect 9826 35264 9831 35320
rect 9489 35262 9831 35264
rect 9489 35259 9555 35262
rect 9765 35259 9831 35262
rect 14825 35322 14891 35325
rect 17309 35322 17375 35325
rect 14825 35320 17375 35322
rect 14825 35264 14830 35320
rect 14886 35264 17314 35320
rect 17370 35264 17375 35320
rect 14825 35262 17375 35264
rect 14825 35259 14891 35262
rect 17309 35259 17375 35262
rect 3049 35186 3115 35189
rect 3509 35186 3575 35189
rect -300 35184 3115 35186
rect -300 35128 3054 35184
rect 3110 35128 3115 35184
rect -300 35126 3115 35128
rect -300 35096 160 35126
rect 3049 35123 3115 35126
rect 3374 35184 3575 35186
rect 3374 35128 3514 35184
rect 3570 35128 3575 35184
rect 3374 35126 3575 35128
rect 1209 35050 1275 35053
rect 798 35048 1275 35050
rect 798 34992 1214 35048
rect 1270 34992 1275 35048
rect 798 34990 1275 34992
rect -300 34914 160 34944
rect 798 34914 858 34990
rect 1209 34987 1275 34990
rect 1485 35048 1551 35053
rect 1485 34992 1490 35048
rect 1546 34992 1551 35048
rect 1485 34987 1551 34992
rect 3049 35050 3115 35053
rect 3374 35050 3434 35126
rect 3509 35123 3575 35126
rect 4061 35186 4127 35189
rect 7649 35186 7715 35189
rect 4061 35184 7715 35186
rect 4061 35128 4066 35184
rect 4122 35128 7654 35184
rect 7710 35128 7715 35184
rect 4061 35126 7715 35128
rect 4061 35123 4127 35126
rect 7649 35123 7715 35126
rect 7925 35186 7991 35189
rect 10317 35186 10383 35189
rect 7925 35184 10383 35186
rect 7925 35128 7930 35184
rect 7986 35128 10322 35184
rect 10378 35128 10383 35184
rect 7925 35126 10383 35128
rect 7925 35123 7991 35126
rect 10317 35123 10383 35126
rect 10869 35186 10935 35189
rect 18413 35186 18479 35189
rect 10869 35184 18479 35186
rect 10869 35128 10874 35184
rect 10930 35128 18418 35184
rect 18474 35128 18479 35184
rect 10869 35126 18479 35128
rect 10869 35123 10935 35126
rect 18413 35123 18479 35126
rect 3049 35048 3434 35050
rect 3049 34992 3054 35048
rect 3110 34992 3434 35048
rect 3049 34990 3434 34992
rect 3509 35050 3575 35053
rect 18229 35050 18295 35053
rect 3509 35048 18295 35050
rect 3509 34992 3514 35048
rect 3570 34992 18234 35048
rect 18290 34992 18295 35048
rect 3509 34990 18295 34992
rect 3049 34987 3115 34990
rect 3509 34987 3575 34990
rect 18229 34987 18295 34990
rect -300 34854 858 34914
rect -300 34824 160 34854
rect -300 34642 160 34672
rect 1488 34642 1548 34987
rect 3233 34914 3299 34917
rect 5993 34916 6059 34917
rect 5942 34914 5948 34916
rect 3233 34912 5948 34914
rect 6012 34912 6059 34916
rect 3233 34856 3238 34912
rect 3294 34856 5948 34912
rect 6054 34856 6059 34912
rect 3233 34854 5948 34856
rect 3233 34851 3299 34854
rect 5942 34852 5948 34854
rect 6012 34852 6059 34856
rect 5993 34851 6059 34852
rect 22185 34914 22251 34917
rect 22840 34914 23300 34944
rect 22185 34912 23300 34914
rect 22185 34856 22190 34912
rect 22246 34856 23300 34912
rect 22185 34854 23300 34856
rect 22185 34851 22251 34854
rect 6144 34848 6460 34849
rect 6144 34784 6150 34848
rect 6214 34784 6230 34848
rect 6294 34784 6310 34848
rect 6374 34784 6390 34848
rect 6454 34784 6460 34848
rect 6144 34783 6460 34784
rect 11342 34848 11658 34849
rect 11342 34784 11348 34848
rect 11412 34784 11428 34848
rect 11492 34784 11508 34848
rect 11572 34784 11588 34848
rect 11652 34784 11658 34848
rect 11342 34783 11658 34784
rect 16540 34848 16856 34849
rect 16540 34784 16546 34848
rect 16610 34784 16626 34848
rect 16690 34784 16706 34848
rect 16770 34784 16786 34848
rect 16850 34784 16856 34848
rect 16540 34783 16856 34784
rect 21738 34848 22054 34849
rect 21738 34784 21744 34848
rect 21808 34784 21824 34848
rect 21888 34784 21904 34848
rect 21968 34784 21984 34848
rect 22048 34784 22054 34848
rect 22840 34824 23300 34854
rect 21738 34783 22054 34784
rect 8201 34778 8267 34781
rect -300 34582 1548 34642
rect 1856 34718 4538 34778
rect -300 34552 160 34582
rect 974 34444 980 34508
rect 1044 34506 1050 34508
rect 1856 34506 1916 34718
rect 2998 34580 3004 34644
rect 3068 34642 3074 34644
rect 3785 34642 3851 34645
rect 4245 34642 4311 34645
rect 3068 34640 3851 34642
rect 3068 34584 3790 34640
rect 3846 34584 3851 34640
rect 3068 34582 3851 34584
rect 3068 34580 3074 34582
rect 3785 34579 3851 34582
rect 4110 34640 4311 34642
rect 4110 34584 4250 34640
rect 4306 34584 4311 34640
rect 4110 34582 4311 34584
rect 4110 34506 4170 34582
rect 4245 34579 4311 34582
rect 1044 34446 1916 34506
rect 2730 34446 4170 34506
rect 4478 34506 4538 34718
rect 6686 34776 8267 34778
rect 6686 34720 8206 34776
rect 8262 34720 8267 34776
rect 6686 34718 8267 34720
rect 4613 34642 4679 34645
rect 6686 34642 6746 34718
rect 8201 34715 8267 34718
rect 8569 34778 8635 34781
rect 8569 34776 11162 34778
rect 8569 34720 8574 34776
rect 8630 34720 11162 34776
rect 8569 34718 11162 34720
rect 8569 34715 8635 34718
rect 4613 34640 6746 34642
rect 4613 34584 4618 34640
rect 4674 34584 6746 34640
rect 4613 34582 6746 34584
rect 6821 34642 6887 34645
rect 9673 34642 9739 34645
rect 6821 34640 9739 34642
rect 6821 34584 6826 34640
rect 6882 34584 9678 34640
rect 9734 34584 9739 34640
rect 6821 34582 9739 34584
rect 4613 34579 4679 34582
rect 6821 34579 6887 34582
rect 9673 34579 9739 34582
rect 9949 34642 10015 34645
rect 10910 34642 10916 34644
rect 9949 34640 10916 34642
rect 9949 34584 9954 34640
rect 10010 34584 10916 34640
rect 9949 34582 10916 34584
rect 9949 34579 10015 34582
rect 10910 34580 10916 34582
rect 10980 34580 10986 34644
rect 11102 34642 11162 34718
rect 11789 34644 11855 34645
rect 11789 34642 11836 34644
rect 11102 34640 11836 34642
rect 11102 34584 11794 34640
rect 11102 34582 11836 34584
rect 11789 34580 11836 34582
rect 11900 34580 11906 34644
rect 11789 34579 11855 34580
rect 10869 34506 10935 34509
rect 4478 34504 10935 34506
rect 4478 34448 10874 34504
rect 10930 34448 10935 34504
rect 4478 34446 10935 34448
rect 1044 34444 1050 34446
rect -300 34370 160 34400
rect 2730 34370 2790 34446
rect 10869 34443 10935 34446
rect 13721 34506 13787 34509
rect 14825 34506 14891 34509
rect 13721 34504 14891 34506
rect 13721 34448 13726 34504
rect 13782 34448 14830 34504
rect 14886 34448 14891 34504
rect 13721 34446 14891 34448
rect 13721 34443 13787 34446
rect 14825 34443 14891 34446
rect 18597 34506 18663 34509
rect 21030 34506 21036 34508
rect 18597 34504 21036 34506
rect 18597 34448 18602 34504
rect 18658 34448 21036 34504
rect 18597 34446 21036 34448
rect 18597 34443 18663 34446
rect 21030 34444 21036 34446
rect 21100 34444 21106 34508
rect -300 34310 2790 34370
rect 21449 34370 21515 34373
rect 22840 34370 23300 34400
rect 21449 34368 23300 34370
rect 21449 34312 21454 34368
rect 21510 34312 23300 34368
rect 21449 34310 23300 34312
rect -300 34280 160 34310
rect 21449 34307 21515 34310
rect 3545 34304 3861 34305
rect 3545 34240 3551 34304
rect 3615 34240 3631 34304
rect 3695 34240 3711 34304
rect 3775 34240 3791 34304
rect 3855 34240 3861 34304
rect 3545 34239 3861 34240
rect 8743 34304 9059 34305
rect 8743 34240 8749 34304
rect 8813 34240 8829 34304
rect 8893 34240 8909 34304
rect 8973 34240 8989 34304
rect 9053 34240 9059 34304
rect 8743 34239 9059 34240
rect 13941 34304 14257 34305
rect 13941 34240 13947 34304
rect 14011 34240 14027 34304
rect 14091 34240 14107 34304
rect 14171 34240 14187 34304
rect 14251 34240 14257 34304
rect 13941 34239 14257 34240
rect 19139 34304 19455 34305
rect 19139 34240 19145 34304
rect 19209 34240 19225 34304
rect 19289 34240 19305 34304
rect 19369 34240 19385 34304
rect 19449 34240 19455 34304
rect 22840 34280 23300 34310
rect 19139 34239 19455 34240
rect 6453 34234 6519 34237
rect 6678 34234 6684 34236
rect 6453 34232 6684 34234
rect 6453 34176 6458 34232
rect 6514 34176 6684 34232
rect 6453 34174 6684 34176
rect 6453 34171 6519 34174
rect 6678 34172 6684 34174
rect 6748 34172 6754 34236
rect -300 34098 160 34128
rect 4061 34098 4127 34101
rect -300 34096 4127 34098
rect -300 34040 4066 34096
rect 4122 34040 4127 34096
rect -300 34038 4127 34040
rect -300 34008 160 34038
rect 4061 34035 4127 34038
rect 5533 34098 5599 34101
rect 9213 34098 9279 34101
rect 11697 34098 11763 34101
rect 5533 34096 9279 34098
rect 5533 34040 5538 34096
rect 5594 34040 9218 34096
rect 9274 34040 9279 34096
rect 5533 34038 9279 34040
rect 5533 34035 5599 34038
rect 9213 34035 9279 34038
rect 11102 34096 11763 34098
rect 11102 34040 11702 34096
rect 11758 34040 11763 34096
rect 11102 34038 11763 34040
rect 1669 33962 1735 33965
rect 3918 33962 3924 33964
rect 1669 33960 3924 33962
rect 1669 33904 1674 33960
rect 1730 33904 3924 33960
rect 1669 33902 3924 33904
rect 1669 33899 1735 33902
rect 3918 33900 3924 33902
rect 3988 33962 3994 33964
rect 8017 33962 8083 33965
rect 3988 33960 8083 33962
rect 3988 33904 8022 33960
rect 8078 33904 8083 33960
rect 3988 33902 8083 33904
rect 3988 33900 3994 33902
rect 8017 33899 8083 33902
rect 8201 33962 8267 33965
rect 11102 33962 11162 34038
rect 11697 34035 11763 34038
rect 11881 34098 11947 34101
rect 18086 34098 18092 34100
rect 11881 34096 18092 34098
rect 11881 34040 11886 34096
rect 11942 34040 18092 34096
rect 11881 34038 18092 34040
rect 11881 34035 11947 34038
rect 18086 34036 18092 34038
rect 18156 34036 18162 34100
rect 22737 34098 22803 34101
rect 18278 34096 22803 34098
rect 18278 34040 22742 34096
rect 22798 34040 22803 34096
rect 18278 34038 22803 34040
rect 8201 33960 11162 33962
rect 8201 33904 8206 33960
rect 8262 33904 11162 33960
rect 8201 33902 11162 33904
rect 11237 33962 11303 33965
rect 18278 33962 18338 34038
rect 22737 34035 22803 34038
rect 11237 33960 18338 33962
rect 11237 33904 11242 33960
rect 11298 33904 18338 33960
rect 11237 33902 18338 33904
rect 8201 33899 8267 33902
rect 11237 33899 11303 33902
rect -300 33826 160 33856
rect 3141 33826 3207 33829
rect -300 33824 3207 33826
rect -300 33768 3146 33824
rect 3202 33768 3207 33824
rect -300 33766 3207 33768
rect -300 33736 160 33766
rect 3141 33763 3207 33766
rect 15837 33828 15903 33829
rect 15837 33824 15884 33828
rect 15948 33826 15954 33828
rect 22185 33826 22251 33829
rect 22840 33826 23300 33856
rect 15837 33768 15842 33824
rect 15837 33764 15884 33768
rect 15948 33766 15994 33826
rect 22185 33824 23300 33826
rect 22185 33768 22190 33824
rect 22246 33768 23300 33824
rect 22185 33766 23300 33768
rect 15948 33764 15954 33766
rect 15837 33763 15903 33764
rect 22185 33763 22251 33766
rect 6144 33760 6460 33761
rect 6144 33696 6150 33760
rect 6214 33696 6230 33760
rect 6294 33696 6310 33760
rect 6374 33696 6390 33760
rect 6454 33696 6460 33760
rect 6144 33695 6460 33696
rect 11342 33760 11658 33761
rect 11342 33696 11348 33760
rect 11412 33696 11428 33760
rect 11492 33696 11508 33760
rect 11572 33696 11588 33760
rect 11652 33696 11658 33760
rect 11342 33695 11658 33696
rect 16540 33760 16856 33761
rect 16540 33696 16546 33760
rect 16610 33696 16626 33760
rect 16690 33696 16706 33760
rect 16770 33696 16786 33760
rect 16850 33696 16856 33760
rect 16540 33695 16856 33696
rect 21738 33760 22054 33761
rect 21738 33696 21744 33760
rect 21808 33696 21824 33760
rect 21888 33696 21904 33760
rect 21968 33696 21984 33760
rect 22048 33696 22054 33760
rect 22840 33736 23300 33766
rect 21738 33695 22054 33696
rect 1853 33690 1919 33693
rect 3182 33690 3188 33692
rect 1853 33688 3188 33690
rect 1853 33632 1858 33688
rect 1914 33632 3188 33688
rect 1853 33630 3188 33632
rect 1853 33627 1919 33630
rect 3182 33628 3188 33630
rect 3252 33628 3258 33692
rect 3877 33690 3943 33693
rect 3374 33688 3943 33690
rect 3374 33632 3882 33688
rect 3938 33632 3943 33688
rect 3374 33630 3943 33632
rect -300 33554 160 33584
rect 3374 33554 3434 33630
rect 3877 33627 3943 33630
rect 11789 33690 11855 33693
rect 11789 33688 15946 33690
rect 11789 33632 11794 33688
rect 11850 33632 15946 33688
rect 11789 33630 15946 33632
rect 11789 33627 11855 33630
rect -300 33494 3434 33554
rect 4613 33554 4679 33557
rect 12750 33554 12756 33556
rect 4613 33552 12756 33554
rect 4613 33496 4618 33552
rect 4674 33496 12756 33552
rect 4613 33494 12756 33496
rect -300 33464 160 33494
rect 4613 33491 4679 33494
rect 12750 33492 12756 33494
rect 12820 33492 12826 33556
rect 12985 33554 13051 33557
rect 15886 33554 15946 33630
rect 17902 33628 17908 33692
rect 17972 33690 17978 33692
rect 21541 33690 21607 33693
rect 17972 33688 21607 33690
rect 17972 33632 21546 33688
rect 21602 33632 21607 33688
rect 17972 33630 21607 33632
rect 17972 33628 17978 33630
rect 21541 33627 21607 33630
rect 19333 33554 19399 33557
rect 12985 33552 14796 33554
rect 12985 33496 12990 33552
rect 13046 33496 14796 33552
rect 12985 33494 14796 33496
rect 15886 33552 19399 33554
rect 15886 33496 19338 33552
rect 19394 33496 19399 33552
rect 15886 33494 19399 33496
rect 12985 33491 13051 33494
rect 1526 33356 1532 33420
rect 1596 33418 1602 33420
rect 10777 33418 10843 33421
rect 1596 33416 10843 33418
rect 1596 33360 10782 33416
rect 10838 33360 10843 33416
rect 1596 33358 10843 33360
rect 1596 33356 1602 33358
rect 10777 33355 10843 33358
rect 11053 33418 11119 33421
rect 14549 33418 14615 33421
rect 11053 33416 14615 33418
rect 11053 33360 11058 33416
rect 11114 33360 14554 33416
rect 14610 33360 14615 33416
rect 11053 33358 14615 33360
rect 14736 33418 14796 33494
rect 19333 33491 19399 33494
rect 17217 33418 17283 33421
rect 14736 33416 17283 33418
rect 14736 33360 17222 33416
rect 17278 33360 17283 33416
rect 14736 33358 17283 33360
rect 11053 33355 11119 33358
rect 14549 33355 14615 33358
rect 17217 33355 17283 33358
rect -300 33282 160 33312
rect 1485 33282 1551 33285
rect -300 33280 1551 33282
rect -300 33224 1490 33280
rect 1546 33224 1551 33280
rect -300 33222 1551 33224
rect -300 33192 160 33222
rect 1485 33219 1551 33222
rect 4797 33282 4863 33285
rect 5022 33282 5028 33284
rect 4797 33280 5028 33282
rect 4797 33224 4802 33280
rect 4858 33224 5028 33280
rect 4797 33222 5028 33224
rect 4797 33219 4863 33222
rect 5022 33220 5028 33222
rect 5092 33220 5098 33284
rect 14549 33282 14615 33285
rect 18321 33282 18387 33285
rect 14549 33280 18387 33282
rect 14549 33224 14554 33280
rect 14610 33224 18326 33280
rect 18382 33224 18387 33280
rect 14549 33222 18387 33224
rect 14549 33219 14615 33222
rect 18321 33219 18387 33222
rect 21265 33282 21331 33285
rect 22840 33282 23300 33312
rect 21265 33280 23300 33282
rect 21265 33224 21270 33280
rect 21326 33224 23300 33280
rect 21265 33222 23300 33224
rect 21265 33219 21331 33222
rect 3545 33216 3861 33217
rect 3545 33152 3551 33216
rect 3615 33152 3631 33216
rect 3695 33152 3711 33216
rect 3775 33152 3791 33216
rect 3855 33152 3861 33216
rect 3545 33151 3861 33152
rect 8743 33216 9059 33217
rect 8743 33152 8749 33216
rect 8813 33152 8829 33216
rect 8893 33152 8909 33216
rect 8973 33152 8989 33216
rect 9053 33152 9059 33216
rect 8743 33151 9059 33152
rect 13941 33216 14257 33217
rect 13941 33152 13947 33216
rect 14011 33152 14027 33216
rect 14091 33152 14107 33216
rect 14171 33152 14187 33216
rect 14251 33152 14257 33216
rect 13941 33151 14257 33152
rect 19139 33216 19455 33217
rect 19139 33152 19145 33216
rect 19209 33152 19225 33216
rect 19289 33152 19305 33216
rect 19369 33152 19385 33216
rect 19449 33152 19455 33216
rect 22840 33192 23300 33222
rect 19139 33151 19455 33152
rect 4838 33146 4844 33148
rect 4800 33084 4844 33146
rect 4908 33146 4914 33148
rect 11789 33146 11855 33149
rect 12014 33146 12020 33148
rect 4908 33086 8402 33146
rect 4908 33084 4914 33086
rect -300 33010 160 33040
rect 3325 33010 3391 33013
rect -300 33008 3391 33010
rect -300 32952 3330 33008
rect 3386 32952 3391 33008
rect -300 32950 3391 32952
rect -300 32920 160 32950
rect 3325 32947 3391 32950
rect 3785 33010 3851 33013
rect 4800 33010 4860 33084
rect 3785 33008 4860 33010
rect 3785 32952 3790 33008
rect 3846 32952 4860 33008
rect 3785 32950 4860 32952
rect 5073 33010 5139 33013
rect 8342 33012 8402 33086
rect 11789 33144 12020 33146
rect 11789 33088 11794 33144
rect 11850 33088 12020 33144
rect 11789 33086 12020 33088
rect 11789 33083 11855 33086
rect 12014 33084 12020 33086
rect 12084 33084 12090 33148
rect 15142 33084 15148 33148
rect 15212 33146 15218 33148
rect 15377 33146 15443 33149
rect 15212 33144 15443 33146
rect 15212 33088 15382 33144
rect 15438 33088 15443 33144
rect 15212 33086 15443 33088
rect 15212 33084 15218 33086
rect 15377 33083 15443 33086
rect 5073 33008 7850 33010
rect 5073 32952 5078 33008
rect 5134 32952 7850 33008
rect 5073 32950 7850 32952
rect 3785 32947 3851 32950
rect 5073 32947 5139 32950
rect 3233 32876 3299 32877
rect 3182 32874 3188 32876
rect 3106 32814 3188 32874
rect 3252 32874 3299 32876
rect 7649 32874 7715 32877
rect 3252 32872 7715 32874
rect 3294 32816 7654 32872
rect 7710 32816 7715 32872
rect 3182 32812 3188 32814
rect 3252 32814 7715 32816
rect 7790 32874 7850 32950
rect 8334 32948 8340 33012
rect 8404 33010 8410 33012
rect 13629 33010 13695 33013
rect 15745 33010 15811 33013
rect 8404 33008 15811 33010
rect 8404 32952 13634 33008
rect 13690 32952 15750 33008
rect 15806 32952 15811 33008
rect 8404 32950 15811 32952
rect 8404 32948 8410 32950
rect 13629 32947 13695 32950
rect 15745 32947 15811 32950
rect 21173 33010 21239 33013
rect 21173 33008 22202 33010
rect 21173 32952 21178 33008
rect 21234 32952 22202 33008
rect 21173 32950 22202 32952
rect 21173 32947 21239 32950
rect 12525 32874 12591 32877
rect 7790 32872 12591 32874
rect 7790 32816 12530 32872
rect 12586 32816 12591 32872
rect 7790 32814 12591 32816
rect 3252 32812 3299 32814
rect 3233 32811 3299 32812
rect 7649 32811 7715 32814
rect 12525 32811 12591 32814
rect 14917 32874 14983 32877
rect 15694 32874 15700 32876
rect 14917 32872 15700 32874
rect 14917 32816 14922 32872
rect 14978 32816 15700 32872
rect 14917 32814 15700 32816
rect 14917 32811 14983 32814
rect 15694 32812 15700 32814
rect 15764 32812 15770 32876
rect 18965 32874 19031 32877
rect 20294 32874 20300 32876
rect 18965 32872 20300 32874
rect 18965 32816 18970 32872
rect 19026 32816 20300 32872
rect 18965 32814 20300 32816
rect 18965 32811 19031 32814
rect 20294 32812 20300 32814
rect 20364 32812 20370 32876
rect -300 32738 160 32768
rect 2957 32738 3023 32741
rect -300 32736 3023 32738
rect -300 32680 2962 32736
rect 3018 32680 3023 32736
rect -300 32678 3023 32680
rect -300 32648 160 32678
rect 2957 32675 3023 32678
rect 8937 32738 9003 32741
rect 11053 32738 11119 32741
rect 8937 32736 11119 32738
rect 8937 32680 8942 32736
rect 8998 32680 11058 32736
rect 11114 32680 11119 32736
rect 8937 32678 11119 32680
rect 8937 32675 9003 32678
rect 11053 32675 11119 32678
rect 11881 32738 11947 32741
rect 14774 32738 14780 32740
rect 11881 32736 14780 32738
rect 11881 32680 11886 32736
rect 11942 32680 14780 32736
rect 11881 32678 14780 32680
rect 11881 32675 11947 32678
rect 14774 32676 14780 32678
rect 14844 32676 14850 32740
rect 22142 32738 22202 32950
rect 22840 32738 23300 32768
rect 22142 32678 23300 32738
rect 6144 32672 6460 32673
rect 6144 32608 6150 32672
rect 6214 32608 6230 32672
rect 6294 32608 6310 32672
rect 6374 32608 6390 32672
rect 6454 32608 6460 32672
rect 6144 32607 6460 32608
rect 11342 32672 11658 32673
rect 11342 32608 11348 32672
rect 11412 32608 11428 32672
rect 11492 32608 11508 32672
rect 11572 32608 11588 32672
rect 11652 32608 11658 32672
rect 11342 32607 11658 32608
rect 16540 32672 16856 32673
rect 16540 32608 16546 32672
rect 16610 32608 16626 32672
rect 16690 32608 16706 32672
rect 16770 32608 16786 32672
rect 16850 32608 16856 32672
rect 16540 32607 16856 32608
rect 21738 32672 22054 32673
rect 21738 32608 21744 32672
rect 21808 32608 21824 32672
rect 21888 32608 21904 32672
rect 21968 32608 21984 32672
rect 22048 32608 22054 32672
rect 22840 32648 23300 32678
rect 21738 32607 22054 32608
rect 12065 32602 12131 32605
rect 14917 32602 14983 32605
rect 11792 32600 14983 32602
rect 11792 32544 12070 32600
rect 12126 32544 14922 32600
rect 14978 32544 14983 32600
rect 11792 32542 14983 32544
rect -300 32466 160 32496
rect 1853 32466 1919 32469
rect -300 32464 1919 32466
rect -300 32408 1858 32464
rect 1914 32408 1919 32464
rect -300 32406 1919 32408
rect -300 32376 160 32406
rect 1853 32403 1919 32406
rect 2221 32466 2287 32469
rect 4061 32466 4127 32469
rect 10685 32466 10751 32469
rect 11792 32466 11852 32542
rect 12065 32539 12131 32542
rect 14917 32539 14983 32542
rect 2221 32464 9690 32466
rect 2221 32408 2226 32464
rect 2282 32408 4066 32464
rect 4122 32408 9690 32464
rect 2221 32406 9690 32408
rect 2221 32403 2287 32406
rect 4061 32403 4127 32406
rect 1761 32330 1827 32333
rect 1894 32330 1900 32332
rect 1761 32328 1900 32330
rect 1761 32272 1766 32328
rect 1822 32272 1900 32328
rect 1761 32270 1900 32272
rect 1761 32267 1827 32270
rect 1894 32268 1900 32270
rect 1964 32268 1970 32332
rect 2957 32330 3023 32333
rect 5993 32330 6059 32333
rect 2957 32328 6059 32330
rect 2957 32272 2962 32328
rect 3018 32272 5998 32328
rect 6054 32272 6059 32328
rect 2957 32270 6059 32272
rect 2957 32267 3023 32270
rect 5993 32267 6059 32270
rect 6821 32332 6887 32333
rect 6821 32328 6868 32332
rect 6932 32330 6938 32332
rect 8569 32330 8635 32333
rect 9630 32330 9690 32406
rect 10685 32464 11852 32466
rect 10685 32408 10690 32464
rect 10746 32408 11852 32464
rect 10685 32406 11852 32408
rect 12157 32466 12223 32469
rect 17861 32466 17927 32469
rect 12157 32464 17927 32466
rect 12157 32408 12162 32464
rect 12218 32408 17866 32464
rect 17922 32408 17927 32464
rect 12157 32406 17927 32408
rect 10685 32403 10751 32406
rect 12157 32403 12223 32406
rect 17861 32403 17927 32406
rect 9765 32330 9831 32333
rect 6821 32272 6826 32328
rect 6821 32268 6868 32272
rect 6932 32270 6978 32330
rect 8569 32328 9322 32330
rect 8569 32272 8574 32328
rect 8630 32272 9322 32328
rect 8569 32270 9322 32272
rect 9630 32328 9831 32330
rect 9630 32272 9770 32328
rect 9826 32272 9831 32328
rect 9630 32270 9831 32272
rect 6932 32268 6938 32270
rect 6821 32267 6887 32268
rect 8569 32267 8635 32270
rect -300 32194 160 32224
rect 1853 32194 1919 32197
rect -300 32192 1919 32194
rect -300 32136 1858 32192
rect 1914 32136 1919 32192
rect -300 32134 1919 32136
rect -300 32104 160 32134
rect 1853 32131 1919 32134
rect 4705 32194 4771 32197
rect 7925 32194 7991 32197
rect 4705 32192 7991 32194
rect 4705 32136 4710 32192
rect 4766 32136 7930 32192
rect 7986 32136 7991 32192
rect 4705 32134 7991 32136
rect 4705 32131 4771 32134
rect 7925 32131 7991 32134
rect 3545 32128 3861 32129
rect 3545 32064 3551 32128
rect 3615 32064 3631 32128
rect 3695 32064 3711 32128
rect 3775 32064 3791 32128
rect 3855 32064 3861 32128
rect 3545 32063 3861 32064
rect 8743 32128 9059 32129
rect 8743 32064 8749 32128
rect 8813 32064 8829 32128
rect 8893 32064 8909 32128
rect 8973 32064 8989 32128
rect 9053 32064 9059 32128
rect 8743 32063 9059 32064
rect 4245 32058 4311 32061
rect 5165 32058 5231 32061
rect 4245 32056 5231 32058
rect 4245 32000 4250 32056
rect 4306 32000 5170 32056
rect 5226 32000 5231 32056
rect 4245 31998 5231 32000
rect 4245 31995 4311 31998
rect 5165 31995 5231 31998
rect 7649 32058 7715 32061
rect 8477 32058 8543 32061
rect 7649 32056 8543 32058
rect 7649 32000 7654 32056
rect 7710 32000 8482 32056
rect 8538 32000 8543 32056
rect 7649 31998 8543 32000
rect 9262 32058 9322 32270
rect 9765 32267 9831 32270
rect 10961 32330 11027 32333
rect 11881 32330 11947 32333
rect 10961 32328 11947 32330
rect 10961 32272 10966 32328
rect 11022 32272 11886 32328
rect 11942 32272 11947 32328
rect 10961 32270 11947 32272
rect 10961 32267 11027 32270
rect 11881 32267 11947 32270
rect 13169 32328 13235 32333
rect 13997 32330 14063 32333
rect 13169 32272 13174 32328
rect 13230 32272 13235 32328
rect 13169 32267 13235 32272
rect 13816 32328 14063 32330
rect 13816 32272 14002 32328
rect 14058 32272 14063 32328
rect 13816 32270 14063 32272
rect 9622 32132 9628 32196
rect 9692 32194 9698 32196
rect 9990 32194 9996 32196
rect 9692 32134 9996 32194
rect 9692 32132 9698 32134
rect 9990 32132 9996 32134
rect 10060 32132 10066 32196
rect 10409 32194 10475 32197
rect 13172 32194 13232 32267
rect 10409 32192 13232 32194
rect 10409 32136 10414 32192
rect 10470 32136 13232 32192
rect 10409 32134 13232 32136
rect 10409 32131 10475 32134
rect 10358 32058 10364 32060
rect 9262 31998 10364 32058
rect 7649 31995 7715 31998
rect 8477 31995 8543 31998
rect 10358 31996 10364 31998
rect 10428 31996 10434 32060
rect 13169 32058 13235 32061
rect 13816 32058 13876 32270
rect 13997 32267 14063 32270
rect 21449 32194 21515 32197
rect 22840 32194 23300 32224
rect 21449 32192 23300 32194
rect 21449 32136 21454 32192
rect 21510 32136 23300 32192
rect 21449 32134 23300 32136
rect 21449 32131 21515 32134
rect 13941 32128 14257 32129
rect 13941 32064 13947 32128
rect 14011 32064 14027 32128
rect 14091 32064 14107 32128
rect 14171 32064 14187 32128
rect 14251 32064 14257 32128
rect 13941 32063 14257 32064
rect 19139 32128 19455 32129
rect 19139 32064 19145 32128
rect 19209 32064 19225 32128
rect 19289 32064 19305 32128
rect 19369 32064 19385 32128
rect 19449 32064 19455 32128
rect 22840 32104 23300 32134
rect 19139 32063 19455 32064
rect 13169 32056 13876 32058
rect 13169 32000 13174 32056
rect 13230 32000 13876 32056
rect 13169 31998 13876 32000
rect 13169 31995 13235 31998
rect -300 31922 160 31952
rect 749 31922 815 31925
rect -300 31920 815 31922
rect -300 31864 754 31920
rect 810 31864 815 31920
rect -300 31862 815 31864
rect -300 31832 160 31862
rect 749 31859 815 31862
rect 1945 31922 2011 31925
rect 2262 31922 2268 31924
rect 1945 31920 2268 31922
rect 1945 31864 1950 31920
rect 2006 31864 2268 31920
rect 1945 31862 2268 31864
rect 1945 31859 2011 31862
rect 2262 31860 2268 31862
rect 2332 31860 2338 31924
rect 2589 31922 2655 31925
rect 4102 31922 4108 31924
rect 2589 31920 4108 31922
rect 2589 31864 2594 31920
rect 2650 31864 4108 31920
rect 2589 31862 4108 31864
rect 2589 31859 2655 31862
rect 4102 31860 4108 31862
rect 4172 31922 4178 31924
rect 4172 31862 4722 31922
rect 4172 31860 4178 31862
rect 1853 31784 1919 31789
rect 2129 31788 2195 31789
rect 2078 31786 2084 31788
rect 1853 31728 1858 31784
rect 1914 31728 1919 31784
rect 1853 31723 1919 31728
rect 2038 31726 2084 31786
rect 2148 31784 2195 31788
rect 2190 31728 2195 31784
rect 2078 31724 2084 31726
rect 2148 31724 2195 31728
rect 2129 31723 2195 31724
rect 4061 31786 4127 31789
rect 4286 31786 4292 31788
rect 4061 31784 4292 31786
rect 4061 31728 4066 31784
rect 4122 31728 4292 31784
rect 4061 31726 4292 31728
rect 4061 31723 4127 31726
rect 4286 31724 4292 31726
rect 4356 31724 4362 31788
rect 4662 31786 4722 31862
rect 9446 31862 13554 31922
rect 5717 31786 5783 31789
rect 7097 31786 7163 31789
rect 4662 31784 5783 31786
rect 4662 31728 5722 31784
rect 5778 31728 5783 31784
rect 4662 31726 5783 31728
rect 5717 31723 5783 31726
rect 5996 31784 7163 31786
rect 5996 31728 7102 31784
rect 7158 31728 7163 31784
rect 5996 31726 7163 31728
rect -300 31650 160 31680
rect 1485 31650 1551 31653
rect -300 31648 1551 31650
rect -300 31592 1490 31648
rect 1546 31592 1551 31648
rect -300 31590 1551 31592
rect 1856 31650 1916 31723
rect 1856 31590 5136 31650
rect -300 31560 160 31590
rect 1485 31587 1551 31590
rect 3233 31514 3299 31517
rect 3693 31514 3759 31517
rect 3233 31512 3759 31514
rect 3233 31456 3238 31512
rect 3294 31456 3698 31512
rect 3754 31456 3759 31512
rect 3233 31454 3759 31456
rect 3233 31451 3299 31454
rect 3693 31451 3759 31454
rect 4245 31514 4311 31517
rect 4654 31514 4660 31516
rect 4245 31512 4660 31514
rect 4245 31456 4250 31512
rect 4306 31456 4660 31512
rect 4245 31454 4660 31456
rect 4245 31451 4311 31454
rect 4654 31452 4660 31454
rect 4724 31452 4730 31516
rect -300 31378 160 31408
rect 3785 31378 3851 31381
rect -300 31376 3851 31378
rect -300 31320 3790 31376
rect 3846 31320 3851 31376
rect -300 31318 3851 31320
rect 5076 31378 5136 31590
rect 5257 31514 5323 31517
rect 5996 31514 6056 31726
rect 7097 31723 7163 31726
rect 8109 31788 8175 31789
rect 8109 31784 8156 31788
rect 8220 31786 8226 31788
rect 8477 31786 8543 31789
rect 9446 31786 9506 31862
rect 8109 31728 8114 31784
rect 8109 31724 8156 31728
rect 8220 31726 8266 31786
rect 8477 31784 9506 31786
rect 8477 31728 8482 31784
rect 8538 31728 9506 31784
rect 8477 31726 9506 31728
rect 9949 31786 10015 31789
rect 13494 31786 13554 31862
rect 13670 31860 13676 31924
rect 13740 31922 13746 31924
rect 13905 31922 13971 31925
rect 20069 31922 20135 31925
rect 13740 31920 13971 31922
rect 13740 31864 13910 31920
rect 13966 31864 13971 31920
rect 13740 31862 13971 31864
rect 13740 31860 13746 31862
rect 13905 31859 13971 31862
rect 14598 31920 20135 31922
rect 14598 31864 20074 31920
rect 20130 31864 20135 31920
rect 14598 31862 20135 31864
rect 14598 31786 14658 31862
rect 20069 31859 20135 31862
rect 20437 31922 20503 31925
rect 21541 31922 21607 31925
rect 20437 31920 21607 31922
rect 20437 31864 20442 31920
rect 20498 31864 21546 31920
rect 21602 31864 21607 31920
rect 20437 31862 21607 31864
rect 20437 31859 20503 31862
rect 21541 31859 21607 31862
rect 9949 31784 12450 31786
rect 9949 31728 9954 31784
rect 10010 31728 12450 31784
rect 9949 31726 12450 31728
rect 13494 31726 14658 31786
rect 14825 31786 14891 31789
rect 14958 31786 14964 31788
rect 14825 31784 14964 31786
rect 14825 31728 14830 31784
rect 14886 31728 14964 31784
rect 14825 31726 14964 31728
rect 8220 31724 8226 31726
rect 8109 31723 8175 31724
rect 8477 31723 8543 31726
rect 9949 31723 10015 31726
rect 12390 31650 12450 31726
rect 14825 31723 14891 31726
rect 14958 31724 14964 31726
rect 15028 31724 15034 31788
rect 15326 31724 15332 31788
rect 15396 31786 15402 31788
rect 15396 31724 15440 31786
rect 15380 31653 15440 31724
rect 12893 31650 12959 31653
rect 12390 31648 12959 31650
rect 12390 31592 12898 31648
rect 12954 31592 12959 31648
rect 12390 31590 12959 31592
rect 12893 31587 12959 31590
rect 15377 31648 15443 31653
rect 15377 31592 15382 31648
rect 15438 31592 15443 31648
rect 15377 31587 15443 31592
rect 22185 31650 22251 31653
rect 22840 31650 23300 31680
rect 22185 31648 23300 31650
rect 22185 31592 22190 31648
rect 22246 31592 23300 31648
rect 22185 31590 23300 31592
rect 22185 31587 22251 31590
rect 6144 31584 6460 31585
rect 6144 31520 6150 31584
rect 6214 31520 6230 31584
rect 6294 31520 6310 31584
rect 6374 31520 6390 31584
rect 6454 31520 6460 31584
rect 6144 31519 6460 31520
rect 11342 31584 11658 31585
rect 11342 31520 11348 31584
rect 11412 31520 11428 31584
rect 11492 31520 11508 31584
rect 11572 31520 11588 31584
rect 11652 31520 11658 31584
rect 11342 31519 11658 31520
rect 16540 31584 16856 31585
rect 16540 31520 16546 31584
rect 16610 31520 16626 31584
rect 16690 31520 16706 31584
rect 16770 31520 16786 31584
rect 16850 31520 16856 31584
rect 16540 31519 16856 31520
rect 21738 31584 22054 31585
rect 21738 31520 21744 31584
rect 21808 31520 21824 31584
rect 21888 31520 21904 31584
rect 21968 31520 21984 31584
rect 22048 31520 22054 31584
rect 22840 31560 23300 31590
rect 21738 31519 22054 31520
rect 5257 31512 6056 31514
rect 5257 31456 5262 31512
rect 5318 31456 6056 31512
rect 5257 31454 6056 31456
rect 13077 31514 13143 31517
rect 13077 31512 15026 31514
rect 13077 31456 13082 31512
rect 13138 31456 15026 31512
rect 13077 31454 15026 31456
rect 5257 31451 5323 31454
rect 13077 31451 13143 31454
rect 5076 31318 5504 31378
rect -300 31288 160 31318
rect 3785 31315 3851 31318
rect 1485 31244 1551 31245
rect 1485 31242 1532 31244
rect 1440 31240 1532 31242
rect 1596 31242 1602 31244
rect 2405 31242 2471 31245
rect 1596 31240 2471 31242
rect 1440 31184 1490 31240
rect 1596 31184 2410 31240
rect 2466 31184 2471 31240
rect 1440 31182 1532 31184
rect 1485 31180 1532 31182
rect 1596 31182 2471 31184
rect 1596 31180 1602 31182
rect 1485 31179 1551 31180
rect 2405 31179 2471 31182
rect 2589 31242 2655 31245
rect 5444 31242 5504 31318
rect 5574 31316 5580 31380
rect 5644 31378 5650 31380
rect 8518 31378 8524 31380
rect 5644 31318 8524 31378
rect 5644 31316 5650 31318
rect 8518 31316 8524 31318
rect 8588 31316 8594 31380
rect 11697 31378 11763 31381
rect 13629 31378 13695 31381
rect 11697 31376 13695 31378
rect 11697 31320 11702 31376
rect 11758 31320 13634 31376
rect 13690 31320 13695 31376
rect 11697 31318 13695 31320
rect 14966 31378 15026 31454
rect 19977 31378 20043 31381
rect 14966 31376 20043 31378
rect 14966 31320 19982 31376
rect 20038 31320 20043 31376
rect 14966 31318 20043 31320
rect 11697 31315 11763 31318
rect 13629 31315 13695 31318
rect 19977 31315 20043 31318
rect 6361 31242 6427 31245
rect 7782 31242 7788 31244
rect 2589 31240 5090 31242
rect 2589 31184 2594 31240
rect 2650 31184 5090 31240
rect 2589 31182 5090 31184
rect 5444 31240 7788 31242
rect 5444 31184 6366 31240
rect 6422 31184 7788 31240
rect 5444 31182 7788 31184
rect 2589 31179 2655 31182
rect -300 31106 160 31136
rect 2681 31106 2747 31109
rect -300 31104 2747 31106
rect -300 31048 2686 31104
rect 2742 31048 2747 31104
rect -300 31046 2747 31048
rect 5030 31106 5090 31182
rect 6361 31179 6427 31182
rect 7782 31180 7788 31182
rect 7852 31242 7858 31244
rect 8477 31242 8543 31245
rect 7852 31240 8543 31242
rect 7852 31184 8482 31240
rect 8538 31184 8543 31240
rect 7852 31182 8543 31184
rect 7852 31180 7858 31182
rect 8477 31179 8543 31182
rect 9765 31242 9831 31245
rect 9765 31240 19626 31242
rect 9765 31184 9770 31240
rect 9826 31184 19626 31240
rect 9765 31182 19626 31184
rect 9765 31179 9831 31182
rect 5165 31106 5231 31109
rect 5030 31104 5231 31106
rect 5030 31048 5170 31104
rect 5226 31048 5231 31104
rect 5030 31046 5231 31048
rect -300 31016 160 31046
rect 2681 31043 2747 31046
rect 5165 31043 5231 31046
rect 5758 31044 5764 31108
rect 5828 31106 5834 31108
rect 7557 31106 7623 31109
rect 5828 31104 7623 31106
rect 5828 31048 7562 31104
rect 7618 31048 7623 31104
rect 5828 31046 7623 31048
rect 5828 31044 5834 31046
rect 7557 31043 7623 31046
rect 9581 31106 9647 31109
rect 11789 31106 11855 31109
rect 9581 31104 11855 31106
rect 9581 31048 9586 31104
rect 9642 31048 11794 31104
rect 11850 31048 11855 31104
rect 9581 31046 11855 31048
rect 9581 31043 9647 31046
rect 11789 31043 11855 31046
rect 14641 31106 14707 31109
rect 15142 31106 15148 31108
rect 14641 31104 15148 31106
rect 14641 31048 14646 31104
rect 14702 31048 15148 31104
rect 14641 31046 15148 31048
rect 14641 31043 14707 31046
rect 15142 31044 15148 31046
rect 15212 31044 15218 31108
rect 3545 31040 3861 31041
rect 3545 30976 3551 31040
rect 3615 30976 3631 31040
rect 3695 30976 3711 31040
rect 3775 30976 3791 31040
rect 3855 30976 3861 31040
rect 3545 30975 3861 30976
rect 8743 31040 9059 31041
rect 8743 30976 8749 31040
rect 8813 30976 8829 31040
rect 8893 30976 8909 31040
rect 8973 30976 8989 31040
rect 9053 30976 9059 31040
rect 8743 30975 9059 30976
rect 13941 31040 14257 31041
rect 13941 30976 13947 31040
rect 14011 30976 14027 31040
rect 14091 30976 14107 31040
rect 14171 30976 14187 31040
rect 14251 30976 14257 31040
rect 13941 30975 14257 30976
rect 19139 31040 19455 31041
rect 19139 30976 19145 31040
rect 19209 30976 19225 31040
rect 19289 30976 19305 31040
rect 19369 30976 19385 31040
rect 19449 30976 19455 31040
rect 19139 30975 19455 30976
rect 5349 30970 5415 30973
rect 7097 30970 7163 30973
rect 5349 30968 7163 30970
rect 5349 30912 5354 30968
rect 5410 30912 7102 30968
rect 7158 30912 7163 30968
rect 5349 30910 7163 30912
rect 5349 30907 5415 30910
rect 7097 30907 7163 30910
rect 10409 30970 10475 30973
rect 10409 30968 12634 30970
rect 10409 30912 10414 30968
rect 10470 30912 12634 30968
rect 10409 30910 12634 30912
rect 10409 30907 10475 30910
rect -300 30834 160 30864
rect 4061 30834 4127 30837
rect -300 30832 4127 30834
rect -300 30776 4066 30832
rect 4122 30776 4127 30832
rect -300 30774 4127 30776
rect -300 30744 160 30774
rect 4061 30771 4127 30774
rect 5165 30834 5231 30837
rect 6085 30834 6151 30837
rect 5165 30832 6151 30834
rect 5165 30776 5170 30832
rect 5226 30776 6090 30832
rect 6146 30776 6151 30832
rect 5165 30774 6151 30776
rect 5165 30771 5231 30774
rect 6085 30771 6151 30774
rect 9622 30772 9628 30836
rect 9692 30834 9698 30836
rect 12433 30834 12499 30837
rect 9692 30832 12499 30834
rect 9692 30776 12438 30832
rect 12494 30776 12499 30832
rect 9692 30774 12499 30776
rect 12574 30834 12634 30910
rect 14774 30908 14780 30972
rect 14844 30970 14850 30972
rect 15193 30970 15259 30973
rect 14844 30968 15259 30970
rect 14844 30912 15198 30968
rect 15254 30912 15259 30968
rect 14844 30910 15259 30912
rect 19566 30970 19626 31182
rect 21449 31106 21515 31109
rect 22840 31106 23300 31136
rect 21449 31104 23300 31106
rect 21449 31048 21454 31104
rect 21510 31048 23300 31104
rect 21449 31046 23300 31048
rect 21449 31043 21515 31046
rect 22840 31016 23300 31046
rect 21265 30970 21331 30973
rect 19566 30968 21331 30970
rect 19566 30912 21270 30968
rect 21326 30912 21331 30968
rect 19566 30910 21331 30912
rect 14844 30908 14850 30910
rect 15193 30907 15259 30910
rect 21265 30907 21331 30910
rect 18873 30834 18939 30837
rect 12574 30832 18939 30834
rect 12574 30776 18878 30832
rect 18934 30776 18939 30832
rect 12574 30774 18939 30776
rect 9692 30772 9698 30774
rect 12433 30771 12499 30774
rect 18873 30771 18939 30774
rect 2078 30636 2084 30700
rect 2148 30698 2154 30700
rect 2589 30698 2655 30701
rect 2148 30696 2655 30698
rect 2148 30640 2594 30696
rect 2650 30640 2655 30696
rect 2148 30638 2655 30640
rect 2148 30636 2154 30638
rect 2589 30635 2655 30638
rect 2865 30698 2931 30701
rect 2865 30696 12956 30698
rect 2865 30640 2870 30696
rect 2926 30640 12956 30696
rect 2865 30638 12956 30640
rect 2865 30635 2931 30638
rect -300 30562 160 30592
rect 1669 30562 1735 30565
rect 5901 30564 5967 30565
rect 5901 30562 5948 30564
rect -300 30560 1735 30562
rect -300 30504 1674 30560
rect 1730 30504 1735 30560
rect -300 30502 1735 30504
rect 5856 30560 5948 30562
rect 5856 30504 5906 30560
rect 5856 30502 5948 30504
rect -300 30472 160 30502
rect 1669 30499 1735 30502
rect 5901 30500 5948 30502
rect 6012 30500 6018 30564
rect 7230 30500 7236 30564
rect 7300 30562 7306 30564
rect 9029 30562 9095 30565
rect 12249 30564 12315 30565
rect 12198 30562 12204 30564
rect 7300 30560 9095 30562
rect 7300 30504 9034 30560
rect 9090 30504 9095 30560
rect 7300 30502 9095 30504
rect 12158 30502 12204 30562
rect 12268 30560 12315 30564
rect 12310 30504 12315 30560
rect 7300 30500 7306 30502
rect 5901 30499 5967 30500
rect 9029 30499 9095 30502
rect 12198 30500 12204 30502
rect 12268 30500 12315 30504
rect 12896 30562 12956 30638
rect 13302 30636 13308 30700
rect 13372 30698 13378 30700
rect 14181 30698 14247 30701
rect 13372 30696 14247 30698
rect 13372 30640 14186 30696
rect 14242 30640 14247 30696
rect 13372 30638 14247 30640
rect 13372 30636 13378 30638
rect 14181 30635 14247 30638
rect 16297 30698 16363 30701
rect 19149 30698 19215 30701
rect 16297 30696 19215 30698
rect 16297 30640 16302 30696
rect 16358 30640 19154 30696
rect 19210 30640 19215 30696
rect 16297 30638 19215 30640
rect 16297 30635 16363 30638
rect 19149 30635 19215 30638
rect 13261 30562 13327 30565
rect 12896 30560 13327 30562
rect 12896 30504 13266 30560
rect 13322 30504 13327 30560
rect 12896 30502 13327 30504
rect 12249 30499 12315 30500
rect 13261 30499 13327 30502
rect 22277 30562 22343 30565
rect 22840 30562 23300 30592
rect 22277 30560 23300 30562
rect 22277 30504 22282 30560
rect 22338 30504 23300 30560
rect 22277 30502 23300 30504
rect 22277 30499 22343 30502
rect 6144 30496 6460 30497
rect 6144 30432 6150 30496
rect 6214 30432 6230 30496
rect 6294 30432 6310 30496
rect 6374 30432 6390 30496
rect 6454 30432 6460 30496
rect 6144 30431 6460 30432
rect 11342 30496 11658 30497
rect 11342 30432 11348 30496
rect 11412 30432 11428 30496
rect 11492 30432 11508 30496
rect 11572 30432 11588 30496
rect 11652 30432 11658 30496
rect 11342 30431 11658 30432
rect 16540 30496 16856 30497
rect 16540 30432 16546 30496
rect 16610 30432 16626 30496
rect 16690 30432 16706 30496
rect 16770 30432 16786 30496
rect 16850 30432 16856 30496
rect 16540 30431 16856 30432
rect 21738 30496 22054 30497
rect 21738 30432 21744 30496
rect 21808 30432 21824 30496
rect 21888 30432 21904 30496
rect 21968 30432 21984 30496
rect 22048 30432 22054 30496
rect 22840 30472 23300 30502
rect 21738 30431 22054 30432
rect 1393 30426 1459 30429
rect 1350 30424 1459 30426
rect 1350 30368 1398 30424
rect 1454 30368 1459 30424
rect 1350 30363 1459 30368
rect 9806 30364 9812 30428
rect 9876 30426 9882 30428
rect 10961 30426 11027 30429
rect 9876 30424 11027 30426
rect 9876 30368 10966 30424
rect 11022 30368 11027 30424
rect 9876 30366 11027 30368
rect 9876 30364 9882 30366
rect 10961 30363 11027 30366
rect 20529 30426 20595 30429
rect 20846 30426 20852 30428
rect 20529 30424 20852 30426
rect 20529 30368 20534 30424
rect 20590 30368 20852 30424
rect 20529 30366 20852 30368
rect 20529 30363 20595 30366
rect 20846 30364 20852 30366
rect 20916 30364 20922 30428
rect -300 30290 160 30320
rect 1350 30290 1410 30363
rect -300 30230 1410 30290
rect -300 30200 160 30230
rect 3182 30228 3188 30292
rect 3252 30290 3258 30292
rect 3601 30290 3667 30293
rect 3252 30288 3667 30290
rect 3252 30232 3606 30288
rect 3662 30232 3667 30288
rect 3252 30230 3667 30232
rect 3252 30228 3258 30230
rect 3601 30227 3667 30230
rect 3877 30290 3943 30293
rect 6085 30290 6151 30293
rect 3877 30288 6151 30290
rect 3877 30232 3882 30288
rect 3938 30232 6090 30288
rect 6146 30232 6151 30288
rect 3877 30230 6151 30232
rect 3877 30227 3943 30230
rect 6085 30227 6151 30230
rect 7189 30290 7255 30293
rect 9857 30290 9923 30293
rect 7189 30288 9923 30290
rect 7189 30232 7194 30288
rect 7250 30232 9862 30288
rect 9918 30232 9923 30288
rect 7189 30230 9923 30232
rect 7189 30227 7255 30230
rect 9857 30227 9923 30230
rect 11605 30290 11671 30293
rect 13261 30290 13327 30293
rect 11605 30288 13327 30290
rect 11605 30232 11610 30288
rect 11666 30232 13266 30288
rect 13322 30232 13327 30288
rect 11605 30230 13327 30232
rect 11605 30227 11671 30230
rect 13261 30227 13327 30230
rect 14641 30290 14707 30293
rect 20253 30290 20319 30293
rect 20529 30290 20595 30293
rect 14641 30288 20595 30290
rect 14641 30232 14646 30288
rect 14702 30232 20258 30288
rect 20314 30232 20534 30288
rect 20590 30232 20595 30288
rect 14641 30230 20595 30232
rect 14641 30227 14707 30230
rect 20253 30227 20319 30230
rect 20529 30227 20595 30230
rect 2497 30154 2563 30157
rect 5165 30156 5231 30157
rect 5165 30154 5212 30156
rect 2497 30152 4170 30154
rect 2497 30096 2502 30152
rect 2558 30096 4170 30152
rect 2497 30094 4170 30096
rect 5120 30152 5212 30154
rect 5120 30096 5170 30152
rect 5120 30094 5212 30096
rect 2497 30091 2563 30094
rect -300 30018 160 30048
rect 749 30018 815 30021
rect -300 30016 815 30018
rect -300 29960 754 30016
rect 810 29960 815 30016
rect -300 29958 815 29960
rect -300 29928 160 29958
rect 749 29955 815 29958
rect 3545 29952 3861 29953
rect 3545 29888 3551 29952
rect 3615 29888 3631 29952
rect 3695 29888 3711 29952
rect 3775 29888 3791 29952
rect 3855 29888 3861 29952
rect 3545 29887 3861 29888
rect 1485 29882 1551 29885
rect 3233 29882 3299 29885
rect 4110 29884 4170 30094
rect 5165 30092 5212 30094
rect 5276 30092 5282 30156
rect 5349 30154 5415 30157
rect 6729 30154 6795 30157
rect 5349 30152 6795 30154
rect 5349 30096 5354 30152
rect 5410 30096 6734 30152
rect 6790 30096 6795 30152
rect 5349 30094 6795 30096
rect 5165 30091 5231 30092
rect 5349 30091 5415 30094
rect 6729 30091 6795 30094
rect 10910 30092 10916 30156
rect 10980 30154 10986 30156
rect 20662 30154 20668 30156
rect 10980 30094 20668 30154
rect 10980 30092 10986 30094
rect 20662 30092 20668 30094
rect 20732 30092 20738 30156
rect 4245 30018 4311 30021
rect 7557 30018 7623 30021
rect 15929 30020 15995 30021
rect 4245 30016 7623 30018
rect 4245 29960 4250 30016
rect 4306 29960 7562 30016
rect 7618 29960 7623 30016
rect 4245 29958 7623 29960
rect 4245 29955 4311 29958
rect 7557 29955 7623 29958
rect 15878 29956 15884 30020
rect 15948 30018 15995 30020
rect 21449 30018 21515 30021
rect 22840 30018 23300 30048
rect 15948 30016 16040 30018
rect 15990 29960 16040 30016
rect 15948 29958 16040 29960
rect 21449 30016 23300 30018
rect 21449 29960 21454 30016
rect 21510 29960 23300 30016
rect 21449 29958 23300 29960
rect 15948 29956 15995 29958
rect 15929 29955 15995 29956
rect 21449 29955 21515 29958
rect 8743 29952 9059 29953
rect 8743 29888 8749 29952
rect 8813 29888 8829 29952
rect 8893 29888 8909 29952
rect 8973 29888 8989 29952
rect 9053 29888 9059 29952
rect 8743 29887 9059 29888
rect 13941 29952 14257 29953
rect 13941 29888 13947 29952
rect 14011 29888 14027 29952
rect 14091 29888 14107 29952
rect 14171 29888 14187 29952
rect 14251 29888 14257 29952
rect 13941 29887 14257 29888
rect 19139 29952 19455 29953
rect 19139 29888 19145 29952
rect 19209 29888 19225 29952
rect 19289 29888 19305 29952
rect 19369 29888 19385 29952
rect 19449 29888 19455 29952
rect 22840 29928 23300 29958
rect 19139 29887 19455 29888
rect 1485 29880 3299 29882
rect 1485 29824 1490 29880
rect 1546 29824 3238 29880
rect 3294 29824 3299 29880
rect 1485 29822 3299 29824
rect 1485 29819 1551 29822
rect 3233 29819 3299 29822
rect 4102 29820 4108 29884
rect 4172 29820 4178 29884
rect 6361 29882 6427 29885
rect 7005 29882 7071 29885
rect 6361 29880 7071 29882
rect 6361 29824 6366 29880
rect 6422 29824 7010 29880
rect 7066 29824 7071 29880
rect 6361 29822 7071 29824
rect 6361 29819 6427 29822
rect 7005 29819 7071 29822
rect 11329 29882 11395 29885
rect 12249 29882 12315 29885
rect 11329 29880 12315 29882
rect 11329 29824 11334 29880
rect 11390 29824 12254 29880
rect 12310 29824 12315 29880
rect 11329 29822 12315 29824
rect 11329 29819 11395 29822
rect 12249 29819 12315 29822
rect -300 29746 160 29776
rect 2773 29746 2839 29749
rect -300 29744 2839 29746
rect -300 29688 2778 29744
rect 2834 29688 2839 29744
rect -300 29686 2839 29688
rect -300 29656 160 29686
rect 2773 29683 2839 29686
rect 3366 29684 3372 29748
rect 3436 29746 3442 29748
rect 13905 29746 13971 29749
rect 3436 29744 13971 29746
rect 3436 29688 13910 29744
rect 13966 29688 13971 29744
rect 3436 29686 13971 29688
rect 3436 29684 3442 29686
rect 13905 29683 13971 29686
rect 289 29610 355 29613
rect 10777 29610 10843 29613
rect 289 29608 10843 29610
rect 289 29552 294 29608
rect 350 29552 10782 29608
rect 10838 29552 10843 29608
rect 289 29550 10843 29552
rect 289 29547 355 29550
rect 10777 29547 10843 29550
rect 13629 29610 13695 29613
rect 15193 29610 15259 29613
rect 13629 29608 15259 29610
rect 13629 29552 13634 29608
rect 13690 29552 15198 29608
rect 15254 29552 15259 29608
rect 13629 29550 15259 29552
rect 13629 29547 13695 29550
rect 15193 29547 15259 29550
rect -300 29474 160 29504
rect 3509 29474 3575 29477
rect 5993 29474 6059 29477
rect -300 29472 3575 29474
rect -300 29416 3514 29472
rect 3570 29416 3575 29472
rect -300 29414 3575 29416
rect -300 29384 160 29414
rect 3509 29411 3575 29414
rect 4478 29472 6059 29474
rect 4478 29416 5998 29472
rect 6054 29416 6059 29472
rect 4478 29414 6059 29416
rect 1945 29338 2011 29341
rect 2221 29338 2287 29341
rect 4478 29338 4538 29414
rect 5993 29411 6059 29414
rect 9438 29412 9444 29476
rect 9508 29412 9514 29476
rect 11789 29474 11855 29477
rect 12341 29474 12407 29477
rect 22185 29474 22251 29477
rect 22840 29474 23300 29504
rect 11789 29472 12407 29474
rect 11789 29416 11794 29472
rect 11850 29416 12346 29472
rect 12402 29416 12407 29472
rect 11789 29414 12407 29416
rect 6144 29408 6460 29409
rect 6144 29344 6150 29408
rect 6214 29344 6230 29408
rect 6294 29344 6310 29408
rect 6374 29344 6390 29408
rect 6454 29344 6460 29408
rect 6144 29343 6460 29344
rect 1945 29336 2287 29338
rect 1945 29280 1950 29336
rect 2006 29280 2226 29336
rect 2282 29280 2287 29336
rect 1945 29278 2287 29280
rect 1945 29275 2011 29278
rect 2221 29275 2287 29278
rect 2730 29278 4538 29338
rect 4613 29338 4679 29341
rect 5022 29338 5028 29340
rect 4613 29336 5028 29338
rect 4613 29280 4618 29336
rect 4674 29280 5028 29336
rect 4613 29278 5028 29280
rect -300 29202 160 29232
rect 1485 29202 1551 29205
rect -300 29200 1551 29202
rect -300 29144 1490 29200
rect 1546 29144 1551 29200
rect -300 29142 1551 29144
rect -300 29112 160 29142
rect 1485 29139 1551 29142
rect 1669 29202 1735 29205
rect 2730 29202 2790 29278
rect 4613 29275 4679 29278
rect 5022 29276 5028 29278
rect 5092 29276 5098 29340
rect 3049 29204 3115 29205
rect 2998 29202 3004 29204
rect 1669 29200 2790 29202
rect 1669 29144 1674 29200
rect 1730 29144 2790 29200
rect 1669 29142 2790 29144
rect 2958 29142 3004 29202
rect 3068 29200 3115 29204
rect 9446 29202 9506 29412
rect 11789 29411 11855 29414
rect 12341 29411 12407 29414
rect 12528 29414 13922 29474
rect 11342 29408 11658 29409
rect 11342 29344 11348 29408
rect 11412 29344 11428 29408
rect 11492 29344 11508 29408
rect 11572 29344 11588 29408
rect 11652 29344 11658 29408
rect 11342 29343 11658 29344
rect 11094 29276 11100 29340
rect 11164 29338 11170 29340
rect 11164 29276 11208 29338
rect 3110 29144 3115 29200
rect 1669 29139 1735 29142
rect 2998 29140 3004 29142
rect 3068 29140 3115 29144
rect 3049 29139 3115 29140
rect 4662 29142 9506 29202
rect 11148 29202 11208 29276
rect 11697 29202 11763 29205
rect 11148 29200 11763 29202
rect 11148 29144 11702 29200
rect 11758 29144 11763 29200
rect 11148 29142 11763 29144
rect 289 29066 355 29069
rect 4662 29066 4722 29142
rect 11697 29139 11763 29142
rect 289 29064 4722 29066
rect 289 29008 294 29064
rect 350 29008 4722 29064
rect 289 29006 4722 29008
rect 289 29003 355 29006
rect 4838 29004 4844 29068
rect 4908 29066 4914 29068
rect 5165 29066 5231 29069
rect 4908 29064 5231 29066
rect 4908 29008 5170 29064
rect 5226 29008 5231 29064
rect 4908 29006 5231 29008
rect 4908 29004 4914 29006
rect 5165 29003 5231 29006
rect 5993 29066 6059 29069
rect 7373 29066 7439 29069
rect 5993 29064 7439 29066
rect 5993 29008 5998 29064
rect 6054 29008 7378 29064
rect 7434 29008 7439 29064
rect 5993 29006 7439 29008
rect 5993 29003 6059 29006
rect 7373 29003 7439 29006
rect 7557 29066 7623 29069
rect 10542 29066 10548 29068
rect 7557 29064 10548 29066
rect 7557 29008 7562 29064
rect 7618 29008 10548 29064
rect 7557 29006 10548 29008
rect 7557 29003 7623 29006
rect 10542 29004 10548 29006
rect 10612 29066 10618 29068
rect 12528 29066 12588 29414
rect 13721 29336 13787 29341
rect 13721 29280 13726 29336
rect 13782 29280 13787 29336
rect 13721 29275 13787 29280
rect 13862 29338 13922 29414
rect 22185 29472 23300 29474
rect 22185 29416 22190 29472
rect 22246 29416 23300 29472
rect 22185 29414 23300 29416
rect 22185 29411 22251 29414
rect 16540 29408 16856 29409
rect 16540 29344 16546 29408
rect 16610 29344 16626 29408
rect 16690 29344 16706 29408
rect 16770 29344 16786 29408
rect 16850 29344 16856 29408
rect 16540 29343 16856 29344
rect 21738 29408 22054 29409
rect 21738 29344 21744 29408
rect 21808 29344 21824 29408
rect 21888 29344 21904 29408
rect 21968 29344 21984 29408
rect 22048 29344 22054 29408
rect 22840 29384 23300 29414
rect 21738 29343 22054 29344
rect 15929 29338 15995 29341
rect 13862 29336 16314 29338
rect 13862 29280 15934 29336
rect 15990 29280 16314 29336
rect 13862 29278 16314 29280
rect 15929 29275 15995 29278
rect 10612 29006 12588 29066
rect 10612 29004 10618 29006
rect -300 28930 160 28960
rect 749 28930 815 28933
rect -300 28928 815 28930
rect -300 28872 754 28928
rect 810 28872 815 28928
rect -300 28870 815 28872
rect -300 28840 160 28870
rect 749 28867 815 28870
rect 4613 28930 4679 28933
rect 8569 28930 8635 28933
rect 4613 28928 8635 28930
rect 4613 28872 4618 28928
rect 4674 28872 8574 28928
rect 8630 28872 8635 28928
rect 4613 28870 8635 28872
rect 4613 28867 4679 28870
rect 8569 28867 8635 28870
rect 9949 28930 10015 28933
rect 10409 28930 10475 28933
rect 13261 28930 13327 28933
rect 9949 28928 10475 28930
rect 9949 28872 9954 28928
rect 10010 28872 10414 28928
rect 10470 28872 10475 28928
rect 9949 28870 10475 28872
rect 9949 28867 10015 28870
rect 10409 28867 10475 28870
rect 10918 28928 13327 28930
rect 10918 28872 13266 28928
rect 13322 28872 13327 28928
rect 10918 28870 13327 28872
rect 3545 28864 3861 28865
rect 3545 28800 3551 28864
rect 3615 28800 3631 28864
rect 3695 28800 3711 28864
rect 3775 28800 3791 28864
rect 3855 28800 3861 28864
rect 3545 28799 3861 28800
rect 8743 28864 9059 28865
rect 8743 28800 8749 28864
rect 8813 28800 8829 28864
rect 8893 28800 8909 28864
rect 8973 28800 8989 28864
rect 9053 28800 9059 28864
rect 8743 28799 9059 28800
rect 5942 28732 5948 28796
rect 6012 28794 6018 28796
rect 6637 28794 6703 28797
rect 6012 28792 6703 28794
rect 6012 28736 6642 28792
rect 6698 28736 6703 28792
rect 6012 28734 6703 28736
rect 6012 28732 6018 28734
rect 6637 28731 6703 28734
rect 8017 28794 8083 28797
rect 8518 28794 8524 28796
rect 8017 28792 8524 28794
rect 8017 28736 8022 28792
rect 8078 28736 8524 28792
rect 8017 28734 8524 28736
rect 8017 28731 8083 28734
rect 8518 28732 8524 28734
rect 8588 28732 8594 28796
rect 9305 28794 9371 28797
rect 10918 28794 10978 28870
rect 13261 28867 13327 28870
rect 13724 28797 13784 29275
rect 16254 29202 16314 29278
rect 16254 29142 17970 29202
rect 16062 29004 16068 29068
rect 16132 29066 16138 29068
rect 17166 29066 17172 29068
rect 16132 29006 17172 29066
rect 16132 29004 16138 29006
rect 17166 29004 17172 29006
rect 17236 29004 17242 29068
rect 17033 28930 17099 28933
rect 17350 28930 17356 28932
rect 17033 28928 17356 28930
rect 17033 28872 17038 28928
rect 17094 28872 17356 28928
rect 17033 28870 17356 28872
rect 17033 28867 17099 28870
rect 17350 28868 17356 28870
rect 17420 28868 17426 28932
rect 17910 28930 17970 29142
rect 18822 29004 18828 29068
rect 18892 29066 18898 29068
rect 20069 29066 20135 29069
rect 18892 29064 20135 29066
rect 18892 29008 20074 29064
rect 20130 29008 20135 29064
rect 18892 29006 20135 29008
rect 18892 29004 18898 29006
rect 20069 29003 20135 29006
rect 18965 28930 19031 28933
rect 17910 28928 19031 28930
rect 17910 28872 18970 28928
rect 19026 28872 19031 28928
rect 17910 28870 19031 28872
rect 18965 28867 19031 28870
rect 21449 28930 21515 28933
rect 22840 28930 23300 28960
rect 21449 28928 23300 28930
rect 21449 28872 21454 28928
rect 21510 28872 23300 28928
rect 21449 28870 23300 28872
rect 21449 28867 21515 28870
rect 13941 28864 14257 28865
rect 13941 28800 13947 28864
rect 14011 28800 14027 28864
rect 14091 28800 14107 28864
rect 14171 28800 14187 28864
rect 14251 28800 14257 28864
rect 13941 28799 14257 28800
rect 19139 28864 19455 28865
rect 19139 28800 19145 28864
rect 19209 28800 19225 28864
rect 19289 28800 19305 28864
rect 19369 28800 19385 28864
rect 19449 28800 19455 28864
rect 22840 28840 23300 28870
rect 19139 28799 19455 28800
rect 9305 28792 10978 28794
rect 9305 28736 9310 28792
rect 9366 28736 10978 28792
rect 9305 28734 10978 28736
rect 11053 28794 11119 28797
rect 13486 28794 13492 28796
rect 11053 28792 13492 28794
rect 11053 28736 11058 28792
rect 11114 28736 13492 28792
rect 11053 28734 13492 28736
rect 9305 28731 9371 28734
rect 11053 28731 11119 28734
rect 13486 28732 13492 28734
rect 13556 28732 13562 28796
rect 13721 28792 13787 28797
rect 13721 28736 13726 28792
rect 13782 28736 13787 28792
rect 13721 28731 13787 28736
rect 14733 28794 14799 28797
rect 16205 28794 16271 28797
rect 14733 28792 16271 28794
rect 14733 28736 14738 28792
rect 14794 28736 16210 28792
rect 16266 28736 16271 28792
rect 14733 28734 16271 28736
rect 14733 28731 14799 28734
rect 16205 28731 16271 28734
rect -300 28658 160 28688
rect 3785 28658 3851 28661
rect -300 28656 3851 28658
rect -300 28600 3790 28656
rect 3846 28600 3851 28656
rect -300 28598 3851 28600
rect -300 28568 160 28598
rect 3785 28595 3851 28598
rect 4153 28658 4219 28661
rect 4286 28658 4292 28660
rect 4153 28656 4292 28658
rect 4153 28600 4158 28656
rect 4214 28600 4292 28656
rect 4153 28598 4292 28600
rect 4153 28595 4219 28598
rect 4286 28596 4292 28598
rect 4356 28596 4362 28660
rect 5257 28658 5323 28661
rect 6678 28658 6684 28660
rect 5257 28656 6684 28658
rect 5257 28600 5262 28656
rect 5318 28600 6684 28656
rect 5257 28598 6684 28600
rect 5257 28595 5323 28598
rect 6678 28596 6684 28598
rect 6748 28658 6754 28660
rect 7833 28658 7899 28661
rect 6748 28656 7899 28658
rect 6748 28600 7838 28656
rect 7894 28600 7899 28656
rect 6748 28598 7899 28600
rect 6748 28596 6754 28598
rect 7833 28595 7899 28598
rect 10174 28596 10180 28660
rect 10244 28658 10250 28660
rect 14590 28658 14596 28660
rect 10244 28598 14596 28658
rect 10244 28596 10250 28598
rect 14590 28596 14596 28598
rect 14660 28596 14666 28660
rect 2262 28460 2268 28524
rect 2332 28522 2338 28524
rect 6913 28522 6979 28525
rect 2332 28520 6979 28522
rect 2332 28464 6918 28520
rect 6974 28464 6979 28520
rect 2332 28462 6979 28464
rect 2332 28460 2338 28462
rect 6913 28459 6979 28462
rect 8477 28522 8543 28525
rect 13118 28522 13124 28524
rect 8477 28520 13124 28522
rect 8477 28464 8482 28520
rect 8538 28464 13124 28520
rect 8477 28462 13124 28464
rect 8477 28459 8543 28462
rect 13118 28460 13124 28462
rect 13188 28460 13194 28524
rect 13997 28522 14063 28525
rect 16205 28522 16271 28525
rect 13997 28520 16271 28522
rect 13997 28464 14002 28520
rect 14058 28464 16210 28520
rect 16266 28464 16271 28520
rect 13997 28462 16271 28464
rect 13997 28459 14063 28462
rect 16205 28459 16271 28462
rect -300 28386 160 28416
rect 1393 28386 1459 28389
rect -300 28384 1459 28386
rect -300 28328 1398 28384
rect 1454 28328 1459 28384
rect -300 28326 1459 28328
rect -300 28296 160 28326
rect 1393 28323 1459 28326
rect 2405 28386 2471 28389
rect 2630 28386 2636 28388
rect 2405 28384 2636 28386
rect 2405 28328 2410 28384
rect 2466 28328 2636 28384
rect 2405 28326 2636 28328
rect 2405 28323 2471 28326
rect 2630 28324 2636 28326
rect 2700 28324 2706 28388
rect 3601 28386 3667 28389
rect 5942 28386 5948 28388
rect 3601 28384 5948 28386
rect 3601 28328 3606 28384
rect 3662 28328 5948 28384
rect 3601 28326 5948 28328
rect 3601 28323 3667 28326
rect 5942 28324 5948 28326
rect 6012 28324 6018 28388
rect 8150 28324 8156 28388
rect 8220 28386 8226 28388
rect 9581 28386 9647 28389
rect 8220 28384 9647 28386
rect 8220 28328 9586 28384
rect 9642 28328 9647 28384
rect 8220 28326 9647 28328
rect 8220 28324 8226 28326
rect 9581 28323 9647 28326
rect 22185 28386 22251 28389
rect 22840 28386 23300 28416
rect 22185 28384 23300 28386
rect 22185 28328 22190 28384
rect 22246 28328 23300 28384
rect 22185 28326 23300 28328
rect 22185 28323 22251 28326
rect 6144 28320 6460 28321
rect 6144 28256 6150 28320
rect 6214 28256 6230 28320
rect 6294 28256 6310 28320
rect 6374 28256 6390 28320
rect 6454 28256 6460 28320
rect 6144 28255 6460 28256
rect 11342 28320 11658 28321
rect 11342 28256 11348 28320
rect 11412 28256 11428 28320
rect 11492 28256 11508 28320
rect 11572 28256 11588 28320
rect 11652 28256 11658 28320
rect 11342 28255 11658 28256
rect 16540 28320 16856 28321
rect 16540 28256 16546 28320
rect 16610 28256 16626 28320
rect 16690 28256 16706 28320
rect 16770 28256 16786 28320
rect 16850 28256 16856 28320
rect 16540 28255 16856 28256
rect 21738 28320 22054 28321
rect 21738 28256 21744 28320
rect 21808 28256 21824 28320
rect 21888 28256 21904 28320
rect 21968 28256 21984 28320
rect 22048 28256 22054 28320
rect 22840 28296 23300 28326
rect 21738 28255 22054 28256
rect 2589 28250 2655 28253
rect 8845 28250 8911 28253
rect 10869 28250 10935 28253
rect 2589 28248 5780 28250
rect 2589 28192 2594 28248
rect 2650 28192 5780 28248
rect 2589 28190 5780 28192
rect 2589 28187 2655 28190
rect -300 28114 160 28144
rect 2957 28114 3023 28117
rect -300 28112 3023 28114
rect -300 28056 2962 28112
rect 3018 28056 3023 28112
rect -300 28054 3023 28056
rect -300 28024 160 28054
rect 2957 28051 3023 28054
rect 3141 28114 3207 28117
rect 5533 28114 5599 28117
rect 3141 28112 5599 28114
rect 3141 28056 3146 28112
rect 3202 28056 5538 28112
rect 5594 28056 5599 28112
rect 3141 28054 5599 28056
rect 5720 28114 5780 28190
rect 8845 28248 10935 28250
rect 8845 28192 8850 28248
rect 8906 28192 10874 28248
rect 10930 28192 10935 28248
rect 8845 28190 10935 28192
rect 8845 28187 8911 28190
rect 10869 28187 10935 28190
rect 8017 28114 8083 28117
rect 5720 28112 8083 28114
rect 5720 28056 8022 28112
rect 8078 28056 8083 28112
rect 5720 28054 8083 28056
rect 3141 28051 3207 28054
rect 5533 28051 5599 28054
rect 8017 28051 8083 28054
rect 8293 28114 8359 28117
rect 12801 28114 12867 28117
rect 8293 28112 12867 28114
rect 8293 28056 8298 28112
rect 8354 28056 12806 28112
rect 12862 28056 12867 28112
rect 8293 28054 12867 28056
rect 8293 28051 8359 28054
rect 12801 28051 12867 28054
rect 1669 27978 1735 27981
rect 4245 27978 4311 27981
rect 4889 27978 4955 27981
rect 1669 27976 4170 27978
rect 1669 27920 1674 27976
rect 1730 27920 4170 27976
rect 1669 27918 4170 27920
rect 1669 27915 1735 27918
rect -300 27842 160 27872
rect 749 27842 815 27845
rect -300 27840 815 27842
rect -300 27784 754 27840
rect 810 27784 815 27840
rect -300 27782 815 27784
rect 4110 27842 4170 27918
rect 4245 27976 4955 27978
rect 4245 27920 4250 27976
rect 4306 27920 4894 27976
rect 4950 27920 4955 27976
rect 4245 27918 4955 27920
rect 4245 27915 4311 27918
rect 4889 27915 4955 27918
rect 5717 27978 5783 27981
rect 7741 27978 7807 27981
rect 5717 27976 7807 27978
rect 5717 27920 5722 27976
rect 5778 27920 7746 27976
rect 7802 27920 7807 27976
rect 5717 27918 7807 27920
rect 5717 27915 5783 27918
rect 7741 27915 7807 27918
rect 8937 27978 9003 27981
rect 9489 27978 9555 27981
rect 8937 27976 9555 27978
rect 8937 27920 8942 27976
rect 8998 27920 9494 27976
rect 9550 27920 9555 27976
rect 8937 27918 9555 27920
rect 8937 27915 9003 27918
rect 9489 27915 9555 27918
rect 11605 27978 11671 27981
rect 14089 27978 14155 27981
rect 11605 27976 14155 27978
rect 11605 27920 11610 27976
rect 11666 27920 14094 27976
rect 14150 27920 14155 27976
rect 11605 27918 14155 27920
rect 11605 27915 11671 27918
rect 14089 27915 14155 27918
rect 14958 27916 14964 27980
rect 15028 27978 15034 27980
rect 17125 27978 17191 27981
rect 19609 27978 19675 27981
rect 15028 27976 17191 27978
rect 15028 27920 17130 27976
rect 17186 27920 17191 27976
rect 15028 27918 17191 27920
rect 15028 27916 15034 27918
rect 17125 27915 17191 27918
rect 17358 27976 19675 27978
rect 17358 27920 19614 27976
rect 19670 27920 19675 27976
rect 17358 27918 19675 27920
rect 7097 27842 7163 27845
rect 4110 27840 7163 27842
rect 4110 27784 7102 27840
rect 7158 27784 7163 27840
rect 4110 27782 7163 27784
rect -300 27752 160 27782
rect 749 27779 815 27782
rect 7097 27779 7163 27782
rect 14457 27842 14523 27845
rect 17358 27842 17418 27918
rect 19609 27915 19675 27918
rect 14457 27840 17418 27842
rect 14457 27784 14462 27840
rect 14518 27784 17418 27840
rect 14457 27782 17418 27784
rect 14457 27779 14523 27782
rect 17534 27780 17540 27844
rect 17604 27842 17610 27844
rect 17677 27842 17743 27845
rect 17604 27840 17743 27842
rect 17604 27784 17682 27840
rect 17738 27784 17743 27840
rect 17604 27782 17743 27784
rect 17604 27780 17610 27782
rect 17677 27779 17743 27782
rect 21081 27842 21147 27845
rect 22840 27842 23300 27872
rect 21081 27840 23300 27842
rect 21081 27784 21086 27840
rect 21142 27784 23300 27840
rect 21081 27782 23300 27784
rect 21081 27779 21147 27782
rect 3545 27776 3861 27777
rect 3545 27712 3551 27776
rect 3615 27712 3631 27776
rect 3695 27712 3711 27776
rect 3775 27712 3791 27776
rect 3855 27712 3861 27776
rect 3545 27711 3861 27712
rect 8743 27776 9059 27777
rect 8743 27712 8749 27776
rect 8813 27712 8829 27776
rect 8893 27712 8909 27776
rect 8973 27712 8989 27776
rect 9053 27712 9059 27776
rect 8743 27711 9059 27712
rect 13941 27776 14257 27777
rect 13941 27712 13947 27776
rect 14011 27712 14027 27776
rect 14091 27712 14107 27776
rect 14171 27712 14187 27776
rect 14251 27712 14257 27776
rect 13941 27711 14257 27712
rect 19139 27776 19455 27777
rect 19139 27712 19145 27776
rect 19209 27712 19225 27776
rect 19289 27712 19305 27776
rect 19369 27712 19385 27776
rect 19449 27712 19455 27776
rect 22840 27752 23300 27782
rect 19139 27711 19455 27712
rect 1209 27706 1275 27709
rect 5073 27708 5139 27709
rect 7281 27708 7347 27709
rect 5022 27706 5028 27708
rect 1209 27704 2790 27706
rect 1209 27648 1214 27704
rect 1270 27648 2790 27704
rect 1209 27646 2790 27648
rect 4982 27646 5028 27706
rect 5092 27704 5139 27708
rect 5134 27648 5139 27704
rect 1209 27643 1275 27646
rect -300 27570 160 27600
rect 1485 27570 1551 27573
rect -300 27568 1551 27570
rect -300 27512 1490 27568
rect 1546 27512 1551 27568
rect -300 27510 1551 27512
rect 2730 27570 2790 27646
rect 5022 27644 5028 27646
rect 5092 27644 5139 27648
rect 7230 27644 7236 27708
rect 7300 27706 7347 27708
rect 7649 27706 7715 27709
rect 7782 27706 7788 27708
rect 7300 27704 7392 27706
rect 7342 27648 7392 27704
rect 7300 27646 7392 27648
rect 7649 27704 7788 27706
rect 7649 27648 7654 27704
rect 7710 27648 7788 27704
rect 7649 27646 7788 27648
rect 7300 27644 7347 27646
rect 5073 27643 5139 27644
rect 7281 27643 7347 27644
rect 7649 27643 7715 27646
rect 7782 27644 7788 27646
rect 7852 27644 7858 27708
rect 14917 27706 14983 27709
rect 16062 27706 16068 27708
rect 14917 27704 16068 27706
rect 14917 27648 14922 27704
rect 14978 27648 16068 27704
rect 14917 27646 16068 27648
rect 14917 27643 14983 27646
rect 16062 27644 16068 27646
rect 16132 27644 16138 27708
rect 9121 27570 9187 27573
rect 2730 27568 9187 27570
rect 2730 27512 9126 27568
rect 9182 27512 9187 27568
rect 2730 27510 9187 27512
rect -300 27480 160 27510
rect 1485 27507 1551 27510
rect 9121 27507 9187 27510
rect 657 27434 723 27437
rect 2814 27434 2820 27436
rect 657 27432 2820 27434
rect 657 27376 662 27432
rect 718 27376 2820 27432
rect 657 27374 2820 27376
rect 657 27371 723 27374
rect 2814 27372 2820 27374
rect 2884 27372 2890 27436
rect 3918 27372 3924 27436
rect 3988 27434 3994 27436
rect 5073 27434 5139 27437
rect 3988 27432 5139 27434
rect 3988 27376 5078 27432
rect 5134 27376 5139 27432
rect 3988 27374 5139 27376
rect 3988 27372 3994 27374
rect 5073 27371 5139 27374
rect 5349 27434 5415 27437
rect 10041 27434 10107 27437
rect 5349 27432 10107 27434
rect 5349 27376 5354 27432
rect 5410 27376 10046 27432
rect 10102 27376 10107 27432
rect 5349 27374 10107 27376
rect 5349 27371 5415 27374
rect 10041 27371 10107 27374
rect 15469 27434 15535 27437
rect 18505 27434 18571 27437
rect 15469 27432 18571 27434
rect 15469 27376 15474 27432
rect 15530 27376 18510 27432
rect 18566 27376 18571 27432
rect 15469 27374 18571 27376
rect 15469 27371 15535 27374
rect 18505 27371 18571 27374
rect -300 27298 160 27328
rect 1301 27298 1367 27301
rect 3141 27300 3207 27301
rect -300 27296 1367 27298
rect -300 27240 1306 27296
rect 1362 27240 1367 27296
rect -300 27238 1367 27240
rect -300 27208 160 27238
rect 1301 27235 1367 27238
rect 1894 27236 1900 27300
rect 1964 27298 1970 27300
rect 1964 27238 2882 27298
rect 1964 27236 1970 27238
rect 1853 27162 1919 27165
rect 2078 27162 2084 27164
rect 1853 27160 2084 27162
rect 1853 27104 1858 27160
rect 1914 27104 2084 27160
rect 1853 27102 2084 27104
rect 1853 27099 1919 27102
rect 2078 27100 2084 27102
rect 2148 27100 2154 27164
rect 2681 27162 2747 27165
rect 2822 27162 2882 27238
rect 3141 27296 3188 27300
rect 3252 27298 3258 27300
rect 4061 27298 4127 27301
rect 4889 27298 4955 27301
rect 3141 27240 3146 27296
rect 3141 27236 3188 27240
rect 3252 27238 3298 27298
rect 4061 27296 4955 27298
rect 4061 27240 4066 27296
rect 4122 27240 4894 27296
rect 4950 27240 4955 27296
rect 4061 27238 4955 27240
rect 3252 27236 3258 27238
rect 3141 27235 3207 27236
rect 4061 27235 4127 27238
rect 4889 27235 4955 27238
rect 12157 27298 12223 27301
rect 12617 27298 12683 27301
rect 12157 27296 12683 27298
rect 12157 27240 12162 27296
rect 12218 27240 12622 27296
rect 12678 27240 12683 27296
rect 12157 27238 12683 27240
rect 12157 27235 12223 27238
rect 12617 27235 12683 27238
rect 22185 27298 22251 27301
rect 22840 27298 23300 27328
rect 22185 27296 23300 27298
rect 22185 27240 22190 27296
rect 22246 27240 23300 27296
rect 22185 27238 23300 27240
rect 22185 27235 22251 27238
rect 6144 27232 6460 27233
rect 6144 27168 6150 27232
rect 6214 27168 6230 27232
rect 6294 27168 6310 27232
rect 6374 27168 6390 27232
rect 6454 27168 6460 27232
rect 6144 27167 6460 27168
rect 11342 27232 11658 27233
rect 11342 27168 11348 27232
rect 11412 27168 11428 27232
rect 11492 27168 11508 27232
rect 11572 27168 11588 27232
rect 11652 27168 11658 27232
rect 11342 27167 11658 27168
rect 16540 27232 16856 27233
rect 16540 27168 16546 27232
rect 16610 27168 16626 27232
rect 16690 27168 16706 27232
rect 16770 27168 16786 27232
rect 16850 27168 16856 27232
rect 16540 27167 16856 27168
rect 21738 27232 22054 27233
rect 21738 27168 21744 27232
rect 21808 27168 21824 27232
rect 21888 27168 21904 27232
rect 21968 27168 21984 27232
rect 22048 27168 22054 27232
rect 22840 27208 23300 27238
rect 21738 27167 22054 27168
rect 3918 27162 3924 27164
rect 2681 27160 3924 27162
rect 2681 27104 2686 27160
rect 2742 27104 3924 27160
rect 2681 27102 3924 27104
rect 2681 27099 2747 27102
rect 3918 27100 3924 27102
rect 3988 27162 3994 27164
rect 4061 27162 4127 27165
rect 3988 27160 4127 27162
rect 3988 27104 4066 27160
rect 4122 27104 4127 27160
rect 3988 27102 4127 27104
rect 3988 27100 3994 27102
rect 4061 27099 4127 27102
rect 4337 27162 4403 27165
rect 8569 27164 8635 27165
rect 4470 27162 4476 27164
rect 4337 27160 4476 27162
rect 4337 27104 4342 27160
rect 4398 27104 4476 27160
rect 4337 27102 4476 27104
rect 4337 27099 4403 27102
rect 4470 27100 4476 27102
rect 4540 27100 4546 27164
rect 8518 27162 8524 27164
rect 8478 27102 8524 27162
rect 8588 27160 8635 27164
rect 8630 27104 8635 27160
rect 8518 27100 8524 27102
rect 8588 27100 8635 27104
rect 9438 27100 9444 27164
rect 9508 27162 9514 27164
rect 10133 27162 10199 27165
rect 10542 27162 10548 27164
rect 9508 27160 10548 27162
rect 9508 27104 10138 27160
rect 10194 27104 10548 27160
rect 9508 27102 10548 27104
rect 9508 27100 9514 27102
rect 8569 27099 8635 27100
rect 10133 27099 10199 27102
rect 10542 27100 10548 27102
rect 10612 27100 10618 27164
rect -300 27026 160 27056
rect 1301 27026 1367 27029
rect -300 27024 1367 27026
rect -300 26968 1306 27024
rect 1362 26968 1367 27024
rect -300 26966 1367 26968
rect -300 26936 160 26966
rect 1301 26963 1367 26966
rect 2957 27026 3023 27029
rect 5533 27026 5599 27029
rect 7373 27026 7439 27029
rect 2957 27024 7439 27026
rect 2957 26968 2962 27024
rect 3018 26968 5538 27024
rect 5594 26968 7378 27024
rect 7434 26968 7439 27024
rect 2957 26966 7439 26968
rect 2957 26963 3023 26966
rect 5533 26963 5599 26966
rect 7373 26963 7439 26966
rect 8518 26964 8524 27028
rect 8588 27026 8594 27028
rect 8661 27026 8727 27029
rect 18045 27026 18111 27029
rect 18873 27026 18939 27029
rect 8588 27024 18939 27026
rect 8588 26968 8666 27024
rect 8722 26968 18050 27024
rect 18106 26968 18878 27024
rect 18934 26968 18939 27024
rect 8588 26966 18939 26968
rect 8588 26964 8594 26966
rect 8661 26963 8727 26966
rect 18045 26963 18111 26966
rect 18873 26963 18939 26966
rect 21449 27024 21515 27029
rect 21449 26968 21454 27024
rect 21510 26968 21515 27024
rect 21449 26963 21515 26968
rect 1393 26890 1459 26893
rect 1526 26890 1532 26892
rect 1393 26888 1532 26890
rect 1393 26832 1398 26888
rect 1454 26832 1532 26888
rect 1393 26830 1532 26832
rect 1393 26827 1459 26830
rect 1526 26828 1532 26830
rect 1596 26828 1602 26892
rect 2497 26890 2563 26893
rect 8661 26890 8727 26893
rect 2497 26888 8727 26890
rect 2497 26832 2502 26888
rect 2558 26832 8666 26888
rect 8722 26832 8727 26888
rect 2497 26830 8727 26832
rect 2497 26827 2563 26830
rect 8661 26827 8727 26830
rect -300 26754 160 26784
rect 1209 26754 1275 26757
rect -300 26752 1275 26754
rect -300 26696 1214 26752
rect 1270 26696 1275 26752
rect -300 26694 1275 26696
rect -300 26664 160 26694
rect 1209 26691 1275 26694
rect 2957 26754 3023 26757
rect 3366 26754 3372 26756
rect 2957 26752 3372 26754
rect 2957 26696 2962 26752
rect 3018 26696 3372 26752
rect 2957 26694 3372 26696
rect 2957 26691 3023 26694
rect 3366 26692 3372 26694
rect 3436 26692 3442 26756
rect 6678 26692 6684 26756
rect 6748 26754 6754 26756
rect 6821 26754 6887 26757
rect 6748 26752 6887 26754
rect 6748 26696 6826 26752
rect 6882 26696 6887 26752
rect 6748 26694 6887 26696
rect 6748 26692 6754 26694
rect 6821 26691 6887 26694
rect 12382 26692 12388 26756
rect 12452 26754 12458 26756
rect 12985 26754 13051 26757
rect 12452 26752 13051 26754
rect 12452 26696 12990 26752
rect 13046 26696 13051 26752
rect 12452 26694 13051 26696
rect 21452 26754 21512 26963
rect 22840 26754 23300 26784
rect 21452 26694 23300 26754
rect 12452 26692 12458 26694
rect 12985 26691 13051 26694
rect 3545 26688 3861 26689
rect 3545 26624 3551 26688
rect 3615 26624 3631 26688
rect 3695 26624 3711 26688
rect 3775 26624 3791 26688
rect 3855 26624 3861 26688
rect 3545 26623 3861 26624
rect 8743 26688 9059 26689
rect 8743 26624 8749 26688
rect 8813 26624 8829 26688
rect 8893 26624 8909 26688
rect 8973 26624 8989 26688
rect 9053 26624 9059 26688
rect 8743 26623 9059 26624
rect 13941 26688 14257 26689
rect 13941 26624 13947 26688
rect 14011 26624 14027 26688
rect 14091 26624 14107 26688
rect 14171 26624 14187 26688
rect 14251 26624 14257 26688
rect 13941 26623 14257 26624
rect 19139 26688 19455 26689
rect 19139 26624 19145 26688
rect 19209 26624 19225 26688
rect 19289 26624 19305 26688
rect 19369 26624 19385 26688
rect 19449 26624 19455 26688
rect 22840 26664 23300 26694
rect 19139 26623 19455 26624
rect 1853 26618 1919 26621
rect 3325 26618 3391 26621
rect 1853 26616 3391 26618
rect 1853 26560 1858 26616
rect 1914 26560 3330 26616
rect 3386 26560 3391 26616
rect 1853 26558 3391 26560
rect 1853 26555 1919 26558
rect 3325 26555 3391 26558
rect 5257 26618 5323 26621
rect 7005 26618 7071 26621
rect 8109 26618 8175 26621
rect 5257 26616 8175 26618
rect 5257 26560 5262 26616
rect 5318 26560 7010 26616
rect 7066 26560 8114 26616
rect 8170 26560 8175 26616
rect 5257 26558 8175 26560
rect 5257 26555 5323 26558
rect 7005 26555 7071 26558
rect 8109 26555 8175 26558
rect -300 26482 160 26512
rect 1761 26482 1827 26485
rect 2037 26482 2103 26485
rect 2497 26484 2563 26485
rect -300 26480 1827 26482
rect -300 26424 1766 26480
rect 1822 26424 1827 26480
rect -300 26422 1827 26424
rect -300 26392 160 26422
rect 1761 26419 1827 26422
rect 1902 26480 2103 26482
rect 1902 26424 2042 26480
rect 2098 26424 2103 26480
rect 1902 26422 2103 26424
rect 1761 26346 1827 26349
rect 1902 26346 1962 26422
rect 2037 26419 2103 26422
rect 2446 26420 2452 26484
rect 2516 26482 2563 26484
rect 3325 26482 3391 26485
rect 14917 26482 14983 26485
rect 2516 26480 2608 26482
rect 2558 26424 2608 26480
rect 2516 26422 2608 26424
rect 3325 26480 14983 26482
rect 3325 26424 3330 26480
rect 3386 26424 14922 26480
rect 14978 26424 14983 26480
rect 3325 26422 14983 26424
rect 2516 26420 2563 26422
rect 2497 26419 2563 26420
rect 3325 26419 3391 26422
rect 14917 26419 14983 26422
rect 1761 26344 1962 26346
rect 1761 26288 1766 26344
rect 1822 26288 1962 26344
rect 1761 26286 1962 26288
rect 3509 26346 3575 26349
rect 6361 26346 6427 26349
rect 6821 26346 6887 26349
rect 3509 26344 6887 26346
rect 3509 26288 3514 26344
rect 3570 26288 6366 26344
rect 6422 26288 6826 26344
rect 6882 26288 6887 26344
rect 3509 26286 6887 26288
rect 1761 26283 1827 26286
rect 3509 26283 3575 26286
rect 6361 26283 6427 26286
rect 6821 26283 6887 26286
rect 7833 26346 7899 26349
rect 8201 26346 8267 26349
rect 10174 26346 10180 26348
rect 7833 26344 10180 26346
rect 7833 26288 7838 26344
rect 7894 26288 8206 26344
rect 8262 26288 10180 26344
rect 7833 26286 10180 26288
rect 7833 26283 7899 26286
rect 8201 26283 8267 26286
rect 10174 26284 10180 26286
rect 10244 26284 10250 26348
rect 10869 26346 10935 26349
rect 13445 26346 13511 26349
rect 10869 26344 13511 26346
rect 10869 26288 10874 26344
rect 10930 26288 13450 26344
rect 13506 26288 13511 26344
rect 10869 26286 13511 26288
rect 10869 26283 10935 26286
rect 13445 26283 13511 26286
rect 15929 26346 15995 26349
rect 19885 26346 19951 26349
rect 15929 26344 19951 26346
rect 15929 26288 15934 26344
rect 15990 26288 19890 26344
rect 19946 26288 19951 26344
rect 15929 26286 19951 26288
rect 15929 26283 15995 26286
rect 19885 26283 19951 26286
rect -300 26210 160 26240
rect 841 26210 907 26213
rect 1342 26210 1348 26212
rect -300 26150 720 26210
rect -300 26120 160 26150
rect 660 26074 720 26150
rect 841 26208 1348 26210
rect 841 26152 846 26208
rect 902 26152 1348 26208
rect 841 26150 1348 26152
rect 841 26147 907 26150
rect 1342 26148 1348 26150
rect 1412 26148 1418 26212
rect 1945 26210 2011 26213
rect 3325 26210 3391 26213
rect 1534 26208 2011 26210
rect 1534 26152 1950 26208
rect 2006 26152 2011 26208
rect 1534 26150 2011 26152
rect 1534 26074 1594 26150
rect 1945 26147 2011 26150
rect 2730 26208 3391 26210
rect 2730 26152 3330 26208
rect 3386 26152 3391 26208
rect 2730 26150 3391 26152
rect 660 26014 1594 26074
rect 1710 26012 1716 26076
rect 1780 26074 1786 26076
rect 2129 26074 2195 26077
rect 1780 26072 2195 26074
rect 1780 26016 2134 26072
rect 2190 26016 2195 26072
rect 1780 26014 2195 26016
rect 1780 26012 1786 26014
rect 2129 26011 2195 26014
rect -300 25938 160 25968
rect 2730 25938 2790 26150
rect 3325 26147 3391 26150
rect 5390 26148 5396 26212
rect 5460 26210 5466 26212
rect 5901 26210 5967 26213
rect 5460 26208 5967 26210
rect 5460 26152 5906 26208
rect 5962 26152 5967 26208
rect 5460 26150 5967 26152
rect 5460 26148 5466 26150
rect 5901 26147 5967 26150
rect 18086 26148 18092 26212
rect 18156 26210 18162 26212
rect 18229 26210 18295 26213
rect 18156 26208 18295 26210
rect 18156 26152 18234 26208
rect 18290 26152 18295 26208
rect 18156 26150 18295 26152
rect 18156 26148 18162 26150
rect 18229 26147 18295 26150
rect 22277 26210 22343 26213
rect 22840 26210 23300 26240
rect 22277 26208 23300 26210
rect 22277 26152 22282 26208
rect 22338 26152 23300 26208
rect 22277 26150 23300 26152
rect 22277 26147 22343 26150
rect 6144 26144 6460 26145
rect 6144 26080 6150 26144
rect 6214 26080 6230 26144
rect 6294 26080 6310 26144
rect 6374 26080 6390 26144
rect 6454 26080 6460 26144
rect 6144 26079 6460 26080
rect 11342 26144 11658 26145
rect 11342 26080 11348 26144
rect 11412 26080 11428 26144
rect 11492 26080 11508 26144
rect 11572 26080 11588 26144
rect 11652 26080 11658 26144
rect 11342 26079 11658 26080
rect 16540 26144 16856 26145
rect 16540 26080 16546 26144
rect 16610 26080 16626 26144
rect 16690 26080 16706 26144
rect 16770 26080 16786 26144
rect 16850 26080 16856 26144
rect 16540 26079 16856 26080
rect 21738 26144 22054 26145
rect 21738 26080 21744 26144
rect 21808 26080 21824 26144
rect 21888 26080 21904 26144
rect 21968 26080 21984 26144
rect 22048 26080 22054 26144
rect 22840 26120 23300 26150
rect 21738 26079 22054 26080
rect 7782 25938 7788 25940
rect -300 25878 2790 25938
rect 4340 25878 7788 25938
rect -300 25848 160 25878
rect 1710 25740 1716 25804
rect 1780 25802 1786 25804
rect 4340 25802 4400 25878
rect 7782 25876 7788 25878
rect 7852 25938 7858 25940
rect 9857 25938 9923 25941
rect 7852 25936 9923 25938
rect 7852 25880 9862 25936
rect 9918 25880 9923 25936
rect 7852 25878 9923 25880
rect 7852 25876 7858 25878
rect 9857 25875 9923 25878
rect 10777 25938 10843 25941
rect 12893 25938 12959 25941
rect 10777 25936 12959 25938
rect 10777 25880 10782 25936
rect 10838 25880 12898 25936
rect 12954 25880 12959 25936
rect 10777 25878 12959 25880
rect 10777 25875 10843 25878
rect 12893 25875 12959 25878
rect 1780 25742 4400 25802
rect 4521 25802 4587 25805
rect 15285 25802 15351 25805
rect 4521 25800 15351 25802
rect 4521 25744 4526 25800
rect 4582 25744 15290 25800
rect 15346 25744 15351 25800
rect 4521 25742 15351 25744
rect 1780 25740 1786 25742
rect 4521 25739 4587 25742
rect 15285 25739 15351 25742
rect -300 25666 160 25696
rect 3049 25666 3115 25669
rect 4521 25668 4587 25669
rect 4470 25666 4476 25668
rect -300 25664 3115 25666
rect -300 25608 3054 25664
rect 3110 25608 3115 25664
rect -300 25606 3115 25608
rect 4430 25606 4476 25666
rect 4540 25664 4587 25668
rect 4582 25608 4587 25664
rect -300 25576 160 25606
rect 3049 25603 3115 25606
rect 4470 25604 4476 25606
rect 4540 25604 4587 25608
rect 5758 25604 5764 25668
rect 5828 25666 5834 25668
rect 6729 25666 6795 25669
rect 5828 25664 6795 25666
rect 5828 25608 6734 25664
rect 6790 25608 6795 25664
rect 5828 25606 6795 25608
rect 5828 25604 5834 25606
rect 4521 25603 4587 25604
rect 6729 25603 6795 25606
rect 7046 25604 7052 25668
rect 7116 25666 7122 25668
rect 7741 25666 7807 25669
rect 7116 25664 7807 25666
rect 7116 25608 7746 25664
rect 7802 25608 7807 25664
rect 7116 25606 7807 25608
rect 7116 25604 7122 25606
rect 7741 25603 7807 25606
rect 21449 25666 21515 25669
rect 22840 25666 23300 25696
rect 21449 25664 23300 25666
rect 21449 25608 21454 25664
rect 21510 25608 23300 25664
rect 21449 25606 23300 25608
rect 21449 25603 21515 25606
rect 3545 25600 3861 25601
rect 3545 25536 3551 25600
rect 3615 25536 3631 25600
rect 3695 25536 3711 25600
rect 3775 25536 3791 25600
rect 3855 25536 3861 25600
rect 3545 25535 3861 25536
rect 8743 25600 9059 25601
rect 8743 25536 8749 25600
rect 8813 25536 8829 25600
rect 8893 25536 8909 25600
rect 8973 25536 8989 25600
rect 9053 25536 9059 25600
rect 8743 25535 9059 25536
rect 13941 25600 14257 25601
rect 13941 25536 13947 25600
rect 14011 25536 14027 25600
rect 14091 25536 14107 25600
rect 14171 25536 14187 25600
rect 14251 25536 14257 25600
rect 13941 25535 14257 25536
rect 19139 25600 19455 25601
rect 19139 25536 19145 25600
rect 19209 25536 19225 25600
rect 19289 25536 19305 25600
rect 19369 25536 19385 25600
rect 19449 25536 19455 25600
rect 22840 25576 23300 25606
rect 19139 25535 19455 25536
rect 2221 25530 2287 25533
rect 6637 25530 6703 25533
rect 6862 25530 6868 25532
rect 2221 25528 3066 25530
rect 2221 25472 2226 25528
rect 2282 25472 3066 25528
rect 2221 25470 3066 25472
rect 2221 25467 2287 25470
rect -300 25394 160 25424
rect 2773 25394 2839 25397
rect 3006 25396 3066 25470
rect 6637 25528 6868 25530
rect 6637 25472 6642 25528
rect 6698 25472 6868 25528
rect 6637 25470 6868 25472
rect 6637 25467 6703 25470
rect 6862 25468 6868 25470
rect 6932 25468 6938 25532
rect 7005 25530 7071 25533
rect 7005 25528 8540 25530
rect 7005 25472 7010 25528
rect 7066 25472 8540 25528
rect 7005 25470 8540 25472
rect 7005 25467 7071 25470
rect -300 25392 2839 25394
rect -300 25336 2778 25392
rect 2834 25336 2839 25392
rect -300 25334 2839 25336
rect -300 25304 160 25334
rect 2773 25331 2839 25334
rect 2998 25332 3004 25396
rect 3068 25332 3074 25396
rect 3601 25394 3667 25397
rect 8293 25394 8359 25397
rect 3601 25392 8359 25394
rect 3601 25336 3606 25392
rect 3662 25336 8298 25392
rect 8354 25336 8359 25392
rect 3601 25334 8359 25336
rect 8480 25394 8540 25470
rect 11881 25394 11947 25397
rect 8480 25392 11947 25394
rect 8480 25336 11886 25392
rect 11942 25336 11947 25392
rect 8480 25334 11947 25336
rect 3601 25331 3667 25334
rect 8293 25331 8359 25334
rect 11881 25331 11947 25334
rect 15929 25394 15995 25397
rect 18270 25394 18276 25396
rect 15929 25392 18276 25394
rect 15929 25336 15934 25392
rect 15990 25336 18276 25392
rect 15929 25334 18276 25336
rect 15929 25331 15995 25334
rect 18270 25332 18276 25334
rect 18340 25332 18346 25396
rect 3182 25196 3188 25260
rect 3252 25258 3258 25260
rect 5073 25258 5139 25261
rect 3252 25256 5139 25258
rect 3252 25200 5078 25256
rect 5134 25200 5139 25256
rect 3252 25198 5139 25200
rect 3252 25196 3258 25198
rect 5073 25195 5139 25198
rect 6545 25258 6611 25261
rect 13302 25258 13308 25260
rect 6545 25256 13308 25258
rect 6545 25200 6550 25256
rect 6606 25200 13308 25256
rect 6545 25198 13308 25200
rect 6545 25195 6611 25198
rect 13302 25196 13308 25198
rect 13372 25258 13378 25260
rect 13629 25258 13695 25261
rect 13372 25256 13695 25258
rect 13372 25200 13634 25256
rect 13690 25200 13695 25256
rect 13372 25198 13695 25200
rect 13372 25196 13378 25198
rect 13629 25195 13695 25198
rect -300 25122 160 25152
rect 1485 25122 1551 25125
rect -300 25120 1551 25122
rect -300 25064 1490 25120
rect 1546 25064 1551 25120
rect -300 25062 1551 25064
rect -300 25032 160 25062
rect 1485 25059 1551 25062
rect 2129 25122 2195 25125
rect 5993 25122 6059 25125
rect 2129 25120 6059 25122
rect 2129 25064 2134 25120
rect 2190 25064 5998 25120
rect 6054 25064 6059 25120
rect 2129 25062 6059 25064
rect 2129 25059 2195 25062
rect 5993 25059 6059 25062
rect 22277 25122 22343 25125
rect 22840 25122 23300 25152
rect 22277 25120 23300 25122
rect 22277 25064 22282 25120
rect 22338 25064 23300 25120
rect 22277 25062 23300 25064
rect 22277 25059 22343 25062
rect 6144 25056 6460 25057
rect 6144 24992 6150 25056
rect 6214 24992 6230 25056
rect 6294 24992 6310 25056
rect 6374 24992 6390 25056
rect 6454 24992 6460 25056
rect 6144 24991 6460 24992
rect 11342 25056 11658 25057
rect 11342 24992 11348 25056
rect 11412 24992 11428 25056
rect 11492 24992 11508 25056
rect 11572 24992 11588 25056
rect 11652 24992 11658 25056
rect 11342 24991 11658 24992
rect 16540 25056 16856 25057
rect 16540 24992 16546 25056
rect 16610 24992 16626 25056
rect 16690 24992 16706 25056
rect 16770 24992 16786 25056
rect 16850 24992 16856 25056
rect 16540 24991 16856 24992
rect 21738 25056 22054 25057
rect 21738 24992 21744 25056
rect 21808 24992 21824 25056
rect 21888 24992 21904 25056
rect 21968 24992 21984 25056
rect 22048 24992 22054 25056
rect 22840 25032 23300 25062
rect 21738 24991 22054 24992
rect 1485 24986 1551 24989
rect 2497 24986 2563 24989
rect 1485 24984 2563 24986
rect 1485 24928 1490 24984
rect 1546 24928 2502 24984
rect 2558 24928 2563 24984
rect 1485 24926 2563 24928
rect 1485 24923 1551 24926
rect 2497 24923 2563 24926
rect 15510 24924 15516 24988
rect 15580 24986 15586 24988
rect 15653 24986 15719 24989
rect 15580 24984 15719 24986
rect 15580 24928 15658 24984
rect 15714 24928 15719 24984
rect 15580 24926 15719 24928
rect 15580 24924 15586 24926
rect 15653 24923 15719 24926
rect -300 24850 160 24880
rect 841 24850 907 24853
rect -300 24848 907 24850
rect -300 24792 846 24848
rect 902 24792 907 24848
rect -300 24790 907 24792
rect -300 24760 160 24790
rect 841 24787 907 24790
rect 5165 24850 5231 24853
rect 9806 24850 9812 24852
rect 5165 24848 9812 24850
rect 5165 24792 5170 24848
rect 5226 24792 9812 24848
rect 5165 24790 9812 24792
rect 5165 24787 5231 24790
rect 9806 24788 9812 24790
rect 9876 24788 9882 24852
rect 11697 24850 11763 24853
rect 12014 24850 12020 24852
rect 11697 24848 12020 24850
rect 11697 24792 11702 24848
rect 11758 24792 12020 24848
rect 11697 24790 12020 24792
rect 11697 24787 11763 24790
rect 12014 24788 12020 24790
rect 12084 24788 12090 24852
rect 12198 24788 12204 24852
rect 12268 24850 12274 24852
rect 12525 24850 12591 24853
rect 12268 24848 12591 24850
rect 12268 24792 12530 24848
rect 12586 24792 12591 24848
rect 12268 24790 12591 24792
rect 12268 24788 12274 24790
rect 12525 24787 12591 24790
rect 16941 24850 17007 24853
rect 18638 24850 18644 24852
rect 16941 24848 18644 24850
rect 16941 24792 16946 24848
rect 17002 24792 18644 24848
rect 16941 24790 18644 24792
rect 16941 24787 17007 24790
rect 18638 24788 18644 24790
rect 18708 24788 18714 24852
rect 1853 24714 1919 24717
rect 1853 24712 3986 24714
rect 1853 24656 1858 24712
rect 1914 24656 3986 24712
rect 1853 24654 3986 24656
rect 1853 24651 1919 24654
rect -300 24578 160 24608
rect 3233 24578 3299 24581
rect -300 24576 3299 24578
rect -300 24520 3238 24576
rect 3294 24520 3299 24576
rect -300 24518 3299 24520
rect 3926 24578 3986 24654
rect 5206 24652 5212 24716
rect 5276 24714 5282 24716
rect 10593 24714 10659 24717
rect 12617 24714 12683 24717
rect 14641 24714 14707 24717
rect 14917 24716 14983 24717
rect 14774 24714 14780 24716
rect 5276 24654 9184 24714
rect 5276 24652 5282 24654
rect 4245 24578 4311 24581
rect 6085 24578 6151 24581
rect 3926 24576 6151 24578
rect 3926 24520 4250 24576
rect 4306 24520 6090 24576
rect 6146 24520 6151 24576
rect 3926 24518 6151 24520
rect 9124 24578 9184 24654
rect 10593 24712 12683 24714
rect 10593 24656 10598 24712
rect 10654 24656 12622 24712
rect 12678 24656 12683 24712
rect 10593 24654 12683 24656
rect 10593 24651 10659 24654
rect 12617 24651 12683 24654
rect 13632 24654 14474 24714
rect 13445 24578 13511 24581
rect 9124 24576 13511 24578
rect 9124 24520 13450 24576
rect 13506 24520 13511 24576
rect 9124 24518 13511 24520
rect -300 24488 160 24518
rect 3233 24515 3299 24518
rect 4245 24515 4311 24518
rect 6085 24515 6151 24518
rect 13445 24515 13511 24518
rect 3545 24512 3861 24513
rect 3545 24448 3551 24512
rect 3615 24448 3631 24512
rect 3695 24448 3711 24512
rect 3775 24448 3791 24512
rect 3855 24448 3861 24512
rect 3545 24447 3861 24448
rect 8743 24512 9059 24513
rect 8743 24448 8749 24512
rect 8813 24448 8829 24512
rect 8893 24448 8909 24512
rect 8973 24448 8989 24512
rect 9053 24448 9059 24512
rect 8743 24447 9059 24448
rect 1393 24442 1459 24445
rect 4245 24444 4311 24445
rect 4245 24442 4292 24444
rect 752 24440 1459 24442
rect 752 24384 1398 24440
rect 1454 24384 1459 24440
rect 752 24382 1459 24384
rect 4200 24440 4292 24442
rect 4200 24384 4250 24440
rect 4200 24382 4292 24384
rect -300 24306 160 24336
rect 752 24306 812 24382
rect 1393 24379 1459 24382
rect 4245 24380 4292 24382
rect 4356 24380 4362 24444
rect 4981 24442 5047 24445
rect 5809 24442 5875 24445
rect 4981 24440 5875 24442
rect 4981 24384 4986 24440
rect 5042 24384 5814 24440
rect 5870 24384 5875 24440
rect 4981 24382 5875 24384
rect 4245 24379 4311 24380
rect 4981 24379 5047 24382
rect 5809 24379 5875 24382
rect 7598 24380 7604 24444
rect 7668 24442 7674 24444
rect 8201 24442 8267 24445
rect 13632 24442 13692 24654
rect 14414 24578 14474 24654
rect 14641 24712 14780 24714
rect 14641 24656 14646 24712
rect 14702 24656 14780 24712
rect 14641 24654 14780 24656
rect 14641 24651 14707 24654
rect 14774 24652 14780 24654
rect 14844 24652 14850 24716
rect 14917 24712 14964 24716
rect 15028 24714 15034 24716
rect 14917 24656 14922 24712
rect 14917 24652 14964 24656
rect 15028 24654 15074 24714
rect 15028 24652 15034 24654
rect 16982 24652 16988 24716
rect 17052 24714 17058 24716
rect 18413 24714 18479 24717
rect 17052 24712 18479 24714
rect 17052 24656 18418 24712
rect 18474 24656 18479 24712
rect 17052 24654 18479 24656
rect 17052 24652 17058 24654
rect 14917 24651 14983 24652
rect 18413 24651 18479 24654
rect 14958 24578 14964 24580
rect 14414 24518 14964 24578
rect 14958 24516 14964 24518
rect 15028 24578 15034 24580
rect 21449 24578 21515 24581
rect 22840 24578 23300 24608
rect 15028 24518 16452 24578
rect 15028 24516 15034 24518
rect 13941 24512 14257 24513
rect 13941 24448 13947 24512
rect 14011 24448 14027 24512
rect 14091 24448 14107 24512
rect 14171 24448 14187 24512
rect 14251 24448 14257 24512
rect 13941 24447 14257 24448
rect 16392 24445 16452 24518
rect 21449 24576 23300 24578
rect 21449 24520 21454 24576
rect 21510 24520 23300 24576
rect 21449 24518 23300 24520
rect 21449 24515 21515 24518
rect 19139 24512 19455 24513
rect 19139 24448 19145 24512
rect 19209 24448 19225 24512
rect 19289 24448 19305 24512
rect 19369 24448 19385 24512
rect 19449 24448 19455 24512
rect 22840 24488 23300 24518
rect 19139 24447 19455 24448
rect 7668 24440 8267 24442
rect 7668 24384 8206 24440
rect 8262 24384 8267 24440
rect 7668 24382 8267 24384
rect 7668 24380 7674 24382
rect 8201 24379 8267 24382
rect 9492 24382 13692 24442
rect 16389 24440 16455 24445
rect 16389 24384 16394 24440
rect 16450 24384 16455 24440
rect -300 24246 812 24306
rect 5809 24306 5875 24309
rect 5942 24306 5948 24308
rect 5809 24304 5948 24306
rect 5809 24248 5814 24304
rect 5870 24248 5948 24304
rect 5809 24246 5948 24248
rect -300 24216 160 24246
rect 5809 24243 5875 24246
rect 5942 24244 5948 24246
rect 6012 24244 6018 24308
rect 7598 24244 7604 24308
rect 7668 24306 7674 24308
rect 7925 24306 7991 24309
rect 7668 24304 7991 24306
rect 7668 24248 7930 24304
rect 7986 24248 7991 24304
rect 7668 24246 7991 24248
rect 7668 24244 7674 24246
rect 7925 24243 7991 24246
rect 4337 24172 4403 24173
rect 4286 24170 4292 24172
rect 4210 24110 4292 24170
rect 4356 24170 4403 24172
rect 7189 24170 7255 24173
rect 9305 24170 9371 24173
rect 9492 24170 9552 24382
rect 16389 24379 16455 24384
rect 10317 24306 10383 24309
rect 20253 24306 20319 24309
rect 10317 24304 20319 24306
rect 10317 24248 10322 24304
rect 10378 24248 20258 24304
rect 20314 24248 20319 24304
rect 10317 24246 20319 24248
rect 10317 24243 10383 24246
rect 20253 24243 20319 24246
rect 4356 24168 6746 24170
rect 4398 24112 6746 24168
rect 4286 24108 4292 24110
rect 4356 24110 6746 24112
rect 4356 24108 4403 24110
rect 4337 24107 4403 24108
rect -300 24034 160 24064
rect 1577 24034 1643 24037
rect -300 24032 1643 24034
rect -300 23976 1582 24032
rect 1638 23976 1643 24032
rect -300 23974 1643 23976
rect -300 23944 160 23974
rect 1577 23971 1643 23974
rect 4797 24034 4863 24037
rect 5022 24034 5028 24036
rect 4797 24032 5028 24034
rect 4797 23976 4802 24032
rect 4858 23976 5028 24032
rect 4797 23974 5028 23976
rect 4797 23971 4863 23974
rect 5022 23972 5028 23974
rect 5092 23972 5098 24036
rect 6686 24034 6746 24110
rect 7189 24168 9552 24170
rect 7189 24112 7194 24168
rect 7250 24112 9310 24168
rect 9366 24112 9552 24168
rect 7189 24110 9552 24112
rect 7189 24107 7255 24110
rect 9305 24107 9371 24110
rect 9622 24108 9628 24172
rect 9692 24170 9698 24172
rect 17350 24170 17356 24172
rect 9692 24110 17356 24170
rect 9692 24108 9698 24110
rect 17350 24108 17356 24110
rect 17420 24108 17426 24172
rect 10041 24034 10107 24037
rect 6686 24032 10107 24034
rect 6686 23976 10046 24032
rect 10102 23976 10107 24032
rect 6686 23974 10107 23976
rect 10041 23971 10107 23974
rect 14457 24034 14523 24037
rect 15142 24034 15148 24036
rect 14457 24032 15148 24034
rect 14457 23976 14462 24032
rect 14518 23976 15148 24032
rect 14457 23974 15148 23976
rect 14457 23971 14523 23974
rect 15142 23972 15148 23974
rect 15212 23972 15218 24036
rect 22185 24034 22251 24037
rect 22840 24034 23300 24064
rect 22185 24032 23300 24034
rect 22185 23976 22190 24032
rect 22246 23976 23300 24032
rect 22185 23974 23300 23976
rect 22185 23971 22251 23974
rect 6144 23968 6460 23969
rect 6144 23904 6150 23968
rect 6214 23904 6230 23968
rect 6294 23904 6310 23968
rect 6374 23904 6390 23968
rect 6454 23904 6460 23968
rect 6144 23903 6460 23904
rect 11342 23968 11658 23969
rect 11342 23904 11348 23968
rect 11412 23904 11428 23968
rect 11492 23904 11508 23968
rect 11572 23904 11588 23968
rect 11652 23904 11658 23968
rect 11342 23903 11658 23904
rect 16540 23968 16856 23969
rect 16540 23904 16546 23968
rect 16610 23904 16626 23968
rect 16690 23904 16706 23968
rect 16770 23904 16786 23968
rect 16850 23904 16856 23968
rect 16540 23903 16856 23904
rect 21738 23968 22054 23969
rect 21738 23904 21744 23968
rect 21808 23904 21824 23968
rect 21888 23904 21904 23968
rect 21968 23904 21984 23968
rect 22048 23904 22054 23968
rect 22840 23944 23300 23974
rect 21738 23903 22054 23904
rect 7046 23836 7052 23900
rect 7116 23898 7122 23900
rect 10317 23898 10383 23901
rect 7116 23896 10383 23898
rect 7116 23840 10322 23896
rect 10378 23840 10383 23896
rect 7116 23838 10383 23840
rect 7116 23836 7122 23838
rect 10317 23835 10383 23838
rect 10501 23900 10567 23901
rect 10501 23896 10548 23900
rect 10612 23898 10618 23900
rect 10501 23840 10506 23896
rect 10501 23836 10548 23840
rect 10612 23838 10658 23898
rect 10612 23836 10618 23838
rect 10501 23835 10567 23836
rect -300 23762 160 23792
rect 749 23762 815 23765
rect -300 23760 815 23762
rect -300 23704 754 23760
rect 810 23704 815 23760
rect -300 23702 815 23704
rect -300 23672 160 23702
rect 749 23699 815 23702
rect 3969 23762 4035 23765
rect 19333 23762 19399 23765
rect 3969 23760 19399 23762
rect 3969 23704 3974 23760
rect 4030 23704 19338 23760
rect 19394 23704 19399 23760
rect 3969 23702 19399 23704
rect 3969 23699 4035 23702
rect 19333 23699 19399 23702
rect 3969 23626 4035 23629
rect 3969 23624 9690 23626
rect 3969 23568 3974 23624
rect 4030 23568 9690 23624
rect 3969 23566 9690 23568
rect 3969 23563 4035 23566
rect -300 23490 160 23520
rect 1393 23490 1459 23493
rect -300 23488 1459 23490
rect -300 23432 1398 23488
rect 1454 23432 1459 23488
rect -300 23430 1459 23432
rect -300 23400 160 23430
rect 1393 23427 1459 23430
rect 2814 23428 2820 23492
rect 2884 23490 2890 23492
rect 2957 23490 3023 23493
rect 2884 23488 3023 23490
rect 2884 23432 2962 23488
rect 3018 23432 3023 23488
rect 2884 23430 3023 23432
rect 2884 23428 2890 23430
rect 2957 23427 3023 23430
rect 3969 23490 4035 23493
rect 4654 23490 4660 23492
rect 3969 23488 4660 23490
rect 3969 23432 3974 23488
rect 4030 23432 4660 23488
rect 3969 23430 4660 23432
rect 3969 23427 4035 23430
rect 4654 23428 4660 23430
rect 4724 23428 4730 23492
rect 5257 23490 5323 23493
rect 8518 23490 8524 23492
rect 5257 23488 8524 23490
rect 5257 23432 5262 23488
rect 5318 23432 8524 23488
rect 5257 23430 8524 23432
rect 5257 23427 5323 23430
rect 8518 23428 8524 23430
rect 8588 23428 8594 23492
rect 9630 23490 9690 23566
rect 11094 23564 11100 23628
rect 11164 23626 11170 23628
rect 11421 23626 11487 23629
rect 11164 23624 11487 23626
rect 11164 23568 11426 23624
rect 11482 23568 11487 23624
rect 11164 23566 11487 23568
rect 11164 23564 11170 23566
rect 11421 23563 11487 23566
rect 13721 23624 13787 23629
rect 13721 23568 13726 23624
rect 13782 23568 13787 23624
rect 13721 23563 13787 23568
rect 10869 23490 10935 23493
rect 13724 23490 13784 23563
rect 9630 23488 13784 23490
rect 9630 23432 10874 23488
rect 10930 23432 13784 23488
rect 9630 23430 13784 23432
rect 10869 23427 10935 23430
rect 16246 23428 16252 23492
rect 16316 23490 16322 23492
rect 17125 23490 17191 23493
rect 16316 23488 17191 23490
rect 16316 23432 17130 23488
rect 17186 23432 17191 23488
rect 16316 23430 17191 23432
rect 16316 23428 16322 23430
rect 17125 23427 17191 23430
rect 19517 23490 19583 23493
rect 19885 23490 19951 23493
rect 19517 23488 19951 23490
rect 19517 23432 19522 23488
rect 19578 23432 19890 23488
rect 19946 23432 19951 23488
rect 19517 23430 19951 23432
rect 19517 23427 19583 23430
rect 19885 23427 19951 23430
rect 20345 23490 20411 23493
rect 21398 23490 21404 23492
rect 20345 23488 21404 23490
rect 20345 23432 20350 23488
rect 20406 23432 21404 23488
rect 20345 23430 21404 23432
rect 20345 23427 20411 23430
rect 21398 23428 21404 23430
rect 21468 23428 21474 23492
rect 21541 23490 21607 23493
rect 22840 23490 23300 23520
rect 21541 23488 23300 23490
rect 21541 23432 21546 23488
rect 21602 23432 23300 23488
rect 21541 23430 23300 23432
rect 21541 23427 21607 23430
rect 3545 23424 3861 23425
rect 3545 23360 3551 23424
rect 3615 23360 3631 23424
rect 3695 23360 3711 23424
rect 3775 23360 3791 23424
rect 3855 23360 3861 23424
rect 3545 23359 3861 23360
rect 8743 23424 9059 23425
rect 8743 23360 8749 23424
rect 8813 23360 8829 23424
rect 8893 23360 8909 23424
rect 8973 23360 8989 23424
rect 9053 23360 9059 23424
rect 8743 23359 9059 23360
rect 13941 23424 14257 23425
rect 13941 23360 13947 23424
rect 14011 23360 14027 23424
rect 14091 23360 14107 23424
rect 14171 23360 14187 23424
rect 14251 23360 14257 23424
rect 13941 23359 14257 23360
rect 19139 23424 19455 23425
rect 19139 23360 19145 23424
rect 19209 23360 19225 23424
rect 19289 23360 19305 23424
rect 19369 23360 19385 23424
rect 19449 23360 19455 23424
rect 22840 23400 23300 23430
rect 19139 23359 19455 23360
rect 5073 23354 5139 23357
rect 9581 23354 9647 23357
rect 12617 23354 12683 23357
rect 5073 23352 7482 23354
rect 5073 23296 5078 23352
rect 5134 23296 7482 23352
rect 5073 23294 7482 23296
rect 5073 23291 5139 23294
rect -300 23218 160 23248
rect 2773 23218 2839 23221
rect -300 23216 2839 23218
rect -300 23160 2778 23216
rect 2834 23160 2839 23216
rect -300 23158 2839 23160
rect -300 23128 160 23158
rect 2773 23155 2839 23158
rect 3601 23218 3667 23221
rect 4245 23218 4311 23221
rect 6545 23218 6611 23221
rect 7281 23220 7347 23221
rect 7230 23218 7236 23220
rect 3601 23216 6611 23218
rect 3601 23160 3606 23216
rect 3662 23160 4250 23216
rect 4306 23160 6550 23216
rect 6606 23160 6611 23216
rect 3601 23158 6611 23160
rect 7190 23158 7236 23218
rect 7300 23216 7347 23220
rect 7342 23160 7347 23216
rect 3601 23155 3667 23158
rect 4245 23155 4311 23158
rect 6545 23155 6611 23158
rect 7230 23156 7236 23158
rect 7300 23156 7347 23160
rect 7422 23218 7482 23294
rect 9581 23352 12683 23354
rect 9581 23296 9586 23352
rect 9642 23296 12622 23352
rect 12678 23296 12683 23352
rect 9581 23294 12683 23296
rect 9581 23291 9647 23294
rect 12617 23291 12683 23294
rect 15377 23354 15443 23357
rect 17401 23354 17467 23357
rect 15377 23352 17467 23354
rect 15377 23296 15382 23352
rect 15438 23296 17406 23352
rect 17462 23296 17467 23352
rect 15377 23294 17467 23296
rect 15377 23291 15443 23294
rect 17401 23291 17467 23294
rect 19517 23354 19583 23357
rect 20621 23354 20687 23357
rect 19517 23352 20687 23354
rect 19517 23296 19522 23352
rect 19578 23296 20626 23352
rect 20682 23296 20687 23352
rect 19517 23294 20687 23296
rect 19517 23291 19583 23294
rect 20621 23291 20687 23294
rect 21214 23292 21220 23356
rect 21284 23292 21290 23356
rect 7422 23158 13370 23218
rect 7281 23155 7347 23156
rect 1577 23082 1643 23085
rect 12893 23082 12959 23085
rect 1577 23080 12959 23082
rect 1577 23024 1582 23080
rect 1638 23024 12898 23080
rect 12954 23024 12959 23080
rect 1577 23022 12959 23024
rect 13310 23082 13370 23158
rect 13486 23156 13492 23220
rect 13556 23218 13562 23220
rect 15469 23218 15535 23221
rect 21222 23218 21282 23292
rect 13556 23216 15535 23218
rect 13556 23160 15474 23216
rect 15530 23160 15535 23216
rect 13556 23158 15535 23160
rect 13556 23156 13562 23158
rect 15469 23155 15535 23158
rect 15702 23158 21282 23218
rect 15377 23082 15443 23085
rect 13310 23080 15443 23082
rect 13310 23024 15382 23080
rect 15438 23024 15443 23080
rect 13310 23022 15443 23024
rect 1577 23019 1643 23022
rect 12893 23019 12959 23022
rect 15377 23019 15443 23022
rect 15561 23082 15627 23085
rect 15702 23082 15762 23158
rect 15561 23080 15762 23082
rect 15561 23024 15566 23080
rect 15622 23024 15762 23080
rect 15561 23022 15762 23024
rect 19333 23082 19399 23085
rect 20345 23082 20411 23085
rect 19333 23080 20411 23082
rect 19333 23024 19338 23080
rect 19394 23024 20350 23080
rect 20406 23024 20411 23080
rect 19333 23022 20411 23024
rect 15561 23019 15627 23022
rect 19333 23019 19399 23022
rect 20345 23019 20411 23022
rect -300 22946 160 22976
rect 1301 22946 1367 22949
rect -300 22944 1367 22946
rect -300 22888 1306 22944
rect 1362 22888 1367 22944
rect -300 22886 1367 22888
rect -300 22856 160 22886
rect 1301 22883 1367 22886
rect 2630 22884 2636 22948
rect 2700 22946 2706 22948
rect 5073 22946 5139 22949
rect 2700 22944 5139 22946
rect 2700 22888 5078 22944
rect 5134 22888 5139 22944
rect 2700 22886 5139 22888
rect 2700 22884 2706 22886
rect 5073 22883 5139 22886
rect 7782 22884 7788 22948
rect 7852 22946 7858 22948
rect 9581 22946 9647 22949
rect 7852 22944 9647 22946
rect 7852 22888 9586 22944
rect 9642 22888 9647 22944
rect 7852 22886 9647 22888
rect 7852 22884 7858 22886
rect 9581 22883 9647 22886
rect 9857 22944 9923 22949
rect 9857 22888 9862 22944
rect 9918 22888 9923 22944
rect 9857 22883 9923 22888
rect 10041 22946 10107 22949
rect 11145 22946 11211 22949
rect 10041 22944 11211 22946
rect 10041 22888 10046 22944
rect 10102 22888 11150 22944
rect 11206 22888 11211 22944
rect 10041 22886 11211 22888
rect 10041 22883 10107 22886
rect 11145 22883 11211 22886
rect 13118 22884 13124 22948
rect 13188 22946 13194 22948
rect 15561 22946 15627 22949
rect 13188 22944 15627 22946
rect 13188 22888 15566 22944
rect 15622 22888 15627 22944
rect 13188 22886 15627 22888
rect 13188 22884 13194 22886
rect 15561 22883 15627 22886
rect 19333 22946 19399 22949
rect 19885 22946 19951 22949
rect 19333 22944 19951 22946
rect 19333 22888 19338 22944
rect 19394 22888 19890 22944
rect 19946 22888 19951 22944
rect 19333 22886 19951 22888
rect 19333 22883 19399 22886
rect 19885 22883 19951 22886
rect 22185 22946 22251 22949
rect 22840 22946 23300 22976
rect 22185 22944 23300 22946
rect 22185 22888 22190 22944
rect 22246 22888 23300 22944
rect 22185 22886 23300 22888
rect 22185 22883 22251 22886
rect 6144 22880 6460 22881
rect 6144 22816 6150 22880
rect 6214 22816 6230 22880
rect 6294 22816 6310 22880
rect 6374 22816 6390 22880
rect 6454 22816 6460 22880
rect 6144 22815 6460 22816
rect 1669 22810 1735 22813
rect 2405 22810 2471 22813
rect 5441 22810 5507 22813
rect 1669 22808 5507 22810
rect 1669 22752 1674 22808
rect 1730 22752 2410 22808
rect 2466 22752 5446 22808
rect 5502 22752 5507 22808
rect 1669 22750 5507 22752
rect 9860 22810 9920 22883
rect 11342 22880 11658 22881
rect 11342 22816 11348 22880
rect 11412 22816 11428 22880
rect 11492 22816 11508 22880
rect 11572 22816 11588 22880
rect 11652 22816 11658 22880
rect 11342 22815 11658 22816
rect 16540 22880 16856 22881
rect 16540 22816 16546 22880
rect 16610 22816 16626 22880
rect 16690 22816 16706 22880
rect 16770 22816 16786 22880
rect 16850 22816 16856 22880
rect 16540 22815 16856 22816
rect 21738 22880 22054 22881
rect 21738 22816 21744 22880
rect 21808 22816 21824 22880
rect 21888 22816 21904 22880
rect 21968 22816 21984 22880
rect 22048 22816 22054 22880
rect 22840 22856 23300 22886
rect 21738 22815 22054 22816
rect 11145 22810 11211 22813
rect 13077 22812 13143 22813
rect 13077 22810 13124 22812
rect 9860 22808 11211 22810
rect 9860 22752 11150 22808
rect 11206 22752 11211 22808
rect 9860 22750 11211 22752
rect 13036 22808 13124 22810
rect 13188 22810 13194 22812
rect 16297 22810 16363 22813
rect 13188 22808 16363 22810
rect 13036 22752 13082 22808
rect 13188 22752 16302 22808
rect 16358 22752 16363 22808
rect 13036 22750 13124 22752
rect 1669 22747 1735 22750
rect 2405 22747 2471 22750
rect 5441 22747 5507 22750
rect 11145 22747 11211 22750
rect 13077 22748 13124 22750
rect 13188 22750 16363 22752
rect 13188 22748 13194 22750
rect 13077 22747 13143 22748
rect 16297 22747 16363 22750
rect 19333 22810 19399 22813
rect 21541 22810 21607 22813
rect 22369 22810 22435 22813
rect 19333 22808 21607 22810
rect 19333 22752 19338 22808
rect 19394 22752 21546 22808
rect 21602 22752 21607 22808
rect 19333 22750 21607 22752
rect 19333 22747 19399 22750
rect 21541 22747 21607 22750
rect 22188 22808 22435 22810
rect 22188 22752 22374 22808
rect 22430 22752 22435 22808
rect 22188 22750 22435 22752
rect -300 22674 160 22704
rect 22188 22677 22248 22750
rect 22369 22747 22435 22750
rect 1117 22674 1183 22677
rect -300 22672 1183 22674
rect -300 22616 1122 22672
rect 1178 22616 1183 22672
rect -300 22614 1183 22616
rect -300 22584 160 22614
rect 1117 22611 1183 22614
rect 2221 22674 2287 22677
rect 10961 22674 11027 22677
rect 2221 22672 11027 22674
rect 2221 22616 2226 22672
rect 2282 22616 10966 22672
rect 11022 22616 11027 22672
rect 2221 22614 11027 22616
rect 2221 22611 2287 22614
rect 10961 22611 11027 22614
rect 11094 22612 11100 22676
rect 11164 22674 11170 22676
rect 20253 22674 20319 22677
rect 11164 22672 20319 22674
rect 11164 22616 20258 22672
rect 20314 22616 20319 22672
rect 11164 22614 20319 22616
rect 11164 22612 11170 22614
rect 20253 22611 20319 22614
rect 22185 22672 22251 22677
rect 22185 22616 22190 22672
rect 22246 22616 22251 22672
rect 22185 22611 22251 22616
rect 1117 22538 1183 22541
rect 4613 22538 4679 22541
rect 1117 22536 4679 22538
rect 1117 22480 1122 22536
rect 1178 22480 4618 22536
rect 4674 22480 4679 22536
rect 1117 22478 4679 22480
rect 1117 22475 1183 22478
rect 4613 22475 4679 22478
rect 5717 22538 5783 22541
rect 15009 22538 15075 22541
rect 5717 22536 15075 22538
rect 5717 22480 5722 22536
rect 5778 22480 15014 22536
rect 15070 22480 15075 22536
rect 5717 22478 15075 22480
rect 5717 22475 5783 22478
rect 15009 22475 15075 22478
rect 19558 22476 19564 22540
rect 19628 22538 19634 22540
rect 22093 22538 22159 22541
rect 19628 22536 22159 22538
rect 19628 22480 22098 22536
rect 22154 22480 22159 22536
rect 19628 22478 22159 22480
rect 19628 22476 19634 22478
rect 22093 22475 22159 22478
rect -300 22402 160 22432
rect 2313 22402 2379 22405
rect -300 22400 2379 22402
rect -300 22344 2318 22400
rect 2374 22344 2379 22400
rect -300 22342 2379 22344
rect -300 22312 160 22342
rect 2313 22339 2379 22342
rect 4654 22340 4660 22404
rect 4724 22402 4730 22404
rect 7782 22402 7788 22404
rect 4724 22342 7788 22402
rect 4724 22340 4730 22342
rect 7782 22340 7788 22342
rect 7852 22340 7858 22404
rect 10174 22340 10180 22404
rect 10244 22402 10250 22404
rect 10317 22402 10383 22405
rect 10244 22400 10383 22402
rect 10244 22344 10322 22400
rect 10378 22344 10383 22400
rect 10244 22342 10383 22344
rect 10244 22340 10250 22342
rect 10317 22339 10383 22342
rect 10961 22402 11027 22405
rect 12934 22402 12940 22404
rect 10961 22400 12940 22402
rect 10961 22344 10966 22400
rect 11022 22344 12940 22400
rect 10961 22342 12940 22344
rect 10961 22339 11027 22342
rect 12934 22340 12940 22342
rect 13004 22340 13010 22404
rect 21449 22402 21515 22405
rect 22840 22402 23300 22432
rect 21449 22400 23300 22402
rect 21449 22344 21454 22400
rect 21510 22344 23300 22400
rect 21449 22342 23300 22344
rect 21449 22339 21515 22342
rect 3545 22336 3861 22337
rect 3545 22272 3551 22336
rect 3615 22272 3631 22336
rect 3695 22272 3711 22336
rect 3775 22272 3791 22336
rect 3855 22272 3861 22336
rect 3545 22271 3861 22272
rect 8743 22336 9059 22337
rect 8743 22272 8749 22336
rect 8813 22272 8829 22336
rect 8893 22272 8909 22336
rect 8973 22272 8989 22336
rect 9053 22272 9059 22336
rect 8743 22271 9059 22272
rect 13941 22336 14257 22337
rect 13941 22272 13947 22336
rect 14011 22272 14027 22336
rect 14091 22272 14107 22336
rect 14171 22272 14187 22336
rect 14251 22272 14257 22336
rect 13941 22271 14257 22272
rect 19139 22336 19455 22337
rect 19139 22272 19145 22336
rect 19209 22272 19225 22336
rect 19289 22272 19305 22336
rect 19369 22272 19385 22336
rect 19449 22272 19455 22336
rect 22840 22312 23300 22342
rect 19139 22271 19455 22272
rect 4337 22266 4403 22269
rect 6453 22266 6519 22269
rect 4337 22264 6519 22266
rect 4337 22208 4342 22264
rect 4398 22208 6458 22264
rect 6514 22208 6519 22264
rect 4337 22206 6519 22208
rect 4337 22203 4403 22206
rect 6453 22203 6519 22206
rect 6862 22204 6868 22268
rect 6932 22266 6938 22268
rect 7557 22266 7623 22269
rect 6932 22264 7623 22266
rect 6932 22208 7562 22264
rect 7618 22208 7623 22264
rect 6932 22206 7623 22208
rect 6932 22204 6938 22206
rect 7557 22203 7623 22206
rect 10910 22204 10916 22268
rect 10980 22266 10986 22268
rect 11145 22266 11211 22269
rect 10980 22264 11211 22266
rect 10980 22208 11150 22264
rect 11206 22208 11211 22264
rect 10980 22206 11211 22208
rect 10980 22204 10986 22206
rect 11145 22203 11211 22206
rect 12433 22264 12499 22269
rect 14825 22268 14891 22269
rect 14774 22266 14780 22268
rect 12433 22208 12438 22264
rect 12494 22208 12499 22264
rect 12433 22203 12499 22208
rect 14734 22206 14780 22266
rect 14844 22264 14891 22268
rect 14886 22208 14891 22264
rect 14774 22204 14780 22206
rect 14844 22204 14891 22208
rect 14825 22203 14891 22204
rect -300 22130 160 22160
rect 1393 22130 1459 22133
rect -300 22128 1459 22130
rect -300 22072 1398 22128
rect 1454 22072 1459 22128
rect -300 22070 1459 22072
rect -300 22040 160 22070
rect 1393 22067 1459 22070
rect 2589 22130 2655 22133
rect 8109 22130 8175 22133
rect 2589 22128 8175 22130
rect 2589 22072 2594 22128
rect 2650 22072 8114 22128
rect 8170 22072 8175 22128
rect 2589 22070 8175 22072
rect 2589 22067 2655 22070
rect 8109 22067 8175 22070
rect 8385 22130 8451 22133
rect 11094 22130 11100 22132
rect 8385 22128 11100 22130
rect 8385 22072 8390 22128
rect 8446 22072 11100 22128
rect 8385 22070 11100 22072
rect 8385 22067 8451 22070
rect 11094 22068 11100 22070
rect 11164 22068 11170 22132
rect 657 21994 723 21997
rect 6269 21994 6335 21997
rect 657 21992 6335 21994
rect 657 21936 662 21992
rect 718 21936 6274 21992
rect 6330 21936 6335 21992
rect 657 21934 6335 21936
rect 657 21931 723 21934
rect 6269 21931 6335 21934
rect 8201 21994 8267 21997
rect 9397 21994 9463 21997
rect 11830 21994 11836 21996
rect 8201 21992 9463 21994
rect 8201 21936 8206 21992
rect 8262 21936 9402 21992
rect 9458 21936 9463 21992
rect 8201 21934 9463 21936
rect 8201 21931 8267 21934
rect 9397 21931 9463 21934
rect 11148 21934 11836 21994
rect -300 21858 160 21888
rect 1209 21858 1275 21861
rect -300 21856 1275 21858
rect -300 21800 1214 21856
rect 1270 21800 1275 21856
rect -300 21798 1275 21800
rect -300 21768 160 21798
rect 1209 21795 1275 21798
rect 2037 21858 2103 21861
rect 4613 21858 4679 21861
rect 11148 21858 11208 21934
rect 11830 21932 11836 21934
rect 11900 21932 11906 21996
rect 12436 21994 12496 22203
rect 13077 22130 13143 22133
rect 13445 22130 13511 22133
rect 13077 22128 13511 22130
rect 13077 22072 13082 22128
rect 13138 22072 13450 22128
rect 13506 22072 13511 22128
rect 13077 22070 13511 22072
rect 13077 22067 13143 22070
rect 13445 22067 13511 22070
rect 19793 22130 19859 22133
rect 19926 22130 19932 22132
rect 19793 22128 19932 22130
rect 19793 22072 19798 22128
rect 19854 22072 19932 22128
rect 19793 22070 19932 22072
rect 19793 22067 19859 22070
rect 19926 22068 19932 22070
rect 19996 22068 20002 22132
rect 21541 22130 21607 22133
rect 22001 22130 22067 22133
rect 21541 22128 22067 22130
rect 21541 22072 21546 22128
rect 21602 22072 22006 22128
rect 22062 22072 22067 22128
rect 21541 22070 22067 22072
rect 21541 22067 21607 22070
rect 22001 22067 22067 22070
rect 12617 21994 12683 21997
rect 12436 21992 12683 21994
rect 12436 21936 12622 21992
rect 12678 21936 12683 21992
rect 12436 21934 12683 21936
rect 2037 21856 4679 21858
rect 2037 21800 2042 21856
rect 2098 21800 4618 21856
rect 4674 21800 4679 21856
rect 2037 21798 4679 21800
rect 2037 21795 2103 21798
rect 4613 21795 4679 21798
rect 9078 21798 11208 21858
rect 11838 21858 11898 21932
rect 12617 21931 12683 21934
rect 18505 21994 18571 21997
rect 22645 21994 22711 21997
rect 18505 21992 22711 21994
rect 18505 21936 18510 21992
rect 18566 21936 22650 21992
rect 22706 21936 22711 21992
rect 18505 21934 22711 21936
rect 18505 21931 18571 21934
rect 22645 21931 22711 21934
rect 13445 21858 13511 21861
rect 11838 21856 13511 21858
rect 11838 21800 13450 21856
rect 13506 21800 13511 21856
rect 11838 21798 13511 21800
rect 6144 21792 6460 21793
rect 6144 21728 6150 21792
rect 6214 21728 6230 21792
rect 6294 21728 6310 21792
rect 6374 21728 6390 21792
rect 6454 21728 6460 21792
rect 6144 21727 6460 21728
rect 1669 21722 1735 21725
rect 4245 21722 4311 21725
rect 1669 21720 4311 21722
rect 1669 21664 1674 21720
rect 1730 21664 4250 21720
rect 4306 21664 4311 21720
rect 1669 21662 4311 21664
rect 1669 21659 1735 21662
rect 4245 21659 4311 21662
rect -300 21586 160 21616
rect 749 21586 815 21589
rect 9078 21586 9138 21798
rect 13445 21795 13511 21798
rect 17033 21858 17099 21861
rect 18137 21858 18203 21861
rect 17033 21856 18203 21858
rect 17033 21800 17038 21856
rect 17094 21800 18142 21856
rect 18198 21800 18203 21856
rect 17033 21798 18203 21800
rect 17033 21795 17099 21798
rect 18137 21795 18203 21798
rect 22185 21858 22251 21861
rect 22840 21858 23300 21888
rect 22185 21856 23300 21858
rect 22185 21800 22190 21856
rect 22246 21800 23300 21856
rect 22185 21798 23300 21800
rect 22185 21795 22251 21798
rect 11342 21792 11658 21793
rect 11342 21728 11348 21792
rect 11412 21728 11428 21792
rect 11492 21728 11508 21792
rect 11572 21728 11588 21792
rect 11652 21728 11658 21792
rect 11342 21727 11658 21728
rect 16540 21792 16856 21793
rect 16540 21728 16546 21792
rect 16610 21728 16626 21792
rect 16690 21728 16706 21792
rect 16770 21728 16786 21792
rect 16850 21728 16856 21792
rect 16540 21727 16856 21728
rect 21738 21792 22054 21793
rect 21738 21728 21744 21792
rect 21808 21728 21824 21792
rect 21888 21728 21904 21792
rect 21968 21728 21984 21792
rect 22048 21728 22054 21792
rect 22840 21768 23300 21798
rect 21738 21727 22054 21728
rect 9949 21722 10015 21725
rect -300 21584 815 21586
rect -300 21528 754 21584
rect 810 21528 815 21584
rect -300 21526 815 21528
rect -300 21496 160 21526
rect 749 21523 815 21526
rect 2730 21526 9138 21586
rect 9216 21720 10015 21722
rect 9216 21664 9954 21720
rect 10010 21664 10015 21720
rect 9216 21662 10015 21664
rect 1761 21450 1827 21453
rect 2730 21450 2790 21526
rect 1761 21448 2790 21450
rect 1761 21392 1766 21448
rect 1822 21392 2790 21448
rect 1761 21390 2790 21392
rect 5533 21450 5599 21453
rect 6862 21450 6868 21452
rect 5533 21448 6868 21450
rect 5533 21392 5538 21448
rect 5594 21392 6868 21448
rect 5533 21390 6868 21392
rect 1761 21387 1827 21390
rect 5533 21387 5599 21390
rect 6862 21388 6868 21390
rect 6932 21388 6938 21452
rect 9216 21450 9276 21662
rect 9949 21659 10015 21662
rect 12198 21660 12204 21724
rect 12268 21722 12274 21724
rect 13169 21722 13235 21725
rect 12268 21720 13235 21722
rect 12268 21664 13174 21720
rect 13230 21664 13235 21720
rect 12268 21662 13235 21664
rect 12268 21660 12274 21662
rect 13169 21659 13235 21662
rect 8572 21390 9276 21450
rect -300 21314 160 21344
rect 1485 21314 1551 21317
rect -300 21312 1551 21314
rect -300 21256 1490 21312
rect 1546 21256 1551 21312
rect -300 21254 1551 21256
rect -300 21224 160 21254
rect 1485 21251 1551 21254
rect 1945 21314 2011 21317
rect 3049 21314 3115 21317
rect 1945 21312 3115 21314
rect 1945 21256 1950 21312
rect 2006 21256 3054 21312
rect 3110 21256 3115 21312
rect 1945 21254 3115 21256
rect 1945 21251 2011 21254
rect 3049 21251 3115 21254
rect 4429 21314 4495 21317
rect 7281 21314 7347 21317
rect 8017 21314 8083 21317
rect 4429 21312 8083 21314
rect 4429 21256 4434 21312
rect 4490 21256 7286 21312
rect 7342 21256 8022 21312
rect 8078 21256 8083 21312
rect 4429 21254 8083 21256
rect 4429 21251 4495 21254
rect 7281 21251 7347 21254
rect 8017 21251 8083 21254
rect 3545 21248 3861 21249
rect 3545 21184 3551 21248
rect 3615 21184 3631 21248
rect 3695 21184 3711 21248
rect 3775 21184 3791 21248
rect 3855 21184 3861 21248
rect 3545 21183 3861 21184
rect 2078 21116 2084 21180
rect 2148 21178 2154 21180
rect 2405 21178 2471 21181
rect 2148 21176 2471 21178
rect 2148 21120 2410 21176
rect 2466 21120 2471 21176
rect 2148 21118 2471 21120
rect 2148 21116 2154 21118
rect 2405 21115 2471 21118
rect 2681 21176 2747 21181
rect 2681 21120 2686 21176
rect 2742 21120 2747 21176
rect 2681 21115 2747 21120
rect 4613 21178 4679 21181
rect 8293 21178 8359 21181
rect 4613 21176 8359 21178
rect 4613 21120 4618 21176
rect 4674 21120 8298 21176
rect 8354 21120 8359 21176
rect 4613 21118 8359 21120
rect 4613 21115 4679 21118
rect 8293 21115 8359 21118
rect -300 21042 160 21072
rect 749 21042 815 21045
rect -300 21040 815 21042
rect -300 20984 754 21040
rect 810 20984 815 21040
rect -300 20982 815 20984
rect 2684 21042 2744 21115
rect 8572 21042 8632 21390
rect 10542 21388 10548 21452
rect 10612 21450 10618 21452
rect 11421 21450 11487 21453
rect 10612 21448 11487 21450
rect 10612 21392 11426 21448
rect 11482 21392 11487 21448
rect 10612 21390 11487 21392
rect 10612 21388 10618 21390
rect 11421 21387 11487 21390
rect 12198 21388 12204 21452
rect 12268 21450 12274 21452
rect 14273 21450 14339 21453
rect 12268 21448 14339 21450
rect 12268 21392 14278 21448
rect 14334 21392 14339 21448
rect 12268 21390 14339 21392
rect 12268 21388 12274 21390
rect 14273 21387 14339 21390
rect 9397 21314 9463 21317
rect 10317 21314 10383 21317
rect 9397 21312 10383 21314
rect 9397 21256 9402 21312
rect 9458 21256 10322 21312
rect 10378 21256 10383 21312
rect 9397 21254 10383 21256
rect 9397 21251 9463 21254
rect 10317 21251 10383 21254
rect 20805 21314 20871 21317
rect 22840 21314 23300 21344
rect 20805 21312 23300 21314
rect 20805 21256 20810 21312
rect 20866 21256 23300 21312
rect 20805 21254 23300 21256
rect 20805 21251 20871 21254
rect 8743 21248 9059 21249
rect 8743 21184 8749 21248
rect 8813 21184 8829 21248
rect 8893 21184 8909 21248
rect 8973 21184 8989 21248
rect 9053 21184 9059 21248
rect 8743 21183 9059 21184
rect 13941 21248 14257 21249
rect 13941 21184 13947 21248
rect 14011 21184 14027 21248
rect 14091 21184 14107 21248
rect 14171 21184 14187 21248
rect 14251 21184 14257 21248
rect 13941 21183 14257 21184
rect 19139 21248 19455 21249
rect 19139 21184 19145 21248
rect 19209 21184 19225 21248
rect 19289 21184 19305 21248
rect 19369 21184 19385 21248
rect 19449 21184 19455 21248
rect 22840 21224 23300 21254
rect 19139 21183 19455 21184
rect 9806 21116 9812 21180
rect 9876 21178 9882 21180
rect 11789 21178 11855 21181
rect 9876 21176 11855 21178
rect 9876 21120 11794 21176
rect 11850 21120 11855 21176
rect 9876 21118 11855 21120
rect 9876 21116 9882 21118
rect 11789 21115 11855 21118
rect 15653 21178 15719 21181
rect 15878 21178 15884 21180
rect 15653 21176 15884 21178
rect 15653 21120 15658 21176
rect 15714 21120 15884 21176
rect 15653 21118 15884 21120
rect 15653 21115 15719 21118
rect 15878 21116 15884 21118
rect 15948 21116 15954 21180
rect 2684 20982 8632 21042
rect 9121 21042 9187 21045
rect 17677 21042 17743 21045
rect 9121 21040 17743 21042
rect 9121 20984 9126 21040
rect 9182 20984 17682 21040
rect 17738 20984 17743 21040
rect 9121 20982 17743 20984
rect -300 20952 160 20982
rect 749 20979 815 20982
rect 9121 20979 9187 20982
rect 17677 20979 17743 20982
rect 2865 20906 2931 20909
rect 4337 20906 4403 20909
rect 2865 20904 4403 20906
rect 2865 20848 2870 20904
rect 2926 20848 4342 20904
rect 4398 20848 4403 20904
rect 2865 20846 4403 20848
rect 2865 20843 2931 20846
rect 4337 20843 4403 20846
rect 6177 20906 6243 20909
rect 10961 20906 11027 20909
rect 6177 20904 11027 20906
rect 6177 20848 6182 20904
rect 6238 20848 10966 20904
rect 11022 20848 11027 20904
rect 6177 20846 11027 20848
rect 6177 20843 6243 20846
rect 10961 20843 11027 20846
rect 12985 20906 13051 20909
rect 13670 20906 13676 20908
rect 12985 20904 13676 20906
rect 12985 20848 12990 20904
rect 13046 20848 13676 20904
rect 12985 20846 13676 20848
rect 12985 20843 13051 20846
rect 13670 20844 13676 20846
rect 13740 20844 13746 20908
rect 13905 20906 13971 20909
rect 15285 20906 15351 20909
rect 13905 20904 15351 20906
rect 13905 20848 13910 20904
rect 13966 20848 15290 20904
rect 15346 20848 15351 20904
rect 13905 20846 15351 20848
rect 13905 20843 13971 20846
rect 15285 20843 15351 20846
rect 19006 20844 19012 20908
rect 19076 20906 19082 20908
rect 19742 20906 19748 20908
rect 19076 20846 19748 20906
rect 19076 20844 19082 20846
rect 19742 20844 19748 20846
rect 19812 20844 19818 20908
rect 22093 20906 22159 20909
rect 22645 20906 22711 20909
rect 22093 20904 22711 20906
rect 22093 20848 22098 20904
rect 22154 20848 22650 20904
rect 22706 20848 22711 20904
rect 22093 20846 22711 20848
rect 22093 20843 22159 20846
rect 22645 20843 22711 20846
rect -300 20770 160 20800
rect 1301 20770 1367 20773
rect 3141 20770 3207 20773
rect 5758 20770 5764 20772
rect -300 20768 1367 20770
rect -300 20712 1306 20768
rect 1362 20712 1367 20768
rect -300 20710 1367 20712
rect -300 20680 160 20710
rect 1301 20707 1367 20710
rect 2316 20710 3066 20770
rect 2316 20637 2376 20710
rect 2313 20632 2379 20637
rect 2589 20636 2655 20637
rect 2589 20634 2636 20636
rect 2313 20576 2318 20632
rect 2374 20576 2379 20632
rect 2313 20571 2379 20576
rect 2544 20632 2636 20634
rect 2544 20576 2594 20632
rect 2544 20574 2636 20576
rect 2589 20572 2636 20574
rect 2700 20572 2706 20636
rect 3006 20634 3066 20710
rect 3141 20768 5764 20770
rect 3141 20712 3146 20768
rect 3202 20712 5764 20768
rect 3141 20710 5764 20712
rect 3141 20707 3207 20710
rect 5758 20708 5764 20710
rect 5828 20708 5834 20772
rect 6913 20770 6979 20773
rect 11053 20770 11119 20773
rect 12566 20770 12572 20772
rect 6913 20768 11119 20770
rect 6913 20712 6918 20768
rect 6974 20712 11058 20768
rect 11114 20712 11119 20768
rect 6913 20710 11119 20712
rect 6913 20707 6979 20710
rect 11053 20707 11119 20710
rect 12390 20710 12572 20770
rect 6144 20704 6460 20705
rect 6144 20640 6150 20704
rect 6214 20640 6230 20704
rect 6294 20640 6310 20704
rect 6374 20640 6390 20704
rect 6454 20640 6460 20704
rect 6144 20639 6460 20640
rect 11342 20704 11658 20705
rect 11342 20640 11348 20704
rect 11412 20640 11428 20704
rect 11492 20640 11508 20704
rect 11572 20640 11588 20704
rect 11652 20640 11658 20704
rect 11342 20639 11658 20640
rect 7281 20634 7347 20637
rect 9438 20634 9444 20636
rect 3006 20574 3434 20634
rect 2589 20571 2655 20572
rect -300 20498 160 20528
rect 3233 20498 3299 20501
rect -300 20496 3299 20498
rect -300 20440 3238 20496
rect 3294 20440 3299 20496
rect -300 20438 3299 20440
rect 3374 20498 3434 20574
rect 7281 20632 9444 20634
rect 7281 20576 7286 20632
rect 7342 20576 9444 20632
rect 7281 20574 9444 20576
rect 7281 20571 7347 20574
rect 9438 20572 9444 20574
rect 9508 20572 9514 20636
rect 10358 20572 10364 20636
rect 10428 20634 10434 20636
rect 11053 20634 11119 20637
rect 10428 20632 11119 20634
rect 10428 20576 11058 20632
rect 11114 20576 11119 20632
rect 10428 20574 11119 20576
rect 10428 20572 10434 20574
rect 11053 20571 11119 20574
rect 3918 20498 3924 20500
rect 3374 20438 3924 20498
rect -300 20408 160 20438
rect 3233 20435 3299 20438
rect 3918 20436 3924 20438
rect 3988 20498 3994 20500
rect 4061 20498 4127 20501
rect 3988 20496 4127 20498
rect 3988 20440 4066 20496
rect 4122 20440 4127 20496
rect 3988 20438 4127 20440
rect 3988 20436 3994 20438
rect 4061 20435 4127 20438
rect 6453 20498 6519 20501
rect 12390 20498 12450 20710
rect 12566 20708 12572 20710
rect 12636 20708 12642 20772
rect 13118 20708 13124 20772
rect 13188 20708 13194 20772
rect 15142 20708 15148 20772
rect 15212 20770 15218 20772
rect 16062 20770 16068 20772
rect 15212 20710 16068 20770
rect 15212 20708 15218 20710
rect 16062 20708 16068 20710
rect 16132 20708 16138 20772
rect 18689 20770 18755 20773
rect 21265 20770 21331 20773
rect 18689 20768 21331 20770
rect 18689 20712 18694 20768
rect 18750 20712 21270 20768
rect 21326 20712 21331 20768
rect 18689 20710 21331 20712
rect 13126 20637 13186 20708
rect 18689 20707 18755 20710
rect 21265 20707 21331 20710
rect 22185 20770 22251 20773
rect 22840 20770 23300 20800
rect 22185 20768 23300 20770
rect 22185 20712 22190 20768
rect 22246 20712 23300 20768
rect 22185 20710 23300 20712
rect 22185 20707 22251 20710
rect 16540 20704 16856 20705
rect 16540 20640 16546 20704
rect 16610 20640 16626 20704
rect 16690 20640 16706 20704
rect 16770 20640 16786 20704
rect 16850 20640 16856 20704
rect 16540 20639 16856 20640
rect 21738 20704 22054 20705
rect 21738 20640 21744 20704
rect 21808 20640 21824 20704
rect 21888 20640 21904 20704
rect 21968 20640 21984 20704
rect 22048 20640 22054 20704
rect 22840 20680 23300 20710
rect 21738 20639 22054 20640
rect 13126 20632 13235 20637
rect 13126 20576 13174 20632
rect 13230 20576 13235 20632
rect 13126 20574 13235 20576
rect 13169 20571 13235 20574
rect 6453 20496 12450 20498
rect 6453 20440 6458 20496
rect 6514 20440 12450 20496
rect 6453 20438 12450 20440
rect 12617 20498 12683 20501
rect 12934 20498 12940 20500
rect 12617 20496 12940 20498
rect 12617 20440 12622 20496
rect 12678 20440 12940 20496
rect 12617 20438 12940 20440
rect 6453 20435 6519 20438
rect 12617 20435 12683 20438
rect 12934 20436 12940 20438
rect 13004 20436 13010 20500
rect 15326 20498 15332 20500
rect 13080 20438 15332 20498
rect 1577 20362 1643 20365
rect 10685 20362 10751 20365
rect 1577 20360 10751 20362
rect 1577 20304 1582 20360
rect 1638 20304 10690 20360
rect 10746 20304 10751 20360
rect 1577 20302 10751 20304
rect 1577 20299 1643 20302
rect 10685 20299 10751 20302
rect 11421 20362 11487 20365
rect 12433 20362 12499 20365
rect 13080 20362 13140 20438
rect 15326 20436 15332 20438
rect 15396 20436 15402 20500
rect 15929 20362 15995 20365
rect 11421 20360 13140 20362
rect 11421 20304 11426 20360
rect 11482 20304 12438 20360
rect 12494 20304 13140 20360
rect 11421 20302 13140 20304
rect 13816 20360 15995 20362
rect 13816 20304 15934 20360
rect 15990 20304 15995 20360
rect 13816 20302 15995 20304
rect 11421 20299 11487 20302
rect 12433 20299 12499 20302
rect -300 20226 160 20256
rect 1485 20226 1551 20229
rect -300 20224 1551 20226
rect -300 20168 1490 20224
rect 1546 20168 1551 20224
rect -300 20166 1551 20168
rect -300 20136 160 20166
rect 1485 20163 1551 20166
rect 4061 20226 4127 20229
rect 8293 20226 8359 20229
rect 4061 20224 8359 20226
rect 4061 20168 4066 20224
rect 4122 20168 8298 20224
rect 8354 20168 8359 20224
rect 4061 20166 8359 20168
rect 4061 20163 4127 20166
rect 8293 20163 8359 20166
rect 10041 20226 10107 20229
rect 13816 20226 13876 20302
rect 15929 20299 15995 20302
rect 16062 20300 16068 20364
rect 16132 20362 16138 20364
rect 17125 20362 17191 20365
rect 16132 20360 17191 20362
rect 16132 20304 17130 20360
rect 17186 20304 17191 20360
rect 16132 20302 17191 20304
rect 16132 20300 16138 20302
rect 17125 20299 17191 20302
rect 10041 20224 13876 20226
rect 10041 20168 10046 20224
rect 10102 20168 13876 20224
rect 10041 20166 13876 20168
rect 21449 20226 21515 20229
rect 22840 20226 23300 20256
rect 21449 20224 23300 20226
rect 21449 20168 21454 20224
rect 21510 20168 23300 20224
rect 21449 20166 23300 20168
rect 10041 20163 10107 20166
rect 21449 20163 21515 20166
rect 3545 20160 3861 20161
rect 3545 20096 3551 20160
rect 3615 20096 3631 20160
rect 3695 20096 3711 20160
rect 3775 20096 3791 20160
rect 3855 20096 3861 20160
rect 3545 20095 3861 20096
rect 8743 20160 9059 20161
rect 8743 20096 8749 20160
rect 8813 20096 8829 20160
rect 8893 20096 8909 20160
rect 8973 20096 8989 20160
rect 9053 20096 9059 20160
rect 8743 20095 9059 20096
rect 13941 20160 14257 20161
rect 13941 20096 13947 20160
rect 14011 20096 14027 20160
rect 14091 20096 14107 20160
rect 14171 20096 14187 20160
rect 14251 20096 14257 20160
rect 13941 20095 14257 20096
rect 19139 20160 19455 20161
rect 19139 20096 19145 20160
rect 19209 20096 19225 20160
rect 19289 20096 19305 20160
rect 19369 20096 19385 20160
rect 19449 20096 19455 20160
rect 22840 20136 23300 20166
rect 19139 20095 19455 20096
rect 4654 20028 4660 20092
rect 4724 20090 4730 20092
rect 7046 20090 7052 20092
rect 4724 20030 7052 20090
rect 4724 20028 4730 20030
rect 7046 20028 7052 20030
rect 7116 20028 7122 20092
rect 8334 20028 8340 20092
rect 8404 20028 8410 20092
rect 16941 20090 17007 20093
rect 17125 20090 17191 20093
rect 14966 20088 17191 20090
rect 14966 20032 16946 20088
rect 17002 20032 17130 20088
rect 17186 20032 17191 20088
rect 14966 20030 17191 20032
rect -300 19954 160 19984
rect 749 19954 815 19957
rect -300 19952 815 19954
rect -300 19896 754 19952
rect 810 19896 815 19952
rect -300 19894 815 19896
rect -300 19864 160 19894
rect 749 19891 815 19894
rect 2313 19954 2379 19957
rect 3233 19954 3299 19957
rect 2313 19952 3299 19954
rect 2313 19896 2318 19952
rect 2374 19896 3238 19952
rect 3294 19896 3299 19952
rect 2313 19894 3299 19896
rect 2313 19891 2379 19894
rect 3233 19891 3299 19894
rect 5349 19954 5415 19957
rect 8342 19954 8402 20028
rect 5349 19952 8402 19954
rect 5349 19896 5354 19952
rect 5410 19896 8402 19952
rect 5349 19894 8402 19896
rect 9397 19954 9463 19957
rect 14089 19954 14155 19957
rect 9397 19952 14155 19954
rect 9397 19896 9402 19952
rect 9458 19896 14094 19952
rect 14150 19896 14155 19952
rect 9397 19894 14155 19896
rect 5349 19891 5415 19894
rect 9397 19891 9463 19894
rect 14089 19891 14155 19894
rect 14273 19954 14339 19957
rect 14966 19954 15026 20030
rect 16941 20027 17007 20030
rect 17125 20027 17191 20030
rect 14273 19952 15026 19954
rect 14273 19896 14278 19952
rect 14334 19896 15026 19952
rect 14273 19894 15026 19896
rect 15101 19954 15167 19957
rect 16757 19954 16823 19957
rect 15101 19952 16823 19954
rect 15101 19896 15106 19952
rect 15162 19896 16762 19952
rect 16818 19896 16823 19952
rect 15101 19894 16823 19896
rect 14273 19891 14339 19894
rect 15101 19891 15167 19894
rect 16757 19891 16823 19894
rect 2313 19818 2379 19821
rect 2446 19818 2452 19820
rect 2313 19816 2452 19818
rect 2313 19760 2318 19816
rect 2374 19760 2452 19816
rect 2313 19758 2452 19760
rect 2313 19755 2379 19758
rect 2446 19756 2452 19758
rect 2516 19756 2522 19820
rect 2589 19818 2655 19821
rect 7373 19818 7439 19821
rect 2589 19816 7439 19818
rect 2589 19760 2594 19816
rect 2650 19760 7378 19816
rect 7434 19760 7439 19816
rect 2589 19758 7439 19760
rect 2589 19755 2655 19758
rect 7373 19755 7439 19758
rect 8518 19756 8524 19820
rect 8588 19818 8594 19820
rect 9305 19818 9371 19821
rect 8588 19816 9371 19818
rect 8588 19760 9310 19816
rect 9366 19760 9371 19816
rect 8588 19758 9371 19760
rect 8588 19756 8594 19758
rect 9305 19755 9371 19758
rect 11237 19818 11303 19821
rect 14406 19818 14412 19820
rect 11237 19816 14412 19818
rect 11237 19760 11242 19816
rect 11298 19760 14412 19816
rect 11237 19758 14412 19760
rect 11237 19755 11303 19758
rect 14406 19756 14412 19758
rect 14476 19756 14482 19820
rect 19558 19756 19564 19820
rect 19628 19818 19634 19820
rect 22093 19818 22159 19821
rect 19628 19816 22159 19818
rect 19628 19760 22098 19816
rect 22154 19760 22159 19816
rect 19628 19758 22159 19760
rect 19628 19756 19634 19758
rect 22093 19755 22159 19758
rect -300 19682 160 19712
rect 1945 19682 2011 19685
rect 5533 19682 5599 19685
rect -300 19622 1824 19682
rect -300 19592 160 19622
rect 1764 19546 1824 19622
rect 1945 19680 5599 19682
rect 1945 19624 1950 19680
rect 2006 19624 5538 19680
rect 5594 19624 5599 19680
rect 1945 19622 5599 19624
rect 1945 19619 2011 19622
rect 5533 19619 5599 19622
rect 7598 19620 7604 19684
rect 7668 19682 7674 19684
rect 9489 19682 9555 19685
rect 7668 19680 9555 19682
rect 7668 19624 9494 19680
rect 9550 19624 9555 19680
rect 7668 19622 9555 19624
rect 7668 19620 7674 19622
rect 9489 19619 9555 19622
rect 14089 19682 14155 19685
rect 15193 19682 15259 19685
rect 14089 19680 15259 19682
rect 14089 19624 14094 19680
rect 14150 19624 15198 19680
rect 15254 19624 15259 19680
rect 14089 19622 15259 19624
rect 14089 19619 14155 19622
rect 15193 19619 15259 19622
rect 18321 19682 18387 19685
rect 20069 19682 20135 19685
rect 18321 19680 20135 19682
rect 18321 19624 18326 19680
rect 18382 19624 20074 19680
rect 20130 19624 20135 19680
rect 18321 19622 20135 19624
rect 18321 19619 18387 19622
rect 20069 19619 20135 19622
rect 22185 19682 22251 19685
rect 22840 19682 23300 19712
rect 22185 19680 23300 19682
rect 22185 19624 22190 19680
rect 22246 19624 23300 19680
rect 22185 19622 23300 19624
rect 22185 19619 22251 19622
rect 6144 19616 6460 19617
rect 6144 19552 6150 19616
rect 6214 19552 6230 19616
rect 6294 19552 6310 19616
rect 6374 19552 6390 19616
rect 6454 19552 6460 19616
rect 6144 19551 6460 19552
rect 11342 19616 11658 19617
rect 11342 19552 11348 19616
rect 11412 19552 11428 19616
rect 11492 19552 11508 19616
rect 11572 19552 11588 19616
rect 11652 19552 11658 19616
rect 11342 19551 11658 19552
rect 16540 19616 16856 19617
rect 16540 19552 16546 19616
rect 16610 19552 16626 19616
rect 16690 19552 16706 19616
rect 16770 19552 16786 19616
rect 16850 19552 16856 19616
rect 16540 19551 16856 19552
rect 21738 19616 22054 19617
rect 21738 19552 21744 19616
rect 21808 19552 21824 19616
rect 21888 19552 21904 19616
rect 21968 19552 21984 19616
rect 22048 19552 22054 19616
rect 22840 19592 23300 19622
rect 21738 19551 22054 19552
rect 2773 19546 2839 19549
rect 1764 19544 2839 19546
rect 1764 19488 2778 19544
rect 2834 19488 2839 19544
rect 1764 19486 2839 19488
rect 2773 19483 2839 19486
rect 2998 19484 3004 19548
rect 3068 19546 3074 19548
rect 3325 19546 3391 19549
rect 3068 19544 3391 19546
rect 3068 19488 3330 19544
rect 3386 19488 3391 19544
rect 3068 19486 3391 19488
rect 3068 19484 3074 19486
rect 3325 19483 3391 19486
rect 4613 19546 4679 19549
rect 5022 19546 5028 19548
rect 4613 19544 5028 19546
rect 4613 19488 4618 19544
rect 4674 19488 5028 19544
rect 4613 19486 5028 19488
rect 4613 19483 4679 19486
rect 5022 19484 5028 19486
rect 5092 19484 5098 19548
rect 5257 19546 5323 19549
rect 9765 19546 9831 19549
rect 11053 19546 11119 19549
rect 5257 19544 5458 19546
rect 5257 19488 5262 19544
rect 5318 19488 5458 19544
rect 5257 19486 5458 19488
rect 5257 19483 5323 19486
rect -300 19410 160 19440
rect 3233 19410 3299 19413
rect -300 19408 3299 19410
rect -300 19352 3238 19408
rect 3294 19352 3299 19408
rect -300 19350 3299 19352
rect -300 19320 160 19350
rect 3233 19347 3299 19350
rect 5206 19348 5212 19412
rect 5276 19348 5282 19412
rect 2405 19274 2471 19277
rect 2405 19272 5090 19274
rect 2405 19216 2410 19272
rect 2466 19216 5090 19272
rect 2405 19214 5090 19216
rect 2405 19211 2471 19214
rect -300 19138 160 19168
rect 2865 19138 2931 19141
rect -300 19136 2931 19138
rect -300 19080 2870 19136
rect 2926 19080 2931 19136
rect -300 19078 2931 19080
rect -300 19048 160 19078
rect 2865 19075 2931 19078
rect 3545 19072 3861 19073
rect 3545 19008 3551 19072
rect 3615 19008 3631 19072
rect 3695 19008 3711 19072
rect 3775 19008 3791 19072
rect 3855 19008 3861 19072
rect 3545 19007 3861 19008
rect 1158 18940 1164 19004
rect 1228 19002 1234 19004
rect 3182 19002 3188 19004
rect 1228 18942 3188 19002
rect 1228 18940 1234 18942
rect 3182 18940 3188 18942
rect 3252 18940 3258 19004
rect 5030 19002 5090 19214
rect 5214 19138 5274 19348
rect 5398 19274 5458 19486
rect 9765 19544 11119 19546
rect 9765 19488 9770 19544
rect 9826 19488 11058 19544
rect 11114 19488 11119 19544
rect 9765 19486 11119 19488
rect 9765 19483 9831 19486
rect 11053 19483 11119 19486
rect 16990 19486 18338 19546
rect 11697 19410 11763 19413
rect 16990 19410 17050 19486
rect 11697 19408 17050 19410
rect 11697 19352 11702 19408
rect 11758 19352 17050 19408
rect 11697 19350 17050 19352
rect 11697 19347 11763 19350
rect 17718 19348 17724 19412
rect 17788 19410 17794 19412
rect 18137 19410 18203 19413
rect 17788 19408 18203 19410
rect 17788 19352 18142 19408
rect 18198 19352 18203 19408
rect 17788 19350 18203 19352
rect 18278 19410 18338 19486
rect 18689 19410 18755 19413
rect 18278 19408 18755 19410
rect 18278 19352 18694 19408
rect 18750 19352 18755 19408
rect 18278 19350 18755 19352
rect 17788 19348 17794 19350
rect 18137 19347 18203 19350
rect 18689 19347 18755 19350
rect 20846 19348 20852 19412
rect 20916 19410 20922 19412
rect 21357 19410 21423 19413
rect 20916 19408 21423 19410
rect 20916 19352 21362 19408
rect 21418 19352 21423 19408
rect 20916 19350 21423 19352
rect 20916 19348 20922 19350
rect 21357 19347 21423 19350
rect 17125 19274 17191 19277
rect 5398 19272 17191 19274
rect 5398 19216 17130 19272
rect 17186 19216 17191 19272
rect 5398 19214 17191 19216
rect 17125 19211 17191 19214
rect 18638 19212 18644 19276
rect 18708 19274 18714 19276
rect 19977 19274 20043 19277
rect 18708 19272 20043 19274
rect 18708 19216 19982 19272
rect 20038 19216 20043 19272
rect 18708 19214 20043 19216
rect 18708 19212 18714 19214
rect 19977 19211 20043 19214
rect 5942 19138 5948 19140
rect 5214 19078 5948 19138
rect 5942 19076 5948 19078
rect 6012 19076 6018 19140
rect 9765 19138 9831 19141
rect 12801 19138 12867 19141
rect 6134 19078 7068 19138
rect 5206 19002 5212 19004
rect 5030 18942 5212 19002
rect 5206 18940 5212 18942
rect 5276 19002 5282 19004
rect 6134 19002 6194 19078
rect 5276 18942 6194 19002
rect 7008 19002 7068 19078
rect 9765 19136 12867 19138
rect 9765 19080 9770 19136
rect 9826 19080 12806 19136
rect 12862 19080 12867 19136
rect 9765 19078 12867 19080
rect 9765 19075 9831 19078
rect 12801 19075 12867 19078
rect 21449 19138 21515 19141
rect 22840 19138 23300 19168
rect 21449 19136 23300 19138
rect 21449 19080 21454 19136
rect 21510 19080 23300 19136
rect 21449 19078 23300 19080
rect 21449 19075 21515 19078
rect 8743 19072 9059 19073
rect 8743 19008 8749 19072
rect 8813 19008 8829 19072
rect 8893 19008 8909 19072
rect 8973 19008 8989 19072
rect 9053 19008 9059 19072
rect 8743 19007 9059 19008
rect 13941 19072 14257 19073
rect 13941 19008 13947 19072
rect 14011 19008 14027 19072
rect 14091 19008 14107 19072
rect 14171 19008 14187 19072
rect 14251 19008 14257 19072
rect 13941 19007 14257 19008
rect 19139 19072 19455 19073
rect 19139 19008 19145 19072
rect 19209 19008 19225 19072
rect 19289 19008 19305 19072
rect 19369 19008 19385 19072
rect 19449 19008 19455 19072
rect 22840 19048 23300 19078
rect 19139 19007 19455 19008
rect 7833 19002 7899 19005
rect 13721 19002 13787 19005
rect 7008 19000 7899 19002
rect 7008 18944 7838 19000
rect 7894 18944 7899 19000
rect 7008 18942 7899 18944
rect 5276 18940 5282 18942
rect 7833 18939 7899 18942
rect 13678 19000 13787 19002
rect 13678 18944 13726 19000
rect 13782 18944 13787 19000
rect 13678 18939 13787 18944
rect -300 18866 160 18896
rect 1669 18866 1735 18869
rect 10225 18866 10291 18869
rect 11881 18866 11947 18869
rect -300 18806 1180 18866
rect -300 18776 160 18806
rect -300 18594 160 18624
rect 933 18594 999 18597
rect -300 18592 999 18594
rect -300 18536 938 18592
rect 994 18536 999 18592
rect -300 18534 999 18536
rect 1120 18594 1180 18806
rect 1669 18864 10291 18866
rect 1669 18808 1674 18864
rect 1730 18808 10230 18864
rect 10286 18808 10291 18864
rect 1669 18806 10291 18808
rect 1669 18803 1735 18806
rect 10225 18803 10291 18806
rect 11102 18864 11947 18866
rect 11102 18808 11886 18864
rect 11942 18808 11947 18864
rect 11102 18806 11947 18808
rect 4286 18668 4292 18732
rect 4356 18730 4362 18732
rect 5257 18730 5323 18733
rect 10869 18730 10935 18733
rect 4356 18728 5323 18730
rect 4356 18672 5262 18728
rect 5318 18672 5323 18728
rect 4356 18670 5323 18672
rect 4356 18668 4362 18670
rect 5257 18667 5323 18670
rect 7238 18728 10935 18730
rect 7238 18672 10874 18728
rect 10930 18672 10935 18728
rect 7238 18670 10935 18672
rect 1669 18594 1735 18597
rect 1120 18592 1735 18594
rect 1120 18536 1674 18592
rect 1730 18536 1735 18592
rect 1120 18534 1735 18536
rect -300 18504 160 18534
rect 933 18531 999 18534
rect 1669 18531 1735 18534
rect 6637 18594 6703 18597
rect 7046 18594 7052 18596
rect 6637 18592 7052 18594
rect 6637 18536 6642 18592
rect 6698 18536 7052 18592
rect 6637 18534 7052 18536
rect 6637 18531 6703 18534
rect 7046 18532 7052 18534
rect 7116 18532 7122 18596
rect 6144 18528 6460 18529
rect 6144 18464 6150 18528
rect 6214 18464 6230 18528
rect 6294 18464 6310 18528
rect 6374 18464 6390 18528
rect 6454 18464 6460 18528
rect 6144 18463 6460 18464
rect 7097 18458 7163 18461
rect 7238 18460 7298 18670
rect 10869 18667 10935 18670
rect 9949 18594 10015 18597
rect 10542 18594 10548 18596
rect 9949 18592 10548 18594
rect 9949 18536 9954 18592
rect 10010 18536 10548 18592
rect 9949 18534 10548 18536
rect 9949 18531 10015 18534
rect 10542 18532 10548 18534
rect 10612 18532 10618 18596
rect 7230 18458 7236 18460
rect 7097 18456 7236 18458
rect 7097 18400 7102 18456
rect 7158 18400 7236 18456
rect 7097 18398 7236 18400
rect 7097 18395 7163 18398
rect 7230 18396 7236 18398
rect 7300 18396 7306 18460
rect 7833 18458 7899 18461
rect 11102 18458 11162 18806
rect 11881 18803 11947 18806
rect 11605 18730 11671 18733
rect 12065 18730 12131 18733
rect 11605 18728 12131 18730
rect 11605 18672 11610 18728
rect 11666 18672 12070 18728
rect 12126 18672 12131 18728
rect 11605 18670 12131 18672
rect 13678 18730 13738 18939
rect 14641 18866 14707 18869
rect 16062 18866 16068 18868
rect 14641 18864 16068 18866
rect 14641 18808 14646 18864
rect 14702 18808 16068 18864
rect 14641 18806 16068 18808
rect 14641 18803 14707 18806
rect 16062 18804 16068 18806
rect 16132 18804 16138 18868
rect 18086 18730 18092 18732
rect 13678 18670 18092 18730
rect 11605 18667 11671 18670
rect 12065 18667 12131 18670
rect 18086 18668 18092 18670
rect 18156 18668 18162 18732
rect 22185 18594 22251 18597
rect 22840 18594 23300 18624
rect 22185 18592 23300 18594
rect 22185 18536 22190 18592
rect 22246 18536 23300 18592
rect 22185 18534 23300 18536
rect 22185 18531 22251 18534
rect 11342 18528 11658 18529
rect 11342 18464 11348 18528
rect 11412 18464 11428 18528
rect 11492 18464 11508 18528
rect 11572 18464 11588 18528
rect 11652 18464 11658 18528
rect 11342 18463 11658 18464
rect 16540 18528 16856 18529
rect 16540 18464 16546 18528
rect 16610 18464 16626 18528
rect 16690 18464 16706 18528
rect 16770 18464 16786 18528
rect 16850 18464 16856 18528
rect 16540 18463 16856 18464
rect 21738 18528 22054 18529
rect 21738 18464 21744 18528
rect 21808 18464 21824 18528
rect 21888 18464 21904 18528
rect 21968 18464 21984 18528
rect 22048 18464 22054 18528
rect 22840 18504 23300 18534
rect 21738 18463 22054 18464
rect 7833 18456 11162 18458
rect 7833 18400 7838 18456
rect 7894 18400 11162 18456
rect 7833 18398 11162 18400
rect 11881 18458 11947 18461
rect 16113 18458 16179 18461
rect 11881 18456 16179 18458
rect 11881 18400 11886 18456
rect 11942 18400 16118 18456
rect 16174 18400 16179 18456
rect 11881 18398 16179 18400
rect 7833 18395 7899 18398
rect 11881 18395 11947 18398
rect 16113 18395 16179 18398
rect -300 18322 160 18352
rect 1853 18322 1919 18325
rect -300 18320 1919 18322
rect -300 18264 1858 18320
rect 1914 18264 1919 18320
rect -300 18262 1919 18264
rect -300 18232 160 18262
rect 1853 18259 1919 18262
rect 4061 18322 4127 18325
rect 7189 18322 7255 18325
rect 4061 18320 7255 18322
rect 4061 18264 4066 18320
rect 4122 18264 7194 18320
rect 7250 18264 7255 18320
rect 4061 18262 7255 18264
rect 4061 18259 4127 18262
rect 7189 18259 7255 18262
rect 8150 18260 8156 18324
rect 8220 18322 8226 18324
rect 12525 18322 12591 18325
rect 8220 18320 12591 18322
rect 8220 18264 12530 18320
rect 12586 18264 12591 18320
rect 8220 18262 12591 18264
rect 8220 18260 8226 18262
rect 12525 18259 12591 18262
rect 13353 18322 13419 18325
rect 17217 18322 17283 18325
rect 13353 18320 17283 18322
rect 13353 18264 13358 18320
rect 13414 18264 17222 18320
rect 17278 18264 17283 18320
rect 13353 18262 17283 18264
rect 13353 18259 13419 18262
rect 17217 18259 17283 18262
rect 2497 18186 2563 18189
rect 5441 18186 5507 18189
rect 2497 18184 5507 18186
rect 2497 18128 2502 18184
rect 2558 18128 5446 18184
rect 5502 18128 5507 18184
rect 2497 18126 5507 18128
rect 2497 18123 2563 18126
rect 5441 18123 5507 18126
rect 5717 18186 5783 18189
rect 7097 18186 7163 18189
rect 11145 18186 11211 18189
rect 5717 18184 6976 18186
rect 5717 18128 5722 18184
rect 5778 18128 6976 18184
rect 5717 18126 6976 18128
rect 5717 18123 5783 18126
rect -300 18050 160 18080
rect 1485 18050 1551 18053
rect -300 18048 1551 18050
rect -300 17992 1490 18048
rect 1546 17992 1551 18048
rect -300 17990 1551 17992
rect -300 17960 160 17990
rect 1485 17987 1551 17990
rect 2773 18050 2839 18053
rect 2773 18048 2882 18050
rect 2773 17992 2778 18048
rect 2834 17992 2882 18048
rect 2773 17987 2882 17992
rect 6678 17988 6684 18052
rect 6748 17988 6754 18052
rect 6916 18050 6976 18126
rect 7097 18184 11211 18186
rect 7097 18128 7102 18184
rect 7158 18128 11150 18184
rect 11206 18128 11211 18184
rect 7097 18126 11211 18128
rect 7097 18123 7163 18126
rect 11145 18123 11211 18126
rect 16205 18186 16271 18189
rect 16982 18186 16988 18188
rect 16205 18184 16988 18186
rect 16205 18128 16210 18184
rect 16266 18128 16988 18184
rect 16205 18126 16988 18128
rect 16205 18123 16271 18126
rect 16982 18124 16988 18126
rect 17052 18124 17058 18188
rect 8569 18050 8635 18053
rect 6916 18048 8635 18050
rect 6916 17992 8574 18048
rect 8630 17992 8635 18048
rect 6916 17990 8635 17992
rect 1577 17914 1643 17917
rect 798 17912 1643 17914
rect 798 17856 1582 17912
rect 1638 17856 1643 17912
rect 798 17854 1643 17856
rect -300 17778 160 17808
rect 798 17778 858 17854
rect 1577 17851 1643 17854
rect 1853 17914 1919 17917
rect 2681 17914 2747 17917
rect 1853 17912 2747 17914
rect 1853 17856 1858 17912
rect 1914 17856 2686 17912
rect 2742 17856 2747 17912
rect 1853 17854 2747 17856
rect 2822 17914 2882 17987
rect 3545 17984 3861 17985
rect 3545 17920 3551 17984
rect 3615 17920 3631 17984
rect 3695 17920 3711 17984
rect 3775 17920 3791 17984
rect 3855 17920 3861 17984
rect 3545 17919 3861 17920
rect 4061 17916 4127 17917
rect 3366 17914 3372 17916
rect 2822 17854 3372 17914
rect 1853 17851 1919 17854
rect 2681 17851 2747 17854
rect 3366 17852 3372 17854
rect 3436 17852 3442 17916
rect 4061 17914 4108 17916
rect 4016 17912 4108 17914
rect 4016 17856 4066 17912
rect 4016 17854 4108 17856
rect 4061 17852 4108 17854
rect 4172 17852 4178 17916
rect 4889 17914 4955 17917
rect 5441 17914 5507 17917
rect 6177 17914 6243 17917
rect 4889 17912 6243 17914
rect 4889 17856 4894 17912
rect 4950 17856 5446 17912
rect 5502 17856 6182 17912
rect 6238 17856 6243 17912
rect 4889 17854 6243 17856
rect 4061 17851 4127 17852
rect 4889 17851 4955 17854
rect 5441 17851 5507 17854
rect 6177 17851 6243 17854
rect -300 17718 858 17778
rect 2773 17778 2839 17781
rect 4337 17778 4403 17781
rect 2773 17776 4403 17778
rect 2773 17720 2778 17776
rect 2834 17720 4342 17776
rect 4398 17720 4403 17776
rect 2773 17718 4403 17720
rect 6686 17778 6746 17988
rect 8569 17987 8635 17990
rect 10685 18050 10751 18053
rect 13721 18050 13787 18053
rect 10685 18048 13787 18050
rect 10685 17992 10690 18048
rect 10746 17992 13726 18048
rect 13782 17992 13787 18048
rect 10685 17990 13787 17992
rect 10685 17987 10751 17990
rect 13721 17987 13787 17990
rect 16246 17988 16252 18052
rect 16316 18050 16322 18052
rect 16982 18050 16988 18052
rect 16316 17990 16988 18050
rect 16316 17988 16322 17990
rect 16982 17988 16988 17990
rect 17052 17988 17058 18052
rect 21449 18050 21515 18053
rect 22840 18050 23300 18080
rect 21449 18048 23300 18050
rect 21449 17992 21454 18048
rect 21510 17992 23300 18048
rect 21449 17990 23300 17992
rect 21449 17987 21515 17990
rect 8743 17984 9059 17985
rect 8743 17920 8749 17984
rect 8813 17920 8829 17984
rect 8893 17920 8909 17984
rect 8973 17920 8989 17984
rect 9053 17920 9059 17984
rect 8743 17919 9059 17920
rect 13941 17984 14257 17985
rect 13941 17920 13947 17984
rect 14011 17920 14027 17984
rect 14091 17920 14107 17984
rect 14171 17920 14187 17984
rect 14251 17920 14257 17984
rect 13941 17919 14257 17920
rect 19139 17984 19455 17985
rect 19139 17920 19145 17984
rect 19209 17920 19225 17984
rect 19289 17920 19305 17984
rect 19369 17920 19385 17984
rect 19449 17920 19455 17984
rect 22840 17960 23300 17990
rect 19139 17919 19455 17920
rect 7005 17914 7071 17917
rect 9213 17914 9279 17917
rect 9438 17914 9444 17916
rect 7005 17912 8632 17914
rect 7005 17856 7010 17912
rect 7066 17856 8632 17912
rect 7005 17854 8632 17856
rect 7005 17851 7071 17854
rect 8385 17778 8451 17781
rect 6686 17776 8451 17778
rect 6686 17720 8390 17776
rect 8446 17720 8451 17776
rect 6686 17718 8451 17720
rect 8572 17778 8632 17854
rect 9213 17912 9444 17914
rect 9213 17856 9218 17912
rect 9274 17856 9444 17912
rect 9213 17854 9444 17856
rect 9213 17851 9279 17854
rect 9438 17852 9444 17854
rect 9508 17852 9514 17916
rect 9581 17778 9647 17781
rect 8572 17776 9647 17778
rect 8572 17720 9586 17776
rect 9642 17720 9647 17776
rect 8572 17718 9647 17720
rect -300 17688 160 17718
rect 2773 17715 2839 17718
rect 4337 17715 4403 17718
rect 8385 17715 8451 17718
rect 9581 17715 9647 17718
rect 12801 17778 12867 17781
rect 12934 17778 12940 17780
rect 12801 17776 12940 17778
rect 12801 17720 12806 17776
rect 12862 17720 12940 17776
rect 12801 17718 12940 17720
rect 12801 17715 12867 17718
rect 12934 17716 12940 17718
rect 13004 17716 13010 17780
rect 15878 17716 15884 17780
rect 15948 17778 15954 17780
rect 19701 17778 19767 17781
rect 15948 17776 19767 17778
rect 15948 17720 19706 17776
rect 19762 17720 19767 17776
rect 15948 17718 19767 17720
rect 15948 17716 15954 17718
rect 19701 17715 19767 17718
rect 473 17642 539 17645
rect 1526 17642 1532 17644
rect 473 17640 1532 17642
rect 473 17584 478 17640
rect 534 17584 1532 17640
rect 473 17582 1532 17584
rect 473 17579 539 17582
rect 1526 17580 1532 17582
rect 1596 17580 1602 17644
rect 2129 17642 2195 17645
rect 3509 17642 3575 17645
rect 7005 17642 7071 17645
rect 8569 17642 8635 17645
rect 11237 17642 11303 17645
rect 2129 17640 6746 17642
rect 2129 17584 2134 17640
rect 2190 17584 3514 17640
rect 3570 17584 6746 17640
rect 2129 17582 6746 17584
rect 2129 17579 2195 17582
rect 3509 17579 3575 17582
rect -300 17506 160 17536
rect 4838 17506 4844 17508
rect -300 17446 858 17506
rect -300 17416 160 17446
rect 798 17370 858 17446
rect 2822 17446 4844 17506
rect 1301 17370 1367 17373
rect 2681 17372 2747 17373
rect 2822 17372 2882 17446
rect 4838 17444 4844 17446
rect 4908 17506 4914 17508
rect 4981 17506 5047 17509
rect 4908 17504 5047 17506
rect 4908 17448 4986 17504
rect 5042 17448 5047 17504
rect 4908 17446 5047 17448
rect 4908 17444 4914 17446
rect 4981 17443 5047 17446
rect 6144 17440 6460 17441
rect 6144 17376 6150 17440
rect 6214 17376 6230 17440
rect 6294 17376 6310 17440
rect 6374 17376 6390 17440
rect 6454 17376 6460 17440
rect 6144 17375 6460 17376
rect 2630 17370 2636 17372
rect 798 17368 1367 17370
rect 798 17312 1306 17368
rect 1362 17312 1367 17368
rect 798 17310 1367 17312
rect 2590 17310 2636 17370
rect 2700 17368 2747 17372
rect 2742 17312 2747 17368
rect 1301 17307 1367 17310
rect 2630 17308 2636 17310
rect 2700 17308 2747 17312
rect 2814 17308 2820 17372
rect 2884 17308 2890 17372
rect 3918 17308 3924 17372
rect 3988 17370 3994 17372
rect 4153 17370 4219 17373
rect 3988 17368 4219 17370
rect 3988 17312 4158 17368
rect 4214 17312 4219 17368
rect 3988 17310 4219 17312
rect 6686 17370 6746 17582
rect 7005 17640 7804 17642
rect 7005 17584 7010 17640
rect 7066 17584 7804 17640
rect 7005 17582 7804 17584
rect 7005 17579 7071 17582
rect 7373 17506 7439 17509
rect 7598 17506 7604 17508
rect 7373 17504 7604 17506
rect 7373 17448 7378 17504
rect 7434 17448 7604 17504
rect 7373 17446 7604 17448
rect 7373 17443 7439 17446
rect 7598 17444 7604 17446
rect 7668 17444 7674 17508
rect 7744 17506 7804 17582
rect 8569 17640 11303 17642
rect 8569 17584 8574 17640
rect 8630 17584 11242 17640
rect 11298 17584 11303 17640
rect 8569 17582 11303 17584
rect 8569 17579 8635 17582
rect 11237 17579 11303 17582
rect 14733 17642 14799 17645
rect 14958 17642 14964 17644
rect 14733 17640 14964 17642
rect 14733 17584 14738 17640
rect 14794 17584 14964 17640
rect 14733 17582 14964 17584
rect 14733 17579 14799 17582
rect 14958 17580 14964 17582
rect 15028 17642 15034 17644
rect 15653 17642 15719 17645
rect 15028 17640 15719 17642
rect 15028 17584 15658 17640
rect 15714 17584 15719 17640
rect 15028 17582 15719 17584
rect 15028 17580 15034 17582
rect 15653 17579 15719 17582
rect 8753 17506 8819 17509
rect 7744 17504 8819 17506
rect 7744 17448 8758 17504
rect 8814 17448 8819 17504
rect 7744 17446 8819 17448
rect 8753 17443 8819 17446
rect 9949 17506 10015 17509
rect 10726 17506 10732 17508
rect 9949 17504 10732 17506
rect 9949 17448 9954 17504
rect 10010 17448 10732 17504
rect 9949 17446 10732 17448
rect 9949 17443 10015 17446
rect 10726 17444 10732 17446
rect 10796 17444 10802 17508
rect 14406 17444 14412 17508
rect 14476 17506 14482 17508
rect 15142 17506 15148 17508
rect 14476 17446 15148 17506
rect 14476 17444 14482 17446
rect 15142 17444 15148 17446
rect 15212 17444 15218 17508
rect 22185 17506 22251 17509
rect 22840 17506 23300 17536
rect 22185 17504 23300 17506
rect 22185 17448 22190 17504
rect 22246 17448 23300 17504
rect 22185 17446 23300 17448
rect 22185 17443 22251 17446
rect 11342 17440 11658 17441
rect 11342 17376 11348 17440
rect 11412 17376 11428 17440
rect 11492 17376 11508 17440
rect 11572 17376 11588 17440
rect 11652 17376 11658 17440
rect 11342 17375 11658 17376
rect 16540 17440 16856 17441
rect 16540 17376 16546 17440
rect 16610 17376 16626 17440
rect 16690 17376 16706 17440
rect 16770 17376 16786 17440
rect 16850 17376 16856 17440
rect 16540 17375 16856 17376
rect 21738 17440 22054 17441
rect 21738 17376 21744 17440
rect 21808 17376 21824 17440
rect 21888 17376 21904 17440
rect 21968 17376 21984 17440
rect 22048 17376 22054 17440
rect 22840 17416 23300 17446
rect 21738 17375 22054 17376
rect 11145 17370 11211 17373
rect 6686 17368 11211 17370
rect 6686 17312 11150 17368
rect 11206 17312 11211 17368
rect 6686 17310 11211 17312
rect 3988 17308 3994 17310
rect 2681 17307 2747 17308
rect 4153 17307 4219 17310
rect 11145 17307 11211 17310
rect 13670 17308 13676 17372
rect 13740 17370 13746 17372
rect 15101 17370 15167 17373
rect 13740 17368 15167 17370
rect 13740 17312 15106 17368
rect 15162 17312 15167 17368
rect 13740 17310 15167 17312
rect 13740 17308 13746 17310
rect 15101 17307 15167 17310
rect -300 17234 160 17264
rect 1945 17234 2011 17237
rect 15009 17234 15075 17237
rect 21265 17236 21331 17237
rect -300 17174 1456 17234
rect -300 17144 160 17174
rect 1396 17098 1456 17174
rect 1945 17232 15075 17234
rect 1945 17176 1950 17232
rect 2006 17176 15014 17232
rect 15070 17176 15075 17232
rect 1945 17174 15075 17176
rect 1945 17171 2011 17174
rect 15009 17171 15075 17174
rect 21214 17172 21220 17236
rect 21284 17234 21331 17236
rect 21284 17232 21376 17234
rect 21326 17176 21376 17232
rect 21284 17174 21376 17176
rect 21284 17172 21331 17174
rect 21265 17171 21331 17172
rect 3877 17098 3943 17101
rect 1396 17096 3943 17098
rect 1396 17040 3882 17096
rect 3938 17040 3943 17096
rect 1396 17038 3943 17040
rect 3877 17035 3943 17038
rect 4061 17098 4127 17101
rect 11145 17098 11211 17101
rect 4061 17096 11211 17098
rect 4061 17040 4066 17096
rect 4122 17040 11150 17096
rect 11206 17040 11211 17096
rect 4061 17038 11211 17040
rect 4061 17035 4127 17038
rect 11145 17035 11211 17038
rect 13486 17036 13492 17100
rect 13556 17098 13562 17100
rect 14733 17098 14799 17101
rect 13556 17096 14799 17098
rect 13556 17040 14738 17096
rect 14794 17040 14799 17096
rect 13556 17038 14799 17040
rect 13556 17036 13562 17038
rect 14733 17035 14799 17038
rect -300 16962 160 16992
rect 1761 16962 1827 16965
rect -300 16960 1827 16962
rect -300 16904 1766 16960
rect 1822 16904 1827 16960
rect -300 16902 1827 16904
rect -300 16872 160 16902
rect 1761 16899 1827 16902
rect 16757 16962 16823 16965
rect 17677 16962 17743 16965
rect 16757 16960 17743 16962
rect 16757 16904 16762 16960
rect 16818 16904 17682 16960
rect 17738 16904 17743 16960
rect 16757 16902 17743 16904
rect 16757 16899 16823 16902
rect 17677 16899 17743 16902
rect 17953 16960 18019 16965
rect 17953 16904 17958 16960
rect 18014 16904 18019 16960
rect 17953 16899 18019 16904
rect 21449 16962 21515 16965
rect 22840 16962 23300 16992
rect 21449 16960 23300 16962
rect 21449 16904 21454 16960
rect 21510 16904 23300 16960
rect 21449 16902 23300 16904
rect 21449 16899 21515 16902
rect 3545 16896 3861 16897
rect 3545 16832 3551 16896
rect 3615 16832 3631 16896
rect 3695 16832 3711 16896
rect 3775 16832 3791 16896
rect 3855 16832 3861 16896
rect 3545 16831 3861 16832
rect 8743 16896 9059 16897
rect 8743 16832 8749 16896
rect 8813 16832 8829 16896
rect 8893 16832 8909 16896
rect 8973 16832 8989 16896
rect 9053 16832 9059 16896
rect 8743 16831 9059 16832
rect 13941 16896 14257 16897
rect 13941 16832 13947 16896
rect 14011 16832 14027 16896
rect 14091 16832 14107 16896
rect 14171 16832 14187 16896
rect 14251 16832 14257 16896
rect 13941 16831 14257 16832
rect 2313 16828 2379 16829
rect 790 16764 796 16828
rect 860 16826 866 16828
rect 1894 16826 1900 16828
rect 860 16766 1900 16826
rect 860 16764 866 16766
rect 1894 16764 1900 16766
rect 1964 16764 1970 16828
rect 2262 16826 2268 16828
rect 2222 16766 2268 16826
rect 2332 16826 2379 16828
rect 3417 16826 3483 16829
rect 2332 16824 3483 16826
rect 2374 16768 3422 16824
rect 3478 16768 3483 16824
rect 2262 16764 2268 16766
rect 2332 16766 3483 16768
rect 2332 16764 2379 16766
rect 2313 16763 2379 16764
rect 3417 16763 3483 16766
rect 4521 16826 4587 16829
rect 10685 16826 10751 16829
rect 10961 16826 11027 16829
rect 4521 16824 8218 16826
rect 4521 16768 4526 16824
rect 4582 16768 8218 16824
rect 4521 16766 8218 16768
rect 4521 16763 4587 16766
rect -300 16690 160 16720
rect 3601 16690 3667 16693
rect -300 16688 3667 16690
rect -300 16632 3606 16688
rect 3662 16632 3667 16688
rect -300 16630 3667 16632
rect -300 16600 160 16630
rect 3601 16627 3667 16630
rect 4102 16628 4108 16692
rect 4172 16690 4178 16692
rect 5901 16690 5967 16693
rect 8158 16692 8218 16766
rect 10685 16824 11027 16826
rect 10685 16768 10690 16824
rect 10746 16768 10966 16824
rect 11022 16768 11027 16824
rect 10685 16766 11027 16768
rect 10685 16763 10751 16766
rect 10961 16763 11027 16766
rect 15285 16826 15351 16829
rect 17956 16826 18016 16899
rect 19139 16896 19455 16897
rect 19139 16832 19145 16896
rect 19209 16832 19225 16896
rect 19289 16832 19305 16896
rect 19369 16832 19385 16896
rect 19449 16832 19455 16896
rect 22840 16872 23300 16902
rect 19139 16831 19455 16832
rect 15285 16824 18016 16826
rect 15285 16768 15290 16824
rect 15346 16768 18016 16824
rect 15285 16766 18016 16768
rect 15285 16763 15351 16766
rect 10501 16692 10567 16693
rect 4172 16688 5967 16690
rect 4172 16632 5906 16688
rect 5962 16632 5967 16688
rect 4172 16630 5967 16632
rect 4172 16628 4178 16630
rect 5901 16627 5967 16630
rect 8150 16628 8156 16692
rect 8220 16628 8226 16692
rect 10501 16688 10548 16692
rect 10612 16690 10618 16692
rect 10501 16632 10506 16688
rect 10501 16628 10548 16632
rect 10612 16630 10658 16690
rect 10612 16628 10618 16630
rect 10910 16628 10916 16692
rect 10980 16690 10986 16692
rect 10980 16628 11024 16690
rect 14590 16628 14596 16692
rect 14660 16690 14666 16692
rect 14733 16690 14799 16693
rect 14660 16688 14799 16690
rect 14660 16632 14738 16688
rect 14794 16632 14799 16688
rect 14660 16630 14799 16632
rect 14660 16628 14666 16630
rect 10501 16627 10567 16628
rect 3366 16492 3372 16556
rect 3436 16554 3442 16556
rect 6862 16554 6868 16556
rect 3436 16494 6868 16554
rect 3436 16492 3442 16494
rect 6862 16492 6868 16494
rect 6932 16492 6938 16556
rect 9673 16554 9739 16557
rect 10174 16554 10180 16556
rect 9673 16552 10180 16554
rect 9673 16496 9678 16552
rect 9734 16496 10180 16552
rect 9673 16494 10180 16496
rect 9673 16491 9739 16494
rect 10174 16492 10180 16494
rect 10244 16492 10250 16556
rect 10964 16554 11024 16628
rect 14733 16627 14799 16630
rect 14774 16554 14780 16556
rect 10964 16494 14780 16554
rect 14774 16492 14780 16494
rect 14844 16492 14850 16556
rect 18781 16554 18847 16557
rect 19793 16554 19859 16557
rect 18781 16552 19859 16554
rect 18781 16496 18786 16552
rect 18842 16496 19798 16552
rect 19854 16496 19859 16552
rect 18781 16494 19859 16496
rect 18781 16491 18847 16494
rect 19793 16491 19859 16494
rect 21449 16554 21515 16557
rect 21449 16552 22202 16554
rect 21449 16496 21454 16552
rect 21510 16496 22202 16552
rect 21449 16494 22202 16496
rect 21449 16491 21515 16494
rect -300 16418 160 16448
rect 3969 16418 4035 16421
rect -300 16416 4035 16418
rect -300 16360 3974 16416
rect 4030 16360 4035 16416
rect -300 16358 4035 16360
rect -300 16328 160 16358
rect 3969 16355 4035 16358
rect 4889 16418 4955 16421
rect 5533 16418 5599 16421
rect 4889 16416 5599 16418
rect 4889 16360 4894 16416
rect 4950 16360 5538 16416
rect 5594 16360 5599 16416
rect 4889 16358 5599 16360
rect 22142 16418 22202 16494
rect 22840 16418 23300 16448
rect 22142 16358 23300 16418
rect 4889 16355 4955 16358
rect 5533 16355 5599 16358
rect 6144 16352 6460 16353
rect 6144 16288 6150 16352
rect 6214 16288 6230 16352
rect 6294 16288 6310 16352
rect 6374 16288 6390 16352
rect 6454 16288 6460 16352
rect 6144 16287 6460 16288
rect 11342 16352 11658 16353
rect 11342 16288 11348 16352
rect 11412 16288 11428 16352
rect 11492 16288 11508 16352
rect 11572 16288 11588 16352
rect 11652 16288 11658 16352
rect 11342 16287 11658 16288
rect 16540 16352 16856 16353
rect 16540 16288 16546 16352
rect 16610 16288 16626 16352
rect 16690 16288 16706 16352
rect 16770 16288 16786 16352
rect 16850 16288 16856 16352
rect 16540 16287 16856 16288
rect 21738 16352 22054 16353
rect 21738 16288 21744 16352
rect 21808 16288 21824 16352
rect 21888 16288 21904 16352
rect 21968 16288 21984 16352
rect 22048 16288 22054 16352
rect 22840 16328 23300 16358
rect 21738 16287 22054 16288
rect 10910 16220 10916 16284
rect 10980 16282 10986 16284
rect 11053 16282 11119 16285
rect 10980 16280 11119 16282
rect 10980 16224 11058 16280
rect 11114 16224 11119 16280
rect 10980 16222 11119 16224
rect 10980 16220 10986 16222
rect 11053 16219 11119 16222
rect -300 16146 160 16176
rect 238 16146 244 16148
rect -300 16086 244 16146
rect -300 16056 160 16086
rect 238 16084 244 16086
rect 308 16084 314 16148
rect 1710 16084 1716 16148
rect 1780 16146 1786 16148
rect 4705 16146 4771 16149
rect 1780 16144 4771 16146
rect 1780 16088 4710 16144
rect 4766 16088 4771 16144
rect 1780 16086 4771 16088
rect 1780 16084 1786 16086
rect 4705 16083 4771 16086
rect 5390 16084 5396 16148
rect 5460 16146 5466 16148
rect 8109 16146 8175 16149
rect 5460 16144 8175 16146
rect 5460 16088 8114 16144
rect 8170 16088 8175 16144
rect 5460 16086 8175 16088
rect 5460 16084 5466 16086
rect 8109 16083 8175 16086
rect 9121 16146 9187 16149
rect 11830 16146 11836 16148
rect 9121 16144 11836 16146
rect 9121 16088 9126 16144
rect 9182 16088 11836 16144
rect 9121 16086 11836 16088
rect 9121 16083 9187 16086
rect 11830 16084 11836 16086
rect 11900 16084 11906 16148
rect 12617 16144 12683 16149
rect 12617 16088 12622 16144
rect 12678 16088 12683 16144
rect 12617 16083 12683 16088
rect 3049 16010 3115 16013
rect 3049 16008 5504 16010
rect 3049 15952 3054 16008
rect 3110 15952 5504 16008
rect 3049 15950 5504 15952
rect 3049 15947 3115 15950
rect -300 15874 160 15904
rect 1577 15874 1643 15877
rect 4889 15876 4955 15877
rect -300 15872 1643 15874
rect -300 15816 1582 15872
rect 1638 15816 1643 15872
rect -300 15814 1643 15816
rect -300 15784 160 15814
rect 1577 15811 1643 15814
rect 4838 15812 4844 15876
rect 4908 15874 4955 15876
rect 4908 15872 5000 15874
rect 4950 15816 5000 15872
rect 4908 15814 5000 15816
rect 4908 15812 4955 15814
rect 4889 15811 4955 15812
rect 3545 15808 3861 15809
rect 3545 15744 3551 15808
rect 3615 15744 3631 15808
rect 3695 15744 3711 15808
rect 3775 15744 3791 15808
rect 3855 15744 3861 15808
rect 3545 15743 3861 15744
rect 1485 15738 1551 15741
rect 982 15736 1551 15738
rect 982 15680 1490 15736
rect 1546 15680 1551 15736
rect 982 15678 1551 15680
rect -300 15602 160 15632
rect 982 15602 1042 15678
rect 1485 15675 1551 15678
rect 4102 15676 4108 15740
rect 4172 15738 4178 15740
rect 4889 15738 4955 15741
rect 4172 15736 4955 15738
rect 4172 15680 4894 15736
rect 4950 15680 4955 15736
rect 4172 15678 4955 15680
rect 5444 15738 5504 15950
rect 7782 15948 7788 16012
rect 7852 16010 7858 16012
rect 12620 16010 12680 16083
rect 7852 15950 12680 16010
rect 7852 15948 7858 15950
rect 19006 15948 19012 16012
rect 19076 16010 19082 16012
rect 19241 16010 19307 16013
rect 19076 16008 19307 16010
rect 19076 15952 19246 16008
rect 19302 15952 19307 16008
rect 19076 15950 19307 15952
rect 19076 15948 19082 15950
rect 19241 15947 19307 15950
rect 9581 15874 9647 15877
rect 13670 15874 13676 15876
rect 9581 15872 13676 15874
rect 9581 15816 9586 15872
rect 9642 15816 13676 15872
rect 9581 15814 13676 15816
rect 9581 15811 9647 15814
rect 13670 15812 13676 15814
rect 13740 15812 13746 15876
rect 21449 15874 21515 15877
rect 22840 15874 23300 15904
rect 21449 15872 23300 15874
rect 21449 15816 21454 15872
rect 21510 15816 23300 15872
rect 21449 15814 23300 15816
rect 21449 15811 21515 15814
rect 8743 15808 9059 15809
rect 8743 15744 8749 15808
rect 8813 15744 8829 15808
rect 8893 15744 8909 15808
rect 8973 15744 8989 15808
rect 9053 15744 9059 15808
rect 8743 15743 9059 15744
rect 13941 15808 14257 15809
rect 13941 15744 13947 15808
rect 14011 15744 14027 15808
rect 14091 15744 14107 15808
rect 14171 15744 14187 15808
rect 14251 15744 14257 15808
rect 13941 15743 14257 15744
rect 19139 15808 19455 15809
rect 19139 15744 19145 15808
rect 19209 15744 19225 15808
rect 19289 15744 19305 15808
rect 19369 15744 19385 15808
rect 19449 15744 19455 15808
rect 22840 15784 23300 15814
rect 19139 15743 19455 15744
rect 6678 15738 6684 15740
rect 5444 15678 6684 15738
rect 4172 15676 4178 15678
rect 4889 15675 4955 15678
rect 6678 15676 6684 15678
rect 6748 15676 6754 15740
rect 4521 15604 4587 15605
rect -300 15542 1042 15602
rect -300 15512 160 15542
rect 4470 15540 4476 15604
rect 4540 15602 4587 15604
rect 4540 15600 4632 15602
rect 4582 15544 4632 15600
rect 4540 15542 4632 15544
rect 4540 15540 4587 15542
rect 7046 15540 7052 15604
rect 7116 15602 7122 15604
rect 7189 15602 7255 15605
rect 16297 15604 16363 15605
rect 7116 15600 7255 15602
rect 7116 15544 7194 15600
rect 7250 15544 7255 15600
rect 7116 15542 7255 15544
rect 7116 15540 7122 15542
rect 4521 15539 4587 15540
rect 7189 15539 7255 15542
rect 10174 15540 10180 15604
rect 10244 15602 10250 15604
rect 16246 15602 16252 15604
rect 10244 15542 16252 15602
rect 16316 15602 16363 15604
rect 16316 15600 16444 15602
rect 16358 15544 16444 15600
rect 10244 15540 10250 15542
rect 16246 15540 16252 15542
rect 16316 15542 16444 15544
rect 16316 15540 16363 15542
rect 16297 15539 16363 15540
rect 1894 15404 1900 15468
rect 1964 15466 1970 15468
rect 5758 15466 5764 15468
rect 1964 15406 5764 15466
rect 1964 15404 1970 15406
rect 5758 15404 5764 15406
rect 5828 15404 5834 15468
rect 12433 15466 12499 15469
rect 13261 15466 13327 15469
rect 18689 15466 18755 15469
rect 12433 15464 18755 15466
rect 12433 15408 12438 15464
rect 12494 15408 13266 15464
rect 13322 15408 18694 15464
rect 18750 15408 18755 15464
rect 12433 15406 18755 15408
rect 12433 15403 12499 15406
rect 13261 15403 13327 15406
rect 18689 15403 18755 15406
rect -300 15330 160 15360
rect 2129 15330 2195 15333
rect 4613 15330 4679 15333
rect 5993 15330 6059 15333
rect -300 15270 1640 15330
rect -300 15240 160 15270
rect 790 15132 796 15196
rect 860 15194 866 15196
rect 1393 15194 1459 15197
rect 860 15192 1459 15194
rect 860 15136 1398 15192
rect 1454 15136 1459 15192
rect 860 15134 1459 15136
rect 860 15132 866 15134
rect 1393 15131 1459 15134
rect -300 15058 160 15088
rect 422 15058 428 15060
rect -300 14998 428 15058
rect -300 14968 160 14998
rect 422 14996 428 14998
rect 492 14996 498 15060
rect 1580 14922 1640 15270
rect 2129 15328 4679 15330
rect 2129 15272 2134 15328
rect 2190 15272 4618 15328
rect 4674 15272 4679 15328
rect 2129 15270 4679 15272
rect 2129 15267 2195 15270
rect 4613 15267 4679 15270
rect 4800 15328 6059 15330
rect 4800 15272 5998 15328
rect 6054 15272 6059 15328
rect 4800 15270 6059 15272
rect 2405 15194 2471 15197
rect 4800 15194 4860 15270
rect 5993 15267 6059 15270
rect 18086 15268 18092 15332
rect 18156 15330 18162 15332
rect 20805 15330 20871 15333
rect 18156 15328 20871 15330
rect 18156 15272 20810 15328
rect 20866 15272 20871 15328
rect 18156 15270 20871 15272
rect 18156 15268 18162 15270
rect 20805 15267 20871 15270
rect 22553 15330 22619 15333
rect 22840 15330 23300 15360
rect 22553 15328 23300 15330
rect 22553 15272 22558 15328
rect 22614 15272 23300 15328
rect 22553 15270 23300 15272
rect 22553 15267 22619 15270
rect 6144 15264 6460 15265
rect 6144 15200 6150 15264
rect 6214 15200 6230 15264
rect 6294 15200 6310 15264
rect 6374 15200 6390 15264
rect 6454 15200 6460 15264
rect 6144 15199 6460 15200
rect 11342 15264 11658 15265
rect 11342 15200 11348 15264
rect 11412 15200 11428 15264
rect 11492 15200 11508 15264
rect 11572 15200 11588 15264
rect 11652 15200 11658 15264
rect 11342 15199 11658 15200
rect 16540 15264 16856 15265
rect 16540 15200 16546 15264
rect 16610 15200 16626 15264
rect 16690 15200 16706 15264
rect 16770 15200 16786 15264
rect 16850 15200 16856 15264
rect 16540 15199 16856 15200
rect 21738 15264 22054 15265
rect 21738 15200 21744 15264
rect 21808 15200 21824 15264
rect 21888 15200 21904 15264
rect 21968 15200 21984 15264
rect 22048 15200 22054 15264
rect 22840 15240 23300 15270
rect 21738 15199 22054 15200
rect 5073 15196 5139 15197
rect 8385 15196 8451 15197
rect 2405 15192 4860 15194
rect 2405 15136 2410 15192
rect 2466 15136 4860 15192
rect 2405 15134 4860 15136
rect 2405 15131 2471 15134
rect 5022 15132 5028 15196
rect 5092 15194 5139 15196
rect 5092 15192 5184 15194
rect 5134 15136 5184 15192
rect 5092 15134 5184 15136
rect 5092 15132 5139 15134
rect 8334 15132 8340 15196
rect 8404 15194 8451 15196
rect 8404 15192 8496 15194
rect 8446 15136 8496 15192
rect 8404 15134 8496 15136
rect 8404 15132 8451 15134
rect 13118 15132 13124 15196
rect 13188 15194 13194 15196
rect 15326 15194 15332 15196
rect 13188 15134 15332 15194
rect 13188 15132 13194 15134
rect 15326 15132 15332 15134
rect 15396 15132 15402 15196
rect 5073 15131 5139 15132
rect 8385 15131 8451 15132
rect 2589 15060 2655 15061
rect 2589 15058 2636 15060
rect 2544 15056 2636 15058
rect 2544 15000 2594 15056
rect 2544 14998 2636 15000
rect 2589 14996 2636 14998
rect 2700 14996 2706 15060
rect 3366 14996 3372 15060
rect 3436 15058 3442 15060
rect 9121 15058 9187 15061
rect 3436 15056 9187 15058
rect 3436 15000 9126 15056
rect 9182 15000 9187 15056
rect 3436 14998 9187 15000
rect 3436 14996 3442 14998
rect 2589 14995 2655 14996
rect 9121 14995 9187 14998
rect 5717 14922 5783 14925
rect 1580 14920 5783 14922
rect 1580 14864 5722 14920
rect 5778 14864 5783 14920
rect 1580 14862 5783 14864
rect 5717 14859 5783 14862
rect 6862 14860 6868 14924
rect 6932 14922 6938 14924
rect 9622 14922 9628 14924
rect 6932 14862 9628 14922
rect 6932 14860 6938 14862
rect 9622 14860 9628 14862
rect 9692 14860 9698 14924
rect 12934 14860 12940 14924
rect 13004 14922 13010 14924
rect 18045 14922 18111 14925
rect 18454 14922 18460 14924
rect 13004 14920 18460 14922
rect 13004 14864 18050 14920
rect 18106 14864 18460 14920
rect 13004 14862 18460 14864
rect 13004 14860 13010 14862
rect 18045 14859 18111 14862
rect 18454 14860 18460 14862
rect 18524 14860 18530 14924
rect 20294 14860 20300 14924
rect 20364 14922 20370 14924
rect 21541 14922 21607 14925
rect 20364 14920 21607 14922
rect 20364 14864 21546 14920
rect 21602 14864 21607 14920
rect 20364 14862 21607 14864
rect 20364 14860 20370 14862
rect 21541 14859 21607 14862
rect -300 14786 160 14816
rect 933 14786 999 14789
rect -300 14784 999 14786
rect -300 14728 938 14784
rect 994 14728 999 14784
rect -300 14726 999 14728
rect -300 14696 160 14726
rect 933 14723 999 14726
rect 4429 14786 4495 14789
rect 6453 14786 6519 14789
rect 7281 14786 7347 14789
rect 4429 14784 4860 14786
rect 4429 14728 4434 14784
rect 4490 14728 4860 14784
rect 4429 14726 4860 14728
rect 4429 14723 4495 14726
rect 3545 14720 3861 14721
rect 3545 14656 3551 14720
rect 3615 14656 3631 14720
rect 3695 14656 3711 14720
rect 3775 14656 3791 14720
rect 3855 14656 3861 14720
rect 3545 14655 3861 14656
rect 657 14650 723 14653
rect 3366 14650 3372 14652
rect 657 14648 3372 14650
rect 657 14592 662 14648
rect 718 14592 3372 14648
rect 657 14590 3372 14592
rect 657 14587 723 14590
rect 3366 14588 3372 14590
rect 3436 14588 3442 14652
rect 4245 14650 4311 14653
rect 4654 14650 4660 14652
rect 4245 14648 4660 14650
rect 4245 14592 4250 14648
rect 4306 14592 4660 14648
rect 4245 14590 4660 14592
rect 4245 14587 4311 14590
rect 4654 14588 4660 14590
rect 4724 14588 4730 14652
rect 4800 14650 4860 14726
rect 6453 14784 7347 14786
rect 6453 14728 6458 14784
rect 6514 14728 7286 14784
rect 7342 14728 7347 14784
rect 6453 14726 7347 14728
rect 6453 14723 6519 14726
rect 7281 14723 7347 14726
rect 21449 14786 21515 14789
rect 22840 14786 23300 14816
rect 21449 14784 23300 14786
rect 21449 14728 21454 14784
rect 21510 14728 23300 14784
rect 21449 14726 23300 14728
rect 21449 14723 21515 14726
rect 8743 14720 9059 14721
rect 8743 14656 8749 14720
rect 8813 14656 8829 14720
rect 8893 14656 8909 14720
rect 8973 14656 8989 14720
rect 9053 14656 9059 14720
rect 8743 14655 9059 14656
rect 13941 14720 14257 14721
rect 13941 14656 13947 14720
rect 14011 14656 14027 14720
rect 14091 14656 14107 14720
rect 14171 14656 14187 14720
rect 14251 14656 14257 14720
rect 13941 14655 14257 14656
rect 19139 14720 19455 14721
rect 19139 14656 19145 14720
rect 19209 14656 19225 14720
rect 19289 14656 19305 14720
rect 19369 14656 19385 14720
rect 19449 14656 19455 14720
rect 22840 14696 23300 14726
rect 19139 14655 19455 14656
rect 8201 14650 8267 14653
rect 4800 14648 8267 14650
rect 4800 14592 8206 14648
rect 8262 14592 8267 14648
rect 4800 14590 8267 14592
rect 8201 14587 8267 14590
rect -300 14514 160 14544
rect 1853 14514 1919 14517
rect -300 14512 1919 14514
rect -300 14456 1858 14512
rect 1914 14456 1919 14512
rect -300 14454 1919 14456
rect -300 14424 160 14454
rect 1853 14451 1919 14454
rect 3877 14514 3943 14517
rect 8293 14514 8359 14517
rect 3877 14512 8359 14514
rect 3877 14456 3882 14512
rect 3938 14456 8298 14512
rect 8354 14456 8359 14512
rect 3877 14454 8359 14456
rect 3877 14451 3943 14454
rect 8293 14451 8359 14454
rect 10777 14514 10843 14517
rect 12709 14514 12775 14517
rect 10777 14512 12775 14514
rect 10777 14456 10782 14512
rect 10838 14456 12714 14512
rect 12770 14456 12775 14512
rect 10777 14454 12775 14456
rect 10777 14451 10843 14454
rect 12709 14451 12775 14454
rect 3233 14378 3299 14381
rect 6729 14378 6795 14381
rect 3233 14376 6795 14378
rect 3233 14320 3238 14376
rect 3294 14320 6734 14376
rect 6790 14320 6795 14376
rect 3233 14318 6795 14320
rect 3233 14315 3299 14318
rect 6729 14315 6795 14318
rect 12198 14316 12204 14380
rect 12268 14378 12274 14380
rect 18045 14378 18111 14381
rect 12268 14376 18111 14378
rect 12268 14320 18050 14376
rect 18106 14320 18111 14376
rect 12268 14318 18111 14320
rect 12268 14316 12274 14318
rect 18045 14315 18111 14318
rect -300 14242 160 14272
rect 1669 14242 1735 14245
rect 3877 14244 3943 14245
rect 3877 14242 3924 14244
rect -300 14240 1735 14242
rect -300 14184 1674 14240
rect 1730 14184 1735 14240
rect -300 14182 1735 14184
rect 3832 14240 3924 14242
rect 3988 14242 3994 14244
rect 5257 14242 5323 14245
rect 3988 14240 5323 14242
rect 3832 14184 3882 14240
rect 3988 14184 5262 14240
rect 5318 14184 5323 14240
rect 3832 14182 3924 14184
rect -300 14152 160 14182
rect 1669 14179 1735 14182
rect 3877 14180 3924 14182
rect 3988 14182 5323 14184
rect 3988 14180 3994 14182
rect 3877 14179 3943 14180
rect 5257 14179 5323 14182
rect 22185 14242 22251 14245
rect 22840 14242 23300 14272
rect 22185 14240 23300 14242
rect 22185 14184 22190 14240
rect 22246 14184 23300 14240
rect 22185 14182 23300 14184
rect 22185 14179 22251 14182
rect 6144 14176 6460 14177
rect 6144 14112 6150 14176
rect 6214 14112 6230 14176
rect 6294 14112 6310 14176
rect 6374 14112 6390 14176
rect 6454 14112 6460 14176
rect 6144 14111 6460 14112
rect 11342 14176 11658 14177
rect 11342 14112 11348 14176
rect 11412 14112 11428 14176
rect 11492 14112 11508 14176
rect 11572 14112 11588 14176
rect 11652 14112 11658 14176
rect 11342 14111 11658 14112
rect 16540 14176 16856 14177
rect 16540 14112 16546 14176
rect 16610 14112 16626 14176
rect 16690 14112 16706 14176
rect 16770 14112 16786 14176
rect 16850 14112 16856 14176
rect 16540 14111 16856 14112
rect 21738 14176 22054 14177
rect 21738 14112 21744 14176
rect 21808 14112 21824 14176
rect 21888 14112 21904 14176
rect 21968 14112 21984 14176
rect 22048 14112 22054 14176
rect 22840 14152 23300 14182
rect 21738 14111 22054 14112
rect 3049 14106 3115 14109
rect 1396 14104 3115 14106
rect 1396 14048 3054 14104
rect 3110 14048 3115 14104
rect 1396 14046 3115 14048
rect -300 13970 160 14000
rect 1396 13970 1456 14046
rect 3049 14043 3115 14046
rect 5073 14106 5139 14109
rect 5942 14106 5948 14108
rect 5073 14104 5948 14106
rect 5073 14048 5078 14104
rect 5134 14048 5948 14104
rect 5073 14046 5948 14048
rect 5073 14043 5139 14046
rect 5942 14044 5948 14046
rect 6012 14044 6018 14108
rect 13302 14044 13308 14108
rect 13372 14106 13378 14108
rect 13372 14046 16130 14106
rect 13372 14044 13378 14046
rect -300 13910 1456 13970
rect 1761 13970 1827 13973
rect 15929 13970 15995 13973
rect 1761 13968 15995 13970
rect 1761 13912 1766 13968
rect 1822 13912 15934 13968
rect 15990 13912 15995 13968
rect 1761 13910 15995 13912
rect 16070 13970 16130 14046
rect 17350 13970 17356 13972
rect 16070 13910 17356 13970
rect -300 13880 160 13910
rect 1761 13907 1827 13910
rect 15929 13907 15995 13910
rect 17350 13908 17356 13910
rect 17420 13908 17426 13972
rect 18822 13908 18828 13972
rect 18892 13970 18898 13972
rect 21173 13970 21239 13973
rect 18892 13968 21239 13970
rect 18892 13912 21178 13968
rect 21234 13912 21239 13968
rect 18892 13910 21239 13912
rect 18892 13908 18898 13910
rect 21173 13907 21239 13910
rect 238 13772 244 13836
rect 308 13834 314 13836
rect 933 13834 999 13837
rect 308 13832 999 13834
rect 308 13776 938 13832
rect 994 13776 999 13832
rect 308 13774 999 13776
rect 308 13772 314 13774
rect 933 13771 999 13774
rect 1393 13834 1459 13837
rect 5574 13834 5580 13836
rect 1393 13832 5580 13834
rect 1393 13776 1398 13832
rect 1454 13776 5580 13832
rect 1393 13774 5580 13776
rect 1393 13771 1459 13774
rect 5574 13772 5580 13774
rect 5644 13772 5650 13836
rect 8201 13834 8267 13837
rect 9765 13834 9831 13837
rect 8201 13832 9831 13834
rect 8201 13776 8206 13832
rect 8262 13776 9770 13832
rect 9826 13776 9831 13832
rect 8201 13774 9831 13776
rect 8201 13771 8267 13774
rect 9765 13771 9831 13774
rect 12341 13834 12407 13837
rect 12341 13832 14474 13834
rect 12341 13776 12346 13832
rect 12402 13776 14474 13832
rect 12341 13774 14474 13776
rect 12341 13771 12407 13774
rect -300 13698 160 13728
rect 2865 13698 2931 13701
rect 2998 13698 3004 13700
rect -300 13638 1042 13698
rect -300 13608 160 13638
rect 982 13562 1042 13638
rect 2865 13696 3004 13698
rect 2865 13640 2870 13696
rect 2926 13640 3004 13696
rect 2865 13638 3004 13640
rect 2865 13635 2931 13638
rect 2998 13636 3004 13638
rect 3068 13636 3074 13700
rect 4521 13698 4587 13701
rect 5022 13698 5028 13700
rect 4521 13696 5028 13698
rect 4521 13640 4526 13696
rect 4582 13640 5028 13696
rect 4521 13638 5028 13640
rect 4521 13635 4587 13638
rect 5022 13636 5028 13638
rect 5092 13636 5098 13700
rect 7230 13636 7236 13700
rect 7300 13698 7306 13700
rect 7833 13698 7899 13701
rect 12525 13700 12591 13701
rect 12525 13698 12572 13700
rect 7300 13696 7899 13698
rect 7300 13640 7838 13696
rect 7894 13640 7899 13696
rect 7300 13638 7899 13640
rect 12480 13696 12572 13698
rect 12480 13640 12530 13696
rect 12480 13638 12572 13640
rect 7300 13636 7306 13638
rect 7833 13635 7899 13638
rect 12525 13636 12572 13638
rect 12636 13636 12642 13700
rect 14414 13698 14474 13774
rect 17953 13700 18019 13701
rect 14414 13638 14658 13698
rect 12525 13635 12591 13636
rect 3545 13632 3861 13633
rect 3545 13568 3551 13632
rect 3615 13568 3631 13632
rect 3695 13568 3711 13632
rect 3775 13568 3791 13632
rect 3855 13568 3861 13632
rect 3545 13567 3861 13568
rect 8743 13632 9059 13633
rect 8743 13568 8749 13632
rect 8813 13568 8829 13632
rect 8893 13568 8909 13632
rect 8973 13568 8989 13632
rect 9053 13568 9059 13632
rect 8743 13567 9059 13568
rect 13941 13632 14257 13633
rect 13941 13568 13947 13632
rect 14011 13568 14027 13632
rect 14091 13568 14107 13632
rect 14171 13568 14187 13632
rect 14251 13568 14257 13632
rect 13941 13567 14257 13568
rect 1761 13562 1827 13565
rect 982 13560 1827 13562
rect 982 13504 1766 13560
rect 1822 13504 1827 13560
rect 982 13502 1827 13504
rect 1761 13499 1827 13502
rect 2589 13562 2655 13565
rect 2814 13562 2820 13564
rect 2589 13560 2820 13562
rect 2589 13504 2594 13560
rect 2650 13504 2820 13560
rect 2589 13502 2820 13504
rect 2589 13499 2655 13502
rect 2814 13500 2820 13502
rect 2884 13500 2890 13564
rect 4889 13562 4955 13565
rect 5901 13562 5967 13565
rect 4889 13560 5967 13562
rect 4889 13504 4894 13560
rect 4950 13504 5906 13560
rect 5962 13504 5967 13560
rect 4889 13502 5967 13504
rect 4889 13499 4955 13502
rect 5901 13499 5967 13502
rect 9438 13500 9444 13564
rect 9508 13562 9514 13564
rect 9581 13562 9647 13565
rect 14598 13564 14658 13638
rect 17902 13636 17908 13700
rect 17972 13698 18019 13700
rect 21449 13698 21515 13701
rect 22840 13698 23300 13728
rect 17972 13696 18064 13698
rect 18014 13640 18064 13696
rect 17972 13638 18064 13640
rect 21449 13696 23300 13698
rect 21449 13640 21454 13696
rect 21510 13640 23300 13696
rect 21449 13638 23300 13640
rect 17972 13636 18019 13638
rect 17953 13635 18019 13636
rect 21449 13635 21515 13638
rect 19139 13632 19455 13633
rect 19139 13568 19145 13632
rect 19209 13568 19225 13632
rect 19289 13568 19305 13632
rect 19369 13568 19385 13632
rect 19449 13568 19455 13632
rect 22840 13608 23300 13638
rect 19139 13567 19455 13568
rect 9508 13560 9647 13562
rect 9508 13504 9586 13560
rect 9642 13504 9647 13560
rect 9508 13502 9647 13504
rect 9508 13500 9514 13502
rect 9581 13499 9647 13502
rect 14590 13500 14596 13564
rect 14660 13500 14666 13564
rect -300 13426 160 13456
rect 4429 13426 4495 13429
rect 6269 13426 6335 13429
rect 15653 13426 15719 13429
rect -300 13424 4495 13426
rect -300 13368 4434 13424
rect 4490 13368 4495 13424
rect -300 13366 4495 13368
rect -300 13336 160 13366
rect 4429 13363 4495 13366
rect 4984 13424 6335 13426
rect 4984 13368 6274 13424
rect 6330 13368 6335 13424
rect 4984 13366 6335 13368
rect 4984 13293 5044 13366
rect 6269 13363 6335 13366
rect 7606 13424 15719 13426
rect 7606 13368 15658 13424
rect 15714 13368 15719 13424
rect 7606 13366 15719 13368
rect 1158 13228 1164 13292
rect 1228 13290 1234 13292
rect 3785 13290 3851 13293
rect 3918 13290 3924 13292
rect 1228 13230 3066 13290
rect 1228 13228 1234 13230
rect -300 13154 160 13184
rect 2865 13154 2931 13157
rect -300 13152 2931 13154
rect -300 13096 2870 13152
rect 2926 13096 2931 13152
rect -300 13094 2931 13096
rect 3006 13154 3066 13230
rect 3785 13288 3924 13290
rect 3785 13232 3790 13288
rect 3846 13232 3924 13288
rect 3785 13230 3924 13232
rect 3785 13227 3851 13230
rect 3918 13228 3924 13230
rect 3988 13228 3994 13292
rect 4613 13290 4679 13293
rect 4838 13290 4844 13292
rect 4613 13288 4844 13290
rect 4613 13232 4618 13288
rect 4674 13232 4844 13288
rect 4613 13230 4844 13232
rect 4613 13227 4679 13230
rect 4838 13228 4844 13230
rect 4908 13228 4914 13292
rect 4981 13288 5047 13293
rect 4981 13232 4986 13288
rect 5042 13232 5047 13288
rect 4981 13227 5047 13232
rect 5349 13290 5415 13293
rect 5717 13290 5783 13293
rect 5349 13288 5783 13290
rect 5349 13232 5354 13288
rect 5410 13232 5722 13288
rect 5778 13232 5783 13288
rect 5349 13230 5783 13232
rect 5349 13227 5415 13230
rect 5717 13227 5783 13230
rect 5942 13228 5948 13292
rect 6012 13228 6018 13292
rect 5950 13154 6010 13228
rect 3006 13094 6010 13154
rect -300 13064 160 13094
rect 2865 13091 2931 13094
rect 6144 13088 6460 13089
rect 6144 13024 6150 13088
rect 6214 13024 6230 13088
rect 6294 13024 6310 13088
rect 6374 13024 6390 13088
rect 6454 13024 6460 13088
rect 6144 13023 6460 13024
rect 422 12956 428 13020
rect 492 13018 498 13020
rect 933 13018 999 13021
rect 492 13016 999 13018
rect 492 12960 938 13016
rect 994 12960 999 13016
rect 492 12958 999 12960
rect 492 12956 498 12958
rect 933 12955 999 12958
rect 1342 12956 1348 13020
rect 1412 13018 1418 13020
rect 2078 13018 2084 13020
rect 1412 12958 2084 13018
rect 1412 12956 1418 12958
rect 2078 12956 2084 12958
rect 2148 12956 2154 13020
rect 7281 13018 7347 13021
rect 6686 13016 7347 13018
rect 6686 12960 7286 13016
rect 7342 12960 7347 13016
rect 6686 12958 7347 12960
rect -300 12882 160 12912
rect 2773 12882 2839 12885
rect -300 12880 2839 12882
rect -300 12824 2778 12880
rect 2834 12824 2839 12880
rect -300 12822 2839 12824
rect -300 12792 160 12822
rect 2773 12819 2839 12822
rect 3049 12882 3115 12885
rect 6686 12882 6746 12958
rect 7281 12955 7347 12958
rect 3049 12880 6746 12882
rect 3049 12824 3054 12880
rect 3110 12824 6746 12880
rect 3049 12822 6746 12824
rect 3049 12819 3115 12822
rect 7230 12820 7236 12884
rect 7300 12882 7306 12884
rect 7373 12882 7439 12885
rect 7300 12880 7439 12882
rect 7300 12824 7378 12880
rect 7434 12824 7439 12880
rect 7300 12822 7439 12824
rect 7300 12820 7306 12822
rect 7373 12819 7439 12822
rect 2589 12746 2655 12749
rect 7606 12746 7666 13366
rect 15653 13363 15719 13366
rect 7741 13290 7807 13293
rect 9438 13290 9444 13292
rect 7741 13288 9444 13290
rect 7741 13232 7746 13288
rect 7802 13232 9444 13288
rect 7741 13230 9444 13232
rect 7741 13227 7807 13230
rect 9438 13228 9444 13230
rect 9508 13228 9514 13292
rect 18321 13290 18387 13293
rect 19926 13290 19932 13292
rect 18321 13288 19932 13290
rect 18321 13232 18326 13288
rect 18382 13232 19932 13288
rect 18321 13230 19932 13232
rect 18321 13227 18387 13230
rect 19926 13228 19932 13230
rect 19996 13228 20002 13292
rect 7925 13154 7991 13157
rect 7925 13152 11208 13154
rect 7925 13096 7930 13152
rect 7986 13096 11208 13152
rect 7925 13094 11208 13096
rect 7925 13091 7991 13094
rect 11148 13021 11208 13094
rect 18822 13092 18828 13156
rect 18892 13154 18898 13156
rect 19977 13154 20043 13157
rect 18892 13152 20043 13154
rect 18892 13096 19982 13152
rect 20038 13096 20043 13152
rect 18892 13094 20043 13096
rect 18892 13092 18898 13094
rect 19977 13091 20043 13094
rect 22185 13154 22251 13157
rect 22840 13154 23300 13184
rect 22185 13152 23300 13154
rect 22185 13096 22190 13152
rect 22246 13096 23300 13152
rect 22185 13094 23300 13096
rect 22185 13091 22251 13094
rect 11342 13088 11658 13089
rect 11342 13024 11348 13088
rect 11412 13024 11428 13088
rect 11492 13024 11508 13088
rect 11572 13024 11588 13088
rect 11652 13024 11658 13088
rect 11342 13023 11658 13024
rect 16540 13088 16856 13089
rect 16540 13024 16546 13088
rect 16610 13024 16626 13088
rect 16690 13024 16706 13088
rect 16770 13024 16786 13088
rect 16850 13024 16856 13088
rect 16540 13023 16856 13024
rect 21738 13088 22054 13089
rect 21738 13024 21744 13088
rect 21808 13024 21824 13088
rect 21888 13024 21904 13088
rect 21968 13024 21984 13088
rect 22048 13024 22054 13088
rect 22840 13064 23300 13094
rect 21738 13023 22054 13024
rect 9857 13018 9923 13021
rect 9814 13016 9923 13018
rect 9814 12960 9862 13016
rect 9918 12960 9923 13016
rect 9814 12955 9923 12960
rect 10225 13018 10291 13021
rect 10593 13018 10659 13021
rect 10225 13016 10659 13018
rect 10225 12960 10230 13016
rect 10286 12960 10598 13016
rect 10654 12960 10659 13016
rect 10225 12958 10659 12960
rect 10225 12955 10291 12958
rect 10593 12955 10659 12958
rect 11145 13016 11211 13021
rect 11145 12960 11150 13016
rect 11206 12960 11211 13016
rect 11145 12955 11211 12960
rect 13169 13018 13235 13021
rect 15561 13018 15627 13021
rect 13169 13016 15627 13018
rect 13169 12960 13174 13016
rect 13230 12960 15566 13016
rect 15622 12960 15627 13016
rect 13169 12958 15627 12960
rect 13169 12955 13235 12958
rect 15561 12955 15627 12958
rect 9814 12749 9874 12955
rect 10225 12882 10291 12885
rect 13813 12882 13879 12885
rect 10225 12880 13879 12882
rect 10225 12824 10230 12880
rect 10286 12824 13818 12880
rect 13874 12824 13879 12880
rect 10225 12822 13879 12824
rect 10225 12819 10291 12822
rect 13813 12819 13879 12822
rect 2589 12744 7666 12746
rect 2589 12688 2594 12744
rect 2650 12688 7666 12744
rect 2589 12686 7666 12688
rect 9029 12746 9095 12749
rect 9029 12744 9690 12746
rect 9029 12688 9034 12744
rect 9090 12688 9690 12744
rect 9029 12686 9690 12688
rect 9814 12744 9923 12749
rect 9814 12688 9862 12744
rect 9918 12688 9923 12744
rect 9814 12686 9923 12688
rect 2589 12683 2655 12686
rect 9029 12683 9095 12686
rect -300 12610 160 12640
rect 3049 12610 3115 12613
rect -300 12608 3115 12610
rect -300 12552 3054 12608
rect 3110 12552 3115 12608
rect -300 12550 3115 12552
rect -300 12520 160 12550
rect 3049 12547 3115 12550
rect 3969 12610 4035 12613
rect 7649 12612 7715 12613
rect 7046 12610 7052 12612
rect 3969 12608 7052 12610
rect 3969 12552 3974 12608
rect 4030 12552 7052 12608
rect 3969 12550 7052 12552
rect 3969 12547 4035 12550
rect 7046 12548 7052 12550
rect 7116 12548 7122 12612
rect 7598 12548 7604 12612
rect 7668 12610 7715 12612
rect 9630 12610 9690 12686
rect 9857 12683 9923 12686
rect 10317 12746 10383 12749
rect 11973 12746 12039 12749
rect 10317 12744 12039 12746
rect 10317 12688 10322 12744
rect 10378 12688 11978 12744
rect 12034 12688 12039 12744
rect 10317 12686 12039 12688
rect 10317 12683 10383 12686
rect 11973 12683 12039 12686
rect 12893 12746 12959 12749
rect 15285 12746 15351 12749
rect 12893 12744 15351 12746
rect 12893 12688 12898 12744
rect 12954 12688 15290 12744
rect 15346 12688 15351 12744
rect 12893 12686 15351 12688
rect 12893 12683 12959 12686
rect 15285 12683 15351 12686
rect 12014 12610 12020 12612
rect 7668 12608 7760 12610
rect 7710 12552 7760 12608
rect 7668 12550 7760 12552
rect 9630 12550 12020 12610
rect 7668 12548 7715 12550
rect 12014 12548 12020 12550
rect 12084 12548 12090 12612
rect 21081 12610 21147 12613
rect 22840 12610 23300 12640
rect 21081 12608 23300 12610
rect 21081 12552 21086 12608
rect 21142 12552 23300 12608
rect 21081 12550 23300 12552
rect 7649 12547 7715 12548
rect 21081 12547 21147 12550
rect 3545 12544 3861 12545
rect 3545 12480 3551 12544
rect 3615 12480 3631 12544
rect 3695 12480 3711 12544
rect 3775 12480 3791 12544
rect 3855 12480 3861 12544
rect 3545 12479 3861 12480
rect 8743 12544 9059 12545
rect 8743 12480 8749 12544
rect 8813 12480 8829 12544
rect 8893 12480 8909 12544
rect 8973 12480 8989 12544
rect 9053 12480 9059 12544
rect 8743 12479 9059 12480
rect 13941 12544 14257 12545
rect 13941 12480 13947 12544
rect 14011 12480 14027 12544
rect 14091 12480 14107 12544
rect 14171 12480 14187 12544
rect 14251 12480 14257 12544
rect 13941 12479 14257 12480
rect 19139 12544 19455 12545
rect 19139 12480 19145 12544
rect 19209 12480 19225 12544
rect 19289 12480 19305 12544
rect 19369 12480 19385 12544
rect 19449 12480 19455 12544
rect 22840 12520 23300 12550
rect 19139 12479 19455 12480
rect 5717 12474 5783 12477
rect 6913 12474 6979 12477
rect 5717 12472 6979 12474
rect 5717 12416 5722 12472
rect 5778 12416 6918 12472
rect 6974 12416 6979 12472
rect 5717 12414 6979 12416
rect 5717 12411 5783 12414
rect 6913 12411 6979 12414
rect 7649 12474 7715 12477
rect 7782 12474 7788 12476
rect 7649 12472 7788 12474
rect 7649 12416 7654 12472
rect 7710 12416 7788 12472
rect 7649 12414 7788 12416
rect 7649 12411 7715 12414
rect 7782 12412 7788 12414
rect 7852 12412 7858 12476
rect 11094 12412 11100 12476
rect 11164 12474 11170 12476
rect 12801 12474 12867 12477
rect 11164 12472 12867 12474
rect 11164 12416 12806 12472
rect 12862 12416 12867 12472
rect 11164 12414 12867 12416
rect 11164 12412 11170 12414
rect 12801 12411 12867 12414
rect 19742 12412 19748 12476
rect 19812 12474 19818 12476
rect 19812 12414 20730 12474
rect 19812 12412 19818 12414
rect -300 12338 160 12368
rect 3969 12338 4035 12341
rect -300 12336 4035 12338
rect -300 12280 3974 12336
rect 4030 12280 4035 12336
rect -300 12278 4035 12280
rect -300 12248 160 12278
rect 3969 12275 4035 12278
rect 4654 12276 4660 12340
rect 4724 12338 4730 12340
rect 5073 12338 5139 12341
rect 4724 12336 5139 12338
rect 4724 12280 5078 12336
rect 5134 12280 5139 12336
rect 4724 12278 5139 12280
rect 4724 12276 4730 12278
rect 5073 12275 5139 12278
rect 6269 12338 6335 12341
rect 7373 12338 7439 12341
rect 15193 12338 15259 12341
rect 19057 12340 19123 12341
rect 6269 12336 7439 12338
rect 6269 12280 6274 12336
rect 6330 12280 7378 12336
rect 7434 12280 7439 12336
rect 6269 12278 7439 12280
rect 6269 12275 6335 12278
rect 7373 12275 7439 12278
rect 7606 12336 15259 12338
rect 7606 12280 15198 12336
rect 15254 12280 15259 12336
rect 7606 12278 15259 12280
rect 1485 12202 1551 12205
rect 7606 12202 7666 12278
rect 15193 12275 15259 12278
rect 19006 12276 19012 12340
rect 19076 12338 19123 12340
rect 20670 12338 20730 12414
rect 20805 12338 20871 12341
rect 19076 12336 19168 12338
rect 19118 12280 19168 12336
rect 19076 12278 19168 12280
rect 20670 12336 20871 12338
rect 20670 12280 20810 12336
rect 20866 12280 20871 12336
rect 20670 12278 20871 12280
rect 19076 12276 19123 12278
rect 19057 12275 19123 12276
rect 20805 12275 20871 12278
rect 1485 12200 7666 12202
rect 1485 12144 1490 12200
rect 1546 12144 7666 12200
rect 1485 12142 7666 12144
rect 11053 12204 11119 12205
rect 11053 12200 11100 12204
rect 11164 12202 11170 12204
rect 11053 12144 11058 12200
rect 1485 12139 1551 12142
rect 11053 12140 11100 12144
rect 11164 12142 11210 12202
rect 11164 12140 11170 12142
rect 11830 12140 11836 12204
rect 11900 12202 11906 12204
rect 13905 12202 13971 12205
rect 18321 12202 18387 12205
rect 11900 12142 12634 12202
rect 11900 12140 11906 12142
rect 11053 12139 11119 12140
rect -300 12066 160 12096
rect 12574 12069 12634 12142
rect 13905 12200 18387 12202
rect 13905 12144 13910 12200
rect 13966 12144 18326 12200
rect 18382 12144 18387 12200
rect 13905 12142 18387 12144
rect 13905 12139 13971 12142
rect 18321 12139 18387 12142
rect 4061 12066 4127 12069
rect 5349 12066 5415 12069
rect -300 12064 4127 12066
rect -300 12008 4066 12064
rect 4122 12008 4127 12064
rect -300 12006 4127 12008
rect -300 11976 160 12006
rect 4061 12003 4127 12006
rect 4478 12064 5415 12066
rect 4478 12008 5354 12064
rect 5410 12008 5415 12064
rect 4478 12006 5415 12008
rect 1577 11930 1643 11933
rect 4153 11932 4219 11933
rect 1577 11928 3112 11930
rect 1577 11872 1582 11928
rect 1638 11872 3112 11928
rect 1577 11870 3112 11872
rect 1577 11867 1643 11870
rect -300 11794 160 11824
rect 1577 11796 1643 11797
rect -300 11734 858 11794
rect -300 11704 160 11734
rect 798 11658 858 11734
rect 1526 11732 1532 11796
rect 1596 11794 1643 11796
rect 1761 11794 1827 11797
rect 1894 11794 1900 11796
rect 1596 11792 1688 11794
rect 1638 11736 1688 11792
rect 1596 11734 1688 11736
rect 1761 11792 1900 11794
rect 1761 11736 1766 11792
rect 1822 11736 1900 11792
rect 1761 11734 1900 11736
rect 1596 11732 1643 11734
rect 1577 11731 1643 11732
rect 1761 11731 1827 11734
rect 1894 11732 1900 11734
rect 1964 11732 1970 11796
rect 3052 11794 3112 11870
rect 3182 11868 3188 11932
rect 3252 11930 3258 11932
rect 3918 11930 3924 11932
rect 3252 11870 3924 11930
rect 3252 11868 3258 11870
rect 3918 11868 3924 11870
rect 3988 11868 3994 11932
rect 4102 11868 4108 11932
rect 4172 11930 4219 11932
rect 4172 11928 4264 11930
rect 4214 11872 4264 11928
rect 4172 11870 4264 11872
rect 4172 11868 4219 11870
rect 4153 11867 4219 11868
rect 4478 11794 4538 12006
rect 5349 12003 5415 12006
rect 5574 12004 5580 12068
rect 5644 12066 5650 12068
rect 5993 12066 6059 12069
rect 5644 12064 6059 12066
rect 5644 12008 5998 12064
rect 6054 12008 6059 12064
rect 5644 12006 6059 12008
rect 5644 12004 5650 12006
rect 5993 12003 6059 12006
rect 7189 12066 7255 12069
rect 7649 12066 7715 12069
rect 9489 12066 9555 12069
rect 7189 12064 9555 12066
rect 7189 12008 7194 12064
rect 7250 12008 7654 12064
rect 7710 12008 9494 12064
rect 9550 12008 9555 12064
rect 7189 12006 9555 12008
rect 12574 12064 12683 12069
rect 12574 12008 12622 12064
rect 12678 12008 12683 12064
rect 12574 12006 12683 12008
rect 7189 12003 7255 12006
rect 7649 12003 7715 12006
rect 9489 12003 9555 12006
rect 12617 12003 12683 12006
rect 17166 12004 17172 12068
rect 17236 12066 17242 12068
rect 17493 12066 17559 12069
rect 17236 12064 17559 12066
rect 17236 12008 17498 12064
rect 17554 12008 17559 12064
rect 17236 12006 17559 12008
rect 17236 12004 17242 12006
rect 17493 12003 17559 12006
rect 22185 12066 22251 12069
rect 22840 12066 23300 12096
rect 22185 12064 23300 12066
rect 22185 12008 22190 12064
rect 22246 12008 23300 12064
rect 22185 12006 23300 12008
rect 22185 12003 22251 12006
rect 6144 12000 6460 12001
rect 6144 11936 6150 12000
rect 6214 11936 6230 12000
rect 6294 11936 6310 12000
rect 6374 11936 6390 12000
rect 6454 11936 6460 12000
rect 6144 11935 6460 11936
rect 11342 12000 11658 12001
rect 11342 11936 11348 12000
rect 11412 11936 11428 12000
rect 11492 11936 11508 12000
rect 11572 11936 11588 12000
rect 11652 11936 11658 12000
rect 11342 11935 11658 11936
rect 16540 12000 16856 12001
rect 16540 11936 16546 12000
rect 16610 11936 16626 12000
rect 16690 11936 16706 12000
rect 16770 11936 16786 12000
rect 16850 11936 16856 12000
rect 16540 11935 16856 11936
rect 21738 12000 22054 12001
rect 21738 11936 21744 12000
rect 21808 11936 21824 12000
rect 21888 11936 21904 12000
rect 21968 11936 21984 12000
rect 22048 11936 22054 12000
rect 22840 11976 23300 12006
rect 21738 11935 22054 11936
rect 7925 11930 7991 11933
rect 10317 11930 10383 11933
rect 12249 11930 12315 11933
rect 7925 11928 10383 11930
rect 7925 11872 7930 11928
rect 7986 11872 10322 11928
rect 10378 11872 10383 11928
rect 7925 11870 10383 11872
rect 7925 11867 7991 11870
rect 10317 11867 10383 11870
rect 11838 11928 12315 11930
rect 11838 11872 12254 11928
rect 12310 11872 12315 11928
rect 11838 11870 12315 11872
rect 3052 11734 4538 11794
rect 5625 11794 5691 11797
rect 10174 11794 10180 11796
rect 5625 11792 10180 11794
rect 5625 11736 5630 11792
rect 5686 11736 10180 11792
rect 5625 11734 10180 11736
rect 5625 11731 5691 11734
rect 10174 11732 10180 11734
rect 10244 11732 10250 11796
rect 10358 11732 10364 11796
rect 10428 11794 10434 11796
rect 11838 11794 11898 11870
rect 12249 11867 12315 11870
rect 16982 11868 16988 11932
rect 17052 11930 17058 11932
rect 17585 11930 17651 11933
rect 17052 11928 17651 11930
rect 17052 11872 17590 11928
rect 17646 11872 17651 11928
rect 17052 11870 17651 11872
rect 17052 11868 17058 11870
rect 17585 11867 17651 11870
rect 10428 11734 11898 11794
rect 13537 11794 13603 11797
rect 16481 11794 16547 11797
rect 13537 11792 16547 11794
rect 13537 11736 13542 11792
rect 13598 11736 16486 11792
rect 16542 11736 16547 11792
rect 13537 11734 16547 11736
rect 10428 11732 10434 11734
rect 13537 11731 13603 11734
rect 16481 11731 16547 11734
rect 18781 11794 18847 11797
rect 22829 11794 22895 11797
rect 18781 11792 22895 11794
rect 18781 11736 18786 11792
rect 18842 11736 22834 11792
rect 22890 11736 22895 11792
rect 18781 11734 22895 11736
rect 18781 11731 18847 11734
rect 22829 11731 22895 11734
rect 1485 11658 1551 11661
rect 798 11656 1551 11658
rect 798 11600 1490 11656
rect 1546 11600 1551 11656
rect 798 11598 1551 11600
rect 1485 11595 1551 11598
rect 2078 11596 2084 11660
rect 2148 11658 2154 11660
rect 2313 11658 2379 11661
rect 2148 11656 2379 11658
rect 2148 11600 2318 11656
rect 2374 11600 2379 11656
rect 2148 11598 2379 11600
rect 2148 11596 2154 11598
rect 2313 11595 2379 11598
rect 2681 11658 2747 11661
rect 8293 11658 8359 11661
rect 20069 11658 20135 11661
rect 2681 11656 20135 11658
rect 2681 11600 2686 11656
rect 2742 11600 8298 11656
rect 8354 11600 20074 11656
rect 20130 11600 20135 11656
rect 2681 11598 20135 11600
rect 2681 11595 2747 11598
rect 8293 11595 8359 11598
rect 20069 11595 20135 11598
rect -300 11522 160 11552
rect 1025 11522 1091 11525
rect -300 11520 1091 11522
rect -300 11464 1030 11520
rect 1086 11464 1091 11520
rect -300 11462 1091 11464
rect -300 11432 160 11462
rect 1025 11459 1091 11462
rect 4981 11522 5047 11525
rect 5206 11522 5212 11524
rect 4981 11520 5212 11522
rect 4981 11464 4986 11520
rect 5042 11464 5212 11520
rect 4981 11462 5212 11464
rect 4981 11459 5047 11462
rect 5206 11460 5212 11462
rect 5276 11460 5282 11524
rect 5349 11522 5415 11525
rect 6361 11522 6427 11525
rect 5349 11520 6427 11522
rect 5349 11464 5354 11520
rect 5410 11464 6366 11520
rect 6422 11464 6427 11520
rect 5349 11462 6427 11464
rect 5349 11459 5415 11462
rect 6361 11459 6427 11462
rect 21081 11522 21147 11525
rect 22840 11522 23300 11552
rect 21081 11520 23300 11522
rect 21081 11464 21086 11520
rect 21142 11464 23300 11520
rect 21081 11462 23300 11464
rect 21081 11459 21147 11462
rect 3545 11456 3861 11457
rect 3545 11392 3551 11456
rect 3615 11392 3631 11456
rect 3695 11392 3711 11456
rect 3775 11392 3791 11456
rect 3855 11392 3861 11456
rect 3545 11391 3861 11392
rect 8743 11456 9059 11457
rect 8743 11392 8749 11456
rect 8813 11392 8829 11456
rect 8893 11392 8909 11456
rect 8973 11392 8989 11456
rect 9053 11392 9059 11456
rect 8743 11391 9059 11392
rect 13941 11456 14257 11457
rect 13941 11392 13947 11456
rect 14011 11392 14027 11456
rect 14091 11392 14107 11456
rect 14171 11392 14187 11456
rect 14251 11392 14257 11456
rect 13941 11391 14257 11392
rect 19139 11456 19455 11457
rect 19139 11392 19145 11456
rect 19209 11392 19225 11456
rect 19289 11392 19305 11456
rect 19369 11392 19385 11456
rect 19449 11392 19455 11456
rect 22840 11432 23300 11462
rect 19139 11391 19455 11392
rect 1669 11386 1735 11389
rect 2589 11386 2655 11389
rect 1669 11384 2655 11386
rect 1669 11328 1674 11384
rect 1730 11328 2594 11384
rect 2650 11328 2655 11384
rect 1669 11326 2655 11328
rect 1669 11323 1735 11326
rect 2589 11323 2655 11326
rect 4102 11324 4108 11388
rect 4172 11386 4178 11388
rect 12065 11386 12131 11389
rect 4172 11326 5642 11386
rect 4172 11324 4178 11326
rect -300 11250 160 11280
rect 2814 11250 2820 11252
rect -300 11190 2820 11250
rect -300 11160 160 11190
rect 2814 11188 2820 11190
rect 2884 11188 2890 11252
rect 3877 11250 3943 11253
rect 5582 11250 5642 11326
rect 9262 11384 12131 11386
rect 9262 11328 12070 11384
rect 12126 11328 12131 11384
rect 9262 11326 12131 11328
rect 9262 11250 9322 11326
rect 12065 11323 12131 11326
rect 16062 11324 16068 11388
rect 16132 11386 16138 11388
rect 16297 11386 16363 11389
rect 16132 11384 16363 11386
rect 16132 11328 16302 11384
rect 16358 11328 16363 11384
rect 16132 11326 16363 11328
rect 16132 11324 16138 11326
rect 16297 11323 16363 11326
rect 21357 11384 21423 11389
rect 21357 11328 21362 11384
rect 21418 11328 21423 11384
rect 21357 11323 21423 11328
rect 3877 11248 4354 11250
rect 3877 11192 3882 11248
rect 3938 11192 4354 11248
rect 3877 11190 4354 11192
rect 5582 11190 9322 11250
rect 9857 11250 9923 11253
rect 11329 11250 11395 11253
rect 20989 11250 21055 11253
rect 9857 11248 21055 11250
rect 9857 11192 9862 11248
rect 9918 11192 11334 11248
rect 11390 11192 20994 11248
rect 21050 11192 21055 11248
rect 9857 11190 21055 11192
rect 3877 11187 3943 11190
rect 2221 11116 2287 11117
rect 2221 11114 2268 11116
rect 2180 11112 2268 11114
rect 2332 11114 2338 11116
rect 2681 11114 2747 11117
rect 2332 11112 2747 11114
rect 2180 11056 2226 11112
rect 2332 11056 2686 11112
rect 2742 11056 2747 11112
rect 2180 11054 2268 11056
rect 2221 11052 2268 11054
rect 2332 11054 2747 11056
rect 4294 11114 4354 11190
rect 9857 11187 9923 11190
rect 11329 11187 11395 11190
rect 20989 11187 21055 11190
rect 13905 11114 13971 11117
rect 4294 11112 13971 11114
rect 4294 11056 13910 11112
rect 13966 11056 13971 11112
rect 4294 11054 13971 11056
rect 2332 11052 2338 11054
rect 2221 11051 2287 11052
rect 2681 11051 2747 11054
rect 13905 11051 13971 11054
rect 15837 11114 15903 11117
rect 21360 11114 21420 11323
rect 15837 11112 21420 11114
rect 15837 11056 15842 11112
rect 15898 11056 21420 11112
rect 15837 11054 21420 11056
rect 15837 11051 15903 11054
rect -300 10978 160 11008
rect 4061 10978 4127 10981
rect 4337 10978 4403 10981
rect -300 10918 3618 10978
rect -300 10888 160 10918
rect 2681 10842 2747 10845
rect 3182 10842 3188 10844
rect 2681 10840 3188 10842
rect 2681 10784 2686 10840
rect 2742 10784 3188 10840
rect 2681 10782 3188 10784
rect 2681 10779 2747 10782
rect 3182 10780 3188 10782
rect 3252 10780 3258 10844
rect 3558 10842 3618 10918
rect 4061 10976 4403 10978
rect 4061 10920 4066 10976
rect 4122 10920 4342 10976
rect 4398 10920 4403 10976
rect 4061 10918 4403 10920
rect 4061 10915 4127 10918
rect 4337 10915 4403 10918
rect 4470 10916 4476 10980
rect 4540 10978 4546 10980
rect 4613 10978 4679 10981
rect 4540 10976 4679 10978
rect 4540 10920 4618 10976
rect 4674 10920 4679 10976
rect 4540 10918 4679 10920
rect 4540 10916 4546 10918
rect 4613 10915 4679 10918
rect 5390 10916 5396 10980
rect 5460 10978 5466 10980
rect 5460 10918 6010 10978
rect 5460 10916 5466 10918
rect 4337 10842 4403 10845
rect 3558 10840 4403 10842
rect 3558 10784 4342 10840
rect 4398 10784 4403 10840
rect 3558 10782 4403 10784
rect 4337 10779 4403 10782
rect 4981 10842 5047 10845
rect 5390 10842 5396 10844
rect 4981 10840 5396 10842
rect 4981 10784 4986 10840
rect 5042 10784 5396 10840
rect 4981 10782 5396 10784
rect 4981 10779 5047 10782
rect 5390 10780 5396 10782
rect 5460 10780 5466 10844
rect -300 10706 160 10736
rect 3969 10706 4035 10709
rect -300 10704 4035 10706
rect -300 10648 3974 10704
rect 4030 10648 4035 10704
rect -300 10646 4035 10648
rect -300 10616 160 10646
rect 3969 10643 4035 10646
rect 4153 10706 4219 10709
rect 5625 10706 5691 10709
rect 4153 10704 5691 10706
rect 4153 10648 4158 10704
rect 4214 10648 5630 10704
rect 5686 10648 5691 10704
rect 4153 10646 5691 10648
rect 5950 10706 6010 10918
rect 6862 10916 6868 10980
rect 6932 10978 6938 10980
rect 7373 10978 7439 10981
rect 10961 10980 11027 10981
rect 10910 10978 10916 10980
rect 6932 10976 7439 10978
rect 6932 10920 7378 10976
rect 7434 10920 7439 10976
rect 6932 10918 7439 10920
rect 10870 10918 10916 10978
rect 10980 10976 11027 10980
rect 11022 10920 11027 10976
rect 6932 10916 6938 10918
rect 7373 10915 7439 10918
rect 10910 10916 10916 10918
rect 10980 10916 11027 10920
rect 10961 10915 11027 10916
rect 15653 10978 15719 10981
rect 16246 10978 16252 10980
rect 15653 10976 16252 10978
rect 15653 10920 15658 10976
rect 15714 10920 16252 10976
rect 15653 10918 16252 10920
rect 15653 10915 15719 10918
rect 16246 10916 16252 10918
rect 16316 10916 16322 10980
rect 22185 10978 22251 10981
rect 22840 10978 23300 11008
rect 22185 10976 23300 10978
rect 22185 10920 22190 10976
rect 22246 10920 23300 10976
rect 22185 10918 23300 10920
rect 22185 10915 22251 10918
rect 6144 10912 6460 10913
rect 6144 10848 6150 10912
rect 6214 10848 6230 10912
rect 6294 10848 6310 10912
rect 6374 10848 6390 10912
rect 6454 10848 6460 10912
rect 6144 10847 6460 10848
rect 11342 10912 11658 10913
rect 11342 10848 11348 10912
rect 11412 10848 11428 10912
rect 11492 10848 11508 10912
rect 11572 10848 11588 10912
rect 11652 10848 11658 10912
rect 11342 10847 11658 10848
rect 16540 10912 16856 10913
rect 16540 10848 16546 10912
rect 16610 10848 16626 10912
rect 16690 10848 16706 10912
rect 16770 10848 16786 10912
rect 16850 10848 16856 10912
rect 16540 10847 16856 10848
rect 21738 10912 22054 10913
rect 21738 10848 21744 10912
rect 21808 10848 21824 10912
rect 21888 10848 21904 10912
rect 21968 10848 21984 10912
rect 22048 10848 22054 10912
rect 22840 10888 23300 10918
rect 21738 10847 22054 10848
rect 8150 10780 8156 10844
rect 8220 10842 8226 10844
rect 10869 10842 10935 10845
rect 8220 10840 10935 10842
rect 8220 10784 10874 10840
rect 10930 10784 10935 10840
rect 8220 10782 10935 10784
rect 8220 10780 8226 10782
rect 10869 10779 10935 10782
rect 6085 10706 6151 10709
rect 5950 10704 6151 10706
rect 5950 10648 6090 10704
rect 6146 10648 6151 10704
rect 5950 10646 6151 10648
rect 4153 10643 4219 10646
rect 5625 10643 5691 10646
rect 6085 10643 6151 10646
rect 6821 10706 6887 10709
rect 11789 10706 11855 10709
rect 6821 10704 11855 10706
rect 6821 10648 6826 10704
rect 6882 10648 11794 10704
rect 11850 10648 11855 10704
rect 6821 10646 11855 10648
rect 6821 10643 6887 10646
rect 11789 10643 11855 10646
rect 14273 10706 14339 10709
rect 19609 10706 19675 10709
rect 14273 10704 19675 10706
rect 14273 10648 14278 10704
rect 14334 10648 19614 10704
rect 19670 10648 19675 10704
rect 14273 10646 19675 10648
rect 14273 10643 14339 10646
rect 19609 10643 19675 10646
rect 21265 10706 21331 10709
rect 21633 10706 21699 10709
rect 21265 10704 21699 10706
rect 21265 10648 21270 10704
rect 21326 10648 21638 10704
rect 21694 10648 21699 10704
rect 21265 10646 21699 10648
rect 21265 10643 21331 10646
rect 21633 10643 21699 10646
rect 2998 10508 3004 10572
rect 3068 10570 3074 10572
rect 4797 10570 4863 10573
rect 9489 10570 9555 10573
rect 10777 10572 10843 10573
rect 3068 10510 4722 10570
rect 3068 10508 3074 10510
rect -300 10434 160 10464
rect 4662 10434 4722 10510
rect 4797 10568 9555 10570
rect 4797 10512 4802 10568
rect 4858 10512 9494 10568
rect 9550 10512 9555 10568
rect 4797 10510 9555 10512
rect 4797 10507 4863 10510
rect 9489 10507 9555 10510
rect 10726 10508 10732 10572
rect 10796 10570 10843 10572
rect 10796 10568 10888 10570
rect 10838 10512 10888 10568
rect 10796 10510 10888 10512
rect 10796 10508 10843 10510
rect 13302 10508 13308 10572
rect 13372 10570 13378 10572
rect 20294 10570 20300 10572
rect 13372 10510 20300 10570
rect 13372 10508 13378 10510
rect 20294 10508 20300 10510
rect 20364 10508 20370 10572
rect 10777 10507 10843 10508
rect 6913 10434 6979 10437
rect -300 10374 3434 10434
rect 4662 10432 6979 10434
rect 4662 10376 6918 10432
rect 6974 10376 6979 10432
rect 4662 10374 6979 10376
rect -300 10344 160 10374
rect 1025 10298 1091 10301
rect 3049 10298 3115 10301
rect 1025 10296 3115 10298
rect 1025 10240 1030 10296
rect 1086 10240 3054 10296
rect 3110 10240 3115 10296
rect 1025 10238 3115 10240
rect 1025 10235 1091 10238
rect 3049 10235 3115 10238
rect -300 10162 160 10192
rect 2773 10162 2839 10165
rect -300 10160 2839 10162
rect -300 10104 2778 10160
rect 2834 10104 2839 10160
rect -300 10102 2839 10104
rect 3374 10162 3434 10374
rect 6913 10371 6979 10374
rect 11237 10434 11303 10437
rect 12198 10434 12204 10436
rect 11237 10432 12204 10434
rect 11237 10376 11242 10432
rect 11298 10376 12204 10432
rect 11237 10374 12204 10376
rect 11237 10371 11303 10374
rect 12198 10372 12204 10374
rect 12268 10372 12274 10436
rect 20897 10434 20963 10437
rect 22840 10434 23300 10464
rect 20897 10432 23300 10434
rect 20897 10376 20902 10432
rect 20958 10376 23300 10432
rect 20897 10374 23300 10376
rect 20897 10371 20963 10374
rect 3545 10368 3861 10369
rect 3545 10304 3551 10368
rect 3615 10304 3631 10368
rect 3695 10304 3711 10368
rect 3775 10304 3791 10368
rect 3855 10304 3861 10368
rect 3545 10303 3861 10304
rect 8743 10368 9059 10369
rect 8743 10304 8749 10368
rect 8813 10304 8829 10368
rect 8893 10304 8909 10368
rect 8973 10304 8989 10368
rect 9053 10304 9059 10368
rect 8743 10303 9059 10304
rect 13941 10368 14257 10369
rect 13941 10304 13947 10368
rect 14011 10304 14027 10368
rect 14091 10304 14107 10368
rect 14171 10304 14187 10368
rect 14251 10304 14257 10368
rect 13941 10303 14257 10304
rect 19139 10368 19455 10369
rect 19139 10304 19145 10368
rect 19209 10304 19225 10368
rect 19289 10304 19305 10368
rect 19369 10304 19385 10368
rect 19449 10304 19455 10368
rect 22840 10344 23300 10374
rect 19139 10303 19455 10304
rect 5390 10236 5396 10300
rect 5460 10298 5466 10300
rect 6545 10298 6611 10301
rect 5460 10296 6611 10298
rect 5460 10240 6550 10296
rect 6606 10240 6611 10296
rect 5460 10238 6611 10240
rect 5460 10236 5466 10238
rect 6545 10235 6611 10238
rect 10961 10298 11027 10301
rect 16297 10298 16363 10301
rect 10961 10296 13738 10298
rect 10961 10240 10966 10296
rect 11022 10240 13738 10296
rect 10961 10238 13738 10240
rect 10961 10235 11027 10238
rect 3969 10162 4035 10165
rect 13537 10162 13603 10165
rect 3374 10160 4035 10162
rect 3374 10104 3974 10160
rect 4030 10104 4035 10160
rect 3374 10102 4035 10104
rect -300 10072 160 10102
rect 2773 10099 2839 10102
rect 3969 10099 4035 10102
rect 4294 10160 13603 10162
rect 4294 10104 13542 10160
rect 13598 10104 13603 10160
rect 4294 10102 13603 10104
rect 13678 10162 13738 10238
rect 14414 10296 16363 10298
rect 14414 10240 16302 10296
rect 16358 10240 16363 10296
rect 14414 10238 16363 10240
rect 14414 10162 14474 10238
rect 16297 10235 16363 10238
rect 13678 10102 14474 10162
rect 14549 10162 14615 10165
rect 16757 10162 16823 10165
rect 14549 10160 16823 10162
rect 14549 10104 14554 10160
rect 14610 10104 16762 10160
rect 16818 10104 16823 10160
rect 14549 10102 16823 10104
rect 4294 10026 4354 10102
rect 13537 10099 13603 10102
rect 14549 10099 14615 10102
rect 16757 10099 16823 10102
rect 2730 9966 4354 10026
rect 4797 10024 4863 10029
rect 4797 9968 4802 10024
rect 4858 9968 4863 10024
rect -300 9890 160 9920
rect 1669 9890 1735 9893
rect -300 9888 1735 9890
rect -300 9832 1674 9888
rect 1730 9832 1735 9888
rect -300 9830 1735 9832
rect -300 9800 160 9830
rect 1669 9827 1735 9830
rect 2221 9754 2287 9757
rect 2730 9754 2790 9966
rect 4797 9963 4863 9968
rect 5073 10026 5139 10029
rect 13486 10026 13492 10028
rect 5073 10024 13492 10026
rect 5073 9968 5078 10024
rect 5134 9968 13492 10024
rect 5073 9966 13492 9968
rect 5073 9963 5139 9966
rect 4800 9890 4860 9963
rect 5073 9892 5139 9893
rect 2221 9752 2790 9754
rect 2221 9696 2226 9752
rect 2282 9696 2790 9752
rect 2221 9694 2790 9696
rect 3558 9830 4860 9890
rect 2221 9691 2287 9694
rect -300 9618 160 9648
rect 3325 9618 3391 9621
rect 3558 9618 3618 9830
rect 5022 9828 5028 9892
rect 5092 9890 5139 9892
rect 5092 9888 5184 9890
rect 5134 9832 5184 9888
rect 5092 9830 5184 9832
rect 5092 9828 5139 9830
rect 5073 9827 5139 9828
rect 6144 9824 6460 9825
rect 6144 9760 6150 9824
rect 6214 9760 6230 9824
rect 6294 9760 6310 9824
rect 6374 9760 6390 9824
rect 6454 9760 6460 9824
rect 6144 9759 6460 9760
rect 11342 9824 11658 9825
rect 11342 9760 11348 9824
rect 11412 9760 11428 9824
rect 11492 9760 11508 9824
rect 11572 9760 11588 9824
rect 11652 9760 11658 9824
rect 11342 9759 11658 9760
rect 12528 9757 12588 9966
rect 13486 9964 13492 9966
rect 13556 9964 13562 10028
rect 13670 9964 13676 10028
rect 13740 10026 13746 10028
rect 14641 10026 14707 10029
rect 13740 10024 14707 10026
rect 13740 9968 14646 10024
rect 14702 9968 14707 10024
rect 13740 9966 14707 9968
rect 13740 9964 13746 9966
rect 14641 9963 14707 9966
rect 17677 10026 17743 10029
rect 18413 10026 18479 10029
rect 17677 10024 18479 10026
rect 17677 9968 17682 10024
rect 17738 9968 18418 10024
rect 18474 9968 18479 10024
rect 17677 9966 18479 9968
rect 17677 9963 17743 9966
rect 18413 9963 18479 9966
rect 12985 9888 13051 9893
rect 12985 9832 12990 9888
rect 13046 9832 13051 9888
rect 12985 9827 13051 9832
rect 22277 9890 22343 9893
rect 22840 9890 23300 9920
rect 22277 9888 23300 9890
rect 22277 9832 22282 9888
rect 22338 9832 23300 9888
rect 22277 9830 23300 9832
rect 22277 9827 22343 9830
rect 3877 9754 3943 9757
rect 5625 9754 5691 9757
rect 7005 9754 7071 9757
rect 8334 9754 8340 9756
rect 3877 9752 5458 9754
rect 3877 9696 3882 9752
rect 3938 9696 5458 9752
rect 3877 9694 5458 9696
rect 3877 9691 3943 9694
rect -300 9616 3391 9618
rect -300 9560 3330 9616
rect 3386 9560 3391 9616
rect -300 9558 3391 9560
rect -300 9528 160 9558
rect 3325 9555 3391 9558
rect 3512 9558 3618 9618
rect 5398 9618 5458 9694
rect 5625 9752 6010 9754
rect 5625 9696 5630 9752
rect 5686 9696 6010 9752
rect 5625 9694 6010 9696
rect 5625 9691 5691 9694
rect 5717 9618 5783 9621
rect 5398 9616 5783 9618
rect 5398 9560 5722 9616
rect 5778 9560 5783 9616
rect 5398 9558 5783 9560
rect 5950 9618 6010 9694
rect 7005 9752 8340 9754
rect 7005 9696 7010 9752
rect 7066 9696 8340 9752
rect 7005 9694 8340 9696
rect 7005 9691 7071 9694
rect 8334 9692 8340 9694
rect 8404 9692 8410 9756
rect 8753 9754 8819 9757
rect 10501 9754 10567 9757
rect 8753 9752 10567 9754
rect 8753 9696 8758 9752
rect 8814 9696 10506 9752
rect 10562 9696 10567 9752
rect 8753 9694 10567 9696
rect 8753 9691 8819 9694
rect 10501 9691 10567 9694
rect 12525 9752 12591 9757
rect 12988 9754 13048 9827
rect 16540 9824 16856 9825
rect 16540 9760 16546 9824
rect 16610 9760 16626 9824
rect 16690 9760 16706 9824
rect 16770 9760 16786 9824
rect 16850 9760 16856 9824
rect 16540 9759 16856 9760
rect 21738 9824 22054 9825
rect 21738 9760 21744 9824
rect 21808 9760 21824 9824
rect 21888 9760 21904 9824
rect 21968 9760 21984 9824
rect 22048 9760 22054 9824
rect 22840 9800 23300 9830
rect 21738 9759 22054 9760
rect 12525 9696 12530 9752
rect 12586 9696 12591 9752
rect 12525 9691 12591 9696
rect 12804 9694 13048 9754
rect 13353 9754 13419 9757
rect 14774 9754 14780 9756
rect 13353 9752 14780 9754
rect 13353 9696 13358 9752
rect 13414 9696 14780 9752
rect 13353 9694 14780 9696
rect 7649 9618 7715 9621
rect 11973 9618 12039 9621
rect 5950 9558 6930 9618
rect 1485 9482 1551 9485
rect 3512 9482 3572 9558
rect 5717 9555 5783 9558
rect 1485 9480 3572 9482
rect 1485 9424 1490 9480
rect 1546 9424 3572 9480
rect 1485 9422 3572 9424
rect 6870 9485 6930 9558
rect 7649 9616 12039 9618
rect 7649 9560 7654 9616
rect 7710 9560 11978 9616
rect 12034 9560 12039 9616
rect 7649 9558 12039 9560
rect 7649 9555 7715 9558
rect 11973 9555 12039 9558
rect 6870 9482 6979 9485
rect 7557 9482 7623 9485
rect 6870 9480 7623 9482
rect 6870 9424 6918 9480
rect 6974 9424 7562 9480
rect 7618 9424 7623 9480
rect 6870 9422 7623 9424
rect 1485 9419 1551 9422
rect 6913 9419 6979 9422
rect 7557 9419 7623 9422
rect 11789 9482 11855 9485
rect 12804 9482 12864 9694
rect 13353 9691 13419 9694
rect 14774 9692 14780 9694
rect 14844 9692 14850 9756
rect 18873 9754 18939 9757
rect 19926 9754 19932 9756
rect 18873 9752 19932 9754
rect 18873 9696 18878 9752
rect 18934 9696 19932 9752
rect 18873 9694 19932 9696
rect 18873 9691 18939 9694
rect 19926 9692 19932 9694
rect 19996 9692 20002 9756
rect 12985 9618 13051 9621
rect 15285 9618 15351 9621
rect 12985 9616 15351 9618
rect 12985 9560 12990 9616
rect 13046 9560 15290 9616
rect 15346 9560 15351 9616
rect 12985 9558 15351 9560
rect 12985 9555 13051 9558
rect 15285 9555 15351 9558
rect 16021 9618 16087 9621
rect 16982 9618 16988 9620
rect 16021 9616 16988 9618
rect 16021 9560 16026 9616
rect 16082 9560 16988 9616
rect 16021 9558 16988 9560
rect 16021 9555 16087 9558
rect 16982 9556 16988 9558
rect 17052 9556 17058 9620
rect 19006 9556 19012 9620
rect 19076 9618 19082 9620
rect 19241 9618 19307 9621
rect 19076 9616 19307 9618
rect 19076 9560 19246 9616
rect 19302 9560 19307 9616
rect 19076 9558 19307 9560
rect 19076 9556 19082 9558
rect 19241 9555 19307 9558
rect 17166 9482 17172 9484
rect 11789 9480 17172 9482
rect 11789 9424 11794 9480
rect 11850 9424 17172 9480
rect 11789 9422 17172 9424
rect 11789 9419 11855 9422
rect 17166 9420 17172 9422
rect 17236 9420 17242 9484
rect 20478 9482 20484 9484
rect 19014 9422 20484 9482
rect -300 9346 160 9376
rect 1577 9346 1643 9349
rect -300 9344 1643 9346
rect -300 9288 1582 9344
rect 1638 9288 1643 9344
rect -300 9286 1643 9288
rect -300 9256 160 9286
rect 1577 9283 1643 9286
rect 2497 9346 2563 9349
rect 2630 9346 2636 9348
rect 2497 9344 2636 9346
rect 2497 9288 2502 9344
rect 2558 9288 2636 9344
rect 2497 9286 2636 9288
rect 2497 9283 2563 9286
rect 2630 9284 2636 9286
rect 2700 9284 2706 9348
rect 4705 9346 4771 9349
rect 5717 9346 5783 9349
rect 4705 9344 5783 9346
rect 4705 9288 4710 9344
rect 4766 9288 5722 9344
rect 5778 9288 5783 9344
rect 4705 9286 5783 9288
rect 4705 9283 4771 9286
rect 5717 9283 5783 9286
rect 11881 9346 11947 9349
rect 12341 9346 12407 9349
rect 13445 9346 13511 9349
rect 11881 9344 13511 9346
rect 11881 9288 11886 9344
rect 11942 9288 12346 9344
rect 12402 9288 13450 9344
rect 13506 9288 13511 9344
rect 11881 9286 13511 9288
rect 11881 9283 11947 9286
rect 12341 9283 12407 9286
rect 13445 9283 13511 9286
rect 15009 9346 15075 9349
rect 19014 9346 19074 9422
rect 20478 9420 20484 9422
rect 20548 9420 20554 9484
rect 15009 9344 19074 9346
rect 15009 9288 15014 9344
rect 15070 9288 19074 9344
rect 15009 9286 19074 9288
rect 21449 9346 21515 9349
rect 22840 9346 23300 9376
rect 21449 9344 23300 9346
rect 21449 9288 21454 9344
rect 21510 9288 23300 9344
rect 21449 9286 23300 9288
rect 15009 9283 15075 9286
rect 21449 9283 21515 9286
rect 3545 9280 3861 9281
rect 3545 9216 3551 9280
rect 3615 9216 3631 9280
rect 3695 9216 3711 9280
rect 3775 9216 3791 9280
rect 3855 9216 3861 9280
rect 3545 9215 3861 9216
rect 8743 9280 9059 9281
rect 8743 9216 8749 9280
rect 8813 9216 8829 9280
rect 8893 9216 8909 9280
rect 8973 9216 8989 9280
rect 9053 9216 9059 9280
rect 8743 9215 9059 9216
rect 13941 9280 14257 9281
rect 13941 9216 13947 9280
rect 14011 9216 14027 9280
rect 14091 9216 14107 9280
rect 14171 9216 14187 9280
rect 14251 9216 14257 9280
rect 13941 9215 14257 9216
rect 19139 9280 19455 9281
rect 19139 9216 19145 9280
rect 19209 9216 19225 9280
rect 19289 9216 19305 9280
rect 19369 9216 19385 9280
rect 19449 9216 19455 9280
rect 22840 9256 23300 9286
rect 19139 9215 19455 9216
rect 3969 9210 4035 9213
rect 4286 9210 4292 9212
rect 3969 9208 4292 9210
rect 3969 9152 3974 9208
rect 4030 9152 4292 9208
rect 3969 9150 4292 9152
rect 3969 9147 4035 9150
rect 4286 9148 4292 9150
rect 4356 9148 4362 9212
rect -300 9074 160 9104
rect 4705 9074 4771 9077
rect -300 9072 4771 9074
rect -300 9016 4710 9072
rect 4766 9016 4771 9072
rect -300 9014 4771 9016
rect -300 8984 160 9014
rect 4705 9011 4771 9014
rect 5758 9012 5764 9076
rect 5828 9074 5834 9076
rect 6453 9074 6519 9077
rect 5828 9072 6519 9074
rect 5828 9016 6458 9072
rect 6514 9016 6519 9072
rect 5828 9014 6519 9016
rect 5828 9012 5834 9014
rect 6453 9011 6519 9014
rect 10041 9074 10107 9077
rect 12341 9074 12407 9077
rect 10041 9072 12407 9074
rect 10041 9016 10046 9072
rect 10102 9016 12346 9072
rect 12402 9016 12407 9072
rect 10041 9014 12407 9016
rect 10041 9011 10107 9014
rect 12341 9011 12407 9014
rect 12709 9074 12775 9077
rect 15837 9074 15903 9077
rect 12709 9072 15903 9074
rect 12709 9016 12714 9072
rect 12770 9016 15842 9072
rect 15898 9016 15903 9072
rect 12709 9014 15903 9016
rect 12709 9011 12775 9014
rect 15837 9011 15903 9014
rect 16246 9012 16252 9076
rect 16316 9074 16322 9076
rect 18597 9074 18663 9077
rect 16316 9072 18663 9074
rect 16316 9016 18602 9072
rect 18658 9016 18663 9072
rect 16316 9014 18663 9016
rect 16316 9012 16322 9014
rect 18597 9011 18663 9014
rect 19057 9074 19123 9077
rect 19057 9072 22202 9074
rect 19057 9016 19062 9072
rect 19118 9016 22202 9072
rect 19057 9014 22202 9016
rect 19057 9011 19123 9014
rect 7649 8938 7715 8941
rect 17125 8938 17191 8941
rect 2730 8936 17191 8938
rect 2730 8880 7654 8936
rect 7710 8880 17130 8936
rect 17186 8880 17191 8936
rect 2730 8878 17191 8880
rect -300 8802 160 8832
rect 1393 8802 1459 8805
rect 2446 8802 2452 8804
rect -300 8800 1459 8802
rect -300 8744 1398 8800
rect 1454 8744 1459 8800
rect -300 8742 1459 8744
rect -300 8712 160 8742
rect 1393 8739 1459 8742
rect 2086 8742 2452 8802
rect 1761 8666 1827 8669
rect 2086 8666 2146 8742
rect 2446 8740 2452 8742
rect 2516 8802 2522 8804
rect 2730 8802 2790 8878
rect 7649 8875 7715 8878
rect 17125 8875 17191 8878
rect 19333 8938 19399 8941
rect 20253 8938 20319 8941
rect 19333 8936 20319 8938
rect 19333 8880 19338 8936
rect 19394 8880 20258 8936
rect 20314 8880 20319 8936
rect 19333 8878 20319 8880
rect 19333 8875 19399 8878
rect 20253 8875 20319 8878
rect 4061 8802 4127 8805
rect 2516 8742 2790 8802
rect 3236 8800 4127 8802
rect 3236 8744 4066 8800
rect 4122 8744 4127 8800
rect 3236 8742 4127 8744
rect 2516 8740 2522 8742
rect 1761 8664 2146 8666
rect 1761 8608 1766 8664
rect 1822 8608 2146 8664
rect 1761 8606 2146 8608
rect 1761 8603 1827 8606
rect 2262 8604 2268 8668
rect 2332 8666 2338 8668
rect 3236 8666 3296 8742
rect 4061 8739 4127 8742
rect 12198 8740 12204 8804
rect 12268 8740 12274 8804
rect 12934 8740 12940 8804
rect 13004 8802 13010 8804
rect 16389 8802 16455 8805
rect 13004 8800 16455 8802
rect 13004 8744 16394 8800
rect 16450 8744 16455 8800
rect 13004 8742 16455 8744
rect 22142 8802 22202 9014
rect 22840 8802 23300 8832
rect 22142 8742 23300 8802
rect 13004 8740 13010 8742
rect 6144 8736 6460 8737
rect 6144 8672 6150 8736
rect 6214 8672 6230 8736
rect 6294 8672 6310 8736
rect 6374 8672 6390 8736
rect 6454 8672 6460 8736
rect 6144 8671 6460 8672
rect 11342 8736 11658 8737
rect 11342 8672 11348 8736
rect 11412 8672 11428 8736
rect 11492 8672 11508 8736
rect 11572 8672 11588 8736
rect 11652 8672 11658 8736
rect 11342 8671 11658 8672
rect 2332 8606 3296 8666
rect 2332 8604 2338 8606
rect 3366 8604 3372 8668
rect 3436 8666 3442 8668
rect 4470 8666 4476 8668
rect 3436 8606 4476 8666
rect 3436 8604 3442 8606
rect 4470 8604 4476 8606
rect 4540 8604 4546 8668
rect 5349 8666 5415 8669
rect 4800 8664 5415 8666
rect 4800 8608 5354 8664
rect 5410 8608 5415 8664
rect 4800 8606 5415 8608
rect -300 8530 160 8560
rect 4800 8530 4860 8606
rect 5349 8603 5415 8606
rect 6862 8604 6868 8668
rect 6932 8666 6938 8668
rect 7005 8666 7071 8669
rect 6932 8664 7071 8666
rect 6932 8608 7010 8664
rect 7066 8608 7071 8664
rect 6932 8606 7071 8608
rect 6932 8604 6938 8606
rect 7005 8603 7071 8606
rect 8569 8666 8635 8669
rect 10041 8666 10107 8669
rect 8569 8664 10107 8666
rect 8569 8608 8574 8664
rect 8630 8608 10046 8664
rect 10102 8608 10107 8664
rect 8569 8606 10107 8608
rect 12206 8666 12266 8740
rect 16389 8739 16455 8742
rect 16540 8736 16856 8737
rect 16540 8672 16546 8736
rect 16610 8672 16626 8736
rect 16690 8672 16706 8736
rect 16770 8672 16786 8736
rect 16850 8672 16856 8736
rect 16540 8671 16856 8672
rect 21738 8736 22054 8737
rect 21738 8672 21744 8736
rect 21808 8672 21824 8736
rect 21888 8672 21904 8736
rect 21968 8672 21984 8736
rect 22048 8672 22054 8736
rect 22840 8712 23300 8742
rect 21738 8671 22054 8672
rect 14181 8666 14247 8669
rect 14733 8666 14799 8669
rect 12206 8664 14799 8666
rect 12206 8608 14186 8664
rect 14242 8608 14738 8664
rect 14794 8608 14799 8664
rect 12206 8606 14799 8608
rect 8569 8603 8635 8606
rect 10041 8603 10107 8606
rect 14181 8603 14247 8606
rect 14733 8603 14799 8606
rect -300 8470 4860 8530
rect -300 8440 160 8470
rect 5022 8468 5028 8532
rect 5092 8530 5098 8532
rect 6269 8530 6335 8533
rect 9622 8530 9628 8532
rect 5092 8528 9628 8530
rect 5092 8472 6274 8528
rect 6330 8472 9628 8528
rect 5092 8470 9628 8472
rect 5092 8468 5098 8470
rect 6269 8467 6335 8470
rect 9622 8468 9628 8470
rect 9692 8530 9698 8532
rect 17953 8530 18019 8533
rect 9692 8528 18019 8530
rect 9692 8472 17958 8528
rect 18014 8472 18019 8528
rect 9692 8470 18019 8472
rect 9692 8468 9698 8470
rect 17953 8467 18019 8470
rect 1393 8394 1459 8397
rect 3182 8394 3188 8396
rect 1393 8392 3188 8394
rect 1393 8336 1398 8392
rect 1454 8336 3188 8392
rect 1393 8334 3188 8336
rect 1393 8331 1459 8334
rect 3182 8332 3188 8334
rect 3252 8332 3258 8396
rect 3366 8332 3372 8396
rect 3436 8394 3442 8396
rect 4521 8394 4587 8397
rect 3436 8392 4587 8394
rect 3436 8336 4526 8392
rect 4582 8336 4587 8392
rect 3436 8334 4587 8336
rect 3436 8332 3442 8334
rect 4521 8331 4587 8334
rect 8017 8394 8083 8397
rect 8334 8394 8340 8396
rect 8017 8392 8340 8394
rect 8017 8336 8022 8392
rect 8078 8336 8340 8392
rect 8017 8334 8340 8336
rect 8017 8331 8083 8334
rect 8334 8332 8340 8334
rect 8404 8332 8410 8396
rect 9438 8332 9444 8396
rect 9508 8394 9514 8396
rect 9581 8394 9647 8397
rect 9508 8392 9647 8394
rect 9508 8336 9586 8392
rect 9642 8336 9647 8392
rect 9508 8334 9647 8336
rect 9508 8332 9514 8334
rect 9581 8331 9647 8334
rect 12433 8394 12499 8397
rect 12934 8394 12940 8396
rect 12433 8392 12940 8394
rect 12433 8336 12438 8392
rect 12494 8336 12940 8392
rect 12433 8334 12940 8336
rect 12433 8331 12499 8334
rect 12934 8332 12940 8334
rect 13004 8332 13010 8396
rect 13118 8332 13124 8396
rect 13188 8394 13194 8396
rect 13261 8394 13327 8397
rect 13188 8392 13327 8394
rect 13188 8336 13266 8392
rect 13322 8336 13327 8392
rect 13188 8334 13327 8336
rect 13188 8332 13194 8334
rect 13261 8331 13327 8334
rect 14733 8394 14799 8397
rect 17534 8394 17540 8396
rect 14733 8392 17540 8394
rect 14733 8336 14738 8392
rect 14794 8336 17540 8392
rect 14733 8334 17540 8336
rect 14733 8331 14799 8334
rect 17534 8332 17540 8334
rect 17604 8332 17610 8396
rect -300 8258 160 8288
rect -300 8198 1410 8258
rect -300 8168 160 8198
rect 1350 8122 1410 8198
rect 2446 8196 2452 8260
rect 2516 8258 2522 8260
rect 3325 8258 3391 8261
rect 5206 8258 5212 8260
rect 2516 8256 3391 8258
rect 2516 8200 3330 8256
rect 3386 8200 3391 8256
rect 2516 8198 3391 8200
rect 2516 8196 2522 8198
rect 3325 8195 3391 8198
rect 4524 8198 5212 8258
rect 3545 8192 3861 8193
rect 3545 8128 3551 8192
rect 3615 8128 3631 8192
rect 3695 8128 3711 8192
rect 3775 8128 3791 8192
rect 3855 8128 3861 8192
rect 3545 8127 3861 8128
rect 4524 8125 4584 8198
rect 5206 8196 5212 8198
rect 5276 8258 5282 8260
rect 10777 8258 10843 8261
rect 14825 8258 14891 8261
rect 18965 8258 19031 8261
rect 22840 8258 23300 8288
rect 5276 8198 8632 8258
rect 5276 8196 5282 8198
rect 2405 8122 2471 8125
rect 1350 8120 2471 8122
rect 1350 8064 2410 8120
rect 2466 8064 2471 8120
rect 1350 8062 2471 8064
rect 2405 8059 2471 8062
rect 4521 8120 4587 8125
rect 4521 8064 4526 8120
rect 4582 8064 4587 8120
rect 4521 8059 4587 8064
rect 5257 8122 5323 8125
rect 7373 8122 7439 8125
rect 5257 8120 7439 8122
rect 5257 8064 5262 8120
rect 5318 8064 7378 8120
rect 7434 8064 7439 8120
rect 5257 8062 7439 8064
rect 5257 8059 5323 8062
rect 7373 8059 7439 8062
rect -300 7986 160 8016
rect 1485 7986 1551 7989
rect 8385 7986 8451 7989
rect -300 7926 1226 7986
rect -300 7896 160 7926
rect 1166 7850 1226 7926
rect 1485 7984 8451 7986
rect 1485 7928 1490 7984
rect 1546 7928 8390 7984
rect 8446 7928 8451 7984
rect 1485 7926 8451 7928
rect 8572 7986 8632 8198
rect 10777 8256 13738 8258
rect 10777 8200 10782 8256
rect 10838 8200 13738 8256
rect 10777 8198 13738 8200
rect 10777 8195 10843 8198
rect 8743 8192 9059 8193
rect 8743 8128 8749 8192
rect 8813 8128 8829 8192
rect 8893 8128 8909 8192
rect 8973 8128 8989 8192
rect 9053 8128 9059 8192
rect 8743 8127 9059 8128
rect 10044 8062 12404 8122
rect 10044 7986 10104 8062
rect 8572 7926 10104 7986
rect 1485 7923 1551 7926
rect 8385 7923 8451 7926
rect 10174 7924 10180 7988
rect 10244 7986 10250 7988
rect 12198 7986 12204 7988
rect 10244 7926 12204 7986
rect 10244 7924 10250 7926
rect 12198 7924 12204 7926
rect 12268 7924 12274 7988
rect 2129 7850 2195 7853
rect 3233 7852 3299 7853
rect 3182 7850 3188 7852
rect 1166 7848 2195 7850
rect 1166 7792 2134 7848
rect 2190 7792 2195 7848
rect 1166 7790 2195 7792
rect 3142 7790 3188 7850
rect 3252 7848 3299 7852
rect 3294 7792 3299 7848
rect 2129 7787 2195 7790
rect 3182 7788 3188 7790
rect 3252 7788 3299 7792
rect 3233 7787 3299 7788
rect 3785 7850 3851 7853
rect 6821 7850 6887 7853
rect 3785 7848 6887 7850
rect 3785 7792 3790 7848
rect 3846 7792 6826 7848
rect 6882 7792 6887 7848
rect 3785 7790 6887 7792
rect 3785 7787 3851 7790
rect 6821 7787 6887 7790
rect 7097 7850 7163 7853
rect 8845 7850 8911 7853
rect 7097 7848 8911 7850
rect 7097 7792 7102 7848
rect 7158 7792 8850 7848
rect 8906 7792 8911 7848
rect 7097 7790 8911 7792
rect 7097 7787 7163 7790
rect 8845 7787 8911 7790
rect 9489 7850 9555 7853
rect 12344 7850 12404 8062
rect 13678 7986 13738 8198
rect 14825 8256 19031 8258
rect 14825 8200 14830 8256
rect 14886 8200 18970 8256
rect 19026 8200 19031 8256
rect 14825 8198 19031 8200
rect 14825 8195 14891 8198
rect 18965 8195 19031 8198
rect 20670 8198 23300 8258
rect 13941 8192 14257 8193
rect 13941 8128 13947 8192
rect 14011 8128 14027 8192
rect 14091 8128 14107 8192
rect 14171 8128 14187 8192
rect 14251 8128 14257 8192
rect 13941 8127 14257 8128
rect 19139 8192 19455 8193
rect 19139 8128 19145 8192
rect 19209 8128 19225 8192
rect 19289 8128 19305 8192
rect 19369 8128 19385 8192
rect 19449 8128 19455 8192
rect 19139 8127 19455 8128
rect 18873 8122 18939 8125
rect 14368 8120 18939 8122
rect 14368 8064 18878 8120
rect 18934 8064 18939 8120
rect 14368 8062 18939 8064
rect 14368 7986 14428 8062
rect 18873 8059 18939 8062
rect 19793 7986 19859 7989
rect 13678 7926 14428 7986
rect 14552 7984 19859 7986
rect 14552 7928 19798 7984
rect 19854 7928 19859 7984
rect 14552 7926 19859 7928
rect 13997 7850 14063 7853
rect 14552 7850 14612 7926
rect 19793 7923 19859 7926
rect 16021 7850 16087 7853
rect 18045 7850 18111 7853
rect 9489 7848 11852 7850
rect 9489 7792 9494 7848
rect 9550 7792 11852 7848
rect 9489 7790 11852 7792
rect 12344 7848 14612 7850
rect 12344 7792 14002 7848
rect 14058 7792 14612 7848
rect 12344 7790 14612 7792
rect 15104 7848 16087 7850
rect 15104 7792 16026 7848
rect 16082 7792 16087 7848
rect 15104 7790 16087 7792
rect 9489 7787 9555 7790
rect -300 7714 160 7744
rect 4153 7714 4219 7717
rect 6729 7714 6795 7717
rect 8753 7714 8819 7717
rect -300 7654 2790 7714
rect -300 7624 160 7654
rect 1485 7578 1551 7581
rect 2078 7578 2084 7580
rect 1485 7576 2084 7578
rect 1485 7520 1490 7576
rect 1546 7520 2084 7576
rect 1485 7518 2084 7520
rect 1485 7515 1551 7518
rect 2078 7516 2084 7518
rect 2148 7516 2154 7580
rect 2730 7578 2790 7654
rect 4153 7712 5826 7714
rect 4153 7656 4158 7712
rect 4214 7656 5826 7712
rect 4153 7654 5826 7656
rect 4153 7651 4219 7654
rect 5766 7580 5826 7654
rect 6729 7712 8819 7714
rect 6729 7656 6734 7712
rect 6790 7656 8758 7712
rect 8814 7656 8819 7712
rect 6729 7654 8819 7656
rect 11792 7714 11852 7790
rect 13997 7787 14063 7790
rect 15104 7714 15164 7790
rect 16021 7787 16087 7790
rect 16254 7848 18111 7850
rect 16254 7792 18050 7848
rect 18106 7792 18111 7848
rect 16254 7790 18111 7792
rect 11792 7654 15164 7714
rect 15285 7714 15351 7717
rect 16254 7714 16314 7790
rect 18045 7787 18111 7790
rect 18413 7850 18479 7853
rect 20670 7850 20730 8198
rect 22840 8168 23300 8198
rect 18413 7848 20730 7850
rect 18413 7792 18418 7848
rect 18474 7792 20730 7848
rect 18413 7790 20730 7792
rect 18413 7787 18479 7790
rect 15285 7712 16314 7714
rect 15285 7656 15290 7712
rect 15346 7656 16314 7712
rect 15285 7654 16314 7656
rect 18781 7716 18847 7717
rect 18781 7712 18828 7716
rect 18892 7714 18898 7716
rect 22840 7714 23300 7744
rect 18781 7656 18786 7712
rect 6729 7651 6795 7654
rect 8753 7651 8819 7654
rect 15285 7651 15351 7654
rect 18781 7652 18828 7656
rect 18892 7654 18938 7714
rect 22142 7654 23300 7714
rect 18892 7652 18898 7654
rect 18781 7651 18847 7652
rect 6144 7648 6460 7649
rect 6144 7584 6150 7648
rect 6214 7584 6230 7648
rect 6294 7584 6310 7648
rect 6374 7584 6390 7648
rect 6454 7584 6460 7648
rect 6144 7583 6460 7584
rect 11342 7648 11658 7649
rect 11342 7584 11348 7648
rect 11412 7584 11428 7648
rect 11492 7584 11508 7648
rect 11572 7584 11588 7648
rect 11652 7584 11658 7648
rect 11342 7583 11658 7584
rect 16540 7648 16856 7649
rect 16540 7584 16546 7648
rect 16610 7584 16626 7648
rect 16690 7584 16706 7648
rect 16770 7584 16786 7648
rect 16850 7584 16856 7648
rect 16540 7583 16856 7584
rect 21738 7648 22054 7649
rect 21738 7584 21744 7648
rect 21808 7584 21824 7648
rect 21888 7584 21904 7648
rect 21968 7584 21984 7648
rect 22048 7584 22054 7648
rect 21738 7583 22054 7584
rect 2730 7518 4354 7578
rect -300 7442 160 7472
rect 4153 7442 4219 7445
rect -300 7440 4219 7442
rect -300 7384 4158 7440
rect 4214 7384 4219 7440
rect -300 7382 4219 7384
rect 4294 7442 4354 7518
rect 4470 7516 4476 7580
rect 4540 7578 4546 7580
rect 5574 7578 5580 7580
rect 4540 7518 5580 7578
rect 4540 7516 4546 7518
rect 5574 7516 5580 7518
rect 5644 7516 5650 7580
rect 5758 7516 5764 7580
rect 5828 7516 5834 7580
rect 12065 7578 12131 7581
rect 13302 7578 13308 7580
rect 12065 7576 13308 7578
rect 12065 7520 12070 7576
rect 12126 7520 13308 7576
rect 12065 7518 13308 7520
rect 12065 7515 12131 7518
rect 13302 7516 13308 7518
rect 13372 7516 13378 7580
rect 14549 7578 14615 7581
rect 16389 7578 16455 7581
rect 14549 7576 16455 7578
rect 14549 7520 14554 7576
rect 14610 7520 16394 7576
rect 16450 7520 16455 7576
rect 14549 7518 16455 7520
rect 14549 7515 14615 7518
rect 16389 7515 16455 7518
rect 4429 7442 4495 7445
rect 4294 7440 4495 7442
rect 4294 7384 4434 7440
rect 4490 7384 4495 7440
rect 4294 7382 4495 7384
rect -300 7352 160 7382
rect 4153 7379 4219 7382
rect 4429 7379 4495 7382
rect 4705 7442 4771 7445
rect 7833 7442 7899 7445
rect 4705 7440 7899 7442
rect 4705 7384 4710 7440
rect 4766 7384 7838 7440
rect 7894 7384 7899 7440
rect 4705 7382 7899 7384
rect 4705 7379 4771 7382
rect 7833 7379 7899 7382
rect 10225 7442 10291 7445
rect 17033 7442 17099 7445
rect 21541 7442 21607 7445
rect 10225 7440 17099 7442
rect 10225 7384 10230 7440
rect 10286 7384 17038 7440
rect 17094 7384 17099 7440
rect 10225 7382 17099 7384
rect 10225 7379 10291 7382
rect 17033 7379 17099 7382
rect 18094 7440 21607 7442
rect 18094 7384 21546 7440
rect 21602 7384 21607 7440
rect 18094 7382 21607 7384
rect 1025 7306 1091 7309
rect 1894 7306 1900 7308
rect 1025 7304 1900 7306
rect 1025 7248 1030 7304
rect 1086 7248 1900 7304
rect 1025 7246 1900 7248
rect 1025 7243 1091 7246
rect 1894 7244 1900 7246
rect 1964 7244 1970 7308
rect 2865 7306 2931 7309
rect 11094 7306 11100 7308
rect 2865 7304 11100 7306
rect 2865 7248 2870 7304
rect 2926 7248 11100 7304
rect 2865 7246 11100 7248
rect 2865 7243 2931 7246
rect 11094 7244 11100 7246
rect 11164 7244 11170 7308
rect 12525 7306 12591 7309
rect 12893 7306 12959 7309
rect 17769 7306 17835 7309
rect 12525 7304 12634 7306
rect 12525 7248 12530 7304
rect 12586 7248 12634 7304
rect 12525 7243 12634 7248
rect 12893 7304 17835 7306
rect 12893 7248 12898 7304
rect 12954 7248 17774 7304
rect 17830 7248 17835 7304
rect 12893 7246 17835 7248
rect 12893 7243 12959 7246
rect 17769 7243 17835 7246
rect -300 7170 160 7200
rect 2221 7172 2287 7173
rect -300 7110 858 7170
rect -300 7080 160 7110
rect 798 7034 858 7110
rect 2221 7168 2268 7172
rect 2332 7170 2338 7172
rect 4521 7170 4587 7173
rect 5441 7170 5507 7173
rect 6085 7170 6151 7173
rect 6913 7170 6979 7173
rect 2221 7112 2226 7168
rect 2221 7108 2268 7112
rect 2332 7110 2378 7170
rect 4294 7168 6979 7170
rect 4294 7112 4526 7168
rect 4582 7112 5446 7168
rect 5502 7112 6090 7168
rect 6146 7112 6918 7168
rect 6974 7112 6979 7168
rect 4294 7110 6979 7112
rect 2332 7108 2338 7110
rect 2221 7107 2287 7108
rect 3545 7104 3861 7105
rect 3545 7040 3551 7104
rect 3615 7040 3631 7104
rect 3695 7040 3711 7104
rect 3775 7040 3791 7104
rect 3855 7040 3861 7104
rect 3545 7039 3861 7040
rect 1761 7034 1827 7037
rect 4294 7036 4354 7110
rect 4521 7107 4587 7110
rect 5441 7107 5507 7110
rect 6085 7107 6151 7110
rect 6913 7107 6979 7110
rect 12341 7170 12407 7173
rect 12574 7170 12634 7243
rect 12341 7168 12634 7170
rect 12341 7112 12346 7168
rect 12402 7112 12634 7168
rect 12341 7110 12634 7112
rect 12341 7107 12407 7110
rect 8743 7104 9059 7105
rect 8743 7040 8749 7104
rect 8813 7040 8829 7104
rect 8893 7040 8909 7104
rect 8973 7040 8989 7104
rect 9053 7040 9059 7104
rect 8743 7039 9059 7040
rect 13941 7104 14257 7105
rect 13941 7040 13947 7104
rect 14011 7040 14027 7104
rect 14091 7040 14107 7104
rect 14171 7040 14187 7104
rect 14251 7040 14257 7104
rect 13941 7039 14257 7040
rect 798 7032 1827 7034
rect 798 6976 1766 7032
rect 1822 6976 1827 7032
rect 798 6974 1827 6976
rect 1761 6971 1827 6974
rect 4286 6972 4292 7036
rect 4356 6972 4362 7036
rect 4654 6972 4660 7036
rect 4724 7034 4730 7036
rect 4981 7034 5047 7037
rect 7046 7034 7052 7036
rect 4724 7032 5047 7034
rect 4724 6976 4986 7032
rect 5042 6976 5047 7032
rect 4724 6974 5047 6976
rect 4724 6972 4730 6974
rect 4981 6971 5047 6974
rect 5582 6974 7052 7034
rect -300 6898 160 6928
rect 4061 6898 4127 6901
rect -300 6896 4127 6898
rect -300 6840 4066 6896
rect 4122 6840 4127 6896
rect -300 6838 4127 6840
rect -300 6808 160 6838
rect 4061 6835 4127 6838
rect 4245 6898 4311 6901
rect 5206 6898 5212 6900
rect 4245 6896 5212 6898
rect 4245 6840 4250 6896
rect 4306 6840 5212 6896
rect 4245 6838 5212 6840
rect 4245 6835 4311 6838
rect 5206 6836 5212 6838
rect 5276 6836 5282 6900
rect 5441 6898 5507 6901
rect 5582 6898 5642 6974
rect 7046 6972 7052 6974
rect 7116 7034 7122 7036
rect 7741 7034 7807 7037
rect 7116 7032 7807 7034
rect 7116 6976 7746 7032
rect 7802 6976 7807 7032
rect 7116 6974 7807 6976
rect 7116 6972 7122 6974
rect 7741 6971 7807 6974
rect 10961 7034 11027 7037
rect 12249 7034 12315 7037
rect 18094 7034 18154 7382
rect 21541 7379 21607 7382
rect 18965 7306 19031 7309
rect 22142 7306 22202 7654
rect 22840 7624 23300 7654
rect 18965 7304 22202 7306
rect 18965 7248 18970 7304
rect 19026 7248 22202 7304
rect 18965 7246 22202 7248
rect 18965 7243 19031 7246
rect 22840 7170 23300 7200
rect 19566 7110 23300 7170
rect 19139 7104 19455 7105
rect 19139 7040 19145 7104
rect 19209 7040 19225 7104
rect 19289 7040 19305 7104
rect 19369 7040 19385 7104
rect 19449 7040 19455 7104
rect 19139 7039 19455 7040
rect 10961 7032 12315 7034
rect 10961 6976 10966 7032
rect 11022 6976 12254 7032
rect 12310 6976 12315 7032
rect 10961 6974 12315 6976
rect 10961 6971 11027 6974
rect 12249 6971 12315 6974
rect 12390 6974 13002 7034
rect 5441 6896 5642 6898
rect 5441 6840 5446 6896
rect 5502 6840 5642 6896
rect 5441 6838 5642 6840
rect 5441 6835 5507 6838
rect 5758 6836 5764 6900
rect 5828 6898 5834 6900
rect 5901 6898 5967 6901
rect 5828 6896 5967 6898
rect 5828 6840 5906 6896
rect 5962 6840 5967 6896
rect 5828 6838 5967 6840
rect 5828 6836 5834 6838
rect 5901 6835 5967 6838
rect 7598 6836 7604 6900
rect 7668 6898 7674 6900
rect 12390 6898 12450 6974
rect 7668 6838 12450 6898
rect 12525 6898 12591 6901
rect 12750 6898 12756 6900
rect 12525 6896 12756 6898
rect 12525 6840 12530 6896
rect 12586 6840 12756 6896
rect 12525 6838 12756 6840
rect 7668 6836 7674 6838
rect 12525 6835 12591 6838
rect 12750 6836 12756 6838
rect 12820 6836 12826 6900
rect 12942 6898 13002 6974
rect 15104 6974 18154 7034
rect 18873 7034 18939 7037
rect 18873 7032 19074 7034
rect 18873 6976 18878 7032
rect 18934 6976 19074 7032
rect 18873 6974 19074 6976
rect 15104 6901 15164 6974
rect 18873 6971 18939 6974
rect 14406 6898 14412 6900
rect 12942 6838 14412 6898
rect 14406 6836 14412 6838
rect 14476 6836 14482 6900
rect 15101 6896 15167 6901
rect 15101 6840 15106 6896
rect 15162 6840 15167 6896
rect 15101 6835 15167 6840
rect 19014 6898 19074 6974
rect 19566 6898 19626 7110
rect 22840 7080 23300 7110
rect 19014 6838 19626 6898
rect 2497 6762 2563 6765
rect 2814 6762 2820 6764
rect 2497 6760 2820 6762
rect 2497 6704 2502 6760
rect 2558 6704 2820 6760
rect 2497 6702 2820 6704
rect 2497 6699 2563 6702
rect 2814 6700 2820 6702
rect 2884 6700 2890 6764
rect 2998 6700 3004 6764
rect 3068 6762 3074 6764
rect 3325 6762 3391 6765
rect 3068 6760 3391 6762
rect 3068 6704 3330 6760
rect 3386 6704 3391 6760
rect 3068 6702 3391 6704
rect 3068 6700 3074 6702
rect 3325 6699 3391 6702
rect 3785 6762 3851 6765
rect 3918 6762 3924 6764
rect 3785 6760 3924 6762
rect 3785 6704 3790 6760
rect 3846 6704 3924 6760
rect 3785 6702 3924 6704
rect 3785 6699 3851 6702
rect 3918 6700 3924 6702
rect 3988 6700 3994 6764
rect 4245 6762 4311 6765
rect 4613 6762 4679 6765
rect 21173 6762 21239 6765
rect 4245 6760 21239 6762
rect 4245 6704 4250 6760
rect 4306 6704 4618 6760
rect 4674 6704 21178 6760
rect 21234 6704 21239 6760
rect 4245 6702 21239 6704
rect 4245 6699 4311 6702
rect 4613 6699 4679 6702
rect 21173 6699 21239 6702
rect 21590 6702 22202 6762
rect -300 6626 160 6656
rect -300 6566 2514 6626
rect -300 6536 160 6566
rect -300 6354 160 6384
rect 2454 6357 2514 6566
rect 2630 6564 2636 6628
rect 2700 6626 2706 6628
rect 4470 6626 4476 6628
rect 2700 6566 4476 6626
rect 2700 6564 2706 6566
rect 4470 6564 4476 6566
rect 4540 6564 4546 6628
rect 4613 6626 4679 6629
rect 5441 6626 5507 6629
rect 4613 6624 5507 6626
rect 4613 6568 4618 6624
rect 4674 6568 5446 6624
rect 5502 6568 5507 6624
rect 4613 6566 5507 6568
rect 4613 6563 4679 6566
rect 5441 6563 5507 6566
rect 7833 6626 7899 6629
rect 10358 6626 10364 6628
rect 7833 6624 10364 6626
rect 7833 6568 7838 6624
rect 7894 6568 10364 6624
rect 7833 6566 10364 6568
rect 7833 6563 7899 6566
rect 10358 6564 10364 6566
rect 10428 6564 10434 6628
rect 14273 6626 14339 6629
rect 12390 6624 14339 6626
rect 12390 6568 14278 6624
rect 14334 6568 14339 6624
rect 12390 6566 14339 6568
rect 3877 6490 3943 6493
rect 4616 6490 4676 6563
rect 6144 6560 6460 6561
rect 6144 6496 6150 6560
rect 6214 6496 6230 6560
rect 6294 6496 6310 6560
rect 6374 6496 6390 6560
rect 6454 6496 6460 6560
rect 6144 6495 6460 6496
rect 11342 6560 11658 6561
rect 11342 6496 11348 6560
rect 11412 6496 11428 6560
rect 11492 6496 11508 6560
rect 11572 6496 11588 6560
rect 11652 6496 11658 6560
rect 11342 6495 11658 6496
rect 3877 6488 4676 6490
rect 3877 6432 3882 6488
rect 3938 6432 4676 6488
rect 3877 6430 4676 6432
rect 3877 6427 3943 6430
rect 1209 6354 1275 6357
rect -300 6352 1275 6354
rect -300 6296 1214 6352
rect 1270 6296 1275 6352
rect -300 6294 1275 6296
rect 2454 6352 2563 6357
rect 2454 6296 2502 6352
rect 2558 6296 2563 6352
rect 2454 6294 2563 6296
rect -300 6264 160 6294
rect 1209 6291 1275 6294
rect 2497 6291 2563 6294
rect 4153 6354 4219 6357
rect 5257 6354 5323 6357
rect 4153 6352 5323 6354
rect 4153 6296 4158 6352
rect 4214 6296 5262 6352
rect 5318 6296 5323 6352
rect 4153 6294 5323 6296
rect 4153 6291 4219 6294
rect 5257 6291 5323 6294
rect 5390 6292 5396 6356
rect 5460 6354 5466 6356
rect 12390 6354 12450 6566
rect 14273 6563 14339 6566
rect 17493 6626 17559 6629
rect 21590 6626 21650 6702
rect 17493 6624 21650 6626
rect 17493 6568 17498 6624
rect 17554 6568 21650 6624
rect 17493 6566 21650 6568
rect 22142 6626 22202 6702
rect 22840 6626 23300 6656
rect 22142 6566 23300 6626
rect 17493 6563 17559 6566
rect 16540 6560 16856 6561
rect 16540 6496 16546 6560
rect 16610 6496 16626 6560
rect 16690 6496 16706 6560
rect 16770 6496 16786 6560
rect 16850 6496 16856 6560
rect 16540 6495 16856 6496
rect 21738 6560 22054 6561
rect 21738 6496 21744 6560
rect 21808 6496 21824 6560
rect 21888 6496 21904 6560
rect 21968 6496 21984 6560
rect 22048 6496 22054 6560
rect 22840 6536 23300 6566
rect 21738 6495 22054 6496
rect 18229 6490 18295 6493
rect 19149 6490 19215 6493
rect 18229 6488 19215 6490
rect 18229 6432 18234 6488
rect 18290 6432 19154 6488
rect 19210 6432 19215 6488
rect 18229 6430 19215 6432
rect 18229 6427 18295 6430
rect 19149 6427 19215 6430
rect 5460 6294 12450 6354
rect 5460 6292 5466 6294
rect 15142 6292 15148 6356
rect 15212 6354 15218 6356
rect 18229 6354 18295 6357
rect 15212 6352 18295 6354
rect 15212 6296 18234 6352
rect 18290 6296 18295 6352
rect 15212 6294 18295 6296
rect 15212 6292 15218 6294
rect 18229 6291 18295 6294
rect 18689 6354 18755 6357
rect 19241 6354 19307 6357
rect 18689 6352 19307 6354
rect 18689 6296 18694 6352
rect 18750 6296 19246 6352
rect 19302 6296 19307 6352
rect 18689 6294 19307 6296
rect 18689 6291 18755 6294
rect 19241 6291 19307 6294
rect 2405 6218 2471 6221
rect 2773 6218 2839 6221
rect 2405 6216 2839 6218
rect 2405 6160 2410 6216
rect 2466 6160 2778 6216
rect 2834 6160 2839 6216
rect 2405 6158 2839 6160
rect 2405 6155 2471 6158
rect 2773 6155 2839 6158
rect 3509 6218 3575 6221
rect 4429 6218 4495 6221
rect 6177 6218 6243 6221
rect 3509 6216 4354 6218
rect 3509 6160 3514 6216
rect 3570 6160 4354 6216
rect 3509 6158 4354 6160
rect 3509 6155 3575 6158
rect -300 6082 160 6112
rect 2814 6082 2820 6084
rect -300 6022 2820 6082
rect -300 5992 160 6022
rect 2814 6020 2820 6022
rect 2884 6020 2890 6084
rect 4294 6082 4354 6158
rect 4429 6216 6243 6218
rect 4429 6160 4434 6216
rect 4490 6160 6182 6216
rect 6238 6160 6243 6216
rect 4429 6158 6243 6160
rect 4429 6155 4495 6158
rect 6177 6155 6243 6158
rect 6637 6218 6703 6221
rect 7373 6218 7439 6221
rect 10174 6218 10180 6220
rect 6637 6216 10180 6218
rect 6637 6160 6642 6216
rect 6698 6160 7378 6216
rect 7434 6160 10180 6216
rect 6637 6158 10180 6160
rect 6637 6155 6703 6158
rect 7373 6155 7439 6158
rect 10174 6156 10180 6158
rect 10244 6156 10250 6220
rect 10777 6218 10843 6221
rect 14549 6218 14615 6221
rect 18086 6218 18092 6220
rect 10777 6216 14428 6218
rect 10777 6160 10782 6216
rect 10838 6160 14428 6216
rect 10777 6158 14428 6160
rect 10777 6155 10843 6158
rect 5993 6082 6059 6085
rect 4294 6080 6059 6082
rect 4294 6024 5998 6080
rect 6054 6024 6059 6080
rect 4294 6022 6059 6024
rect 5993 6019 6059 6022
rect 6269 6082 6335 6085
rect 8385 6082 8451 6085
rect 6269 6080 8451 6082
rect 6269 6024 6274 6080
rect 6330 6024 8390 6080
rect 8446 6024 8451 6080
rect 6269 6022 8451 6024
rect 6269 6019 6335 6022
rect 8385 6019 8451 6022
rect 9765 6082 9831 6085
rect 12801 6082 12867 6085
rect 9765 6080 12867 6082
rect 9765 6024 9770 6080
rect 9826 6024 12806 6080
rect 12862 6024 12867 6080
rect 9765 6022 12867 6024
rect 14368 6082 14428 6158
rect 14549 6216 18092 6218
rect 14549 6160 14554 6216
rect 14610 6160 18092 6216
rect 14549 6158 18092 6160
rect 14549 6155 14615 6158
rect 18086 6156 18092 6158
rect 18156 6156 18162 6220
rect 18600 6158 19626 6218
rect 18600 6085 18660 6158
rect 14368 6022 15808 6082
rect 9765 6019 9831 6022
rect 12801 6019 12867 6022
rect 3545 6016 3861 6017
rect 3545 5952 3551 6016
rect 3615 5952 3631 6016
rect 3695 5952 3711 6016
rect 3775 5952 3791 6016
rect 3855 5952 3861 6016
rect 3545 5951 3861 5952
rect 8743 6016 9059 6017
rect 8743 5952 8749 6016
rect 8813 5952 8829 6016
rect 8893 5952 8909 6016
rect 8973 5952 8989 6016
rect 9053 5952 9059 6016
rect 8743 5951 9059 5952
rect 13941 6016 14257 6017
rect 13941 5952 13947 6016
rect 14011 5952 14027 6016
rect 14091 5952 14107 6016
rect 14171 5952 14187 6016
rect 14251 5952 14257 6016
rect 13941 5951 14257 5952
rect 15748 5949 15808 6022
rect 18597 6080 18663 6085
rect 18597 6024 18602 6080
rect 18658 6024 18663 6080
rect 18597 6019 18663 6024
rect 19566 6082 19626 6158
rect 22840 6082 23300 6112
rect 19566 6022 23300 6082
rect 19139 6016 19455 6017
rect 19139 5952 19145 6016
rect 19209 5952 19225 6016
rect 19289 5952 19305 6016
rect 19369 5952 19385 6016
rect 19449 5952 19455 6016
rect 22840 5992 23300 6022
rect 19139 5951 19455 5952
rect 15745 5946 15811 5949
rect 18689 5946 18755 5949
rect 15745 5944 18755 5946
rect 15745 5888 15750 5944
rect 15806 5888 18694 5944
rect 18750 5888 18755 5944
rect 15745 5886 18755 5888
rect 15745 5883 15811 5886
rect 18689 5883 18755 5886
rect -300 5810 160 5840
rect 4061 5810 4127 5813
rect -300 5808 4127 5810
rect -300 5752 4066 5808
rect 4122 5752 4127 5808
rect -300 5750 4127 5752
rect -300 5720 160 5750
rect 4061 5747 4127 5750
rect 4470 5748 4476 5812
rect 4540 5810 4546 5812
rect 15101 5810 15167 5813
rect 20161 5810 20227 5813
rect 20989 5810 21055 5813
rect 4540 5750 12450 5810
rect 4540 5748 4546 5750
rect 2497 5674 2563 5677
rect 3325 5674 3391 5677
rect 2497 5672 3391 5674
rect 2497 5616 2502 5672
rect 2558 5616 3330 5672
rect 3386 5616 3391 5672
rect 2497 5614 3391 5616
rect 2497 5611 2563 5614
rect 3325 5611 3391 5614
rect 4153 5674 4219 5677
rect 8937 5674 9003 5677
rect 4153 5672 9003 5674
rect 4153 5616 4158 5672
rect 4214 5616 8942 5672
rect 8998 5616 9003 5672
rect 4153 5614 9003 5616
rect 4153 5611 4219 5614
rect 8937 5611 9003 5614
rect 9622 5612 9628 5676
rect 9692 5674 9698 5676
rect 10961 5674 11027 5677
rect 9692 5672 11027 5674
rect 9692 5616 10966 5672
rect 11022 5616 11027 5672
rect 9692 5614 11027 5616
rect 12390 5674 12450 5750
rect 15101 5808 21055 5810
rect 15101 5752 15106 5808
rect 15162 5752 20166 5808
rect 20222 5752 20994 5808
rect 21050 5752 21055 5808
rect 15101 5750 21055 5752
rect 15101 5747 15167 5750
rect 20161 5747 20227 5750
rect 20989 5747 21055 5750
rect 18321 5674 18387 5677
rect 12390 5672 18387 5674
rect 12390 5616 18326 5672
rect 18382 5616 18387 5672
rect 12390 5614 18387 5616
rect 9692 5612 9698 5614
rect 10961 5611 11027 5614
rect 18321 5611 18387 5614
rect 18781 5674 18847 5677
rect 19006 5674 19012 5676
rect 18781 5672 19012 5674
rect 18781 5616 18786 5672
rect 18842 5616 19012 5672
rect 18781 5614 19012 5616
rect 18781 5611 18847 5614
rect 19006 5612 19012 5614
rect 19076 5674 19082 5676
rect 19149 5674 19215 5677
rect 22369 5674 22435 5677
rect 19076 5672 19215 5674
rect 19076 5616 19154 5672
rect 19210 5616 19215 5672
rect 19076 5614 19215 5616
rect 19076 5612 19082 5614
rect 19149 5611 19215 5614
rect 21590 5672 22435 5674
rect 21590 5616 22374 5672
rect 22430 5616 22435 5672
rect 21590 5614 22435 5616
rect -300 5538 160 5568
rect 4061 5538 4127 5541
rect -300 5536 4127 5538
rect -300 5480 4066 5536
rect 4122 5480 4127 5536
rect -300 5478 4127 5480
rect -300 5448 160 5478
rect 4061 5475 4127 5478
rect 12157 5538 12223 5541
rect 15561 5538 15627 5541
rect 12157 5536 15627 5538
rect 12157 5480 12162 5536
rect 12218 5480 15566 5536
rect 15622 5480 15627 5536
rect 12157 5478 15627 5480
rect 12157 5475 12223 5478
rect 15561 5475 15627 5478
rect 18413 5540 18479 5541
rect 18413 5536 18460 5540
rect 18524 5538 18530 5540
rect 21590 5538 21650 5614
rect 22369 5611 22435 5614
rect 22840 5538 23300 5568
rect 18413 5480 18418 5536
rect 18413 5476 18460 5480
rect 18524 5478 18570 5538
rect 19382 5478 21650 5538
rect 22142 5478 23300 5538
rect 18524 5476 18530 5478
rect 18413 5475 18479 5476
rect 6144 5472 6460 5473
rect 6144 5408 6150 5472
rect 6214 5408 6230 5472
rect 6294 5408 6310 5472
rect 6374 5408 6390 5472
rect 6454 5408 6460 5472
rect 6144 5407 6460 5408
rect 11342 5472 11658 5473
rect 11342 5408 11348 5472
rect 11412 5408 11428 5472
rect 11492 5408 11508 5472
rect 11572 5408 11588 5472
rect 11652 5408 11658 5472
rect 11342 5407 11658 5408
rect 16540 5472 16856 5473
rect 16540 5408 16546 5472
rect 16610 5408 16626 5472
rect 16690 5408 16706 5472
rect 16770 5408 16786 5472
rect 16850 5408 16856 5472
rect 16540 5407 16856 5408
rect 1485 5402 1551 5405
rect 3366 5402 3372 5404
rect 1485 5400 3372 5402
rect 1485 5344 1490 5400
rect 1546 5344 3372 5400
rect 1485 5342 3372 5344
rect 1485 5339 1551 5342
rect 3366 5340 3372 5342
rect 3436 5340 3442 5404
rect 17718 5340 17724 5404
rect 17788 5402 17794 5404
rect 19382 5402 19442 5478
rect 21738 5472 22054 5473
rect 21738 5408 21744 5472
rect 21808 5408 21824 5472
rect 21888 5408 21904 5472
rect 21968 5408 21984 5472
rect 22048 5408 22054 5472
rect 21738 5407 22054 5408
rect 17788 5342 19442 5402
rect 17788 5340 17794 5342
rect -300 5266 160 5296
rect 4061 5266 4127 5269
rect -300 5264 4127 5266
rect -300 5208 4066 5264
rect 4122 5208 4127 5264
rect -300 5206 4127 5208
rect -300 5176 160 5206
rect 4061 5203 4127 5206
rect 5993 5266 6059 5269
rect 12249 5266 12315 5269
rect 13169 5266 13235 5269
rect 5993 5264 12315 5266
rect 5993 5208 5998 5264
rect 6054 5208 12254 5264
rect 12310 5208 12315 5264
rect 5993 5206 12315 5208
rect 5993 5203 6059 5206
rect 12249 5203 12315 5206
rect 12390 5264 13235 5266
rect 12390 5208 13174 5264
rect 13230 5208 13235 5264
rect 12390 5206 13235 5208
rect 1853 5130 1919 5133
rect 3049 5130 3115 5133
rect 5022 5130 5028 5132
rect 1853 5128 2790 5130
rect 1853 5072 1858 5128
rect 1914 5072 2790 5128
rect 1853 5070 2790 5072
rect 1853 5067 1919 5070
rect -300 4994 160 5024
rect -300 4934 674 4994
rect -300 4904 160 4934
rect 614 4722 674 4934
rect 1301 4722 1367 4725
rect 614 4720 1367 4722
rect 614 4664 1306 4720
rect 1362 4664 1367 4720
rect 614 4662 1367 4664
rect 2730 4722 2790 5070
rect 3049 5128 5028 5130
rect 3049 5072 3054 5128
rect 3110 5072 5028 5128
rect 3049 5070 5028 5072
rect 3049 5067 3115 5070
rect 5022 5068 5028 5070
rect 5092 5068 5098 5132
rect 5206 5068 5212 5132
rect 5276 5130 5282 5132
rect 12390 5130 12450 5206
rect 13169 5203 13235 5206
rect 14549 5266 14615 5269
rect 22142 5266 22202 5478
rect 22840 5448 23300 5478
rect 14549 5264 22202 5266
rect 14549 5208 14554 5264
rect 14610 5208 22202 5264
rect 14549 5206 22202 5208
rect 14549 5203 14615 5206
rect 5276 5070 12450 5130
rect 15377 5130 15443 5133
rect 15377 5128 19626 5130
rect 15377 5072 15382 5128
rect 15438 5072 19626 5128
rect 15377 5070 19626 5072
rect 5276 5068 5282 5070
rect 15377 5067 15443 5070
rect 4889 4994 4955 4997
rect 7373 4994 7439 4997
rect 4889 4992 7439 4994
rect 4889 4936 4894 4992
rect 4950 4936 7378 4992
rect 7434 4936 7439 4992
rect 4889 4934 7439 4936
rect 4889 4931 4955 4934
rect 7373 4931 7439 4934
rect 15929 4994 15995 4997
rect 18413 4994 18479 4997
rect 15929 4992 18479 4994
rect 15929 4936 15934 4992
rect 15990 4936 18418 4992
rect 18474 4936 18479 4992
rect 15929 4934 18479 4936
rect 19566 4994 19626 5070
rect 22840 4994 23300 5024
rect 19566 4934 23300 4994
rect 15929 4931 15995 4934
rect 18413 4931 18479 4934
rect 3545 4928 3861 4929
rect 3545 4864 3551 4928
rect 3615 4864 3631 4928
rect 3695 4864 3711 4928
rect 3775 4864 3791 4928
rect 3855 4864 3861 4928
rect 3545 4863 3861 4864
rect 8743 4928 9059 4929
rect 8743 4864 8749 4928
rect 8813 4864 8829 4928
rect 8893 4864 8909 4928
rect 8973 4864 8989 4928
rect 9053 4864 9059 4928
rect 8743 4863 9059 4864
rect 13941 4928 14257 4929
rect 13941 4864 13947 4928
rect 14011 4864 14027 4928
rect 14091 4864 14107 4928
rect 14171 4864 14187 4928
rect 14251 4864 14257 4928
rect 13941 4863 14257 4864
rect 19139 4928 19455 4929
rect 19139 4864 19145 4928
rect 19209 4864 19225 4928
rect 19289 4864 19305 4928
rect 19369 4864 19385 4928
rect 19449 4864 19455 4928
rect 22840 4904 23300 4934
rect 19139 4863 19455 4864
rect 14917 4858 14983 4861
rect 18597 4858 18663 4861
rect 14917 4856 18663 4858
rect 14917 4800 14922 4856
rect 14978 4800 18602 4856
rect 18658 4800 18663 4856
rect 14917 4798 18663 4800
rect 14917 4795 14983 4798
rect 18597 4795 18663 4798
rect 9213 4722 9279 4725
rect 2730 4720 9279 4722
rect 2730 4664 9218 4720
rect 9274 4664 9279 4720
rect 2730 4662 9279 4664
rect 1301 4659 1367 4662
rect 9213 4659 9279 4662
rect 15561 4722 15627 4725
rect 21081 4722 21147 4725
rect 15561 4720 21147 4722
rect 15561 4664 15566 4720
rect 15622 4664 21086 4720
rect 21142 4664 21147 4720
rect 15561 4662 21147 4664
rect 15561 4659 15627 4662
rect 21081 4659 21147 4662
rect 2446 4524 2452 4588
rect 2516 4586 2522 4588
rect 2681 4586 2747 4589
rect 2516 4584 2747 4586
rect 2516 4528 2686 4584
rect 2742 4528 2747 4584
rect 2516 4526 2747 4528
rect 2516 4524 2522 4526
rect 2681 4523 2747 4526
rect 3601 4586 3667 4589
rect 4337 4588 4403 4589
rect 4102 4586 4108 4588
rect 3601 4584 4108 4586
rect 3601 4528 3606 4584
rect 3662 4528 4108 4584
rect 3601 4526 4108 4528
rect 3601 4523 3667 4526
rect 4102 4524 4108 4526
rect 4172 4524 4178 4588
rect 4286 4524 4292 4588
rect 4356 4586 4403 4588
rect 4981 4586 5047 4589
rect 4356 4584 4448 4586
rect 4398 4528 4448 4584
rect 4356 4526 4448 4528
rect 4981 4584 6746 4586
rect 4981 4528 4986 4584
rect 5042 4528 6746 4584
rect 4981 4526 6746 4528
rect 4356 4524 4403 4526
rect 4337 4523 4403 4524
rect 4981 4523 5047 4526
rect 3693 4450 3759 4453
rect 4654 4450 4660 4452
rect 3693 4448 4660 4450
rect 3693 4392 3698 4448
rect 3754 4392 4660 4448
rect 3693 4390 4660 4392
rect 3693 4387 3759 4390
rect 4654 4388 4660 4390
rect 4724 4388 4730 4452
rect 6686 4450 6746 4526
rect 8150 4524 8156 4588
rect 8220 4586 8226 4588
rect 12566 4586 12572 4588
rect 8220 4526 12572 4586
rect 8220 4524 8226 4526
rect 12566 4524 12572 4526
rect 12636 4524 12642 4588
rect 16113 4586 16179 4589
rect 19517 4586 19583 4589
rect 16113 4584 19583 4586
rect 16113 4528 16118 4584
rect 16174 4528 19522 4584
rect 19578 4528 19583 4584
rect 16113 4526 19583 4528
rect 16113 4523 16179 4526
rect 19517 4523 19583 4526
rect 21590 4526 22202 4586
rect 10542 4450 10548 4452
rect 6686 4390 10548 4450
rect 10542 4388 10548 4390
rect 10612 4388 10618 4452
rect 13629 4450 13695 4453
rect 16297 4450 16363 4453
rect 13629 4448 16363 4450
rect 13629 4392 13634 4448
rect 13690 4392 16302 4448
rect 16358 4392 16363 4448
rect 13629 4390 16363 4392
rect 13629 4387 13695 4390
rect 16297 4387 16363 4390
rect 17217 4450 17283 4453
rect 18229 4450 18295 4453
rect 17217 4448 18295 4450
rect 17217 4392 17222 4448
rect 17278 4392 18234 4448
rect 18290 4392 18295 4448
rect 17217 4390 18295 4392
rect 17217 4387 17283 4390
rect 18229 4387 18295 4390
rect 18638 4388 18644 4452
rect 18708 4450 18714 4452
rect 21590 4450 21650 4526
rect 18708 4390 21650 4450
rect 22142 4450 22202 4526
rect 22840 4450 23300 4480
rect 22142 4390 23300 4450
rect 18708 4388 18714 4390
rect 6144 4384 6460 4385
rect 6144 4320 6150 4384
rect 6214 4320 6230 4384
rect 6294 4320 6310 4384
rect 6374 4320 6390 4384
rect 6454 4320 6460 4384
rect 6144 4319 6460 4320
rect 11342 4384 11658 4385
rect 11342 4320 11348 4384
rect 11412 4320 11428 4384
rect 11492 4320 11508 4384
rect 11572 4320 11588 4384
rect 11652 4320 11658 4384
rect 11342 4319 11658 4320
rect 16540 4384 16856 4385
rect 16540 4320 16546 4384
rect 16610 4320 16626 4384
rect 16690 4320 16706 4384
rect 16770 4320 16786 4384
rect 16850 4320 16856 4384
rect 16540 4319 16856 4320
rect 21738 4384 22054 4385
rect 21738 4320 21744 4384
rect 21808 4320 21824 4384
rect 21888 4320 21904 4384
rect 21968 4320 21984 4384
rect 22048 4320 22054 4384
rect 22840 4360 23300 4390
rect 21738 4319 22054 4320
rect 14590 4314 14596 4316
rect 12390 4254 14596 4314
rect 4102 4116 4108 4180
rect 4172 4178 4178 4180
rect 12390 4178 12450 4254
rect 14590 4252 14596 4254
rect 14660 4252 14666 4316
rect 18229 4314 18295 4317
rect 20069 4314 20135 4317
rect 18229 4312 20135 4314
rect 18229 4256 18234 4312
rect 18290 4256 20074 4312
rect 20130 4256 20135 4312
rect 18229 4254 20135 4256
rect 18229 4251 18295 4254
rect 20069 4251 20135 4254
rect 4172 4118 12450 4178
rect 14733 4178 14799 4181
rect 21357 4178 21423 4181
rect 14733 4176 21423 4178
rect 14733 4120 14738 4176
rect 14794 4120 21362 4176
rect 21418 4120 21423 4176
rect 14733 4118 21423 4120
rect 4172 4116 4178 4118
rect 14733 4115 14799 4118
rect 21357 4115 21423 4118
rect 5165 4042 5231 4045
rect 7465 4042 7531 4045
rect 5165 4040 7531 4042
rect 5165 3984 5170 4040
rect 5226 3984 7470 4040
rect 7526 3984 7531 4040
rect 5165 3982 7531 3984
rect 5165 3979 5231 3982
rect 7465 3979 7531 3982
rect 15653 4044 15719 4045
rect 15653 4040 15700 4044
rect 15764 4042 15770 4044
rect 18045 4042 18111 4045
rect 15653 3984 15658 4040
rect 15653 3980 15700 3984
rect 15764 3982 15810 4042
rect 15886 4040 18111 4042
rect 15886 3984 18050 4040
rect 18106 3984 18111 4040
rect 15886 3982 18111 3984
rect 15764 3980 15770 3982
rect 15653 3979 15719 3980
rect 5574 3844 5580 3908
rect 5644 3906 5650 3908
rect 7281 3906 7347 3909
rect 5644 3904 7347 3906
rect 5644 3848 7286 3904
rect 7342 3848 7347 3904
rect 5644 3846 7347 3848
rect 5644 3844 5650 3846
rect 7281 3843 7347 3846
rect 14641 3906 14707 3909
rect 15886 3906 15946 3982
rect 18045 3979 18111 3982
rect 18229 4044 18295 4045
rect 18229 4040 18276 4044
rect 18340 4042 18346 4044
rect 19241 4042 19307 4045
rect 20069 4044 20135 4045
rect 20069 4042 20116 4044
rect 18229 3984 18234 4040
rect 18229 3980 18276 3984
rect 18340 3982 18386 4042
rect 19241 4040 19810 4042
rect 19241 3984 19246 4040
rect 19302 3984 19810 4040
rect 19241 3982 19810 3984
rect 20024 4040 20116 4042
rect 20024 3984 20074 4040
rect 20024 3982 20116 3984
rect 18340 3980 18346 3982
rect 18229 3979 18295 3980
rect 19241 3979 19307 3982
rect 14641 3904 15946 3906
rect 14641 3848 14646 3904
rect 14702 3848 15946 3904
rect 14641 3846 15946 3848
rect 16021 3906 16087 3909
rect 18873 3906 18939 3909
rect 16021 3904 18939 3906
rect 16021 3848 16026 3904
rect 16082 3848 18878 3904
rect 18934 3848 18939 3904
rect 16021 3846 18939 3848
rect 14641 3843 14707 3846
rect 16021 3843 16087 3846
rect 18873 3843 18939 3846
rect 3545 3840 3861 3841
rect 3545 3776 3551 3840
rect 3615 3776 3631 3840
rect 3695 3776 3711 3840
rect 3775 3776 3791 3840
rect 3855 3776 3861 3840
rect 3545 3775 3861 3776
rect 8743 3840 9059 3841
rect 8743 3776 8749 3840
rect 8813 3776 8829 3840
rect 8893 3776 8909 3840
rect 8973 3776 8989 3840
rect 9053 3776 9059 3840
rect 8743 3775 9059 3776
rect 13941 3840 14257 3841
rect 13941 3776 13947 3840
rect 14011 3776 14027 3840
rect 14091 3776 14107 3840
rect 14171 3776 14187 3840
rect 14251 3776 14257 3840
rect 13941 3775 14257 3776
rect 19139 3840 19455 3841
rect 19139 3776 19145 3840
rect 19209 3776 19225 3840
rect 19289 3776 19305 3840
rect 19369 3776 19385 3840
rect 19449 3776 19455 3840
rect 19139 3775 19455 3776
rect 14365 3770 14431 3773
rect 18413 3770 18479 3773
rect 14365 3768 18479 3770
rect 14365 3712 14370 3768
rect 14426 3712 18418 3768
rect 18474 3712 18479 3768
rect 14365 3710 18479 3712
rect 19750 3770 19810 3982
rect 20069 3980 20116 3982
rect 20180 3980 20186 4044
rect 20069 3979 20135 3980
rect 20161 3906 20227 3909
rect 22840 3906 23300 3936
rect 20161 3904 23300 3906
rect 20161 3848 20166 3904
rect 20222 3848 23300 3904
rect 20161 3846 23300 3848
rect 20161 3843 20227 3846
rect 22840 3816 23300 3846
rect 19750 3710 22202 3770
rect 14365 3707 14431 3710
rect 18413 3707 18479 3710
rect 933 3634 999 3637
rect 4153 3634 4219 3637
rect 933 3632 4219 3634
rect 933 3576 938 3632
rect 994 3576 4158 3632
rect 4214 3576 4219 3632
rect 933 3574 4219 3576
rect 933 3571 999 3574
rect 4153 3571 4219 3574
rect 5257 3634 5323 3637
rect 7966 3634 7972 3636
rect 5257 3632 7972 3634
rect 5257 3576 5262 3632
rect 5318 3576 7972 3632
rect 5257 3574 7972 3576
rect 5257 3571 5323 3574
rect 7966 3572 7972 3574
rect 8036 3572 8042 3636
rect 14089 3634 14155 3637
rect 15469 3636 15535 3637
rect 15142 3634 15148 3636
rect 14089 3632 15148 3634
rect 14089 3576 14094 3632
rect 14150 3576 15148 3632
rect 14089 3574 15148 3576
rect 14089 3571 14155 3574
rect 15142 3572 15148 3574
rect 15212 3572 15218 3636
rect 15469 3632 15516 3636
rect 15580 3634 15586 3636
rect 15745 3634 15811 3637
rect 20713 3634 20779 3637
rect 15469 3576 15474 3632
rect 15469 3572 15516 3576
rect 15580 3574 15626 3634
rect 15745 3632 20779 3634
rect 15745 3576 15750 3632
rect 15806 3576 20718 3632
rect 20774 3576 20779 3632
rect 15745 3574 20779 3576
rect 15580 3572 15586 3574
rect 15469 3571 15535 3572
rect 15745 3571 15811 3574
rect 20713 3571 20779 3574
rect 10501 3498 10567 3501
rect 2730 3496 10567 3498
rect 2730 3440 10506 3496
rect 10562 3440 10567 3496
rect 2730 3438 10567 3440
rect 1485 3362 1551 3365
rect 2730 3362 2790 3438
rect 10501 3435 10567 3438
rect 16297 3498 16363 3501
rect 20805 3498 20871 3501
rect 16297 3496 20871 3498
rect 16297 3440 16302 3496
rect 16358 3440 20810 3496
rect 20866 3440 20871 3496
rect 16297 3438 20871 3440
rect 16297 3435 16363 3438
rect 20805 3435 20871 3438
rect 1485 3360 2790 3362
rect 1485 3304 1490 3360
rect 1546 3304 2790 3360
rect 1485 3302 2790 3304
rect 2865 3362 2931 3365
rect 5717 3362 5783 3365
rect 16297 3364 16363 3365
rect 16246 3362 16252 3364
rect 2865 3360 5783 3362
rect 2865 3304 2870 3360
rect 2926 3304 5722 3360
rect 5778 3304 5783 3360
rect 2865 3302 5783 3304
rect 16206 3302 16252 3362
rect 16316 3360 16363 3364
rect 16358 3304 16363 3360
rect 1485 3299 1551 3302
rect 2865 3299 2931 3302
rect 5717 3299 5783 3302
rect 16246 3300 16252 3302
rect 16316 3300 16363 3304
rect 16297 3299 16363 3300
rect 17401 3362 17467 3365
rect 18045 3364 18111 3365
rect 17718 3362 17724 3364
rect 17401 3360 17724 3362
rect 17401 3304 17406 3360
rect 17462 3304 17724 3360
rect 17401 3302 17724 3304
rect 17401 3299 17467 3302
rect 17718 3300 17724 3302
rect 17788 3300 17794 3364
rect 18045 3360 18092 3364
rect 18156 3362 18162 3364
rect 18321 3362 18387 3365
rect 18822 3362 18828 3364
rect 18045 3304 18050 3360
rect 18045 3300 18092 3304
rect 18156 3302 18202 3362
rect 18321 3360 18828 3362
rect 18321 3304 18326 3360
rect 18382 3304 18828 3360
rect 18321 3302 18828 3304
rect 18156 3300 18162 3302
rect 18045 3299 18111 3300
rect 18321 3299 18387 3302
rect 18822 3300 18828 3302
rect 18892 3300 18898 3364
rect 22142 3362 22202 3710
rect 22840 3362 23300 3392
rect 22142 3302 23300 3362
rect 6144 3296 6460 3297
rect 6144 3232 6150 3296
rect 6214 3232 6230 3296
rect 6294 3232 6310 3296
rect 6374 3232 6390 3296
rect 6454 3232 6460 3296
rect 6144 3231 6460 3232
rect 11342 3296 11658 3297
rect 11342 3232 11348 3296
rect 11412 3232 11428 3296
rect 11492 3232 11508 3296
rect 11572 3232 11588 3296
rect 11652 3232 11658 3296
rect 11342 3231 11658 3232
rect 16540 3296 16856 3297
rect 16540 3232 16546 3296
rect 16610 3232 16626 3296
rect 16690 3232 16706 3296
rect 16770 3232 16786 3296
rect 16850 3232 16856 3296
rect 16540 3231 16856 3232
rect 21738 3296 22054 3297
rect 21738 3232 21744 3296
rect 21808 3232 21824 3296
rect 21888 3232 21904 3296
rect 21968 3232 21984 3296
rect 22048 3232 22054 3296
rect 22840 3272 23300 3302
rect 21738 3231 22054 3232
rect 2037 3226 2103 3229
rect 5441 3226 5507 3229
rect 2037 3224 5507 3226
rect 2037 3168 2042 3224
rect 2098 3168 5446 3224
rect 5502 3168 5507 3224
rect 2037 3166 5507 3168
rect 2037 3163 2103 3166
rect 5441 3163 5507 3166
rect 8334 3164 8340 3228
rect 8404 3164 8410 3228
rect 8518 3164 8524 3228
rect 8588 3226 8594 3228
rect 8753 3226 8819 3229
rect 8588 3224 8819 3226
rect 8588 3168 8758 3224
rect 8814 3168 8819 3224
rect 8588 3166 8819 3168
rect 8588 3164 8594 3166
rect 5441 3090 5507 3093
rect 8342 3090 8402 3164
rect 8753 3163 8819 3166
rect 9213 3226 9279 3229
rect 9806 3226 9812 3228
rect 9213 3224 9812 3226
rect 9213 3168 9218 3224
rect 9274 3168 9812 3224
rect 9213 3166 9812 3168
rect 9213 3163 9279 3166
rect 9806 3164 9812 3166
rect 9876 3164 9882 3228
rect 15101 3226 15167 3229
rect 15837 3226 15903 3229
rect 15101 3224 15903 3226
rect 15101 3168 15106 3224
rect 15162 3168 15842 3224
rect 15898 3168 15903 3224
rect 15101 3166 15903 3168
rect 15101 3163 15167 3166
rect 15837 3163 15903 3166
rect 18597 3226 18663 3229
rect 19006 3226 19012 3228
rect 18597 3224 19012 3226
rect 18597 3168 18602 3224
rect 18658 3168 19012 3224
rect 18597 3166 19012 3168
rect 18597 3163 18663 3166
rect 19006 3164 19012 3166
rect 19076 3164 19082 3228
rect 8569 3090 8635 3093
rect 5441 3088 8402 3090
rect 5441 3032 5446 3088
rect 5502 3032 8402 3088
rect 5441 3030 8402 3032
rect 8526 3088 8635 3090
rect 8526 3032 8574 3088
rect 8630 3032 8635 3088
rect 5441 3027 5507 3030
rect 8526 3027 8635 3032
rect 9489 3090 9555 3093
rect 12014 3090 12020 3092
rect 9489 3088 12020 3090
rect 9489 3032 9494 3088
rect 9550 3032 12020 3088
rect 9489 3030 12020 3032
rect 9489 3027 9555 3030
rect 12014 3028 12020 3030
rect 12084 3028 12090 3092
rect 14365 3090 14431 3093
rect 20989 3090 21055 3093
rect 14365 3088 21055 3090
rect 14365 3032 14370 3088
rect 14426 3032 20994 3088
rect 21050 3032 21055 3088
rect 14365 3030 21055 3032
rect 14365 3027 14431 3030
rect 20989 3027 21055 3030
rect 4061 2954 4127 2957
rect 8201 2954 8267 2957
rect 4061 2952 8267 2954
rect 4061 2896 4066 2952
rect 4122 2896 8206 2952
rect 8262 2896 8267 2952
rect 4061 2894 8267 2896
rect 4061 2891 4127 2894
rect 8201 2891 8267 2894
rect 5942 2756 5948 2820
rect 6012 2818 6018 2820
rect 8526 2818 8586 3027
rect 13813 2954 13879 2957
rect 14733 2954 14799 2957
rect 17953 2954 18019 2957
rect 13813 2952 14474 2954
rect 13813 2896 13818 2952
rect 13874 2896 14474 2952
rect 13813 2894 14474 2896
rect 13813 2891 13879 2894
rect 6012 2758 6930 2818
rect 6012 2756 6018 2758
rect 3545 2752 3861 2753
rect 3545 2688 3551 2752
rect 3615 2688 3631 2752
rect 3695 2688 3711 2752
rect 3775 2688 3791 2752
rect 3855 2688 3861 2752
rect 3545 2687 3861 2688
rect 6870 2682 6930 2758
rect 8342 2758 8586 2818
rect 7189 2682 7255 2685
rect 6870 2680 7255 2682
rect 6870 2624 7194 2680
rect 7250 2624 7255 2680
rect 6870 2622 7255 2624
rect 7189 2619 7255 2622
rect 7925 2682 7991 2685
rect 8150 2682 8156 2684
rect 7925 2680 8156 2682
rect 7925 2624 7930 2680
rect 7986 2624 8156 2680
rect 7925 2622 8156 2624
rect 7925 2619 7991 2622
rect 8150 2620 8156 2622
rect 8220 2620 8226 2684
rect 2865 2548 2931 2549
rect 2814 2484 2820 2548
rect 2884 2546 2931 2548
rect 4153 2546 4219 2549
rect 5625 2546 5691 2549
rect 2884 2544 2976 2546
rect 2926 2488 2976 2544
rect 2884 2486 2976 2488
rect 4153 2544 5691 2546
rect 4153 2488 4158 2544
rect 4214 2488 5630 2544
rect 5686 2488 5691 2544
rect 4153 2486 5691 2488
rect 2884 2484 2931 2486
rect 2865 2483 2931 2484
rect 4153 2483 4219 2486
rect 5625 2483 5691 2486
rect 6545 2546 6611 2549
rect 7598 2546 7604 2548
rect 6545 2544 7604 2546
rect 6545 2488 6550 2544
rect 6606 2488 7604 2544
rect 6545 2486 7604 2488
rect 6545 2483 6611 2486
rect 7598 2484 7604 2486
rect 7668 2484 7674 2548
rect 6269 2410 6335 2413
rect 6862 2410 6868 2412
rect 6269 2408 6868 2410
rect 6269 2352 6274 2408
rect 6330 2352 6868 2408
rect 6269 2350 6868 2352
rect 6269 2347 6335 2350
rect 6862 2348 6868 2350
rect 6932 2348 6938 2412
rect 790 2212 796 2276
rect 860 2212 866 2276
rect 4797 2274 4863 2277
rect 5441 2276 5507 2277
rect 5206 2274 5212 2276
rect 4797 2272 5212 2274
rect 4797 2216 4802 2272
rect 4858 2216 5212 2272
rect 4797 2214 5212 2216
rect 798 2138 858 2212
rect 4797 2211 4863 2214
rect 5206 2212 5212 2214
rect 5276 2212 5282 2276
rect 5390 2212 5396 2276
rect 5460 2274 5507 2276
rect 8201 2274 8267 2277
rect 8342 2274 8402 2758
rect 9254 2756 9260 2820
rect 9324 2756 9330 2820
rect 8743 2752 9059 2753
rect 8743 2688 8749 2752
rect 8813 2688 8829 2752
rect 8893 2688 8909 2752
rect 8973 2688 8989 2752
rect 9053 2688 9059 2752
rect 8743 2687 9059 2688
rect 8753 2546 8819 2549
rect 9262 2546 9322 2756
rect 13941 2752 14257 2753
rect 13941 2688 13947 2752
rect 14011 2688 14027 2752
rect 14091 2688 14107 2752
rect 14171 2688 14187 2752
rect 14251 2688 14257 2752
rect 13941 2687 14257 2688
rect 8753 2544 9322 2546
rect 8753 2488 8758 2544
rect 8814 2488 9322 2544
rect 8753 2486 9322 2488
rect 14414 2546 14474 2894
rect 14733 2952 18019 2954
rect 14733 2896 14738 2952
rect 14794 2896 17958 2952
rect 18014 2896 18019 2952
rect 14733 2894 18019 2896
rect 14733 2891 14799 2894
rect 17953 2891 18019 2894
rect 16113 2818 16179 2821
rect 18597 2818 18663 2821
rect 16113 2816 18663 2818
rect 16113 2760 16118 2816
rect 16174 2760 18602 2816
rect 18658 2760 18663 2816
rect 16113 2758 18663 2760
rect 16113 2755 16179 2758
rect 18597 2755 18663 2758
rect 21081 2818 21147 2821
rect 22840 2818 23300 2848
rect 21081 2816 23300 2818
rect 21081 2760 21086 2816
rect 21142 2760 23300 2816
rect 21081 2758 23300 2760
rect 21081 2755 21147 2758
rect 19139 2752 19455 2753
rect 19139 2688 19145 2752
rect 19209 2688 19225 2752
rect 19289 2688 19305 2752
rect 19369 2688 19385 2752
rect 19449 2688 19455 2752
rect 22840 2728 23300 2758
rect 19139 2687 19455 2688
rect 14549 2682 14615 2685
rect 16113 2682 16179 2685
rect 14549 2680 16179 2682
rect 14549 2624 14554 2680
rect 14610 2624 16118 2680
rect 16174 2624 16179 2680
rect 14549 2622 16179 2624
rect 14549 2619 14615 2622
rect 16113 2619 16179 2622
rect 16573 2682 16639 2685
rect 17350 2682 17356 2684
rect 16573 2680 17356 2682
rect 16573 2624 16578 2680
rect 16634 2624 17356 2680
rect 16573 2622 17356 2624
rect 16573 2619 16639 2622
rect 17350 2620 17356 2622
rect 17420 2620 17426 2684
rect 17902 2620 17908 2684
rect 17972 2682 17978 2684
rect 18505 2682 18571 2685
rect 17972 2680 18571 2682
rect 17972 2624 18510 2680
rect 18566 2624 18571 2680
rect 17972 2622 18571 2624
rect 17972 2620 17978 2622
rect 18505 2619 18571 2622
rect 14414 2486 17234 2546
rect 8753 2483 8819 2486
rect 14365 2410 14431 2413
rect 17174 2410 17234 2486
rect 17350 2484 17356 2548
rect 17420 2546 17426 2548
rect 17585 2546 17651 2549
rect 17420 2544 17651 2546
rect 17420 2488 17590 2544
rect 17646 2488 17651 2544
rect 17420 2486 17651 2488
rect 17420 2484 17426 2486
rect 17585 2483 17651 2486
rect 18689 2546 18755 2549
rect 18689 2544 22386 2546
rect 18689 2488 18694 2544
rect 18750 2488 22386 2544
rect 18689 2486 22386 2488
rect 18689 2483 18755 2486
rect 18689 2410 18755 2413
rect 14365 2408 17050 2410
rect 14365 2352 14370 2408
rect 14426 2352 17050 2408
rect 14365 2350 17050 2352
rect 17174 2408 18755 2410
rect 17174 2352 18694 2408
rect 18750 2352 18755 2408
rect 17174 2350 18755 2352
rect 14365 2347 14431 2350
rect 5460 2272 5552 2274
rect 5502 2216 5552 2272
rect 5460 2214 5552 2216
rect 8201 2272 8402 2274
rect 8201 2216 8206 2272
rect 8262 2216 8402 2272
rect 8201 2214 8402 2216
rect 16990 2274 17050 2350
rect 18689 2347 18755 2350
rect 20713 2274 20779 2277
rect 20989 2276 21055 2277
rect 21357 2276 21423 2277
rect 20989 2274 21036 2276
rect 16990 2272 20779 2274
rect 16990 2216 20718 2272
rect 20774 2216 20779 2272
rect 16990 2214 20779 2216
rect 20944 2272 21036 2274
rect 20944 2216 20994 2272
rect 20944 2214 21036 2216
rect 5460 2212 5507 2214
rect 5441 2211 5507 2212
rect 8201 2211 8267 2214
rect 20713 2211 20779 2214
rect 20989 2212 21036 2214
rect 21100 2212 21106 2276
rect 21357 2274 21404 2276
rect 21312 2272 21404 2274
rect 21312 2216 21362 2272
rect 21312 2214 21404 2216
rect 21357 2212 21404 2214
rect 21468 2212 21474 2276
rect 22326 2274 22386 2486
rect 22840 2274 23300 2304
rect 22326 2214 23300 2274
rect 20989 2211 21055 2212
rect 21357 2211 21423 2212
rect 6144 2208 6460 2209
rect 6144 2144 6150 2208
rect 6214 2144 6230 2208
rect 6294 2144 6310 2208
rect 6374 2144 6390 2208
rect 6454 2144 6460 2208
rect 6144 2143 6460 2144
rect 11342 2208 11658 2209
rect 11342 2144 11348 2208
rect 11412 2144 11428 2208
rect 11492 2144 11508 2208
rect 11572 2144 11588 2208
rect 11652 2144 11658 2208
rect 11342 2143 11658 2144
rect 16540 2208 16856 2209
rect 16540 2144 16546 2208
rect 16610 2144 16626 2208
rect 16690 2144 16706 2208
rect 16770 2144 16786 2208
rect 16850 2144 16856 2208
rect 16540 2143 16856 2144
rect 21738 2208 22054 2209
rect 21738 2144 21744 2208
rect 21808 2144 21824 2208
rect 21888 2144 21904 2208
rect 21968 2144 21984 2208
rect 22048 2144 22054 2208
rect 22840 2184 23300 2214
rect 21738 2143 22054 2144
rect 5717 2138 5783 2141
rect 21541 2138 21607 2141
rect 798 2136 5783 2138
rect 798 2080 5722 2136
rect 5778 2080 5783 2136
rect 798 2078 5783 2080
rect 5717 2075 5783 2078
rect 16990 2136 21607 2138
rect 16990 2080 21546 2136
rect 21602 2080 21607 2136
rect 16990 2078 21607 2080
rect 974 1940 980 2004
rect 1044 2002 1050 2004
rect 9765 2002 9831 2005
rect 1044 2000 9831 2002
rect 1044 1944 9770 2000
rect 9826 1944 9831 2000
rect 1044 1942 9831 1944
rect 1044 1940 1050 1942
rect 9765 1939 9831 1942
rect 10133 2002 10199 2005
rect 11973 2002 12039 2005
rect 10133 2000 12039 2002
rect 10133 1944 10138 2000
rect 10194 1944 11978 2000
rect 12034 1944 12039 2000
rect 10133 1942 12039 1944
rect 10133 1939 10199 1942
rect 11973 1939 12039 1942
rect 12709 2002 12775 2005
rect 13445 2002 13511 2005
rect 16990 2002 17050 2078
rect 21541 2075 21607 2078
rect 12709 2000 13370 2002
rect 12709 1944 12714 2000
rect 12770 1944 13370 2000
rect 12709 1942 13370 1944
rect 12709 1939 12775 1942
rect 606 1804 612 1868
rect 676 1866 682 1868
rect 7005 1866 7071 1869
rect 676 1864 7071 1866
rect 676 1808 7010 1864
rect 7066 1808 7071 1864
rect 676 1806 7071 1808
rect 676 1804 682 1806
rect 7005 1803 7071 1806
rect 7414 1804 7420 1868
rect 7484 1866 7490 1868
rect 7649 1866 7715 1869
rect 7484 1864 7715 1866
rect 7484 1808 7654 1864
rect 7710 1808 7715 1864
rect 7484 1806 7715 1808
rect 13310 1866 13370 1942
rect 13445 2000 17050 2002
rect 13445 1944 13450 2000
rect 13506 1944 17050 2000
rect 13445 1942 17050 1944
rect 18965 2002 19031 2005
rect 18965 2000 20960 2002
rect 18965 1944 18970 2000
rect 19026 1944 20960 2000
rect 18965 1942 20960 1944
rect 13445 1939 13511 1942
rect 18965 1939 19031 1942
rect 18638 1866 18644 1868
rect 13310 1806 18644 1866
rect 7484 1804 7490 1806
rect 7649 1803 7715 1806
rect 18638 1804 18644 1806
rect 18708 1804 18714 1868
rect 14549 1730 14615 1733
rect 17033 1732 17099 1733
rect 14549 1728 16866 1730
rect 14549 1672 14554 1728
rect 14610 1672 16866 1728
rect 14549 1670 16866 1672
rect 14549 1667 14615 1670
rect 3545 1664 3861 1665
rect 3545 1600 3551 1664
rect 3615 1600 3631 1664
rect 3695 1600 3711 1664
rect 3775 1600 3791 1664
rect 3855 1600 3861 1664
rect 3545 1599 3861 1600
rect 8743 1664 9059 1665
rect 8743 1600 8749 1664
rect 8813 1600 8829 1664
rect 8893 1600 8909 1664
rect 8973 1600 8989 1664
rect 9053 1600 9059 1664
rect 8743 1599 9059 1600
rect 13941 1664 14257 1665
rect 13941 1600 13947 1664
rect 14011 1600 14027 1664
rect 14091 1600 14107 1664
rect 14171 1600 14187 1664
rect 14251 1600 14257 1664
rect 13941 1599 14257 1600
rect 14917 1594 14983 1597
rect 15745 1594 15811 1597
rect 14917 1592 15811 1594
rect 14917 1536 14922 1592
rect 14978 1536 15750 1592
rect 15806 1536 15811 1592
rect 14917 1534 15811 1536
rect 16806 1594 16866 1670
rect 16982 1668 16988 1732
rect 17052 1730 17099 1732
rect 20900 1730 20960 1942
rect 22840 1730 23300 1760
rect 17052 1728 17144 1730
rect 17094 1672 17144 1728
rect 17052 1670 17144 1672
rect 20900 1670 23300 1730
rect 17052 1668 17099 1670
rect 17033 1667 17099 1668
rect 19139 1664 19455 1665
rect 19139 1600 19145 1664
rect 19209 1600 19225 1664
rect 19289 1600 19305 1664
rect 19369 1600 19385 1664
rect 19449 1600 19455 1664
rect 22840 1640 23300 1670
rect 19139 1599 19455 1600
rect 18137 1594 18203 1597
rect 16806 1592 18203 1594
rect 16806 1536 18142 1592
rect 18198 1536 18203 1592
rect 16806 1534 18203 1536
rect 14917 1531 14983 1534
rect 15745 1531 15811 1534
rect 18137 1531 18203 1534
rect 749 1458 815 1461
rect 7189 1458 7255 1461
rect 749 1456 7255 1458
rect 749 1400 754 1456
rect 810 1400 7194 1456
rect 7250 1400 7255 1456
rect 749 1398 7255 1400
rect 749 1395 815 1398
rect 7189 1395 7255 1398
rect 8201 1458 8267 1461
rect 9397 1458 9463 1461
rect 8201 1456 9463 1458
rect 8201 1400 8206 1456
rect 8262 1400 9402 1456
rect 9458 1400 9463 1456
rect 8201 1398 9463 1400
rect 8201 1395 8267 1398
rect 9397 1395 9463 1398
rect 14365 1458 14431 1461
rect 16849 1458 16915 1461
rect 14365 1456 16915 1458
rect 14365 1400 14370 1456
rect 14426 1400 16854 1456
rect 16910 1400 16915 1456
rect 14365 1398 16915 1400
rect 14365 1395 14431 1398
rect 16849 1395 16915 1398
rect 1158 1260 1164 1324
rect 1228 1322 1234 1324
rect 3509 1322 3575 1325
rect 1228 1320 3575 1322
rect 1228 1264 3514 1320
rect 3570 1264 3575 1320
rect 1228 1262 3575 1264
rect 1228 1260 1234 1262
rect 3509 1259 3575 1262
rect 4102 1260 4108 1324
rect 4172 1260 4178 1324
rect 7230 1260 7236 1324
rect 7300 1322 7306 1324
rect 7373 1322 7439 1325
rect 9857 1324 9923 1325
rect 7300 1320 7439 1322
rect 7300 1264 7378 1320
rect 7434 1264 7439 1320
rect 7300 1262 7439 1264
rect 7300 1260 7306 1262
rect 3325 1186 3391 1189
rect 4110 1186 4170 1260
rect 7373 1259 7439 1262
rect 9806 1260 9812 1324
rect 9876 1322 9923 1324
rect 9876 1320 9968 1322
rect 9918 1264 9968 1320
rect 9876 1262 9968 1264
rect 19014 1262 22202 1322
rect 9876 1260 9923 1262
rect 9857 1259 9923 1260
rect 19014 1188 19074 1262
rect 3325 1184 4170 1186
rect 3325 1128 3330 1184
rect 3386 1128 4170 1184
rect 3325 1126 4170 1128
rect 3325 1123 3391 1126
rect 19006 1124 19012 1188
rect 19076 1124 19082 1188
rect 22142 1186 22202 1262
rect 22840 1186 23300 1216
rect 22142 1126 23300 1186
rect 6144 1120 6460 1121
rect 6144 1056 6150 1120
rect 6214 1056 6230 1120
rect 6294 1056 6310 1120
rect 6374 1056 6390 1120
rect 6454 1056 6460 1120
rect 6144 1055 6460 1056
rect 11342 1120 11658 1121
rect 11342 1056 11348 1120
rect 11412 1056 11428 1120
rect 11492 1056 11508 1120
rect 11572 1056 11588 1120
rect 11652 1056 11658 1120
rect 11342 1055 11658 1056
rect 16540 1120 16856 1121
rect 16540 1056 16546 1120
rect 16610 1056 16626 1120
rect 16690 1056 16706 1120
rect 16770 1056 16786 1120
rect 16850 1056 16856 1120
rect 16540 1055 16856 1056
rect 21738 1120 22054 1121
rect 21738 1056 21744 1120
rect 21808 1056 21824 1120
rect 21888 1056 21904 1120
rect 21968 1056 21984 1120
rect 22048 1056 22054 1120
rect 22840 1096 23300 1126
rect 21738 1055 22054 1056
rect 9622 914 9628 916
rect 2730 854 9628 914
rect 1485 778 1551 781
rect 2730 778 2790 854
rect 9622 852 9628 854
rect 9692 852 9698 916
rect 15377 914 15443 917
rect 19926 914 19932 916
rect 15377 912 19932 914
rect 15377 856 15382 912
rect 15438 856 19932 912
rect 15377 854 19932 856
rect 15377 851 15443 854
rect 19926 852 19932 854
rect 19996 852 20002 916
rect 20662 852 20668 916
rect 20732 852 20738 916
rect 1485 776 2790 778
rect 1485 720 1490 776
rect 1546 720 2790 776
rect 1485 718 2790 720
rect 4797 778 4863 781
rect 20670 778 20730 852
rect 4797 776 20730 778
rect 4797 720 4802 776
rect 4858 720 20730 776
rect 4797 718 20730 720
rect 1485 715 1551 718
rect 4797 715 4863 718
rect 18822 580 18828 644
rect 18892 642 18898 644
rect 22840 642 23300 672
rect 18892 582 23300 642
rect 18892 580 18898 582
rect 22840 552 23300 582
rect 8518 36 8524 100
rect 8588 98 8594 100
rect 8937 98 9003 101
rect 8588 96 9003 98
rect 8588 40 8942 96
rect 8998 40 9003 96
rect 8588 38 9003 40
rect 8588 36 8594 38
rect 8937 35 9003 38
<< via3 >>
rect 6150 43548 6214 43552
rect 6150 43492 6154 43548
rect 6154 43492 6210 43548
rect 6210 43492 6214 43548
rect 6150 43488 6214 43492
rect 6230 43548 6294 43552
rect 6230 43492 6234 43548
rect 6234 43492 6290 43548
rect 6290 43492 6294 43548
rect 6230 43488 6294 43492
rect 6310 43548 6374 43552
rect 6310 43492 6314 43548
rect 6314 43492 6370 43548
rect 6370 43492 6374 43548
rect 6310 43488 6374 43492
rect 6390 43548 6454 43552
rect 6390 43492 6394 43548
rect 6394 43492 6450 43548
rect 6450 43492 6454 43548
rect 6390 43488 6454 43492
rect 11348 43548 11412 43552
rect 11348 43492 11352 43548
rect 11352 43492 11408 43548
rect 11408 43492 11412 43548
rect 11348 43488 11412 43492
rect 11428 43548 11492 43552
rect 11428 43492 11432 43548
rect 11432 43492 11488 43548
rect 11488 43492 11492 43548
rect 11428 43488 11492 43492
rect 11508 43548 11572 43552
rect 11508 43492 11512 43548
rect 11512 43492 11568 43548
rect 11568 43492 11572 43548
rect 11508 43488 11572 43492
rect 11588 43548 11652 43552
rect 11588 43492 11592 43548
rect 11592 43492 11648 43548
rect 11648 43492 11652 43548
rect 11588 43488 11652 43492
rect 16546 43548 16610 43552
rect 16546 43492 16550 43548
rect 16550 43492 16606 43548
rect 16606 43492 16610 43548
rect 16546 43488 16610 43492
rect 16626 43548 16690 43552
rect 16626 43492 16630 43548
rect 16630 43492 16686 43548
rect 16686 43492 16690 43548
rect 16626 43488 16690 43492
rect 16706 43548 16770 43552
rect 16706 43492 16710 43548
rect 16710 43492 16766 43548
rect 16766 43492 16770 43548
rect 16706 43488 16770 43492
rect 16786 43548 16850 43552
rect 16786 43492 16790 43548
rect 16790 43492 16846 43548
rect 16846 43492 16850 43548
rect 16786 43488 16850 43492
rect 21744 43548 21808 43552
rect 21744 43492 21748 43548
rect 21748 43492 21804 43548
rect 21804 43492 21808 43548
rect 21744 43488 21808 43492
rect 21824 43548 21888 43552
rect 21824 43492 21828 43548
rect 21828 43492 21884 43548
rect 21884 43492 21888 43548
rect 21824 43488 21888 43492
rect 21904 43548 21968 43552
rect 21904 43492 21908 43548
rect 21908 43492 21964 43548
rect 21964 43492 21968 43548
rect 21904 43488 21968 43492
rect 21984 43548 22048 43552
rect 21984 43492 21988 43548
rect 21988 43492 22044 43548
rect 22044 43492 22048 43548
rect 21984 43488 22048 43492
rect 11836 43148 11900 43212
rect 3551 43004 3615 43008
rect 3551 42948 3555 43004
rect 3555 42948 3611 43004
rect 3611 42948 3615 43004
rect 3551 42944 3615 42948
rect 3631 43004 3695 43008
rect 3631 42948 3635 43004
rect 3635 42948 3691 43004
rect 3691 42948 3695 43004
rect 3631 42944 3695 42948
rect 3711 43004 3775 43008
rect 3711 42948 3715 43004
rect 3715 42948 3771 43004
rect 3771 42948 3775 43004
rect 3711 42944 3775 42948
rect 3791 43004 3855 43008
rect 3791 42948 3795 43004
rect 3795 42948 3851 43004
rect 3851 42948 3855 43004
rect 3791 42944 3855 42948
rect 8749 43004 8813 43008
rect 8749 42948 8753 43004
rect 8753 42948 8809 43004
rect 8809 42948 8813 43004
rect 8749 42944 8813 42948
rect 8829 43004 8893 43008
rect 8829 42948 8833 43004
rect 8833 42948 8889 43004
rect 8889 42948 8893 43004
rect 8829 42944 8893 42948
rect 8909 43004 8973 43008
rect 8909 42948 8913 43004
rect 8913 42948 8969 43004
rect 8969 42948 8973 43004
rect 8909 42944 8973 42948
rect 8989 43004 9053 43008
rect 8989 42948 8993 43004
rect 8993 42948 9049 43004
rect 9049 42948 9053 43004
rect 8989 42944 9053 42948
rect 5028 42876 5092 42940
rect 13947 43004 14011 43008
rect 13947 42948 13951 43004
rect 13951 42948 14007 43004
rect 14007 42948 14011 43004
rect 13947 42944 14011 42948
rect 14027 43004 14091 43008
rect 14027 42948 14031 43004
rect 14031 42948 14087 43004
rect 14087 42948 14091 43004
rect 14027 42944 14091 42948
rect 14107 43004 14171 43008
rect 14107 42948 14111 43004
rect 14111 42948 14167 43004
rect 14167 42948 14171 43004
rect 14107 42944 14171 42948
rect 14187 43004 14251 43008
rect 14187 42948 14191 43004
rect 14191 42948 14247 43004
rect 14247 42948 14251 43004
rect 14187 42944 14251 42948
rect 19145 43004 19209 43008
rect 19145 42948 19149 43004
rect 19149 42948 19205 43004
rect 19205 42948 19209 43004
rect 19145 42944 19209 42948
rect 19225 43004 19289 43008
rect 19225 42948 19229 43004
rect 19229 42948 19285 43004
rect 19285 42948 19289 43004
rect 19225 42944 19289 42948
rect 19305 43004 19369 43008
rect 19305 42948 19309 43004
rect 19309 42948 19365 43004
rect 19365 42948 19369 43004
rect 19305 42944 19369 42948
rect 19385 43004 19449 43008
rect 19385 42948 19389 43004
rect 19389 42948 19445 43004
rect 19445 42948 19449 43004
rect 19385 42944 19449 42948
rect 13124 42936 13188 42940
rect 13124 42880 13138 42936
rect 13138 42880 13188 42936
rect 13124 42876 13188 42880
rect 6684 42468 6748 42532
rect 6150 42460 6214 42464
rect 6150 42404 6154 42460
rect 6154 42404 6210 42460
rect 6210 42404 6214 42460
rect 6150 42400 6214 42404
rect 6230 42460 6294 42464
rect 6230 42404 6234 42460
rect 6234 42404 6290 42460
rect 6290 42404 6294 42460
rect 6230 42400 6294 42404
rect 6310 42460 6374 42464
rect 6310 42404 6314 42460
rect 6314 42404 6370 42460
rect 6370 42404 6374 42460
rect 6310 42400 6374 42404
rect 6390 42460 6454 42464
rect 6390 42404 6394 42460
rect 6394 42404 6450 42460
rect 6450 42404 6454 42460
rect 6390 42400 6454 42404
rect 11348 42460 11412 42464
rect 11348 42404 11352 42460
rect 11352 42404 11408 42460
rect 11408 42404 11412 42460
rect 11348 42400 11412 42404
rect 11428 42460 11492 42464
rect 11428 42404 11432 42460
rect 11432 42404 11488 42460
rect 11488 42404 11492 42460
rect 11428 42400 11492 42404
rect 11508 42460 11572 42464
rect 11508 42404 11512 42460
rect 11512 42404 11568 42460
rect 11568 42404 11572 42460
rect 11508 42400 11572 42404
rect 11588 42460 11652 42464
rect 11588 42404 11592 42460
rect 11592 42404 11648 42460
rect 11648 42404 11652 42460
rect 11588 42400 11652 42404
rect 9260 42332 9324 42396
rect 9444 42332 9508 42396
rect 17908 42876 17972 42940
rect 16546 42460 16610 42464
rect 16546 42404 16550 42460
rect 16550 42404 16606 42460
rect 16606 42404 16610 42460
rect 16546 42400 16610 42404
rect 16626 42460 16690 42464
rect 16626 42404 16630 42460
rect 16630 42404 16686 42460
rect 16686 42404 16690 42460
rect 16626 42400 16690 42404
rect 16706 42460 16770 42464
rect 16706 42404 16710 42460
rect 16710 42404 16766 42460
rect 16766 42404 16770 42460
rect 16706 42400 16770 42404
rect 16786 42460 16850 42464
rect 16786 42404 16790 42460
rect 16790 42404 16846 42460
rect 16846 42404 16850 42460
rect 16786 42400 16850 42404
rect 21744 42460 21808 42464
rect 21744 42404 21748 42460
rect 21748 42404 21804 42460
rect 21804 42404 21808 42460
rect 21744 42400 21808 42404
rect 21824 42460 21888 42464
rect 21824 42404 21828 42460
rect 21828 42404 21884 42460
rect 21884 42404 21888 42460
rect 21824 42400 21888 42404
rect 21904 42460 21968 42464
rect 21904 42404 21908 42460
rect 21908 42404 21964 42460
rect 21964 42404 21968 42460
rect 21904 42400 21968 42404
rect 21984 42460 22048 42464
rect 21984 42404 21988 42460
rect 21988 42404 22044 42460
rect 22044 42404 22048 42460
rect 21984 42400 22048 42404
rect 19748 42332 19812 42396
rect 8340 42196 8404 42260
rect 10180 41924 10244 41988
rect 3551 41916 3615 41920
rect 3551 41860 3555 41916
rect 3555 41860 3611 41916
rect 3611 41860 3615 41916
rect 3551 41856 3615 41860
rect 3631 41916 3695 41920
rect 3631 41860 3635 41916
rect 3635 41860 3691 41916
rect 3691 41860 3695 41916
rect 3631 41856 3695 41860
rect 3711 41916 3775 41920
rect 3711 41860 3715 41916
rect 3715 41860 3771 41916
rect 3771 41860 3775 41916
rect 3711 41856 3775 41860
rect 3791 41916 3855 41920
rect 3791 41860 3795 41916
rect 3795 41860 3851 41916
rect 3851 41860 3855 41916
rect 3791 41856 3855 41860
rect 8749 41916 8813 41920
rect 8749 41860 8753 41916
rect 8753 41860 8809 41916
rect 8809 41860 8813 41916
rect 8749 41856 8813 41860
rect 8829 41916 8893 41920
rect 8829 41860 8833 41916
rect 8833 41860 8889 41916
rect 8889 41860 8893 41916
rect 8829 41856 8893 41860
rect 8909 41916 8973 41920
rect 8909 41860 8913 41916
rect 8913 41860 8969 41916
rect 8969 41860 8973 41916
rect 8909 41856 8973 41860
rect 8989 41916 9053 41920
rect 8989 41860 8993 41916
rect 8993 41860 9049 41916
rect 9049 41860 9053 41916
rect 8989 41856 9053 41860
rect 13947 41916 14011 41920
rect 13947 41860 13951 41916
rect 13951 41860 14007 41916
rect 14007 41860 14011 41916
rect 13947 41856 14011 41860
rect 14027 41916 14091 41920
rect 14027 41860 14031 41916
rect 14031 41860 14087 41916
rect 14087 41860 14091 41916
rect 14027 41856 14091 41860
rect 14107 41916 14171 41920
rect 14107 41860 14111 41916
rect 14111 41860 14167 41916
rect 14167 41860 14171 41916
rect 14107 41856 14171 41860
rect 14187 41916 14251 41920
rect 14187 41860 14191 41916
rect 14191 41860 14247 41916
rect 14247 41860 14251 41916
rect 14187 41856 14251 41860
rect 796 41652 860 41716
rect 20484 42196 20548 42260
rect 17724 42060 17788 42124
rect 19145 41916 19209 41920
rect 19145 41860 19149 41916
rect 19149 41860 19205 41916
rect 19205 41860 19209 41916
rect 19145 41856 19209 41860
rect 19225 41916 19289 41920
rect 19225 41860 19229 41916
rect 19229 41860 19285 41916
rect 19285 41860 19289 41916
rect 19225 41856 19289 41860
rect 19305 41916 19369 41920
rect 19305 41860 19309 41916
rect 19309 41860 19365 41916
rect 19365 41860 19369 41916
rect 19305 41856 19369 41860
rect 19385 41916 19449 41920
rect 19385 41860 19389 41916
rect 19389 41860 19445 41916
rect 19445 41860 19449 41916
rect 19385 41856 19449 41860
rect 18092 41788 18156 41852
rect 15148 41712 15212 41716
rect 15148 41656 15198 41712
rect 15198 41656 15212 41712
rect 15148 41652 15212 41656
rect 16068 41652 16132 41716
rect 4660 41516 4724 41580
rect 7420 41576 7484 41580
rect 7420 41520 7434 41576
rect 7434 41520 7484 41576
rect 7420 41516 7484 41520
rect 15332 41380 15396 41444
rect 17356 41516 17420 41580
rect 6150 41372 6214 41376
rect 6150 41316 6154 41372
rect 6154 41316 6210 41372
rect 6210 41316 6214 41372
rect 6150 41312 6214 41316
rect 6230 41372 6294 41376
rect 6230 41316 6234 41372
rect 6234 41316 6290 41372
rect 6290 41316 6294 41372
rect 6230 41312 6294 41316
rect 6310 41372 6374 41376
rect 6310 41316 6314 41372
rect 6314 41316 6370 41372
rect 6370 41316 6374 41372
rect 6310 41312 6374 41316
rect 6390 41372 6454 41376
rect 6390 41316 6394 41372
rect 6394 41316 6450 41372
rect 6450 41316 6454 41372
rect 6390 41312 6454 41316
rect 11348 41372 11412 41376
rect 11348 41316 11352 41372
rect 11352 41316 11408 41372
rect 11408 41316 11412 41372
rect 11348 41312 11412 41316
rect 11428 41372 11492 41376
rect 11428 41316 11432 41372
rect 11432 41316 11488 41372
rect 11488 41316 11492 41372
rect 11428 41312 11492 41316
rect 11508 41372 11572 41376
rect 11508 41316 11512 41372
rect 11512 41316 11568 41372
rect 11568 41316 11572 41372
rect 11508 41312 11572 41316
rect 11588 41372 11652 41376
rect 11588 41316 11592 41372
rect 11592 41316 11648 41372
rect 11648 41316 11652 41372
rect 11588 41312 11652 41316
rect 16546 41372 16610 41376
rect 16546 41316 16550 41372
rect 16550 41316 16606 41372
rect 16606 41316 16610 41372
rect 16546 41312 16610 41316
rect 16626 41372 16690 41376
rect 16626 41316 16630 41372
rect 16630 41316 16686 41372
rect 16686 41316 16690 41372
rect 16626 41312 16690 41316
rect 16706 41372 16770 41376
rect 16706 41316 16710 41372
rect 16710 41316 16766 41372
rect 16766 41316 16770 41372
rect 16706 41312 16770 41316
rect 16786 41372 16850 41376
rect 16786 41316 16790 41372
rect 16790 41316 16846 41372
rect 16846 41316 16850 41372
rect 16786 41312 16850 41316
rect 18276 41304 18340 41308
rect 18276 41248 18326 41304
rect 18326 41248 18340 41304
rect 18276 41244 18340 41248
rect 21744 41372 21808 41376
rect 21744 41316 21748 41372
rect 21748 41316 21804 41372
rect 21804 41316 21808 41372
rect 21744 41312 21808 41316
rect 21824 41372 21888 41376
rect 21824 41316 21828 41372
rect 21828 41316 21884 41372
rect 21884 41316 21888 41372
rect 21824 41312 21888 41316
rect 21904 41372 21968 41376
rect 21904 41316 21908 41372
rect 21908 41316 21964 41372
rect 21964 41316 21968 41372
rect 21904 41312 21968 41316
rect 21984 41372 22048 41376
rect 21984 41316 21988 41372
rect 21988 41316 22044 41372
rect 22044 41316 22048 41372
rect 21984 41312 22048 41316
rect 17724 40836 17788 40900
rect 3551 40828 3615 40832
rect 3551 40772 3555 40828
rect 3555 40772 3611 40828
rect 3611 40772 3615 40828
rect 3551 40768 3615 40772
rect 3631 40828 3695 40832
rect 3631 40772 3635 40828
rect 3635 40772 3691 40828
rect 3691 40772 3695 40828
rect 3631 40768 3695 40772
rect 3711 40828 3775 40832
rect 3711 40772 3715 40828
rect 3715 40772 3771 40828
rect 3771 40772 3775 40828
rect 3711 40768 3775 40772
rect 3791 40828 3855 40832
rect 3791 40772 3795 40828
rect 3795 40772 3851 40828
rect 3851 40772 3855 40828
rect 3791 40768 3855 40772
rect 8749 40828 8813 40832
rect 8749 40772 8753 40828
rect 8753 40772 8809 40828
rect 8809 40772 8813 40828
rect 8749 40768 8813 40772
rect 8829 40828 8893 40832
rect 8829 40772 8833 40828
rect 8833 40772 8889 40828
rect 8889 40772 8893 40828
rect 8829 40768 8893 40772
rect 8909 40828 8973 40832
rect 8909 40772 8913 40828
rect 8913 40772 8969 40828
rect 8969 40772 8973 40828
rect 8909 40768 8973 40772
rect 8989 40828 9053 40832
rect 8989 40772 8993 40828
rect 8993 40772 9049 40828
rect 9049 40772 9053 40828
rect 8989 40768 9053 40772
rect 13947 40828 14011 40832
rect 13947 40772 13951 40828
rect 13951 40772 14007 40828
rect 14007 40772 14011 40828
rect 13947 40768 14011 40772
rect 14027 40828 14091 40832
rect 14027 40772 14031 40828
rect 14031 40772 14087 40828
rect 14087 40772 14091 40828
rect 14027 40768 14091 40772
rect 14107 40828 14171 40832
rect 14107 40772 14111 40828
rect 14111 40772 14167 40828
rect 14167 40772 14171 40828
rect 14107 40768 14171 40772
rect 14187 40828 14251 40832
rect 14187 40772 14191 40828
rect 14191 40772 14247 40828
rect 14247 40772 14251 40828
rect 14187 40768 14251 40772
rect 19145 40828 19209 40832
rect 19145 40772 19149 40828
rect 19149 40772 19205 40828
rect 19205 40772 19209 40828
rect 19145 40768 19209 40772
rect 19225 40828 19289 40832
rect 19225 40772 19229 40828
rect 19229 40772 19285 40828
rect 19285 40772 19289 40828
rect 19225 40768 19289 40772
rect 19305 40828 19369 40832
rect 19305 40772 19309 40828
rect 19309 40772 19365 40828
rect 19365 40772 19369 40828
rect 19305 40768 19369 40772
rect 19385 40828 19449 40832
rect 19385 40772 19389 40828
rect 19389 40772 19445 40828
rect 19445 40772 19449 40828
rect 19385 40768 19449 40772
rect 19932 40700 19996 40764
rect 612 40564 676 40628
rect 17908 40564 17972 40628
rect 19748 40428 19812 40492
rect 6150 40284 6214 40288
rect 6150 40228 6154 40284
rect 6154 40228 6210 40284
rect 6210 40228 6214 40284
rect 6150 40224 6214 40228
rect 6230 40284 6294 40288
rect 6230 40228 6234 40284
rect 6234 40228 6290 40284
rect 6290 40228 6294 40284
rect 6230 40224 6294 40228
rect 6310 40284 6374 40288
rect 6310 40228 6314 40284
rect 6314 40228 6370 40284
rect 6370 40228 6374 40284
rect 6310 40224 6374 40228
rect 6390 40284 6454 40288
rect 6390 40228 6394 40284
rect 6394 40228 6450 40284
rect 6450 40228 6454 40284
rect 6390 40224 6454 40228
rect 11348 40284 11412 40288
rect 11348 40228 11352 40284
rect 11352 40228 11408 40284
rect 11408 40228 11412 40284
rect 11348 40224 11412 40228
rect 11428 40284 11492 40288
rect 11428 40228 11432 40284
rect 11432 40228 11488 40284
rect 11488 40228 11492 40284
rect 11428 40224 11492 40228
rect 11508 40284 11572 40288
rect 11508 40228 11512 40284
rect 11512 40228 11568 40284
rect 11568 40228 11572 40284
rect 11508 40224 11572 40228
rect 11588 40284 11652 40288
rect 11588 40228 11592 40284
rect 11592 40228 11648 40284
rect 11648 40228 11652 40284
rect 11588 40224 11652 40228
rect 16546 40284 16610 40288
rect 16546 40228 16550 40284
rect 16550 40228 16606 40284
rect 16606 40228 16610 40284
rect 16546 40224 16610 40228
rect 16626 40284 16690 40288
rect 16626 40228 16630 40284
rect 16630 40228 16686 40284
rect 16686 40228 16690 40284
rect 16626 40224 16690 40228
rect 16706 40284 16770 40288
rect 16706 40228 16710 40284
rect 16710 40228 16766 40284
rect 16766 40228 16770 40284
rect 16706 40224 16770 40228
rect 16786 40284 16850 40288
rect 16786 40228 16790 40284
rect 16790 40228 16846 40284
rect 16846 40228 16850 40284
rect 16786 40224 16850 40228
rect 21744 40284 21808 40288
rect 21744 40228 21748 40284
rect 21748 40228 21804 40284
rect 21804 40228 21808 40284
rect 21744 40224 21808 40228
rect 21824 40284 21888 40288
rect 21824 40228 21828 40284
rect 21828 40228 21884 40284
rect 21884 40228 21888 40284
rect 21824 40224 21888 40228
rect 21904 40284 21968 40288
rect 21904 40228 21908 40284
rect 21908 40228 21964 40284
rect 21964 40228 21968 40284
rect 21904 40224 21968 40228
rect 21984 40284 22048 40288
rect 21984 40228 21988 40284
rect 21988 40228 22044 40284
rect 22044 40228 22048 40284
rect 21984 40224 22048 40228
rect 5396 40156 5460 40220
rect 19012 40080 19076 40084
rect 19012 40024 19062 40080
rect 19062 40024 19076 40080
rect 19012 40020 19076 40024
rect 19564 40020 19628 40084
rect 5028 39884 5092 39948
rect 19932 39884 19996 39948
rect 3551 39740 3615 39744
rect 3551 39684 3555 39740
rect 3555 39684 3611 39740
rect 3611 39684 3615 39740
rect 3551 39680 3615 39684
rect 3631 39740 3695 39744
rect 3631 39684 3635 39740
rect 3635 39684 3691 39740
rect 3691 39684 3695 39740
rect 3631 39680 3695 39684
rect 3711 39740 3775 39744
rect 3711 39684 3715 39740
rect 3715 39684 3771 39740
rect 3771 39684 3775 39740
rect 3711 39680 3775 39684
rect 3791 39740 3855 39744
rect 3791 39684 3795 39740
rect 3795 39684 3851 39740
rect 3851 39684 3855 39740
rect 3791 39680 3855 39684
rect 8749 39740 8813 39744
rect 8749 39684 8753 39740
rect 8753 39684 8809 39740
rect 8809 39684 8813 39740
rect 8749 39680 8813 39684
rect 8829 39740 8893 39744
rect 8829 39684 8833 39740
rect 8833 39684 8889 39740
rect 8889 39684 8893 39740
rect 8829 39680 8893 39684
rect 8909 39740 8973 39744
rect 8909 39684 8913 39740
rect 8913 39684 8969 39740
rect 8969 39684 8973 39740
rect 8909 39680 8973 39684
rect 8989 39740 9053 39744
rect 8989 39684 8993 39740
rect 8993 39684 9049 39740
rect 9049 39684 9053 39740
rect 8989 39680 9053 39684
rect 13947 39740 14011 39744
rect 13947 39684 13951 39740
rect 13951 39684 14007 39740
rect 14007 39684 14011 39740
rect 13947 39680 14011 39684
rect 14027 39740 14091 39744
rect 14027 39684 14031 39740
rect 14031 39684 14087 39740
rect 14087 39684 14091 39740
rect 14027 39680 14091 39684
rect 14107 39740 14171 39744
rect 14107 39684 14111 39740
rect 14111 39684 14167 39740
rect 14167 39684 14171 39740
rect 14107 39680 14171 39684
rect 14187 39740 14251 39744
rect 14187 39684 14191 39740
rect 14191 39684 14247 39740
rect 14247 39684 14251 39740
rect 14187 39680 14251 39684
rect 19145 39740 19209 39744
rect 19145 39684 19149 39740
rect 19149 39684 19205 39740
rect 19205 39684 19209 39740
rect 19145 39680 19209 39684
rect 19225 39740 19289 39744
rect 19225 39684 19229 39740
rect 19229 39684 19285 39740
rect 19285 39684 19289 39740
rect 19225 39680 19289 39684
rect 19305 39740 19369 39744
rect 19305 39684 19309 39740
rect 19309 39684 19365 39740
rect 19365 39684 19369 39740
rect 19305 39680 19369 39684
rect 19385 39740 19449 39744
rect 19385 39684 19389 39740
rect 19389 39684 19445 39740
rect 19445 39684 19449 39740
rect 19385 39680 19449 39684
rect 6150 39196 6214 39200
rect 6150 39140 6154 39196
rect 6154 39140 6210 39196
rect 6210 39140 6214 39196
rect 6150 39136 6214 39140
rect 6230 39196 6294 39200
rect 6230 39140 6234 39196
rect 6234 39140 6290 39196
rect 6290 39140 6294 39196
rect 6230 39136 6294 39140
rect 6310 39196 6374 39200
rect 6310 39140 6314 39196
rect 6314 39140 6370 39196
rect 6370 39140 6374 39196
rect 6310 39136 6374 39140
rect 6390 39196 6454 39200
rect 6390 39140 6394 39196
rect 6394 39140 6450 39196
rect 6450 39140 6454 39196
rect 6390 39136 6454 39140
rect 11348 39196 11412 39200
rect 11348 39140 11352 39196
rect 11352 39140 11408 39196
rect 11408 39140 11412 39196
rect 11348 39136 11412 39140
rect 11428 39196 11492 39200
rect 11428 39140 11432 39196
rect 11432 39140 11488 39196
rect 11488 39140 11492 39196
rect 11428 39136 11492 39140
rect 11508 39196 11572 39200
rect 11508 39140 11512 39196
rect 11512 39140 11568 39196
rect 11568 39140 11572 39196
rect 11508 39136 11572 39140
rect 11588 39196 11652 39200
rect 11588 39140 11592 39196
rect 11592 39140 11648 39196
rect 11648 39140 11652 39196
rect 11588 39136 11652 39140
rect 16546 39196 16610 39200
rect 16546 39140 16550 39196
rect 16550 39140 16606 39196
rect 16606 39140 16610 39196
rect 16546 39136 16610 39140
rect 16626 39196 16690 39200
rect 16626 39140 16630 39196
rect 16630 39140 16686 39196
rect 16686 39140 16690 39196
rect 16626 39136 16690 39140
rect 16706 39196 16770 39200
rect 16706 39140 16710 39196
rect 16710 39140 16766 39196
rect 16766 39140 16770 39196
rect 16706 39136 16770 39140
rect 16786 39196 16850 39200
rect 16786 39140 16790 39196
rect 16790 39140 16846 39196
rect 16846 39140 16850 39196
rect 16786 39136 16850 39140
rect 21744 39196 21808 39200
rect 21744 39140 21748 39196
rect 21748 39140 21804 39196
rect 21804 39140 21808 39196
rect 21744 39136 21808 39140
rect 21824 39196 21888 39200
rect 21824 39140 21828 39196
rect 21828 39140 21884 39196
rect 21884 39140 21888 39196
rect 21824 39136 21888 39140
rect 21904 39196 21968 39200
rect 21904 39140 21908 39196
rect 21908 39140 21964 39196
rect 21964 39140 21968 39196
rect 21904 39136 21968 39140
rect 21984 39196 22048 39200
rect 21984 39140 21988 39196
rect 21988 39140 22044 39196
rect 22044 39140 22048 39196
rect 21984 39136 22048 39140
rect 18092 38932 18156 38996
rect 2268 38660 2332 38724
rect 15332 38660 15396 38724
rect 18276 38660 18340 38724
rect 20116 38660 20180 38724
rect 3551 38652 3615 38656
rect 3551 38596 3555 38652
rect 3555 38596 3611 38652
rect 3611 38596 3615 38652
rect 3551 38592 3615 38596
rect 3631 38652 3695 38656
rect 3631 38596 3635 38652
rect 3635 38596 3691 38652
rect 3691 38596 3695 38652
rect 3631 38592 3695 38596
rect 3711 38652 3775 38656
rect 3711 38596 3715 38652
rect 3715 38596 3771 38652
rect 3771 38596 3775 38652
rect 3711 38592 3775 38596
rect 3791 38652 3855 38656
rect 3791 38596 3795 38652
rect 3795 38596 3851 38652
rect 3851 38596 3855 38652
rect 3791 38592 3855 38596
rect 8749 38652 8813 38656
rect 8749 38596 8753 38652
rect 8753 38596 8809 38652
rect 8809 38596 8813 38652
rect 8749 38592 8813 38596
rect 8829 38652 8893 38656
rect 8829 38596 8833 38652
rect 8833 38596 8889 38652
rect 8889 38596 8893 38652
rect 8829 38592 8893 38596
rect 8909 38652 8973 38656
rect 8909 38596 8913 38652
rect 8913 38596 8969 38652
rect 8969 38596 8973 38652
rect 8909 38592 8973 38596
rect 8989 38652 9053 38656
rect 8989 38596 8993 38652
rect 8993 38596 9049 38652
rect 9049 38596 9053 38652
rect 8989 38592 9053 38596
rect 13947 38652 14011 38656
rect 13947 38596 13951 38652
rect 13951 38596 14007 38652
rect 14007 38596 14011 38652
rect 13947 38592 14011 38596
rect 14027 38652 14091 38656
rect 14027 38596 14031 38652
rect 14031 38596 14087 38652
rect 14087 38596 14091 38652
rect 14027 38592 14091 38596
rect 14107 38652 14171 38656
rect 14107 38596 14111 38652
rect 14111 38596 14167 38652
rect 14167 38596 14171 38652
rect 14107 38592 14171 38596
rect 14187 38652 14251 38656
rect 14187 38596 14191 38652
rect 14191 38596 14247 38652
rect 14247 38596 14251 38652
rect 14187 38592 14251 38596
rect 19145 38652 19209 38656
rect 19145 38596 19149 38652
rect 19149 38596 19205 38652
rect 19205 38596 19209 38652
rect 19145 38592 19209 38596
rect 19225 38652 19289 38656
rect 19225 38596 19229 38652
rect 19229 38596 19285 38652
rect 19285 38596 19289 38652
rect 19225 38592 19289 38596
rect 19305 38652 19369 38656
rect 19305 38596 19309 38652
rect 19309 38596 19365 38652
rect 19365 38596 19369 38652
rect 19305 38592 19369 38596
rect 19385 38652 19449 38656
rect 19385 38596 19389 38652
rect 19389 38596 19445 38652
rect 19445 38596 19449 38652
rect 19385 38592 19449 38596
rect 8156 38388 8220 38452
rect 12572 38388 12636 38452
rect 6150 38108 6214 38112
rect 6150 38052 6154 38108
rect 6154 38052 6210 38108
rect 6210 38052 6214 38108
rect 6150 38048 6214 38052
rect 6230 38108 6294 38112
rect 6230 38052 6234 38108
rect 6234 38052 6290 38108
rect 6290 38052 6294 38108
rect 6230 38048 6294 38052
rect 6310 38108 6374 38112
rect 6310 38052 6314 38108
rect 6314 38052 6370 38108
rect 6370 38052 6374 38108
rect 6310 38048 6374 38052
rect 6390 38108 6454 38112
rect 6390 38052 6394 38108
rect 6394 38052 6450 38108
rect 6450 38052 6454 38108
rect 6390 38048 6454 38052
rect 11348 38108 11412 38112
rect 11348 38052 11352 38108
rect 11352 38052 11408 38108
rect 11408 38052 11412 38108
rect 11348 38048 11412 38052
rect 11428 38108 11492 38112
rect 11428 38052 11432 38108
rect 11432 38052 11488 38108
rect 11488 38052 11492 38108
rect 11428 38048 11492 38052
rect 11508 38108 11572 38112
rect 11508 38052 11512 38108
rect 11512 38052 11568 38108
rect 11568 38052 11572 38108
rect 11508 38048 11572 38052
rect 11588 38108 11652 38112
rect 11588 38052 11592 38108
rect 11592 38052 11648 38108
rect 11648 38052 11652 38108
rect 11588 38048 11652 38052
rect 16546 38108 16610 38112
rect 16546 38052 16550 38108
rect 16550 38052 16606 38108
rect 16606 38052 16610 38108
rect 16546 38048 16610 38052
rect 16626 38108 16690 38112
rect 16626 38052 16630 38108
rect 16630 38052 16686 38108
rect 16686 38052 16690 38108
rect 16626 38048 16690 38052
rect 16706 38108 16770 38112
rect 16706 38052 16710 38108
rect 16710 38052 16766 38108
rect 16766 38052 16770 38108
rect 16706 38048 16770 38052
rect 16786 38108 16850 38112
rect 16786 38052 16790 38108
rect 16790 38052 16846 38108
rect 16846 38052 16850 38108
rect 16786 38048 16850 38052
rect 21744 38108 21808 38112
rect 21744 38052 21748 38108
rect 21748 38052 21804 38108
rect 21804 38052 21808 38108
rect 21744 38048 21808 38052
rect 21824 38108 21888 38112
rect 21824 38052 21828 38108
rect 21828 38052 21884 38108
rect 21884 38052 21888 38108
rect 21824 38048 21888 38052
rect 21904 38108 21968 38112
rect 21904 38052 21908 38108
rect 21908 38052 21964 38108
rect 21964 38052 21968 38108
rect 21904 38048 21968 38052
rect 21984 38108 22048 38112
rect 21984 38052 21988 38108
rect 21988 38052 22044 38108
rect 22044 38052 22048 38108
rect 21984 38048 22048 38052
rect 9812 37708 9876 37772
rect 4844 37632 4908 37636
rect 4844 37576 4894 37632
rect 4894 37576 4908 37632
rect 4844 37572 4908 37576
rect 3551 37564 3615 37568
rect 3551 37508 3555 37564
rect 3555 37508 3611 37564
rect 3611 37508 3615 37564
rect 3551 37504 3615 37508
rect 3631 37564 3695 37568
rect 3631 37508 3635 37564
rect 3635 37508 3691 37564
rect 3691 37508 3695 37564
rect 3631 37504 3695 37508
rect 3711 37564 3775 37568
rect 3711 37508 3715 37564
rect 3715 37508 3771 37564
rect 3771 37508 3775 37564
rect 3711 37504 3775 37508
rect 3791 37564 3855 37568
rect 3791 37508 3795 37564
rect 3795 37508 3851 37564
rect 3851 37508 3855 37564
rect 3791 37504 3855 37508
rect 8749 37564 8813 37568
rect 8749 37508 8753 37564
rect 8753 37508 8809 37564
rect 8809 37508 8813 37564
rect 8749 37504 8813 37508
rect 8829 37564 8893 37568
rect 8829 37508 8833 37564
rect 8833 37508 8889 37564
rect 8889 37508 8893 37564
rect 8829 37504 8893 37508
rect 8909 37564 8973 37568
rect 8909 37508 8913 37564
rect 8913 37508 8969 37564
rect 8969 37508 8973 37564
rect 8909 37504 8973 37508
rect 8989 37564 9053 37568
rect 8989 37508 8993 37564
rect 8993 37508 9049 37564
rect 9049 37508 9053 37564
rect 8989 37504 9053 37508
rect 13947 37564 14011 37568
rect 13947 37508 13951 37564
rect 13951 37508 14007 37564
rect 14007 37508 14011 37564
rect 13947 37504 14011 37508
rect 14027 37564 14091 37568
rect 14027 37508 14031 37564
rect 14031 37508 14087 37564
rect 14087 37508 14091 37564
rect 14027 37504 14091 37508
rect 14107 37564 14171 37568
rect 14107 37508 14111 37564
rect 14111 37508 14167 37564
rect 14167 37508 14171 37564
rect 14107 37504 14171 37508
rect 14187 37564 14251 37568
rect 14187 37508 14191 37564
rect 14191 37508 14247 37564
rect 14247 37508 14251 37564
rect 14187 37504 14251 37508
rect 19145 37564 19209 37568
rect 19145 37508 19149 37564
rect 19149 37508 19205 37564
rect 19205 37508 19209 37564
rect 19145 37504 19209 37508
rect 19225 37564 19289 37568
rect 19225 37508 19229 37564
rect 19229 37508 19285 37564
rect 19285 37508 19289 37564
rect 19225 37504 19289 37508
rect 19305 37564 19369 37568
rect 19305 37508 19309 37564
rect 19309 37508 19365 37564
rect 19365 37508 19369 37564
rect 19305 37504 19369 37508
rect 19385 37564 19449 37568
rect 19385 37508 19389 37564
rect 19389 37508 19445 37564
rect 19445 37508 19449 37564
rect 19385 37504 19449 37508
rect 7972 37300 8036 37364
rect 8524 37164 8588 37228
rect 14412 37164 14476 37228
rect 7788 37088 7852 37092
rect 7788 37032 7802 37088
rect 7802 37032 7852 37088
rect 7788 37028 7852 37032
rect 6150 37020 6214 37024
rect 6150 36964 6154 37020
rect 6154 36964 6210 37020
rect 6210 36964 6214 37020
rect 6150 36960 6214 36964
rect 6230 37020 6294 37024
rect 6230 36964 6234 37020
rect 6234 36964 6290 37020
rect 6290 36964 6294 37020
rect 6230 36960 6294 36964
rect 6310 37020 6374 37024
rect 6310 36964 6314 37020
rect 6314 36964 6370 37020
rect 6370 36964 6374 37020
rect 6310 36960 6374 36964
rect 6390 37020 6454 37024
rect 6390 36964 6394 37020
rect 6394 36964 6450 37020
rect 6450 36964 6454 37020
rect 6390 36960 6454 36964
rect 11348 37020 11412 37024
rect 11348 36964 11352 37020
rect 11352 36964 11408 37020
rect 11408 36964 11412 37020
rect 11348 36960 11412 36964
rect 11428 37020 11492 37024
rect 11428 36964 11432 37020
rect 11432 36964 11488 37020
rect 11488 36964 11492 37020
rect 11428 36960 11492 36964
rect 11508 37020 11572 37024
rect 11508 36964 11512 37020
rect 11512 36964 11568 37020
rect 11568 36964 11572 37020
rect 11508 36960 11572 36964
rect 11588 37020 11652 37024
rect 11588 36964 11592 37020
rect 11592 36964 11648 37020
rect 11648 36964 11652 37020
rect 11588 36960 11652 36964
rect 16546 37020 16610 37024
rect 16546 36964 16550 37020
rect 16550 36964 16606 37020
rect 16606 36964 16610 37020
rect 16546 36960 16610 36964
rect 16626 37020 16690 37024
rect 16626 36964 16630 37020
rect 16630 36964 16686 37020
rect 16686 36964 16690 37020
rect 16626 36960 16690 36964
rect 16706 37020 16770 37024
rect 16706 36964 16710 37020
rect 16710 36964 16766 37020
rect 16766 36964 16770 37020
rect 16706 36960 16770 36964
rect 16786 37020 16850 37024
rect 16786 36964 16790 37020
rect 16790 36964 16846 37020
rect 16846 36964 16850 37020
rect 16786 36960 16850 36964
rect 21744 37020 21808 37024
rect 21744 36964 21748 37020
rect 21748 36964 21804 37020
rect 21804 36964 21808 37020
rect 21744 36960 21808 36964
rect 21824 37020 21888 37024
rect 21824 36964 21828 37020
rect 21828 36964 21884 37020
rect 21884 36964 21888 37020
rect 21824 36960 21888 36964
rect 21904 37020 21968 37024
rect 21904 36964 21908 37020
rect 21908 36964 21964 37020
rect 21964 36964 21968 37020
rect 21904 36960 21968 36964
rect 21984 37020 22048 37024
rect 21984 36964 21988 37020
rect 21988 36964 22044 37020
rect 22044 36964 22048 37020
rect 21984 36960 22048 36964
rect 6684 36756 6748 36820
rect 6868 36816 6932 36820
rect 6868 36760 6918 36816
rect 6918 36760 6932 36816
rect 6868 36756 6932 36760
rect 2268 36620 2332 36684
rect 7236 36620 7300 36684
rect 14780 36620 14844 36684
rect 5028 36484 5092 36548
rect 3551 36476 3615 36480
rect 3551 36420 3555 36476
rect 3555 36420 3611 36476
rect 3611 36420 3615 36476
rect 3551 36416 3615 36420
rect 3631 36476 3695 36480
rect 3631 36420 3635 36476
rect 3635 36420 3691 36476
rect 3691 36420 3695 36476
rect 3631 36416 3695 36420
rect 3711 36476 3775 36480
rect 3711 36420 3715 36476
rect 3715 36420 3771 36476
rect 3771 36420 3775 36476
rect 3711 36416 3775 36420
rect 3791 36476 3855 36480
rect 3791 36420 3795 36476
rect 3795 36420 3851 36476
rect 3851 36420 3855 36476
rect 3791 36416 3855 36420
rect 8749 36476 8813 36480
rect 8749 36420 8753 36476
rect 8753 36420 8809 36476
rect 8809 36420 8813 36476
rect 8749 36416 8813 36420
rect 8829 36476 8893 36480
rect 8829 36420 8833 36476
rect 8833 36420 8889 36476
rect 8889 36420 8893 36476
rect 8829 36416 8893 36420
rect 8909 36476 8973 36480
rect 8909 36420 8913 36476
rect 8913 36420 8969 36476
rect 8969 36420 8973 36476
rect 8909 36416 8973 36420
rect 8989 36476 9053 36480
rect 8989 36420 8993 36476
rect 8993 36420 9049 36476
rect 9049 36420 9053 36476
rect 8989 36416 9053 36420
rect 13947 36476 14011 36480
rect 13947 36420 13951 36476
rect 13951 36420 14007 36476
rect 14007 36420 14011 36476
rect 13947 36416 14011 36420
rect 14027 36476 14091 36480
rect 14027 36420 14031 36476
rect 14031 36420 14087 36476
rect 14087 36420 14091 36476
rect 14027 36416 14091 36420
rect 14107 36476 14171 36480
rect 14107 36420 14111 36476
rect 14111 36420 14167 36476
rect 14167 36420 14171 36476
rect 14107 36416 14171 36420
rect 14187 36476 14251 36480
rect 14187 36420 14191 36476
rect 14191 36420 14247 36476
rect 14247 36420 14251 36476
rect 14187 36416 14251 36420
rect 19145 36476 19209 36480
rect 19145 36420 19149 36476
rect 19149 36420 19205 36476
rect 19205 36420 19209 36476
rect 19145 36416 19209 36420
rect 19225 36476 19289 36480
rect 19225 36420 19229 36476
rect 19229 36420 19285 36476
rect 19285 36420 19289 36476
rect 19225 36416 19289 36420
rect 19305 36476 19369 36480
rect 19305 36420 19309 36476
rect 19309 36420 19365 36476
rect 19365 36420 19369 36476
rect 19305 36416 19369 36420
rect 19385 36476 19449 36480
rect 19385 36420 19389 36476
rect 19389 36420 19445 36476
rect 19445 36420 19449 36476
rect 19385 36416 19449 36420
rect 15516 36212 15580 36276
rect 17724 36212 17788 36276
rect 7604 35940 7668 36004
rect 9996 35940 10060 36004
rect 10732 35940 10796 36004
rect 6150 35932 6214 35936
rect 6150 35876 6154 35932
rect 6154 35876 6210 35932
rect 6210 35876 6214 35932
rect 6150 35872 6214 35876
rect 6230 35932 6294 35936
rect 6230 35876 6234 35932
rect 6234 35876 6290 35932
rect 6290 35876 6294 35932
rect 6230 35872 6294 35876
rect 6310 35932 6374 35936
rect 6310 35876 6314 35932
rect 6314 35876 6370 35932
rect 6370 35876 6374 35932
rect 6310 35872 6374 35876
rect 6390 35932 6454 35936
rect 6390 35876 6394 35932
rect 6394 35876 6450 35932
rect 6450 35876 6454 35932
rect 6390 35872 6454 35876
rect 11348 35932 11412 35936
rect 11348 35876 11352 35932
rect 11352 35876 11408 35932
rect 11408 35876 11412 35932
rect 11348 35872 11412 35876
rect 11428 35932 11492 35936
rect 11428 35876 11432 35932
rect 11432 35876 11488 35932
rect 11488 35876 11492 35932
rect 11428 35872 11492 35876
rect 11508 35932 11572 35936
rect 11508 35876 11512 35932
rect 11512 35876 11568 35932
rect 11568 35876 11572 35932
rect 11508 35872 11572 35876
rect 11588 35932 11652 35936
rect 11588 35876 11592 35932
rect 11592 35876 11648 35932
rect 11648 35876 11652 35932
rect 11588 35872 11652 35876
rect 16546 35932 16610 35936
rect 16546 35876 16550 35932
rect 16550 35876 16606 35932
rect 16606 35876 16610 35932
rect 16546 35872 16610 35876
rect 16626 35932 16690 35936
rect 16626 35876 16630 35932
rect 16630 35876 16686 35932
rect 16686 35876 16690 35932
rect 16626 35872 16690 35876
rect 16706 35932 16770 35936
rect 16706 35876 16710 35932
rect 16710 35876 16766 35932
rect 16766 35876 16770 35932
rect 16706 35872 16770 35876
rect 16786 35932 16850 35936
rect 16786 35876 16790 35932
rect 16790 35876 16846 35932
rect 16846 35876 16850 35932
rect 16786 35872 16850 35876
rect 21744 35932 21808 35936
rect 21744 35876 21748 35932
rect 21748 35876 21804 35932
rect 21804 35876 21808 35932
rect 21744 35872 21808 35876
rect 21824 35932 21888 35936
rect 21824 35876 21828 35932
rect 21828 35876 21884 35932
rect 21884 35876 21888 35932
rect 21824 35872 21888 35876
rect 21904 35932 21968 35936
rect 21904 35876 21908 35932
rect 21908 35876 21964 35932
rect 21964 35876 21968 35932
rect 21904 35872 21968 35876
rect 21984 35932 22048 35936
rect 21984 35876 21988 35932
rect 21988 35876 22044 35932
rect 22044 35876 22048 35932
rect 21984 35872 22048 35876
rect 5764 35804 5828 35868
rect 8340 35804 8404 35868
rect 11100 35804 11164 35868
rect 15332 35532 15396 35596
rect 5396 35396 5460 35460
rect 9444 35456 9508 35460
rect 9444 35400 9458 35456
rect 9458 35400 9508 35456
rect 9444 35396 9508 35400
rect 3551 35388 3615 35392
rect 3551 35332 3555 35388
rect 3555 35332 3611 35388
rect 3611 35332 3615 35388
rect 3551 35328 3615 35332
rect 3631 35388 3695 35392
rect 3631 35332 3635 35388
rect 3635 35332 3691 35388
rect 3691 35332 3695 35388
rect 3631 35328 3695 35332
rect 3711 35388 3775 35392
rect 3711 35332 3715 35388
rect 3715 35332 3771 35388
rect 3771 35332 3775 35388
rect 3711 35328 3775 35332
rect 3791 35388 3855 35392
rect 3791 35332 3795 35388
rect 3795 35332 3851 35388
rect 3851 35332 3855 35388
rect 3791 35328 3855 35332
rect 8749 35388 8813 35392
rect 8749 35332 8753 35388
rect 8753 35332 8809 35388
rect 8809 35332 8813 35388
rect 8749 35328 8813 35332
rect 8829 35388 8893 35392
rect 8829 35332 8833 35388
rect 8833 35332 8889 35388
rect 8889 35332 8893 35388
rect 8829 35328 8893 35332
rect 8909 35388 8973 35392
rect 8909 35332 8913 35388
rect 8913 35332 8969 35388
rect 8969 35332 8973 35388
rect 8909 35328 8973 35332
rect 8989 35388 9053 35392
rect 8989 35332 8993 35388
rect 8993 35332 9049 35388
rect 9049 35332 9053 35388
rect 8989 35328 9053 35332
rect 13947 35388 14011 35392
rect 13947 35332 13951 35388
rect 13951 35332 14007 35388
rect 14007 35332 14011 35388
rect 13947 35328 14011 35332
rect 14027 35388 14091 35392
rect 14027 35332 14031 35388
rect 14031 35332 14087 35388
rect 14087 35332 14091 35388
rect 14027 35328 14091 35332
rect 14107 35388 14171 35392
rect 14107 35332 14111 35388
rect 14111 35332 14167 35388
rect 14167 35332 14171 35388
rect 14107 35328 14171 35332
rect 14187 35388 14251 35392
rect 14187 35332 14191 35388
rect 14191 35332 14247 35388
rect 14247 35332 14251 35388
rect 14187 35328 14251 35332
rect 19145 35388 19209 35392
rect 19145 35332 19149 35388
rect 19149 35332 19205 35388
rect 19205 35332 19209 35388
rect 19145 35328 19209 35332
rect 19225 35388 19289 35392
rect 19225 35332 19229 35388
rect 19229 35332 19285 35388
rect 19285 35332 19289 35388
rect 19225 35328 19289 35332
rect 19305 35388 19369 35392
rect 19305 35332 19309 35388
rect 19309 35332 19365 35388
rect 19365 35332 19369 35388
rect 19305 35328 19369 35332
rect 19385 35388 19449 35392
rect 19385 35332 19389 35388
rect 19389 35332 19445 35388
rect 19445 35332 19449 35388
rect 19385 35328 19449 35332
rect 1716 35320 1780 35324
rect 1716 35264 1730 35320
rect 1730 35264 1780 35320
rect 1716 35260 1780 35264
rect 2452 35260 2516 35324
rect 5948 34912 6012 34916
rect 5948 34856 5998 34912
rect 5998 34856 6012 34912
rect 5948 34852 6012 34856
rect 6150 34844 6214 34848
rect 6150 34788 6154 34844
rect 6154 34788 6210 34844
rect 6210 34788 6214 34844
rect 6150 34784 6214 34788
rect 6230 34844 6294 34848
rect 6230 34788 6234 34844
rect 6234 34788 6290 34844
rect 6290 34788 6294 34844
rect 6230 34784 6294 34788
rect 6310 34844 6374 34848
rect 6310 34788 6314 34844
rect 6314 34788 6370 34844
rect 6370 34788 6374 34844
rect 6310 34784 6374 34788
rect 6390 34844 6454 34848
rect 6390 34788 6394 34844
rect 6394 34788 6450 34844
rect 6450 34788 6454 34844
rect 6390 34784 6454 34788
rect 11348 34844 11412 34848
rect 11348 34788 11352 34844
rect 11352 34788 11408 34844
rect 11408 34788 11412 34844
rect 11348 34784 11412 34788
rect 11428 34844 11492 34848
rect 11428 34788 11432 34844
rect 11432 34788 11488 34844
rect 11488 34788 11492 34844
rect 11428 34784 11492 34788
rect 11508 34844 11572 34848
rect 11508 34788 11512 34844
rect 11512 34788 11568 34844
rect 11568 34788 11572 34844
rect 11508 34784 11572 34788
rect 11588 34844 11652 34848
rect 11588 34788 11592 34844
rect 11592 34788 11648 34844
rect 11648 34788 11652 34844
rect 11588 34784 11652 34788
rect 16546 34844 16610 34848
rect 16546 34788 16550 34844
rect 16550 34788 16606 34844
rect 16606 34788 16610 34844
rect 16546 34784 16610 34788
rect 16626 34844 16690 34848
rect 16626 34788 16630 34844
rect 16630 34788 16686 34844
rect 16686 34788 16690 34844
rect 16626 34784 16690 34788
rect 16706 34844 16770 34848
rect 16706 34788 16710 34844
rect 16710 34788 16766 34844
rect 16766 34788 16770 34844
rect 16706 34784 16770 34788
rect 16786 34844 16850 34848
rect 16786 34788 16790 34844
rect 16790 34788 16846 34844
rect 16846 34788 16850 34844
rect 16786 34784 16850 34788
rect 21744 34844 21808 34848
rect 21744 34788 21748 34844
rect 21748 34788 21804 34844
rect 21804 34788 21808 34844
rect 21744 34784 21808 34788
rect 21824 34844 21888 34848
rect 21824 34788 21828 34844
rect 21828 34788 21884 34844
rect 21884 34788 21888 34844
rect 21824 34784 21888 34788
rect 21904 34844 21968 34848
rect 21904 34788 21908 34844
rect 21908 34788 21964 34844
rect 21964 34788 21968 34844
rect 21904 34784 21968 34788
rect 21984 34844 22048 34848
rect 21984 34788 21988 34844
rect 21988 34788 22044 34844
rect 22044 34788 22048 34844
rect 21984 34784 22048 34788
rect 980 34444 1044 34508
rect 3004 34580 3068 34644
rect 10916 34580 10980 34644
rect 11836 34640 11900 34644
rect 11836 34584 11850 34640
rect 11850 34584 11900 34640
rect 11836 34580 11900 34584
rect 21036 34444 21100 34508
rect 3551 34300 3615 34304
rect 3551 34244 3555 34300
rect 3555 34244 3611 34300
rect 3611 34244 3615 34300
rect 3551 34240 3615 34244
rect 3631 34300 3695 34304
rect 3631 34244 3635 34300
rect 3635 34244 3691 34300
rect 3691 34244 3695 34300
rect 3631 34240 3695 34244
rect 3711 34300 3775 34304
rect 3711 34244 3715 34300
rect 3715 34244 3771 34300
rect 3771 34244 3775 34300
rect 3711 34240 3775 34244
rect 3791 34300 3855 34304
rect 3791 34244 3795 34300
rect 3795 34244 3851 34300
rect 3851 34244 3855 34300
rect 3791 34240 3855 34244
rect 8749 34300 8813 34304
rect 8749 34244 8753 34300
rect 8753 34244 8809 34300
rect 8809 34244 8813 34300
rect 8749 34240 8813 34244
rect 8829 34300 8893 34304
rect 8829 34244 8833 34300
rect 8833 34244 8889 34300
rect 8889 34244 8893 34300
rect 8829 34240 8893 34244
rect 8909 34300 8973 34304
rect 8909 34244 8913 34300
rect 8913 34244 8969 34300
rect 8969 34244 8973 34300
rect 8909 34240 8973 34244
rect 8989 34300 9053 34304
rect 8989 34244 8993 34300
rect 8993 34244 9049 34300
rect 9049 34244 9053 34300
rect 8989 34240 9053 34244
rect 13947 34300 14011 34304
rect 13947 34244 13951 34300
rect 13951 34244 14007 34300
rect 14007 34244 14011 34300
rect 13947 34240 14011 34244
rect 14027 34300 14091 34304
rect 14027 34244 14031 34300
rect 14031 34244 14087 34300
rect 14087 34244 14091 34300
rect 14027 34240 14091 34244
rect 14107 34300 14171 34304
rect 14107 34244 14111 34300
rect 14111 34244 14167 34300
rect 14167 34244 14171 34300
rect 14107 34240 14171 34244
rect 14187 34300 14251 34304
rect 14187 34244 14191 34300
rect 14191 34244 14247 34300
rect 14247 34244 14251 34300
rect 14187 34240 14251 34244
rect 19145 34300 19209 34304
rect 19145 34244 19149 34300
rect 19149 34244 19205 34300
rect 19205 34244 19209 34300
rect 19145 34240 19209 34244
rect 19225 34300 19289 34304
rect 19225 34244 19229 34300
rect 19229 34244 19285 34300
rect 19285 34244 19289 34300
rect 19225 34240 19289 34244
rect 19305 34300 19369 34304
rect 19305 34244 19309 34300
rect 19309 34244 19365 34300
rect 19365 34244 19369 34300
rect 19305 34240 19369 34244
rect 19385 34300 19449 34304
rect 19385 34244 19389 34300
rect 19389 34244 19445 34300
rect 19445 34244 19449 34300
rect 19385 34240 19449 34244
rect 6684 34172 6748 34236
rect 3924 33900 3988 33964
rect 18092 34036 18156 34100
rect 15884 33824 15948 33828
rect 15884 33768 15898 33824
rect 15898 33768 15948 33824
rect 15884 33764 15948 33768
rect 6150 33756 6214 33760
rect 6150 33700 6154 33756
rect 6154 33700 6210 33756
rect 6210 33700 6214 33756
rect 6150 33696 6214 33700
rect 6230 33756 6294 33760
rect 6230 33700 6234 33756
rect 6234 33700 6290 33756
rect 6290 33700 6294 33756
rect 6230 33696 6294 33700
rect 6310 33756 6374 33760
rect 6310 33700 6314 33756
rect 6314 33700 6370 33756
rect 6370 33700 6374 33756
rect 6310 33696 6374 33700
rect 6390 33756 6454 33760
rect 6390 33700 6394 33756
rect 6394 33700 6450 33756
rect 6450 33700 6454 33756
rect 6390 33696 6454 33700
rect 11348 33756 11412 33760
rect 11348 33700 11352 33756
rect 11352 33700 11408 33756
rect 11408 33700 11412 33756
rect 11348 33696 11412 33700
rect 11428 33756 11492 33760
rect 11428 33700 11432 33756
rect 11432 33700 11488 33756
rect 11488 33700 11492 33756
rect 11428 33696 11492 33700
rect 11508 33756 11572 33760
rect 11508 33700 11512 33756
rect 11512 33700 11568 33756
rect 11568 33700 11572 33756
rect 11508 33696 11572 33700
rect 11588 33756 11652 33760
rect 11588 33700 11592 33756
rect 11592 33700 11648 33756
rect 11648 33700 11652 33756
rect 11588 33696 11652 33700
rect 16546 33756 16610 33760
rect 16546 33700 16550 33756
rect 16550 33700 16606 33756
rect 16606 33700 16610 33756
rect 16546 33696 16610 33700
rect 16626 33756 16690 33760
rect 16626 33700 16630 33756
rect 16630 33700 16686 33756
rect 16686 33700 16690 33756
rect 16626 33696 16690 33700
rect 16706 33756 16770 33760
rect 16706 33700 16710 33756
rect 16710 33700 16766 33756
rect 16766 33700 16770 33756
rect 16706 33696 16770 33700
rect 16786 33756 16850 33760
rect 16786 33700 16790 33756
rect 16790 33700 16846 33756
rect 16846 33700 16850 33756
rect 16786 33696 16850 33700
rect 21744 33756 21808 33760
rect 21744 33700 21748 33756
rect 21748 33700 21804 33756
rect 21804 33700 21808 33756
rect 21744 33696 21808 33700
rect 21824 33756 21888 33760
rect 21824 33700 21828 33756
rect 21828 33700 21884 33756
rect 21884 33700 21888 33756
rect 21824 33696 21888 33700
rect 21904 33756 21968 33760
rect 21904 33700 21908 33756
rect 21908 33700 21964 33756
rect 21964 33700 21968 33756
rect 21904 33696 21968 33700
rect 21984 33756 22048 33760
rect 21984 33700 21988 33756
rect 21988 33700 22044 33756
rect 22044 33700 22048 33756
rect 21984 33696 22048 33700
rect 3188 33628 3252 33692
rect 12756 33492 12820 33556
rect 17908 33628 17972 33692
rect 1532 33356 1596 33420
rect 5028 33220 5092 33284
rect 3551 33212 3615 33216
rect 3551 33156 3555 33212
rect 3555 33156 3611 33212
rect 3611 33156 3615 33212
rect 3551 33152 3615 33156
rect 3631 33212 3695 33216
rect 3631 33156 3635 33212
rect 3635 33156 3691 33212
rect 3691 33156 3695 33212
rect 3631 33152 3695 33156
rect 3711 33212 3775 33216
rect 3711 33156 3715 33212
rect 3715 33156 3771 33212
rect 3771 33156 3775 33212
rect 3711 33152 3775 33156
rect 3791 33212 3855 33216
rect 3791 33156 3795 33212
rect 3795 33156 3851 33212
rect 3851 33156 3855 33212
rect 3791 33152 3855 33156
rect 8749 33212 8813 33216
rect 8749 33156 8753 33212
rect 8753 33156 8809 33212
rect 8809 33156 8813 33212
rect 8749 33152 8813 33156
rect 8829 33212 8893 33216
rect 8829 33156 8833 33212
rect 8833 33156 8889 33212
rect 8889 33156 8893 33212
rect 8829 33152 8893 33156
rect 8909 33212 8973 33216
rect 8909 33156 8913 33212
rect 8913 33156 8969 33212
rect 8969 33156 8973 33212
rect 8909 33152 8973 33156
rect 8989 33212 9053 33216
rect 8989 33156 8993 33212
rect 8993 33156 9049 33212
rect 9049 33156 9053 33212
rect 8989 33152 9053 33156
rect 13947 33212 14011 33216
rect 13947 33156 13951 33212
rect 13951 33156 14007 33212
rect 14007 33156 14011 33212
rect 13947 33152 14011 33156
rect 14027 33212 14091 33216
rect 14027 33156 14031 33212
rect 14031 33156 14087 33212
rect 14087 33156 14091 33212
rect 14027 33152 14091 33156
rect 14107 33212 14171 33216
rect 14107 33156 14111 33212
rect 14111 33156 14167 33212
rect 14167 33156 14171 33212
rect 14107 33152 14171 33156
rect 14187 33212 14251 33216
rect 14187 33156 14191 33212
rect 14191 33156 14247 33212
rect 14247 33156 14251 33212
rect 14187 33152 14251 33156
rect 19145 33212 19209 33216
rect 19145 33156 19149 33212
rect 19149 33156 19205 33212
rect 19205 33156 19209 33212
rect 19145 33152 19209 33156
rect 19225 33212 19289 33216
rect 19225 33156 19229 33212
rect 19229 33156 19285 33212
rect 19285 33156 19289 33212
rect 19225 33152 19289 33156
rect 19305 33212 19369 33216
rect 19305 33156 19309 33212
rect 19309 33156 19365 33212
rect 19365 33156 19369 33212
rect 19305 33152 19369 33156
rect 19385 33212 19449 33216
rect 19385 33156 19389 33212
rect 19389 33156 19445 33212
rect 19445 33156 19449 33212
rect 19385 33152 19449 33156
rect 4844 33084 4908 33148
rect 12020 33084 12084 33148
rect 15148 33084 15212 33148
rect 3188 32872 3252 32876
rect 3188 32816 3238 32872
rect 3238 32816 3252 32872
rect 3188 32812 3252 32816
rect 8340 32948 8404 33012
rect 15700 32812 15764 32876
rect 20300 32812 20364 32876
rect 14780 32676 14844 32740
rect 6150 32668 6214 32672
rect 6150 32612 6154 32668
rect 6154 32612 6210 32668
rect 6210 32612 6214 32668
rect 6150 32608 6214 32612
rect 6230 32668 6294 32672
rect 6230 32612 6234 32668
rect 6234 32612 6290 32668
rect 6290 32612 6294 32668
rect 6230 32608 6294 32612
rect 6310 32668 6374 32672
rect 6310 32612 6314 32668
rect 6314 32612 6370 32668
rect 6370 32612 6374 32668
rect 6310 32608 6374 32612
rect 6390 32668 6454 32672
rect 6390 32612 6394 32668
rect 6394 32612 6450 32668
rect 6450 32612 6454 32668
rect 6390 32608 6454 32612
rect 11348 32668 11412 32672
rect 11348 32612 11352 32668
rect 11352 32612 11408 32668
rect 11408 32612 11412 32668
rect 11348 32608 11412 32612
rect 11428 32668 11492 32672
rect 11428 32612 11432 32668
rect 11432 32612 11488 32668
rect 11488 32612 11492 32668
rect 11428 32608 11492 32612
rect 11508 32668 11572 32672
rect 11508 32612 11512 32668
rect 11512 32612 11568 32668
rect 11568 32612 11572 32668
rect 11508 32608 11572 32612
rect 11588 32668 11652 32672
rect 11588 32612 11592 32668
rect 11592 32612 11648 32668
rect 11648 32612 11652 32668
rect 11588 32608 11652 32612
rect 16546 32668 16610 32672
rect 16546 32612 16550 32668
rect 16550 32612 16606 32668
rect 16606 32612 16610 32668
rect 16546 32608 16610 32612
rect 16626 32668 16690 32672
rect 16626 32612 16630 32668
rect 16630 32612 16686 32668
rect 16686 32612 16690 32668
rect 16626 32608 16690 32612
rect 16706 32668 16770 32672
rect 16706 32612 16710 32668
rect 16710 32612 16766 32668
rect 16766 32612 16770 32668
rect 16706 32608 16770 32612
rect 16786 32668 16850 32672
rect 16786 32612 16790 32668
rect 16790 32612 16846 32668
rect 16846 32612 16850 32668
rect 16786 32608 16850 32612
rect 21744 32668 21808 32672
rect 21744 32612 21748 32668
rect 21748 32612 21804 32668
rect 21804 32612 21808 32668
rect 21744 32608 21808 32612
rect 21824 32668 21888 32672
rect 21824 32612 21828 32668
rect 21828 32612 21884 32668
rect 21884 32612 21888 32668
rect 21824 32608 21888 32612
rect 21904 32668 21968 32672
rect 21904 32612 21908 32668
rect 21908 32612 21964 32668
rect 21964 32612 21968 32668
rect 21904 32608 21968 32612
rect 21984 32668 22048 32672
rect 21984 32612 21988 32668
rect 21988 32612 22044 32668
rect 22044 32612 22048 32668
rect 21984 32608 22048 32612
rect 1900 32268 1964 32332
rect 6868 32328 6932 32332
rect 6868 32272 6882 32328
rect 6882 32272 6932 32328
rect 6868 32268 6932 32272
rect 3551 32124 3615 32128
rect 3551 32068 3555 32124
rect 3555 32068 3611 32124
rect 3611 32068 3615 32124
rect 3551 32064 3615 32068
rect 3631 32124 3695 32128
rect 3631 32068 3635 32124
rect 3635 32068 3691 32124
rect 3691 32068 3695 32124
rect 3631 32064 3695 32068
rect 3711 32124 3775 32128
rect 3711 32068 3715 32124
rect 3715 32068 3771 32124
rect 3771 32068 3775 32124
rect 3711 32064 3775 32068
rect 3791 32124 3855 32128
rect 3791 32068 3795 32124
rect 3795 32068 3851 32124
rect 3851 32068 3855 32124
rect 3791 32064 3855 32068
rect 8749 32124 8813 32128
rect 8749 32068 8753 32124
rect 8753 32068 8809 32124
rect 8809 32068 8813 32124
rect 8749 32064 8813 32068
rect 8829 32124 8893 32128
rect 8829 32068 8833 32124
rect 8833 32068 8889 32124
rect 8889 32068 8893 32124
rect 8829 32064 8893 32068
rect 8909 32124 8973 32128
rect 8909 32068 8913 32124
rect 8913 32068 8969 32124
rect 8969 32068 8973 32124
rect 8909 32064 8973 32068
rect 8989 32124 9053 32128
rect 8989 32068 8993 32124
rect 8993 32068 9049 32124
rect 9049 32068 9053 32124
rect 8989 32064 9053 32068
rect 9628 32132 9692 32196
rect 9996 32132 10060 32196
rect 10364 31996 10428 32060
rect 13947 32124 14011 32128
rect 13947 32068 13951 32124
rect 13951 32068 14007 32124
rect 14007 32068 14011 32124
rect 13947 32064 14011 32068
rect 14027 32124 14091 32128
rect 14027 32068 14031 32124
rect 14031 32068 14087 32124
rect 14087 32068 14091 32124
rect 14027 32064 14091 32068
rect 14107 32124 14171 32128
rect 14107 32068 14111 32124
rect 14111 32068 14167 32124
rect 14167 32068 14171 32124
rect 14107 32064 14171 32068
rect 14187 32124 14251 32128
rect 14187 32068 14191 32124
rect 14191 32068 14247 32124
rect 14247 32068 14251 32124
rect 14187 32064 14251 32068
rect 19145 32124 19209 32128
rect 19145 32068 19149 32124
rect 19149 32068 19205 32124
rect 19205 32068 19209 32124
rect 19145 32064 19209 32068
rect 19225 32124 19289 32128
rect 19225 32068 19229 32124
rect 19229 32068 19285 32124
rect 19285 32068 19289 32124
rect 19225 32064 19289 32068
rect 19305 32124 19369 32128
rect 19305 32068 19309 32124
rect 19309 32068 19365 32124
rect 19365 32068 19369 32124
rect 19305 32064 19369 32068
rect 19385 32124 19449 32128
rect 19385 32068 19389 32124
rect 19389 32068 19445 32124
rect 19445 32068 19449 32124
rect 19385 32064 19449 32068
rect 2268 31860 2332 31924
rect 4108 31860 4172 31924
rect 2084 31784 2148 31788
rect 2084 31728 2134 31784
rect 2134 31728 2148 31784
rect 2084 31724 2148 31728
rect 4292 31724 4356 31788
rect 4660 31452 4724 31516
rect 8156 31784 8220 31788
rect 8156 31728 8170 31784
rect 8170 31728 8220 31784
rect 8156 31724 8220 31728
rect 13676 31860 13740 31924
rect 14964 31724 15028 31788
rect 15332 31724 15396 31788
rect 6150 31580 6214 31584
rect 6150 31524 6154 31580
rect 6154 31524 6210 31580
rect 6210 31524 6214 31580
rect 6150 31520 6214 31524
rect 6230 31580 6294 31584
rect 6230 31524 6234 31580
rect 6234 31524 6290 31580
rect 6290 31524 6294 31580
rect 6230 31520 6294 31524
rect 6310 31580 6374 31584
rect 6310 31524 6314 31580
rect 6314 31524 6370 31580
rect 6370 31524 6374 31580
rect 6310 31520 6374 31524
rect 6390 31580 6454 31584
rect 6390 31524 6394 31580
rect 6394 31524 6450 31580
rect 6450 31524 6454 31580
rect 6390 31520 6454 31524
rect 11348 31580 11412 31584
rect 11348 31524 11352 31580
rect 11352 31524 11408 31580
rect 11408 31524 11412 31580
rect 11348 31520 11412 31524
rect 11428 31580 11492 31584
rect 11428 31524 11432 31580
rect 11432 31524 11488 31580
rect 11488 31524 11492 31580
rect 11428 31520 11492 31524
rect 11508 31580 11572 31584
rect 11508 31524 11512 31580
rect 11512 31524 11568 31580
rect 11568 31524 11572 31580
rect 11508 31520 11572 31524
rect 11588 31580 11652 31584
rect 11588 31524 11592 31580
rect 11592 31524 11648 31580
rect 11648 31524 11652 31580
rect 11588 31520 11652 31524
rect 16546 31580 16610 31584
rect 16546 31524 16550 31580
rect 16550 31524 16606 31580
rect 16606 31524 16610 31580
rect 16546 31520 16610 31524
rect 16626 31580 16690 31584
rect 16626 31524 16630 31580
rect 16630 31524 16686 31580
rect 16686 31524 16690 31580
rect 16626 31520 16690 31524
rect 16706 31580 16770 31584
rect 16706 31524 16710 31580
rect 16710 31524 16766 31580
rect 16766 31524 16770 31580
rect 16706 31520 16770 31524
rect 16786 31580 16850 31584
rect 16786 31524 16790 31580
rect 16790 31524 16846 31580
rect 16846 31524 16850 31580
rect 16786 31520 16850 31524
rect 21744 31580 21808 31584
rect 21744 31524 21748 31580
rect 21748 31524 21804 31580
rect 21804 31524 21808 31580
rect 21744 31520 21808 31524
rect 21824 31580 21888 31584
rect 21824 31524 21828 31580
rect 21828 31524 21884 31580
rect 21884 31524 21888 31580
rect 21824 31520 21888 31524
rect 21904 31580 21968 31584
rect 21904 31524 21908 31580
rect 21908 31524 21964 31580
rect 21964 31524 21968 31580
rect 21904 31520 21968 31524
rect 21984 31580 22048 31584
rect 21984 31524 21988 31580
rect 21988 31524 22044 31580
rect 22044 31524 22048 31580
rect 21984 31520 22048 31524
rect 1532 31240 1596 31244
rect 1532 31184 1546 31240
rect 1546 31184 1596 31240
rect 1532 31180 1596 31184
rect 5580 31316 5644 31380
rect 8524 31316 8588 31380
rect 7788 31180 7852 31244
rect 5764 31044 5828 31108
rect 15148 31044 15212 31108
rect 3551 31036 3615 31040
rect 3551 30980 3555 31036
rect 3555 30980 3611 31036
rect 3611 30980 3615 31036
rect 3551 30976 3615 30980
rect 3631 31036 3695 31040
rect 3631 30980 3635 31036
rect 3635 30980 3691 31036
rect 3691 30980 3695 31036
rect 3631 30976 3695 30980
rect 3711 31036 3775 31040
rect 3711 30980 3715 31036
rect 3715 30980 3771 31036
rect 3771 30980 3775 31036
rect 3711 30976 3775 30980
rect 3791 31036 3855 31040
rect 3791 30980 3795 31036
rect 3795 30980 3851 31036
rect 3851 30980 3855 31036
rect 3791 30976 3855 30980
rect 8749 31036 8813 31040
rect 8749 30980 8753 31036
rect 8753 30980 8809 31036
rect 8809 30980 8813 31036
rect 8749 30976 8813 30980
rect 8829 31036 8893 31040
rect 8829 30980 8833 31036
rect 8833 30980 8889 31036
rect 8889 30980 8893 31036
rect 8829 30976 8893 30980
rect 8909 31036 8973 31040
rect 8909 30980 8913 31036
rect 8913 30980 8969 31036
rect 8969 30980 8973 31036
rect 8909 30976 8973 30980
rect 8989 31036 9053 31040
rect 8989 30980 8993 31036
rect 8993 30980 9049 31036
rect 9049 30980 9053 31036
rect 8989 30976 9053 30980
rect 13947 31036 14011 31040
rect 13947 30980 13951 31036
rect 13951 30980 14007 31036
rect 14007 30980 14011 31036
rect 13947 30976 14011 30980
rect 14027 31036 14091 31040
rect 14027 30980 14031 31036
rect 14031 30980 14087 31036
rect 14087 30980 14091 31036
rect 14027 30976 14091 30980
rect 14107 31036 14171 31040
rect 14107 30980 14111 31036
rect 14111 30980 14167 31036
rect 14167 30980 14171 31036
rect 14107 30976 14171 30980
rect 14187 31036 14251 31040
rect 14187 30980 14191 31036
rect 14191 30980 14247 31036
rect 14247 30980 14251 31036
rect 14187 30976 14251 30980
rect 19145 31036 19209 31040
rect 19145 30980 19149 31036
rect 19149 30980 19205 31036
rect 19205 30980 19209 31036
rect 19145 30976 19209 30980
rect 19225 31036 19289 31040
rect 19225 30980 19229 31036
rect 19229 30980 19285 31036
rect 19285 30980 19289 31036
rect 19225 30976 19289 30980
rect 19305 31036 19369 31040
rect 19305 30980 19309 31036
rect 19309 30980 19365 31036
rect 19365 30980 19369 31036
rect 19305 30976 19369 30980
rect 19385 31036 19449 31040
rect 19385 30980 19389 31036
rect 19389 30980 19445 31036
rect 19445 30980 19449 31036
rect 19385 30976 19449 30980
rect 9628 30772 9692 30836
rect 14780 30908 14844 30972
rect 2084 30636 2148 30700
rect 5948 30560 6012 30564
rect 5948 30504 5962 30560
rect 5962 30504 6012 30560
rect 5948 30500 6012 30504
rect 7236 30500 7300 30564
rect 12204 30560 12268 30564
rect 12204 30504 12254 30560
rect 12254 30504 12268 30560
rect 12204 30500 12268 30504
rect 13308 30636 13372 30700
rect 6150 30492 6214 30496
rect 6150 30436 6154 30492
rect 6154 30436 6210 30492
rect 6210 30436 6214 30492
rect 6150 30432 6214 30436
rect 6230 30492 6294 30496
rect 6230 30436 6234 30492
rect 6234 30436 6290 30492
rect 6290 30436 6294 30492
rect 6230 30432 6294 30436
rect 6310 30492 6374 30496
rect 6310 30436 6314 30492
rect 6314 30436 6370 30492
rect 6370 30436 6374 30492
rect 6310 30432 6374 30436
rect 6390 30492 6454 30496
rect 6390 30436 6394 30492
rect 6394 30436 6450 30492
rect 6450 30436 6454 30492
rect 6390 30432 6454 30436
rect 11348 30492 11412 30496
rect 11348 30436 11352 30492
rect 11352 30436 11408 30492
rect 11408 30436 11412 30492
rect 11348 30432 11412 30436
rect 11428 30492 11492 30496
rect 11428 30436 11432 30492
rect 11432 30436 11488 30492
rect 11488 30436 11492 30492
rect 11428 30432 11492 30436
rect 11508 30492 11572 30496
rect 11508 30436 11512 30492
rect 11512 30436 11568 30492
rect 11568 30436 11572 30492
rect 11508 30432 11572 30436
rect 11588 30492 11652 30496
rect 11588 30436 11592 30492
rect 11592 30436 11648 30492
rect 11648 30436 11652 30492
rect 11588 30432 11652 30436
rect 16546 30492 16610 30496
rect 16546 30436 16550 30492
rect 16550 30436 16606 30492
rect 16606 30436 16610 30492
rect 16546 30432 16610 30436
rect 16626 30492 16690 30496
rect 16626 30436 16630 30492
rect 16630 30436 16686 30492
rect 16686 30436 16690 30492
rect 16626 30432 16690 30436
rect 16706 30492 16770 30496
rect 16706 30436 16710 30492
rect 16710 30436 16766 30492
rect 16766 30436 16770 30492
rect 16706 30432 16770 30436
rect 16786 30492 16850 30496
rect 16786 30436 16790 30492
rect 16790 30436 16846 30492
rect 16846 30436 16850 30492
rect 16786 30432 16850 30436
rect 21744 30492 21808 30496
rect 21744 30436 21748 30492
rect 21748 30436 21804 30492
rect 21804 30436 21808 30492
rect 21744 30432 21808 30436
rect 21824 30492 21888 30496
rect 21824 30436 21828 30492
rect 21828 30436 21884 30492
rect 21884 30436 21888 30492
rect 21824 30432 21888 30436
rect 21904 30492 21968 30496
rect 21904 30436 21908 30492
rect 21908 30436 21964 30492
rect 21964 30436 21968 30492
rect 21904 30432 21968 30436
rect 21984 30492 22048 30496
rect 21984 30436 21988 30492
rect 21988 30436 22044 30492
rect 22044 30436 22048 30492
rect 21984 30432 22048 30436
rect 9812 30364 9876 30428
rect 20852 30364 20916 30428
rect 3188 30228 3252 30292
rect 5212 30152 5276 30156
rect 5212 30096 5226 30152
rect 5226 30096 5276 30152
rect 3551 29948 3615 29952
rect 3551 29892 3555 29948
rect 3555 29892 3611 29948
rect 3611 29892 3615 29948
rect 3551 29888 3615 29892
rect 3631 29948 3695 29952
rect 3631 29892 3635 29948
rect 3635 29892 3691 29948
rect 3691 29892 3695 29948
rect 3631 29888 3695 29892
rect 3711 29948 3775 29952
rect 3711 29892 3715 29948
rect 3715 29892 3771 29948
rect 3771 29892 3775 29948
rect 3711 29888 3775 29892
rect 3791 29948 3855 29952
rect 3791 29892 3795 29948
rect 3795 29892 3851 29948
rect 3851 29892 3855 29948
rect 3791 29888 3855 29892
rect 5212 30092 5276 30096
rect 10916 30092 10980 30156
rect 20668 30092 20732 30156
rect 15884 30016 15948 30020
rect 15884 29960 15934 30016
rect 15934 29960 15948 30016
rect 15884 29956 15948 29960
rect 8749 29948 8813 29952
rect 8749 29892 8753 29948
rect 8753 29892 8809 29948
rect 8809 29892 8813 29948
rect 8749 29888 8813 29892
rect 8829 29948 8893 29952
rect 8829 29892 8833 29948
rect 8833 29892 8889 29948
rect 8889 29892 8893 29948
rect 8829 29888 8893 29892
rect 8909 29948 8973 29952
rect 8909 29892 8913 29948
rect 8913 29892 8969 29948
rect 8969 29892 8973 29948
rect 8909 29888 8973 29892
rect 8989 29948 9053 29952
rect 8989 29892 8993 29948
rect 8993 29892 9049 29948
rect 9049 29892 9053 29948
rect 8989 29888 9053 29892
rect 13947 29948 14011 29952
rect 13947 29892 13951 29948
rect 13951 29892 14007 29948
rect 14007 29892 14011 29948
rect 13947 29888 14011 29892
rect 14027 29948 14091 29952
rect 14027 29892 14031 29948
rect 14031 29892 14087 29948
rect 14087 29892 14091 29948
rect 14027 29888 14091 29892
rect 14107 29948 14171 29952
rect 14107 29892 14111 29948
rect 14111 29892 14167 29948
rect 14167 29892 14171 29948
rect 14107 29888 14171 29892
rect 14187 29948 14251 29952
rect 14187 29892 14191 29948
rect 14191 29892 14247 29948
rect 14247 29892 14251 29948
rect 14187 29888 14251 29892
rect 19145 29948 19209 29952
rect 19145 29892 19149 29948
rect 19149 29892 19205 29948
rect 19205 29892 19209 29948
rect 19145 29888 19209 29892
rect 19225 29948 19289 29952
rect 19225 29892 19229 29948
rect 19229 29892 19285 29948
rect 19285 29892 19289 29948
rect 19225 29888 19289 29892
rect 19305 29948 19369 29952
rect 19305 29892 19309 29948
rect 19309 29892 19365 29948
rect 19365 29892 19369 29948
rect 19305 29888 19369 29892
rect 19385 29948 19449 29952
rect 19385 29892 19389 29948
rect 19389 29892 19445 29948
rect 19445 29892 19449 29948
rect 19385 29888 19449 29892
rect 4108 29820 4172 29884
rect 3372 29684 3436 29748
rect 9444 29412 9508 29476
rect 6150 29404 6214 29408
rect 6150 29348 6154 29404
rect 6154 29348 6210 29404
rect 6210 29348 6214 29404
rect 6150 29344 6214 29348
rect 6230 29404 6294 29408
rect 6230 29348 6234 29404
rect 6234 29348 6290 29404
rect 6290 29348 6294 29404
rect 6230 29344 6294 29348
rect 6310 29404 6374 29408
rect 6310 29348 6314 29404
rect 6314 29348 6370 29404
rect 6370 29348 6374 29404
rect 6310 29344 6374 29348
rect 6390 29404 6454 29408
rect 6390 29348 6394 29404
rect 6394 29348 6450 29404
rect 6450 29348 6454 29404
rect 6390 29344 6454 29348
rect 5028 29276 5092 29340
rect 3004 29200 3068 29204
rect 11348 29404 11412 29408
rect 11348 29348 11352 29404
rect 11352 29348 11408 29404
rect 11408 29348 11412 29404
rect 11348 29344 11412 29348
rect 11428 29404 11492 29408
rect 11428 29348 11432 29404
rect 11432 29348 11488 29404
rect 11488 29348 11492 29404
rect 11428 29344 11492 29348
rect 11508 29404 11572 29408
rect 11508 29348 11512 29404
rect 11512 29348 11568 29404
rect 11568 29348 11572 29404
rect 11508 29344 11572 29348
rect 11588 29404 11652 29408
rect 11588 29348 11592 29404
rect 11592 29348 11648 29404
rect 11648 29348 11652 29404
rect 11588 29344 11652 29348
rect 11100 29276 11164 29340
rect 3004 29144 3054 29200
rect 3054 29144 3068 29200
rect 3004 29140 3068 29144
rect 4844 29004 4908 29068
rect 10548 29004 10612 29068
rect 16546 29404 16610 29408
rect 16546 29348 16550 29404
rect 16550 29348 16606 29404
rect 16606 29348 16610 29404
rect 16546 29344 16610 29348
rect 16626 29404 16690 29408
rect 16626 29348 16630 29404
rect 16630 29348 16686 29404
rect 16686 29348 16690 29404
rect 16626 29344 16690 29348
rect 16706 29404 16770 29408
rect 16706 29348 16710 29404
rect 16710 29348 16766 29404
rect 16766 29348 16770 29404
rect 16706 29344 16770 29348
rect 16786 29404 16850 29408
rect 16786 29348 16790 29404
rect 16790 29348 16846 29404
rect 16846 29348 16850 29404
rect 16786 29344 16850 29348
rect 21744 29404 21808 29408
rect 21744 29348 21748 29404
rect 21748 29348 21804 29404
rect 21804 29348 21808 29404
rect 21744 29344 21808 29348
rect 21824 29404 21888 29408
rect 21824 29348 21828 29404
rect 21828 29348 21884 29404
rect 21884 29348 21888 29404
rect 21824 29344 21888 29348
rect 21904 29404 21968 29408
rect 21904 29348 21908 29404
rect 21908 29348 21964 29404
rect 21964 29348 21968 29404
rect 21904 29344 21968 29348
rect 21984 29404 22048 29408
rect 21984 29348 21988 29404
rect 21988 29348 22044 29404
rect 22044 29348 22048 29404
rect 21984 29344 22048 29348
rect 3551 28860 3615 28864
rect 3551 28804 3555 28860
rect 3555 28804 3611 28860
rect 3611 28804 3615 28860
rect 3551 28800 3615 28804
rect 3631 28860 3695 28864
rect 3631 28804 3635 28860
rect 3635 28804 3691 28860
rect 3691 28804 3695 28860
rect 3631 28800 3695 28804
rect 3711 28860 3775 28864
rect 3711 28804 3715 28860
rect 3715 28804 3771 28860
rect 3771 28804 3775 28860
rect 3711 28800 3775 28804
rect 3791 28860 3855 28864
rect 3791 28804 3795 28860
rect 3795 28804 3851 28860
rect 3851 28804 3855 28860
rect 3791 28800 3855 28804
rect 8749 28860 8813 28864
rect 8749 28804 8753 28860
rect 8753 28804 8809 28860
rect 8809 28804 8813 28860
rect 8749 28800 8813 28804
rect 8829 28860 8893 28864
rect 8829 28804 8833 28860
rect 8833 28804 8889 28860
rect 8889 28804 8893 28860
rect 8829 28800 8893 28804
rect 8909 28860 8973 28864
rect 8909 28804 8913 28860
rect 8913 28804 8969 28860
rect 8969 28804 8973 28860
rect 8909 28800 8973 28804
rect 8989 28860 9053 28864
rect 8989 28804 8993 28860
rect 8993 28804 9049 28860
rect 9049 28804 9053 28860
rect 8989 28800 9053 28804
rect 5948 28732 6012 28796
rect 8524 28732 8588 28796
rect 16068 29004 16132 29068
rect 17172 29004 17236 29068
rect 17356 28868 17420 28932
rect 18828 29004 18892 29068
rect 13947 28860 14011 28864
rect 13947 28804 13951 28860
rect 13951 28804 14007 28860
rect 14007 28804 14011 28860
rect 13947 28800 14011 28804
rect 14027 28860 14091 28864
rect 14027 28804 14031 28860
rect 14031 28804 14087 28860
rect 14087 28804 14091 28860
rect 14027 28800 14091 28804
rect 14107 28860 14171 28864
rect 14107 28804 14111 28860
rect 14111 28804 14167 28860
rect 14167 28804 14171 28860
rect 14107 28800 14171 28804
rect 14187 28860 14251 28864
rect 14187 28804 14191 28860
rect 14191 28804 14247 28860
rect 14247 28804 14251 28860
rect 14187 28800 14251 28804
rect 19145 28860 19209 28864
rect 19145 28804 19149 28860
rect 19149 28804 19205 28860
rect 19205 28804 19209 28860
rect 19145 28800 19209 28804
rect 19225 28860 19289 28864
rect 19225 28804 19229 28860
rect 19229 28804 19285 28860
rect 19285 28804 19289 28860
rect 19225 28800 19289 28804
rect 19305 28860 19369 28864
rect 19305 28804 19309 28860
rect 19309 28804 19365 28860
rect 19365 28804 19369 28860
rect 19305 28800 19369 28804
rect 19385 28860 19449 28864
rect 19385 28804 19389 28860
rect 19389 28804 19445 28860
rect 19445 28804 19449 28860
rect 19385 28800 19449 28804
rect 13492 28732 13556 28796
rect 4292 28596 4356 28660
rect 6684 28596 6748 28660
rect 10180 28596 10244 28660
rect 14596 28596 14660 28660
rect 2268 28460 2332 28524
rect 13124 28460 13188 28524
rect 2636 28324 2700 28388
rect 5948 28324 6012 28388
rect 8156 28324 8220 28388
rect 6150 28316 6214 28320
rect 6150 28260 6154 28316
rect 6154 28260 6210 28316
rect 6210 28260 6214 28316
rect 6150 28256 6214 28260
rect 6230 28316 6294 28320
rect 6230 28260 6234 28316
rect 6234 28260 6290 28316
rect 6290 28260 6294 28316
rect 6230 28256 6294 28260
rect 6310 28316 6374 28320
rect 6310 28260 6314 28316
rect 6314 28260 6370 28316
rect 6370 28260 6374 28316
rect 6310 28256 6374 28260
rect 6390 28316 6454 28320
rect 6390 28260 6394 28316
rect 6394 28260 6450 28316
rect 6450 28260 6454 28316
rect 6390 28256 6454 28260
rect 11348 28316 11412 28320
rect 11348 28260 11352 28316
rect 11352 28260 11408 28316
rect 11408 28260 11412 28316
rect 11348 28256 11412 28260
rect 11428 28316 11492 28320
rect 11428 28260 11432 28316
rect 11432 28260 11488 28316
rect 11488 28260 11492 28316
rect 11428 28256 11492 28260
rect 11508 28316 11572 28320
rect 11508 28260 11512 28316
rect 11512 28260 11568 28316
rect 11568 28260 11572 28316
rect 11508 28256 11572 28260
rect 11588 28316 11652 28320
rect 11588 28260 11592 28316
rect 11592 28260 11648 28316
rect 11648 28260 11652 28316
rect 11588 28256 11652 28260
rect 16546 28316 16610 28320
rect 16546 28260 16550 28316
rect 16550 28260 16606 28316
rect 16606 28260 16610 28316
rect 16546 28256 16610 28260
rect 16626 28316 16690 28320
rect 16626 28260 16630 28316
rect 16630 28260 16686 28316
rect 16686 28260 16690 28316
rect 16626 28256 16690 28260
rect 16706 28316 16770 28320
rect 16706 28260 16710 28316
rect 16710 28260 16766 28316
rect 16766 28260 16770 28316
rect 16706 28256 16770 28260
rect 16786 28316 16850 28320
rect 16786 28260 16790 28316
rect 16790 28260 16846 28316
rect 16846 28260 16850 28316
rect 16786 28256 16850 28260
rect 21744 28316 21808 28320
rect 21744 28260 21748 28316
rect 21748 28260 21804 28316
rect 21804 28260 21808 28316
rect 21744 28256 21808 28260
rect 21824 28316 21888 28320
rect 21824 28260 21828 28316
rect 21828 28260 21884 28316
rect 21884 28260 21888 28316
rect 21824 28256 21888 28260
rect 21904 28316 21968 28320
rect 21904 28260 21908 28316
rect 21908 28260 21964 28316
rect 21964 28260 21968 28316
rect 21904 28256 21968 28260
rect 21984 28316 22048 28320
rect 21984 28260 21988 28316
rect 21988 28260 22044 28316
rect 22044 28260 22048 28316
rect 21984 28256 22048 28260
rect 14964 27916 15028 27980
rect 17540 27780 17604 27844
rect 3551 27772 3615 27776
rect 3551 27716 3555 27772
rect 3555 27716 3611 27772
rect 3611 27716 3615 27772
rect 3551 27712 3615 27716
rect 3631 27772 3695 27776
rect 3631 27716 3635 27772
rect 3635 27716 3691 27772
rect 3691 27716 3695 27772
rect 3631 27712 3695 27716
rect 3711 27772 3775 27776
rect 3711 27716 3715 27772
rect 3715 27716 3771 27772
rect 3771 27716 3775 27772
rect 3711 27712 3775 27716
rect 3791 27772 3855 27776
rect 3791 27716 3795 27772
rect 3795 27716 3851 27772
rect 3851 27716 3855 27772
rect 3791 27712 3855 27716
rect 8749 27772 8813 27776
rect 8749 27716 8753 27772
rect 8753 27716 8809 27772
rect 8809 27716 8813 27772
rect 8749 27712 8813 27716
rect 8829 27772 8893 27776
rect 8829 27716 8833 27772
rect 8833 27716 8889 27772
rect 8889 27716 8893 27772
rect 8829 27712 8893 27716
rect 8909 27772 8973 27776
rect 8909 27716 8913 27772
rect 8913 27716 8969 27772
rect 8969 27716 8973 27772
rect 8909 27712 8973 27716
rect 8989 27772 9053 27776
rect 8989 27716 8993 27772
rect 8993 27716 9049 27772
rect 9049 27716 9053 27772
rect 8989 27712 9053 27716
rect 13947 27772 14011 27776
rect 13947 27716 13951 27772
rect 13951 27716 14007 27772
rect 14007 27716 14011 27772
rect 13947 27712 14011 27716
rect 14027 27772 14091 27776
rect 14027 27716 14031 27772
rect 14031 27716 14087 27772
rect 14087 27716 14091 27772
rect 14027 27712 14091 27716
rect 14107 27772 14171 27776
rect 14107 27716 14111 27772
rect 14111 27716 14167 27772
rect 14167 27716 14171 27772
rect 14107 27712 14171 27716
rect 14187 27772 14251 27776
rect 14187 27716 14191 27772
rect 14191 27716 14247 27772
rect 14247 27716 14251 27772
rect 14187 27712 14251 27716
rect 19145 27772 19209 27776
rect 19145 27716 19149 27772
rect 19149 27716 19205 27772
rect 19205 27716 19209 27772
rect 19145 27712 19209 27716
rect 19225 27772 19289 27776
rect 19225 27716 19229 27772
rect 19229 27716 19285 27772
rect 19285 27716 19289 27772
rect 19225 27712 19289 27716
rect 19305 27772 19369 27776
rect 19305 27716 19309 27772
rect 19309 27716 19365 27772
rect 19365 27716 19369 27772
rect 19305 27712 19369 27716
rect 19385 27772 19449 27776
rect 19385 27716 19389 27772
rect 19389 27716 19445 27772
rect 19445 27716 19449 27772
rect 19385 27712 19449 27716
rect 5028 27704 5092 27708
rect 5028 27648 5078 27704
rect 5078 27648 5092 27704
rect 5028 27644 5092 27648
rect 7236 27704 7300 27708
rect 7236 27648 7286 27704
rect 7286 27648 7300 27704
rect 7236 27644 7300 27648
rect 7788 27644 7852 27708
rect 16068 27644 16132 27708
rect 2820 27372 2884 27436
rect 3924 27372 3988 27436
rect 1900 27236 1964 27300
rect 2084 27100 2148 27164
rect 3188 27296 3252 27300
rect 3188 27240 3202 27296
rect 3202 27240 3252 27296
rect 3188 27236 3252 27240
rect 6150 27228 6214 27232
rect 6150 27172 6154 27228
rect 6154 27172 6210 27228
rect 6210 27172 6214 27228
rect 6150 27168 6214 27172
rect 6230 27228 6294 27232
rect 6230 27172 6234 27228
rect 6234 27172 6290 27228
rect 6290 27172 6294 27228
rect 6230 27168 6294 27172
rect 6310 27228 6374 27232
rect 6310 27172 6314 27228
rect 6314 27172 6370 27228
rect 6370 27172 6374 27228
rect 6310 27168 6374 27172
rect 6390 27228 6454 27232
rect 6390 27172 6394 27228
rect 6394 27172 6450 27228
rect 6450 27172 6454 27228
rect 6390 27168 6454 27172
rect 11348 27228 11412 27232
rect 11348 27172 11352 27228
rect 11352 27172 11408 27228
rect 11408 27172 11412 27228
rect 11348 27168 11412 27172
rect 11428 27228 11492 27232
rect 11428 27172 11432 27228
rect 11432 27172 11488 27228
rect 11488 27172 11492 27228
rect 11428 27168 11492 27172
rect 11508 27228 11572 27232
rect 11508 27172 11512 27228
rect 11512 27172 11568 27228
rect 11568 27172 11572 27228
rect 11508 27168 11572 27172
rect 11588 27228 11652 27232
rect 11588 27172 11592 27228
rect 11592 27172 11648 27228
rect 11648 27172 11652 27228
rect 11588 27168 11652 27172
rect 16546 27228 16610 27232
rect 16546 27172 16550 27228
rect 16550 27172 16606 27228
rect 16606 27172 16610 27228
rect 16546 27168 16610 27172
rect 16626 27228 16690 27232
rect 16626 27172 16630 27228
rect 16630 27172 16686 27228
rect 16686 27172 16690 27228
rect 16626 27168 16690 27172
rect 16706 27228 16770 27232
rect 16706 27172 16710 27228
rect 16710 27172 16766 27228
rect 16766 27172 16770 27228
rect 16706 27168 16770 27172
rect 16786 27228 16850 27232
rect 16786 27172 16790 27228
rect 16790 27172 16846 27228
rect 16846 27172 16850 27228
rect 16786 27168 16850 27172
rect 21744 27228 21808 27232
rect 21744 27172 21748 27228
rect 21748 27172 21804 27228
rect 21804 27172 21808 27228
rect 21744 27168 21808 27172
rect 21824 27228 21888 27232
rect 21824 27172 21828 27228
rect 21828 27172 21884 27228
rect 21884 27172 21888 27228
rect 21824 27168 21888 27172
rect 21904 27228 21968 27232
rect 21904 27172 21908 27228
rect 21908 27172 21964 27228
rect 21964 27172 21968 27228
rect 21904 27168 21968 27172
rect 21984 27228 22048 27232
rect 21984 27172 21988 27228
rect 21988 27172 22044 27228
rect 22044 27172 22048 27228
rect 21984 27168 22048 27172
rect 3924 27100 3988 27164
rect 4476 27100 4540 27164
rect 8524 27160 8588 27164
rect 8524 27104 8574 27160
rect 8574 27104 8588 27160
rect 8524 27100 8588 27104
rect 9444 27100 9508 27164
rect 10548 27100 10612 27164
rect 8524 26964 8588 27028
rect 1532 26828 1596 26892
rect 3372 26692 3436 26756
rect 6684 26692 6748 26756
rect 12388 26692 12452 26756
rect 3551 26684 3615 26688
rect 3551 26628 3555 26684
rect 3555 26628 3611 26684
rect 3611 26628 3615 26684
rect 3551 26624 3615 26628
rect 3631 26684 3695 26688
rect 3631 26628 3635 26684
rect 3635 26628 3691 26684
rect 3691 26628 3695 26684
rect 3631 26624 3695 26628
rect 3711 26684 3775 26688
rect 3711 26628 3715 26684
rect 3715 26628 3771 26684
rect 3771 26628 3775 26684
rect 3711 26624 3775 26628
rect 3791 26684 3855 26688
rect 3791 26628 3795 26684
rect 3795 26628 3851 26684
rect 3851 26628 3855 26684
rect 3791 26624 3855 26628
rect 8749 26684 8813 26688
rect 8749 26628 8753 26684
rect 8753 26628 8809 26684
rect 8809 26628 8813 26684
rect 8749 26624 8813 26628
rect 8829 26684 8893 26688
rect 8829 26628 8833 26684
rect 8833 26628 8889 26684
rect 8889 26628 8893 26684
rect 8829 26624 8893 26628
rect 8909 26684 8973 26688
rect 8909 26628 8913 26684
rect 8913 26628 8969 26684
rect 8969 26628 8973 26684
rect 8909 26624 8973 26628
rect 8989 26684 9053 26688
rect 8989 26628 8993 26684
rect 8993 26628 9049 26684
rect 9049 26628 9053 26684
rect 8989 26624 9053 26628
rect 13947 26684 14011 26688
rect 13947 26628 13951 26684
rect 13951 26628 14007 26684
rect 14007 26628 14011 26684
rect 13947 26624 14011 26628
rect 14027 26684 14091 26688
rect 14027 26628 14031 26684
rect 14031 26628 14087 26684
rect 14087 26628 14091 26684
rect 14027 26624 14091 26628
rect 14107 26684 14171 26688
rect 14107 26628 14111 26684
rect 14111 26628 14167 26684
rect 14167 26628 14171 26684
rect 14107 26624 14171 26628
rect 14187 26684 14251 26688
rect 14187 26628 14191 26684
rect 14191 26628 14247 26684
rect 14247 26628 14251 26684
rect 14187 26624 14251 26628
rect 19145 26684 19209 26688
rect 19145 26628 19149 26684
rect 19149 26628 19205 26684
rect 19205 26628 19209 26684
rect 19145 26624 19209 26628
rect 19225 26684 19289 26688
rect 19225 26628 19229 26684
rect 19229 26628 19285 26684
rect 19285 26628 19289 26684
rect 19225 26624 19289 26628
rect 19305 26684 19369 26688
rect 19305 26628 19309 26684
rect 19309 26628 19365 26684
rect 19365 26628 19369 26684
rect 19305 26624 19369 26628
rect 19385 26684 19449 26688
rect 19385 26628 19389 26684
rect 19389 26628 19445 26684
rect 19445 26628 19449 26684
rect 19385 26624 19449 26628
rect 2452 26480 2516 26484
rect 2452 26424 2502 26480
rect 2502 26424 2516 26480
rect 2452 26420 2516 26424
rect 10180 26284 10244 26348
rect 1348 26148 1412 26212
rect 1716 26012 1780 26076
rect 5396 26148 5460 26212
rect 18092 26148 18156 26212
rect 6150 26140 6214 26144
rect 6150 26084 6154 26140
rect 6154 26084 6210 26140
rect 6210 26084 6214 26140
rect 6150 26080 6214 26084
rect 6230 26140 6294 26144
rect 6230 26084 6234 26140
rect 6234 26084 6290 26140
rect 6290 26084 6294 26140
rect 6230 26080 6294 26084
rect 6310 26140 6374 26144
rect 6310 26084 6314 26140
rect 6314 26084 6370 26140
rect 6370 26084 6374 26140
rect 6310 26080 6374 26084
rect 6390 26140 6454 26144
rect 6390 26084 6394 26140
rect 6394 26084 6450 26140
rect 6450 26084 6454 26140
rect 6390 26080 6454 26084
rect 11348 26140 11412 26144
rect 11348 26084 11352 26140
rect 11352 26084 11408 26140
rect 11408 26084 11412 26140
rect 11348 26080 11412 26084
rect 11428 26140 11492 26144
rect 11428 26084 11432 26140
rect 11432 26084 11488 26140
rect 11488 26084 11492 26140
rect 11428 26080 11492 26084
rect 11508 26140 11572 26144
rect 11508 26084 11512 26140
rect 11512 26084 11568 26140
rect 11568 26084 11572 26140
rect 11508 26080 11572 26084
rect 11588 26140 11652 26144
rect 11588 26084 11592 26140
rect 11592 26084 11648 26140
rect 11648 26084 11652 26140
rect 11588 26080 11652 26084
rect 16546 26140 16610 26144
rect 16546 26084 16550 26140
rect 16550 26084 16606 26140
rect 16606 26084 16610 26140
rect 16546 26080 16610 26084
rect 16626 26140 16690 26144
rect 16626 26084 16630 26140
rect 16630 26084 16686 26140
rect 16686 26084 16690 26140
rect 16626 26080 16690 26084
rect 16706 26140 16770 26144
rect 16706 26084 16710 26140
rect 16710 26084 16766 26140
rect 16766 26084 16770 26140
rect 16706 26080 16770 26084
rect 16786 26140 16850 26144
rect 16786 26084 16790 26140
rect 16790 26084 16846 26140
rect 16846 26084 16850 26140
rect 16786 26080 16850 26084
rect 21744 26140 21808 26144
rect 21744 26084 21748 26140
rect 21748 26084 21804 26140
rect 21804 26084 21808 26140
rect 21744 26080 21808 26084
rect 21824 26140 21888 26144
rect 21824 26084 21828 26140
rect 21828 26084 21884 26140
rect 21884 26084 21888 26140
rect 21824 26080 21888 26084
rect 21904 26140 21968 26144
rect 21904 26084 21908 26140
rect 21908 26084 21964 26140
rect 21964 26084 21968 26140
rect 21904 26080 21968 26084
rect 21984 26140 22048 26144
rect 21984 26084 21988 26140
rect 21988 26084 22044 26140
rect 22044 26084 22048 26140
rect 21984 26080 22048 26084
rect 1716 25740 1780 25804
rect 7788 25876 7852 25940
rect 4476 25664 4540 25668
rect 4476 25608 4526 25664
rect 4526 25608 4540 25664
rect 4476 25604 4540 25608
rect 5764 25604 5828 25668
rect 7052 25604 7116 25668
rect 3551 25596 3615 25600
rect 3551 25540 3555 25596
rect 3555 25540 3611 25596
rect 3611 25540 3615 25596
rect 3551 25536 3615 25540
rect 3631 25596 3695 25600
rect 3631 25540 3635 25596
rect 3635 25540 3691 25596
rect 3691 25540 3695 25596
rect 3631 25536 3695 25540
rect 3711 25596 3775 25600
rect 3711 25540 3715 25596
rect 3715 25540 3771 25596
rect 3771 25540 3775 25596
rect 3711 25536 3775 25540
rect 3791 25596 3855 25600
rect 3791 25540 3795 25596
rect 3795 25540 3851 25596
rect 3851 25540 3855 25596
rect 3791 25536 3855 25540
rect 8749 25596 8813 25600
rect 8749 25540 8753 25596
rect 8753 25540 8809 25596
rect 8809 25540 8813 25596
rect 8749 25536 8813 25540
rect 8829 25596 8893 25600
rect 8829 25540 8833 25596
rect 8833 25540 8889 25596
rect 8889 25540 8893 25596
rect 8829 25536 8893 25540
rect 8909 25596 8973 25600
rect 8909 25540 8913 25596
rect 8913 25540 8969 25596
rect 8969 25540 8973 25596
rect 8909 25536 8973 25540
rect 8989 25596 9053 25600
rect 8989 25540 8993 25596
rect 8993 25540 9049 25596
rect 9049 25540 9053 25596
rect 8989 25536 9053 25540
rect 13947 25596 14011 25600
rect 13947 25540 13951 25596
rect 13951 25540 14007 25596
rect 14007 25540 14011 25596
rect 13947 25536 14011 25540
rect 14027 25596 14091 25600
rect 14027 25540 14031 25596
rect 14031 25540 14087 25596
rect 14087 25540 14091 25596
rect 14027 25536 14091 25540
rect 14107 25596 14171 25600
rect 14107 25540 14111 25596
rect 14111 25540 14167 25596
rect 14167 25540 14171 25596
rect 14107 25536 14171 25540
rect 14187 25596 14251 25600
rect 14187 25540 14191 25596
rect 14191 25540 14247 25596
rect 14247 25540 14251 25596
rect 14187 25536 14251 25540
rect 19145 25596 19209 25600
rect 19145 25540 19149 25596
rect 19149 25540 19205 25596
rect 19205 25540 19209 25596
rect 19145 25536 19209 25540
rect 19225 25596 19289 25600
rect 19225 25540 19229 25596
rect 19229 25540 19285 25596
rect 19285 25540 19289 25596
rect 19225 25536 19289 25540
rect 19305 25596 19369 25600
rect 19305 25540 19309 25596
rect 19309 25540 19365 25596
rect 19365 25540 19369 25596
rect 19305 25536 19369 25540
rect 19385 25596 19449 25600
rect 19385 25540 19389 25596
rect 19389 25540 19445 25596
rect 19445 25540 19449 25596
rect 19385 25536 19449 25540
rect 6868 25468 6932 25532
rect 3004 25332 3068 25396
rect 18276 25332 18340 25396
rect 3188 25196 3252 25260
rect 13308 25196 13372 25260
rect 6150 25052 6214 25056
rect 6150 24996 6154 25052
rect 6154 24996 6210 25052
rect 6210 24996 6214 25052
rect 6150 24992 6214 24996
rect 6230 25052 6294 25056
rect 6230 24996 6234 25052
rect 6234 24996 6290 25052
rect 6290 24996 6294 25052
rect 6230 24992 6294 24996
rect 6310 25052 6374 25056
rect 6310 24996 6314 25052
rect 6314 24996 6370 25052
rect 6370 24996 6374 25052
rect 6310 24992 6374 24996
rect 6390 25052 6454 25056
rect 6390 24996 6394 25052
rect 6394 24996 6450 25052
rect 6450 24996 6454 25052
rect 6390 24992 6454 24996
rect 11348 25052 11412 25056
rect 11348 24996 11352 25052
rect 11352 24996 11408 25052
rect 11408 24996 11412 25052
rect 11348 24992 11412 24996
rect 11428 25052 11492 25056
rect 11428 24996 11432 25052
rect 11432 24996 11488 25052
rect 11488 24996 11492 25052
rect 11428 24992 11492 24996
rect 11508 25052 11572 25056
rect 11508 24996 11512 25052
rect 11512 24996 11568 25052
rect 11568 24996 11572 25052
rect 11508 24992 11572 24996
rect 11588 25052 11652 25056
rect 11588 24996 11592 25052
rect 11592 24996 11648 25052
rect 11648 24996 11652 25052
rect 11588 24992 11652 24996
rect 16546 25052 16610 25056
rect 16546 24996 16550 25052
rect 16550 24996 16606 25052
rect 16606 24996 16610 25052
rect 16546 24992 16610 24996
rect 16626 25052 16690 25056
rect 16626 24996 16630 25052
rect 16630 24996 16686 25052
rect 16686 24996 16690 25052
rect 16626 24992 16690 24996
rect 16706 25052 16770 25056
rect 16706 24996 16710 25052
rect 16710 24996 16766 25052
rect 16766 24996 16770 25052
rect 16706 24992 16770 24996
rect 16786 25052 16850 25056
rect 16786 24996 16790 25052
rect 16790 24996 16846 25052
rect 16846 24996 16850 25052
rect 16786 24992 16850 24996
rect 21744 25052 21808 25056
rect 21744 24996 21748 25052
rect 21748 24996 21804 25052
rect 21804 24996 21808 25052
rect 21744 24992 21808 24996
rect 21824 25052 21888 25056
rect 21824 24996 21828 25052
rect 21828 24996 21884 25052
rect 21884 24996 21888 25052
rect 21824 24992 21888 24996
rect 21904 25052 21968 25056
rect 21904 24996 21908 25052
rect 21908 24996 21964 25052
rect 21964 24996 21968 25052
rect 21904 24992 21968 24996
rect 21984 25052 22048 25056
rect 21984 24996 21988 25052
rect 21988 24996 22044 25052
rect 22044 24996 22048 25052
rect 21984 24992 22048 24996
rect 15516 24924 15580 24988
rect 9812 24788 9876 24852
rect 12020 24788 12084 24852
rect 12204 24788 12268 24852
rect 18644 24788 18708 24852
rect 5212 24652 5276 24716
rect 3551 24508 3615 24512
rect 3551 24452 3555 24508
rect 3555 24452 3611 24508
rect 3611 24452 3615 24508
rect 3551 24448 3615 24452
rect 3631 24508 3695 24512
rect 3631 24452 3635 24508
rect 3635 24452 3691 24508
rect 3691 24452 3695 24508
rect 3631 24448 3695 24452
rect 3711 24508 3775 24512
rect 3711 24452 3715 24508
rect 3715 24452 3771 24508
rect 3771 24452 3775 24508
rect 3711 24448 3775 24452
rect 3791 24508 3855 24512
rect 3791 24452 3795 24508
rect 3795 24452 3851 24508
rect 3851 24452 3855 24508
rect 3791 24448 3855 24452
rect 8749 24508 8813 24512
rect 8749 24452 8753 24508
rect 8753 24452 8809 24508
rect 8809 24452 8813 24508
rect 8749 24448 8813 24452
rect 8829 24508 8893 24512
rect 8829 24452 8833 24508
rect 8833 24452 8889 24508
rect 8889 24452 8893 24508
rect 8829 24448 8893 24452
rect 8909 24508 8973 24512
rect 8909 24452 8913 24508
rect 8913 24452 8969 24508
rect 8969 24452 8973 24508
rect 8909 24448 8973 24452
rect 8989 24508 9053 24512
rect 8989 24452 8993 24508
rect 8993 24452 9049 24508
rect 9049 24452 9053 24508
rect 8989 24448 9053 24452
rect 4292 24440 4356 24444
rect 4292 24384 4306 24440
rect 4306 24384 4356 24440
rect 4292 24380 4356 24384
rect 7604 24380 7668 24444
rect 14780 24652 14844 24716
rect 14964 24712 15028 24716
rect 14964 24656 14978 24712
rect 14978 24656 15028 24712
rect 14964 24652 15028 24656
rect 16988 24652 17052 24716
rect 14964 24516 15028 24580
rect 13947 24508 14011 24512
rect 13947 24452 13951 24508
rect 13951 24452 14007 24508
rect 14007 24452 14011 24508
rect 13947 24448 14011 24452
rect 14027 24508 14091 24512
rect 14027 24452 14031 24508
rect 14031 24452 14087 24508
rect 14087 24452 14091 24508
rect 14027 24448 14091 24452
rect 14107 24508 14171 24512
rect 14107 24452 14111 24508
rect 14111 24452 14167 24508
rect 14167 24452 14171 24508
rect 14107 24448 14171 24452
rect 14187 24508 14251 24512
rect 14187 24452 14191 24508
rect 14191 24452 14247 24508
rect 14247 24452 14251 24508
rect 14187 24448 14251 24452
rect 19145 24508 19209 24512
rect 19145 24452 19149 24508
rect 19149 24452 19205 24508
rect 19205 24452 19209 24508
rect 19145 24448 19209 24452
rect 19225 24508 19289 24512
rect 19225 24452 19229 24508
rect 19229 24452 19285 24508
rect 19285 24452 19289 24508
rect 19225 24448 19289 24452
rect 19305 24508 19369 24512
rect 19305 24452 19309 24508
rect 19309 24452 19365 24508
rect 19365 24452 19369 24508
rect 19305 24448 19369 24452
rect 19385 24508 19449 24512
rect 19385 24452 19389 24508
rect 19389 24452 19445 24508
rect 19445 24452 19449 24508
rect 19385 24448 19449 24452
rect 5948 24244 6012 24308
rect 7604 24244 7668 24308
rect 4292 24168 4356 24172
rect 4292 24112 4342 24168
rect 4342 24112 4356 24168
rect 4292 24108 4356 24112
rect 5028 23972 5092 24036
rect 9628 24108 9692 24172
rect 17356 24108 17420 24172
rect 15148 23972 15212 24036
rect 6150 23964 6214 23968
rect 6150 23908 6154 23964
rect 6154 23908 6210 23964
rect 6210 23908 6214 23964
rect 6150 23904 6214 23908
rect 6230 23964 6294 23968
rect 6230 23908 6234 23964
rect 6234 23908 6290 23964
rect 6290 23908 6294 23964
rect 6230 23904 6294 23908
rect 6310 23964 6374 23968
rect 6310 23908 6314 23964
rect 6314 23908 6370 23964
rect 6370 23908 6374 23964
rect 6310 23904 6374 23908
rect 6390 23964 6454 23968
rect 6390 23908 6394 23964
rect 6394 23908 6450 23964
rect 6450 23908 6454 23964
rect 6390 23904 6454 23908
rect 11348 23964 11412 23968
rect 11348 23908 11352 23964
rect 11352 23908 11408 23964
rect 11408 23908 11412 23964
rect 11348 23904 11412 23908
rect 11428 23964 11492 23968
rect 11428 23908 11432 23964
rect 11432 23908 11488 23964
rect 11488 23908 11492 23964
rect 11428 23904 11492 23908
rect 11508 23964 11572 23968
rect 11508 23908 11512 23964
rect 11512 23908 11568 23964
rect 11568 23908 11572 23964
rect 11508 23904 11572 23908
rect 11588 23964 11652 23968
rect 11588 23908 11592 23964
rect 11592 23908 11648 23964
rect 11648 23908 11652 23964
rect 11588 23904 11652 23908
rect 16546 23964 16610 23968
rect 16546 23908 16550 23964
rect 16550 23908 16606 23964
rect 16606 23908 16610 23964
rect 16546 23904 16610 23908
rect 16626 23964 16690 23968
rect 16626 23908 16630 23964
rect 16630 23908 16686 23964
rect 16686 23908 16690 23964
rect 16626 23904 16690 23908
rect 16706 23964 16770 23968
rect 16706 23908 16710 23964
rect 16710 23908 16766 23964
rect 16766 23908 16770 23964
rect 16706 23904 16770 23908
rect 16786 23964 16850 23968
rect 16786 23908 16790 23964
rect 16790 23908 16846 23964
rect 16846 23908 16850 23964
rect 16786 23904 16850 23908
rect 21744 23964 21808 23968
rect 21744 23908 21748 23964
rect 21748 23908 21804 23964
rect 21804 23908 21808 23964
rect 21744 23904 21808 23908
rect 21824 23964 21888 23968
rect 21824 23908 21828 23964
rect 21828 23908 21884 23964
rect 21884 23908 21888 23964
rect 21824 23904 21888 23908
rect 21904 23964 21968 23968
rect 21904 23908 21908 23964
rect 21908 23908 21964 23964
rect 21964 23908 21968 23964
rect 21904 23904 21968 23908
rect 21984 23964 22048 23968
rect 21984 23908 21988 23964
rect 21988 23908 22044 23964
rect 22044 23908 22048 23964
rect 21984 23904 22048 23908
rect 7052 23836 7116 23900
rect 10548 23896 10612 23900
rect 10548 23840 10562 23896
rect 10562 23840 10612 23896
rect 10548 23836 10612 23840
rect 2820 23428 2884 23492
rect 4660 23428 4724 23492
rect 8524 23428 8588 23492
rect 11100 23564 11164 23628
rect 16252 23428 16316 23492
rect 21404 23428 21468 23492
rect 3551 23420 3615 23424
rect 3551 23364 3555 23420
rect 3555 23364 3611 23420
rect 3611 23364 3615 23420
rect 3551 23360 3615 23364
rect 3631 23420 3695 23424
rect 3631 23364 3635 23420
rect 3635 23364 3691 23420
rect 3691 23364 3695 23420
rect 3631 23360 3695 23364
rect 3711 23420 3775 23424
rect 3711 23364 3715 23420
rect 3715 23364 3771 23420
rect 3771 23364 3775 23420
rect 3711 23360 3775 23364
rect 3791 23420 3855 23424
rect 3791 23364 3795 23420
rect 3795 23364 3851 23420
rect 3851 23364 3855 23420
rect 3791 23360 3855 23364
rect 8749 23420 8813 23424
rect 8749 23364 8753 23420
rect 8753 23364 8809 23420
rect 8809 23364 8813 23420
rect 8749 23360 8813 23364
rect 8829 23420 8893 23424
rect 8829 23364 8833 23420
rect 8833 23364 8889 23420
rect 8889 23364 8893 23420
rect 8829 23360 8893 23364
rect 8909 23420 8973 23424
rect 8909 23364 8913 23420
rect 8913 23364 8969 23420
rect 8969 23364 8973 23420
rect 8909 23360 8973 23364
rect 8989 23420 9053 23424
rect 8989 23364 8993 23420
rect 8993 23364 9049 23420
rect 9049 23364 9053 23420
rect 8989 23360 9053 23364
rect 13947 23420 14011 23424
rect 13947 23364 13951 23420
rect 13951 23364 14007 23420
rect 14007 23364 14011 23420
rect 13947 23360 14011 23364
rect 14027 23420 14091 23424
rect 14027 23364 14031 23420
rect 14031 23364 14087 23420
rect 14087 23364 14091 23420
rect 14027 23360 14091 23364
rect 14107 23420 14171 23424
rect 14107 23364 14111 23420
rect 14111 23364 14167 23420
rect 14167 23364 14171 23420
rect 14107 23360 14171 23364
rect 14187 23420 14251 23424
rect 14187 23364 14191 23420
rect 14191 23364 14247 23420
rect 14247 23364 14251 23420
rect 14187 23360 14251 23364
rect 19145 23420 19209 23424
rect 19145 23364 19149 23420
rect 19149 23364 19205 23420
rect 19205 23364 19209 23420
rect 19145 23360 19209 23364
rect 19225 23420 19289 23424
rect 19225 23364 19229 23420
rect 19229 23364 19285 23420
rect 19285 23364 19289 23420
rect 19225 23360 19289 23364
rect 19305 23420 19369 23424
rect 19305 23364 19309 23420
rect 19309 23364 19365 23420
rect 19365 23364 19369 23420
rect 19305 23360 19369 23364
rect 19385 23420 19449 23424
rect 19385 23364 19389 23420
rect 19389 23364 19445 23420
rect 19445 23364 19449 23420
rect 19385 23360 19449 23364
rect 7236 23216 7300 23220
rect 7236 23160 7286 23216
rect 7286 23160 7300 23216
rect 7236 23156 7300 23160
rect 21220 23292 21284 23356
rect 13492 23156 13556 23220
rect 2636 22884 2700 22948
rect 7788 22884 7852 22948
rect 13124 22884 13188 22948
rect 6150 22876 6214 22880
rect 6150 22820 6154 22876
rect 6154 22820 6210 22876
rect 6210 22820 6214 22876
rect 6150 22816 6214 22820
rect 6230 22876 6294 22880
rect 6230 22820 6234 22876
rect 6234 22820 6290 22876
rect 6290 22820 6294 22876
rect 6230 22816 6294 22820
rect 6310 22876 6374 22880
rect 6310 22820 6314 22876
rect 6314 22820 6370 22876
rect 6370 22820 6374 22876
rect 6310 22816 6374 22820
rect 6390 22876 6454 22880
rect 6390 22820 6394 22876
rect 6394 22820 6450 22876
rect 6450 22820 6454 22876
rect 6390 22816 6454 22820
rect 11348 22876 11412 22880
rect 11348 22820 11352 22876
rect 11352 22820 11408 22876
rect 11408 22820 11412 22876
rect 11348 22816 11412 22820
rect 11428 22876 11492 22880
rect 11428 22820 11432 22876
rect 11432 22820 11488 22876
rect 11488 22820 11492 22876
rect 11428 22816 11492 22820
rect 11508 22876 11572 22880
rect 11508 22820 11512 22876
rect 11512 22820 11568 22876
rect 11568 22820 11572 22876
rect 11508 22816 11572 22820
rect 11588 22876 11652 22880
rect 11588 22820 11592 22876
rect 11592 22820 11648 22876
rect 11648 22820 11652 22876
rect 11588 22816 11652 22820
rect 16546 22876 16610 22880
rect 16546 22820 16550 22876
rect 16550 22820 16606 22876
rect 16606 22820 16610 22876
rect 16546 22816 16610 22820
rect 16626 22876 16690 22880
rect 16626 22820 16630 22876
rect 16630 22820 16686 22876
rect 16686 22820 16690 22876
rect 16626 22816 16690 22820
rect 16706 22876 16770 22880
rect 16706 22820 16710 22876
rect 16710 22820 16766 22876
rect 16766 22820 16770 22876
rect 16706 22816 16770 22820
rect 16786 22876 16850 22880
rect 16786 22820 16790 22876
rect 16790 22820 16846 22876
rect 16846 22820 16850 22876
rect 16786 22816 16850 22820
rect 21744 22876 21808 22880
rect 21744 22820 21748 22876
rect 21748 22820 21804 22876
rect 21804 22820 21808 22876
rect 21744 22816 21808 22820
rect 21824 22876 21888 22880
rect 21824 22820 21828 22876
rect 21828 22820 21884 22876
rect 21884 22820 21888 22876
rect 21824 22816 21888 22820
rect 21904 22876 21968 22880
rect 21904 22820 21908 22876
rect 21908 22820 21964 22876
rect 21964 22820 21968 22876
rect 21904 22816 21968 22820
rect 21984 22876 22048 22880
rect 21984 22820 21988 22876
rect 21988 22820 22044 22876
rect 22044 22820 22048 22876
rect 21984 22816 22048 22820
rect 13124 22808 13188 22812
rect 13124 22752 13138 22808
rect 13138 22752 13188 22808
rect 13124 22748 13188 22752
rect 11100 22612 11164 22676
rect 19564 22476 19628 22540
rect 4660 22340 4724 22404
rect 7788 22340 7852 22404
rect 10180 22340 10244 22404
rect 12940 22340 13004 22404
rect 3551 22332 3615 22336
rect 3551 22276 3555 22332
rect 3555 22276 3611 22332
rect 3611 22276 3615 22332
rect 3551 22272 3615 22276
rect 3631 22332 3695 22336
rect 3631 22276 3635 22332
rect 3635 22276 3691 22332
rect 3691 22276 3695 22332
rect 3631 22272 3695 22276
rect 3711 22332 3775 22336
rect 3711 22276 3715 22332
rect 3715 22276 3771 22332
rect 3771 22276 3775 22332
rect 3711 22272 3775 22276
rect 3791 22332 3855 22336
rect 3791 22276 3795 22332
rect 3795 22276 3851 22332
rect 3851 22276 3855 22332
rect 3791 22272 3855 22276
rect 8749 22332 8813 22336
rect 8749 22276 8753 22332
rect 8753 22276 8809 22332
rect 8809 22276 8813 22332
rect 8749 22272 8813 22276
rect 8829 22332 8893 22336
rect 8829 22276 8833 22332
rect 8833 22276 8889 22332
rect 8889 22276 8893 22332
rect 8829 22272 8893 22276
rect 8909 22332 8973 22336
rect 8909 22276 8913 22332
rect 8913 22276 8969 22332
rect 8969 22276 8973 22332
rect 8909 22272 8973 22276
rect 8989 22332 9053 22336
rect 8989 22276 8993 22332
rect 8993 22276 9049 22332
rect 9049 22276 9053 22332
rect 8989 22272 9053 22276
rect 13947 22332 14011 22336
rect 13947 22276 13951 22332
rect 13951 22276 14007 22332
rect 14007 22276 14011 22332
rect 13947 22272 14011 22276
rect 14027 22332 14091 22336
rect 14027 22276 14031 22332
rect 14031 22276 14087 22332
rect 14087 22276 14091 22332
rect 14027 22272 14091 22276
rect 14107 22332 14171 22336
rect 14107 22276 14111 22332
rect 14111 22276 14167 22332
rect 14167 22276 14171 22332
rect 14107 22272 14171 22276
rect 14187 22332 14251 22336
rect 14187 22276 14191 22332
rect 14191 22276 14247 22332
rect 14247 22276 14251 22332
rect 14187 22272 14251 22276
rect 19145 22332 19209 22336
rect 19145 22276 19149 22332
rect 19149 22276 19205 22332
rect 19205 22276 19209 22332
rect 19145 22272 19209 22276
rect 19225 22332 19289 22336
rect 19225 22276 19229 22332
rect 19229 22276 19285 22332
rect 19285 22276 19289 22332
rect 19225 22272 19289 22276
rect 19305 22332 19369 22336
rect 19305 22276 19309 22332
rect 19309 22276 19365 22332
rect 19365 22276 19369 22332
rect 19305 22272 19369 22276
rect 19385 22332 19449 22336
rect 19385 22276 19389 22332
rect 19389 22276 19445 22332
rect 19445 22276 19449 22332
rect 19385 22272 19449 22276
rect 6868 22204 6932 22268
rect 10916 22204 10980 22268
rect 14780 22264 14844 22268
rect 14780 22208 14830 22264
rect 14830 22208 14844 22264
rect 14780 22204 14844 22208
rect 11100 22068 11164 22132
rect 11836 21932 11900 21996
rect 19932 22068 19996 22132
rect 6150 21788 6214 21792
rect 6150 21732 6154 21788
rect 6154 21732 6210 21788
rect 6210 21732 6214 21788
rect 6150 21728 6214 21732
rect 6230 21788 6294 21792
rect 6230 21732 6234 21788
rect 6234 21732 6290 21788
rect 6290 21732 6294 21788
rect 6230 21728 6294 21732
rect 6310 21788 6374 21792
rect 6310 21732 6314 21788
rect 6314 21732 6370 21788
rect 6370 21732 6374 21788
rect 6310 21728 6374 21732
rect 6390 21788 6454 21792
rect 6390 21732 6394 21788
rect 6394 21732 6450 21788
rect 6450 21732 6454 21788
rect 6390 21728 6454 21732
rect 11348 21788 11412 21792
rect 11348 21732 11352 21788
rect 11352 21732 11408 21788
rect 11408 21732 11412 21788
rect 11348 21728 11412 21732
rect 11428 21788 11492 21792
rect 11428 21732 11432 21788
rect 11432 21732 11488 21788
rect 11488 21732 11492 21788
rect 11428 21728 11492 21732
rect 11508 21788 11572 21792
rect 11508 21732 11512 21788
rect 11512 21732 11568 21788
rect 11568 21732 11572 21788
rect 11508 21728 11572 21732
rect 11588 21788 11652 21792
rect 11588 21732 11592 21788
rect 11592 21732 11648 21788
rect 11648 21732 11652 21788
rect 11588 21728 11652 21732
rect 16546 21788 16610 21792
rect 16546 21732 16550 21788
rect 16550 21732 16606 21788
rect 16606 21732 16610 21788
rect 16546 21728 16610 21732
rect 16626 21788 16690 21792
rect 16626 21732 16630 21788
rect 16630 21732 16686 21788
rect 16686 21732 16690 21788
rect 16626 21728 16690 21732
rect 16706 21788 16770 21792
rect 16706 21732 16710 21788
rect 16710 21732 16766 21788
rect 16766 21732 16770 21788
rect 16706 21728 16770 21732
rect 16786 21788 16850 21792
rect 16786 21732 16790 21788
rect 16790 21732 16846 21788
rect 16846 21732 16850 21788
rect 16786 21728 16850 21732
rect 21744 21788 21808 21792
rect 21744 21732 21748 21788
rect 21748 21732 21804 21788
rect 21804 21732 21808 21788
rect 21744 21728 21808 21732
rect 21824 21788 21888 21792
rect 21824 21732 21828 21788
rect 21828 21732 21884 21788
rect 21884 21732 21888 21788
rect 21824 21728 21888 21732
rect 21904 21788 21968 21792
rect 21904 21732 21908 21788
rect 21908 21732 21964 21788
rect 21964 21732 21968 21788
rect 21904 21728 21968 21732
rect 21984 21788 22048 21792
rect 21984 21732 21988 21788
rect 21988 21732 22044 21788
rect 22044 21732 22048 21788
rect 21984 21728 22048 21732
rect 6868 21388 6932 21452
rect 12204 21660 12268 21724
rect 3551 21244 3615 21248
rect 3551 21188 3555 21244
rect 3555 21188 3611 21244
rect 3611 21188 3615 21244
rect 3551 21184 3615 21188
rect 3631 21244 3695 21248
rect 3631 21188 3635 21244
rect 3635 21188 3691 21244
rect 3691 21188 3695 21244
rect 3631 21184 3695 21188
rect 3711 21244 3775 21248
rect 3711 21188 3715 21244
rect 3715 21188 3771 21244
rect 3771 21188 3775 21244
rect 3711 21184 3775 21188
rect 3791 21244 3855 21248
rect 3791 21188 3795 21244
rect 3795 21188 3851 21244
rect 3851 21188 3855 21244
rect 3791 21184 3855 21188
rect 2084 21116 2148 21180
rect 10548 21388 10612 21452
rect 12204 21388 12268 21452
rect 8749 21244 8813 21248
rect 8749 21188 8753 21244
rect 8753 21188 8809 21244
rect 8809 21188 8813 21244
rect 8749 21184 8813 21188
rect 8829 21244 8893 21248
rect 8829 21188 8833 21244
rect 8833 21188 8889 21244
rect 8889 21188 8893 21244
rect 8829 21184 8893 21188
rect 8909 21244 8973 21248
rect 8909 21188 8913 21244
rect 8913 21188 8969 21244
rect 8969 21188 8973 21244
rect 8909 21184 8973 21188
rect 8989 21244 9053 21248
rect 8989 21188 8993 21244
rect 8993 21188 9049 21244
rect 9049 21188 9053 21244
rect 8989 21184 9053 21188
rect 13947 21244 14011 21248
rect 13947 21188 13951 21244
rect 13951 21188 14007 21244
rect 14007 21188 14011 21244
rect 13947 21184 14011 21188
rect 14027 21244 14091 21248
rect 14027 21188 14031 21244
rect 14031 21188 14087 21244
rect 14087 21188 14091 21244
rect 14027 21184 14091 21188
rect 14107 21244 14171 21248
rect 14107 21188 14111 21244
rect 14111 21188 14167 21244
rect 14167 21188 14171 21244
rect 14107 21184 14171 21188
rect 14187 21244 14251 21248
rect 14187 21188 14191 21244
rect 14191 21188 14247 21244
rect 14247 21188 14251 21244
rect 14187 21184 14251 21188
rect 19145 21244 19209 21248
rect 19145 21188 19149 21244
rect 19149 21188 19205 21244
rect 19205 21188 19209 21244
rect 19145 21184 19209 21188
rect 19225 21244 19289 21248
rect 19225 21188 19229 21244
rect 19229 21188 19285 21244
rect 19285 21188 19289 21244
rect 19225 21184 19289 21188
rect 19305 21244 19369 21248
rect 19305 21188 19309 21244
rect 19309 21188 19365 21244
rect 19365 21188 19369 21244
rect 19305 21184 19369 21188
rect 19385 21244 19449 21248
rect 19385 21188 19389 21244
rect 19389 21188 19445 21244
rect 19445 21188 19449 21244
rect 19385 21184 19449 21188
rect 9812 21116 9876 21180
rect 15884 21116 15948 21180
rect 13676 20844 13740 20908
rect 19012 20844 19076 20908
rect 19748 20844 19812 20908
rect 2636 20632 2700 20636
rect 2636 20576 2650 20632
rect 2650 20576 2700 20632
rect 2636 20572 2700 20576
rect 5764 20708 5828 20772
rect 6150 20700 6214 20704
rect 6150 20644 6154 20700
rect 6154 20644 6210 20700
rect 6210 20644 6214 20700
rect 6150 20640 6214 20644
rect 6230 20700 6294 20704
rect 6230 20644 6234 20700
rect 6234 20644 6290 20700
rect 6290 20644 6294 20700
rect 6230 20640 6294 20644
rect 6310 20700 6374 20704
rect 6310 20644 6314 20700
rect 6314 20644 6370 20700
rect 6370 20644 6374 20700
rect 6310 20640 6374 20644
rect 6390 20700 6454 20704
rect 6390 20644 6394 20700
rect 6394 20644 6450 20700
rect 6450 20644 6454 20700
rect 6390 20640 6454 20644
rect 11348 20700 11412 20704
rect 11348 20644 11352 20700
rect 11352 20644 11408 20700
rect 11408 20644 11412 20700
rect 11348 20640 11412 20644
rect 11428 20700 11492 20704
rect 11428 20644 11432 20700
rect 11432 20644 11488 20700
rect 11488 20644 11492 20700
rect 11428 20640 11492 20644
rect 11508 20700 11572 20704
rect 11508 20644 11512 20700
rect 11512 20644 11568 20700
rect 11568 20644 11572 20700
rect 11508 20640 11572 20644
rect 11588 20700 11652 20704
rect 11588 20644 11592 20700
rect 11592 20644 11648 20700
rect 11648 20644 11652 20700
rect 11588 20640 11652 20644
rect 9444 20572 9508 20636
rect 10364 20572 10428 20636
rect 3924 20436 3988 20500
rect 12572 20708 12636 20772
rect 13124 20708 13188 20772
rect 15148 20708 15212 20772
rect 16068 20708 16132 20772
rect 16546 20700 16610 20704
rect 16546 20644 16550 20700
rect 16550 20644 16606 20700
rect 16606 20644 16610 20700
rect 16546 20640 16610 20644
rect 16626 20700 16690 20704
rect 16626 20644 16630 20700
rect 16630 20644 16686 20700
rect 16686 20644 16690 20700
rect 16626 20640 16690 20644
rect 16706 20700 16770 20704
rect 16706 20644 16710 20700
rect 16710 20644 16766 20700
rect 16766 20644 16770 20700
rect 16706 20640 16770 20644
rect 16786 20700 16850 20704
rect 16786 20644 16790 20700
rect 16790 20644 16846 20700
rect 16846 20644 16850 20700
rect 16786 20640 16850 20644
rect 21744 20700 21808 20704
rect 21744 20644 21748 20700
rect 21748 20644 21804 20700
rect 21804 20644 21808 20700
rect 21744 20640 21808 20644
rect 21824 20700 21888 20704
rect 21824 20644 21828 20700
rect 21828 20644 21884 20700
rect 21884 20644 21888 20700
rect 21824 20640 21888 20644
rect 21904 20700 21968 20704
rect 21904 20644 21908 20700
rect 21908 20644 21964 20700
rect 21964 20644 21968 20700
rect 21904 20640 21968 20644
rect 21984 20700 22048 20704
rect 21984 20644 21988 20700
rect 21988 20644 22044 20700
rect 22044 20644 22048 20700
rect 21984 20640 22048 20644
rect 12940 20436 13004 20500
rect 15332 20436 15396 20500
rect 16068 20300 16132 20364
rect 3551 20156 3615 20160
rect 3551 20100 3555 20156
rect 3555 20100 3611 20156
rect 3611 20100 3615 20156
rect 3551 20096 3615 20100
rect 3631 20156 3695 20160
rect 3631 20100 3635 20156
rect 3635 20100 3691 20156
rect 3691 20100 3695 20156
rect 3631 20096 3695 20100
rect 3711 20156 3775 20160
rect 3711 20100 3715 20156
rect 3715 20100 3771 20156
rect 3771 20100 3775 20156
rect 3711 20096 3775 20100
rect 3791 20156 3855 20160
rect 3791 20100 3795 20156
rect 3795 20100 3851 20156
rect 3851 20100 3855 20156
rect 3791 20096 3855 20100
rect 8749 20156 8813 20160
rect 8749 20100 8753 20156
rect 8753 20100 8809 20156
rect 8809 20100 8813 20156
rect 8749 20096 8813 20100
rect 8829 20156 8893 20160
rect 8829 20100 8833 20156
rect 8833 20100 8889 20156
rect 8889 20100 8893 20156
rect 8829 20096 8893 20100
rect 8909 20156 8973 20160
rect 8909 20100 8913 20156
rect 8913 20100 8969 20156
rect 8969 20100 8973 20156
rect 8909 20096 8973 20100
rect 8989 20156 9053 20160
rect 8989 20100 8993 20156
rect 8993 20100 9049 20156
rect 9049 20100 9053 20156
rect 8989 20096 9053 20100
rect 13947 20156 14011 20160
rect 13947 20100 13951 20156
rect 13951 20100 14007 20156
rect 14007 20100 14011 20156
rect 13947 20096 14011 20100
rect 14027 20156 14091 20160
rect 14027 20100 14031 20156
rect 14031 20100 14087 20156
rect 14087 20100 14091 20156
rect 14027 20096 14091 20100
rect 14107 20156 14171 20160
rect 14107 20100 14111 20156
rect 14111 20100 14167 20156
rect 14167 20100 14171 20156
rect 14107 20096 14171 20100
rect 14187 20156 14251 20160
rect 14187 20100 14191 20156
rect 14191 20100 14247 20156
rect 14247 20100 14251 20156
rect 14187 20096 14251 20100
rect 19145 20156 19209 20160
rect 19145 20100 19149 20156
rect 19149 20100 19205 20156
rect 19205 20100 19209 20156
rect 19145 20096 19209 20100
rect 19225 20156 19289 20160
rect 19225 20100 19229 20156
rect 19229 20100 19285 20156
rect 19285 20100 19289 20156
rect 19225 20096 19289 20100
rect 19305 20156 19369 20160
rect 19305 20100 19309 20156
rect 19309 20100 19365 20156
rect 19365 20100 19369 20156
rect 19305 20096 19369 20100
rect 19385 20156 19449 20160
rect 19385 20100 19389 20156
rect 19389 20100 19445 20156
rect 19445 20100 19449 20156
rect 19385 20096 19449 20100
rect 4660 20028 4724 20092
rect 7052 20028 7116 20092
rect 8340 20028 8404 20092
rect 2452 19756 2516 19820
rect 8524 19756 8588 19820
rect 14412 19756 14476 19820
rect 19564 19756 19628 19820
rect 7604 19620 7668 19684
rect 6150 19612 6214 19616
rect 6150 19556 6154 19612
rect 6154 19556 6210 19612
rect 6210 19556 6214 19612
rect 6150 19552 6214 19556
rect 6230 19612 6294 19616
rect 6230 19556 6234 19612
rect 6234 19556 6290 19612
rect 6290 19556 6294 19612
rect 6230 19552 6294 19556
rect 6310 19612 6374 19616
rect 6310 19556 6314 19612
rect 6314 19556 6370 19612
rect 6370 19556 6374 19612
rect 6310 19552 6374 19556
rect 6390 19612 6454 19616
rect 6390 19556 6394 19612
rect 6394 19556 6450 19612
rect 6450 19556 6454 19612
rect 6390 19552 6454 19556
rect 11348 19612 11412 19616
rect 11348 19556 11352 19612
rect 11352 19556 11408 19612
rect 11408 19556 11412 19612
rect 11348 19552 11412 19556
rect 11428 19612 11492 19616
rect 11428 19556 11432 19612
rect 11432 19556 11488 19612
rect 11488 19556 11492 19612
rect 11428 19552 11492 19556
rect 11508 19612 11572 19616
rect 11508 19556 11512 19612
rect 11512 19556 11568 19612
rect 11568 19556 11572 19612
rect 11508 19552 11572 19556
rect 11588 19612 11652 19616
rect 11588 19556 11592 19612
rect 11592 19556 11648 19612
rect 11648 19556 11652 19612
rect 11588 19552 11652 19556
rect 16546 19612 16610 19616
rect 16546 19556 16550 19612
rect 16550 19556 16606 19612
rect 16606 19556 16610 19612
rect 16546 19552 16610 19556
rect 16626 19612 16690 19616
rect 16626 19556 16630 19612
rect 16630 19556 16686 19612
rect 16686 19556 16690 19612
rect 16626 19552 16690 19556
rect 16706 19612 16770 19616
rect 16706 19556 16710 19612
rect 16710 19556 16766 19612
rect 16766 19556 16770 19612
rect 16706 19552 16770 19556
rect 16786 19612 16850 19616
rect 16786 19556 16790 19612
rect 16790 19556 16846 19612
rect 16846 19556 16850 19612
rect 16786 19552 16850 19556
rect 21744 19612 21808 19616
rect 21744 19556 21748 19612
rect 21748 19556 21804 19612
rect 21804 19556 21808 19612
rect 21744 19552 21808 19556
rect 21824 19612 21888 19616
rect 21824 19556 21828 19612
rect 21828 19556 21884 19612
rect 21884 19556 21888 19612
rect 21824 19552 21888 19556
rect 21904 19612 21968 19616
rect 21904 19556 21908 19612
rect 21908 19556 21964 19612
rect 21964 19556 21968 19612
rect 21904 19552 21968 19556
rect 21984 19612 22048 19616
rect 21984 19556 21988 19612
rect 21988 19556 22044 19612
rect 22044 19556 22048 19612
rect 21984 19552 22048 19556
rect 3004 19484 3068 19548
rect 5028 19484 5092 19548
rect 5212 19348 5276 19412
rect 3551 19068 3615 19072
rect 3551 19012 3555 19068
rect 3555 19012 3611 19068
rect 3611 19012 3615 19068
rect 3551 19008 3615 19012
rect 3631 19068 3695 19072
rect 3631 19012 3635 19068
rect 3635 19012 3691 19068
rect 3691 19012 3695 19068
rect 3631 19008 3695 19012
rect 3711 19068 3775 19072
rect 3711 19012 3715 19068
rect 3715 19012 3771 19068
rect 3771 19012 3775 19068
rect 3711 19008 3775 19012
rect 3791 19068 3855 19072
rect 3791 19012 3795 19068
rect 3795 19012 3851 19068
rect 3851 19012 3855 19068
rect 3791 19008 3855 19012
rect 1164 18940 1228 19004
rect 3188 18940 3252 19004
rect 17724 19348 17788 19412
rect 20852 19348 20916 19412
rect 18644 19212 18708 19276
rect 5948 19076 6012 19140
rect 5212 18940 5276 19004
rect 8749 19068 8813 19072
rect 8749 19012 8753 19068
rect 8753 19012 8809 19068
rect 8809 19012 8813 19068
rect 8749 19008 8813 19012
rect 8829 19068 8893 19072
rect 8829 19012 8833 19068
rect 8833 19012 8889 19068
rect 8889 19012 8893 19068
rect 8829 19008 8893 19012
rect 8909 19068 8973 19072
rect 8909 19012 8913 19068
rect 8913 19012 8969 19068
rect 8969 19012 8973 19068
rect 8909 19008 8973 19012
rect 8989 19068 9053 19072
rect 8989 19012 8993 19068
rect 8993 19012 9049 19068
rect 9049 19012 9053 19068
rect 8989 19008 9053 19012
rect 13947 19068 14011 19072
rect 13947 19012 13951 19068
rect 13951 19012 14007 19068
rect 14007 19012 14011 19068
rect 13947 19008 14011 19012
rect 14027 19068 14091 19072
rect 14027 19012 14031 19068
rect 14031 19012 14087 19068
rect 14087 19012 14091 19068
rect 14027 19008 14091 19012
rect 14107 19068 14171 19072
rect 14107 19012 14111 19068
rect 14111 19012 14167 19068
rect 14167 19012 14171 19068
rect 14107 19008 14171 19012
rect 14187 19068 14251 19072
rect 14187 19012 14191 19068
rect 14191 19012 14247 19068
rect 14247 19012 14251 19068
rect 14187 19008 14251 19012
rect 19145 19068 19209 19072
rect 19145 19012 19149 19068
rect 19149 19012 19205 19068
rect 19205 19012 19209 19068
rect 19145 19008 19209 19012
rect 19225 19068 19289 19072
rect 19225 19012 19229 19068
rect 19229 19012 19285 19068
rect 19285 19012 19289 19068
rect 19225 19008 19289 19012
rect 19305 19068 19369 19072
rect 19305 19012 19309 19068
rect 19309 19012 19365 19068
rect 19365 19012 19369 19068
rect 19305 19008 19369 19012
rect 19385 19068 19449 19072
rect 19385 19012 19389 19068
rect 19389 19012 19445 19068
rect 19445 19012 19449 19068
rect 19385 19008 19449 19012
rect 4292 18668 4356 18732
rect 7052 18532 7116 18596
rect 6150 18524 6214 18528
rect 6150 18468 6154 18524
rect 6154 18468 6210 18524
rect 6210 18468 6214 18524
rect 6150 18464 6214 18468
rect 6230 18524 6294 18528
rect 6230 18468 6234 18524
rect 6234 18468 6290 18524
rect 6290 18468 6294 18524
rect 6230 18464 6294 18468
rect 6310 18524 6374 18528
rect 6310 18468 6314 18524
rect 6314 18468 6370 18524
rect 6370 18468 6374 18524
rect 6310 18464 6374 18468
rect 6390 18524 6454 18528
rect 6390 18468 6394 18524
rect 6394 18468 6450 18524
rect 6450 18468 6454 18524
rect 6390 18464 6454 18468
rect 10548 18532 10612 18596
rect 7236 18396 7300 18460
rect 16068 18804 16132 18868
rect 18092 18668 18156 18732
rect 11348 18524 11412 18528
rect 11348 18468 11352 18524
rect 11352 18468 11408 18524
rect 11408 18468 11412 18524
rect 11348 18464 11412 18468
rect 11428 18524 11492 18528
rect 11428 18468 11432 18524
rect 11432 18468 11488 18524
rect 11488 18468 11492 18524
rect 11428 18464 11492 18468
rect 11508 18524 11572 18528
rect 11508 18468 11512 18524
rect 11512 18468 11568 18524
rect 11568 18468 11572 18524
rect 11508 18464 11572 18468
rect 11588 18524 11652 18528
rect 11588 18468 11592 18524
rect 11592 18468 11648 18524
rect 11648 18468 11652 18524
rect 11588 18464 11652 18468
rect 16546 18524 16610 18528
rect 16546 18468 16550 18524
rect 16550 18468 16606 18524
rect 16606 18468 16610 18524
rect 16546 18464 16610 18468
rect 16626 18524 16690 18528
rect 16626 18468 16630 18524
rect 16630 18468 16686 18524
rect 16686 18468 16690 18524
rect 16626 18464 16690 18468
rect 16706 18524 16770 18528
rect 16706 18468 16710 18524
rect 16710 18468 16766 18524
rect 16766 18468 16770 18524
rect 16706 18464 16770 18468
rect 16786 18524 16850 18528
rect 16786 18468 16790 18524
rect 16790 18468 16846 18524
rect 16846 18468 16850 18524
rect 16786 18464 16850 18468
rect 21744 18524 21808 18528
rect 21744 18468 21748 18524
rect 21748 18468 21804 18524
rect 21804 18468 21808 18524
rect 21744 18464 21808 18468
rect 21824 18524 21888 18528
rect 21824 18468 21828 18524
rect 21828 18468 21884 18524
rect 21884 18468 21888 18524
rect 21824 18464 21888 18468
rect 21904 18524 21968 18528
rect 21904 18468 21908 18524
rect 21908 18468 21964 18524
rect 21964 18468 21968 18524
rect 21904 18464 21968 18468
rect 21984 18524 22048 18528
rect 21984 18468 21988 18524
rect 21988 18468 22044 18524
rect 22044 18468 22048 18524
rect 21984 18464 22048 18468
rect 8156 18260 8220 18324
rect 6684 17988 6748 18052
rect 16988 18124 17052 18188
rect 3551 17980 3615 17984
rect 3551 17924 3555 17980
rect 3555 17924 3611 17980
rect 3611 17924 3615 17980
rect 3551 17920 3615 17924
rect 3631 17980 3695 17984
rect 3631 17924 3635 17980
rect 3635 17924 3691 17980
rect 3691 17924 3695 17980
rect 3631 17920 3695 17924
rect 3711 17980 3775 17984
rect 3711 17924 3715 17980
rect 3715 17924 3771 17980
rect 3771 17924 3775 17980
rect 3711 17920 3775 17924
rect 3791 17980 3855 17984
rect 3791 17924 3795 17980
rect 3795 17924 3851 17980
rect 3851 17924 3855 17980
rect 3791 17920 3855 17924
rect 3372 17852 3436 17916
rect 4108 17912 4172 17916
rect 4108 17856 4122 17912
rect 4122 17856 4172 17912
rect 4108 17852 4172 17856
rect 16252 17988 16316 18052
rect 16988 17988 17052 18052
rect 8749 17980 8813 17984
rect 8749 17924 8753 17980
rect 8753 17924 8809 17980
rect 8809 17924 8813 17980
rect 8749 17920 8813 17924
rect 8829 17980 8893 17984
rect 8829 17924 8833 17980
rect 8833 17924 8889 17980
rect 8889 17924 8893 17980
rect 8829 17920 8893 17924
rect 8909 17980 8973 17984
rect 8909 17924 8913 17980
rect 8913 17924 8969 17980
rect 8969 17924 8973 17980
rect 8909 17920 8973 17924
rect 8989 17980 9053 17984
rect 8989 17924 8993 17980
rect 8993 17924 9049 17980
rect 9049 17924 9053 17980
rect 8989 17920 9053 17924
rect 13947 17980 14011 17984
rect 13947 17924 13951 17980
rect 13951 17924 14007 17980
rect 14007 17924 14011 17980
rect 13947 17920 14011 17924
rect 14027 17980 14091 17984
rect 14027 17924 14031 17980
rect 14031 17924 14087 17980
rect 14087 17924 14091 17980
rect 14027 17920 14091 17924
rect 14107 17980 14171 17984
rect 14107 17924 14111 17980
rect 14111 17924 14167 17980
rect 14167 17924 14171 17980
rect 14107 17920 14171 17924
rect 14187 17980 14251 17984
rect 14187 17924 14191 17980
rect 14191 17924 14247 17980
rect 14247 17924 14251 17980
rect 14187 17920 14251 17924
rect 19145 17980 19209 17984
rect 19145 17924 19149 17980
rect 19149 17924 19205 17980
rect 19205 17924 19209 17980
rect 19145 17920 19209 17924
rect 19225 17980 19289 17984
rect 19225 17924 19229 17980
rect 19229 17924 19285 17980
rect 19285 17924 19289 17980
rect 19225 17920 19289 17924
rect 19305 17980 19369 17984
rect 19305 17924 19309 17980
rect 19309 17924 19365 17980
rect 19365 17924 19369 17980
rect 19305 17920 19369 17924
rect 19385 17980 19449 17984
rect 19385 17924 19389 17980
rect 19389 17924 19445 17980
rect 19445 17924 19449 17980
rect 19385 17920 19449 17924
rect 9444 17852 9508 17916
rect 12940 17716 13004 17780
rect 15884 17716 15948 17780
rect 1532 17580 1596 17644
rect 4844 17444 4908 17508
rect 6150 17436 6214 17440
rect 6150 17380 6154 17436
rect 6154 17380 6210 17436
rect 6210 17380 6214 17436
rect 6150 17376 6214 17380
rect 6230 17436 6294 17440
rect 6230 17380 6234 17436
rect 6234 17380 6290 17436
rect 6290 17380 6294 17436
rect 6230 17376 6294 17380
rect 6310 17436 6374 17440
rect 6310 17380 6314 17436
rect 6314 17380 6370 17436
rect 6370 17380 6374 17436
rect 6310 17376 6374 17380
rect 6390 17436 6454 17440
rect 6390 17380 6394 17436
rect 6394 17380 6450 17436
rect 6450 17380 6454 17436
rect 6390 17376 6454 17380
rect 2636 17368 2700 17372
rect 2636 17312 2686 17368
rect 2686 17312 2700 17368
rect 2636 17308 2700 17312
rect 2820 17308 2884 17372
rect 3924 17308 3988 17372
rect 7604 17444 7668 17508
rect 14964 17580 15028 17644
rect 10732 17444 10796 17508
rect 14412 17444 14476 17508
rect 15148 17444 15212 17508
rect 11348 17436 11412 17440
rect 11348 17380 11352 17436
rect 11352 17380 11408 17436
rect 11408 17380 11412 17436
rect 11348 17376 11412 17380
rect 11428 17436 11492 17440
rect 11428 17380 11432 17436
rect 11432 17380 11488 17436
rect 11488 17380 11492 17436
rect 11428 17376 11492 17380
rect 11508 17436 11572 17440
rect 11508 17380 11512 17436
rect 11512 17380 11568 17436
rect 11568 17380 11572 17436
rect 11508 17376 11572 17380
rect 11588 17436 11652 17440
rect 11588 17380 11592 17436
rect 11592 17380 11648 17436
rect 11648 17380 11652 17436
rect 11588 17376 11652 17380
rect 16546 17436 16610 17440
rect 16546 17380 16550 17436
rect 16550 17380 16606 17436
rect 16606 17380 16610 17436
rect 16546 17376 16610 17380
rect 16626 17436 16690 17440
rect 16626 17380 16630 17436
rect 16630 17380 16686 17436
rect 16686 17380 16690 17436
rect 16626 17376 16690 17380
rect 16706 17436 16770 17440
rect 16706 17380 16710 17436
rect 16710 17380 16766 17436
rect 16766 17380 16770 17436
rect 16706 17376 16770 17380
rect 16786 17436 16850 17440
rect 16786 17380 16790 17436
rect 16790 17380 16846 17436
rect 16846 17380 16850 17436
rect 16786 17376 16850 17380
rect 21744 17436 21808 17440
rect 21744 17380 21748 17436
rect 21748 17380 21804 17436
rect 21804 17380 21808 17436
rect 21744 17376 21808 17380
rect 21824 17436 21888 17440
rect 21824 17380 21828 17436
rect 21828 17380 21884 17436
rect 21884 17380 21888 17436
rect 21824 17376 21888 17380
rect 21904 17436 21968 17440
rect 21904 17380 21908 17436
rect 21908 17380 21964 17436
rect 21964 17380 21968 17436
rect 21904 17376 21968 17380
rect 21984 17436 22048 17440
rect 21984 17380 21988 17436
rect 21988 17380 22044 17436
rect 22044 17380 22048 17436
rect 21984 17376 22048 17380
rect 13676 17308 13740 17372
rect 21220 17232 21284 17236
rect 21220 17176 21270 17232
rect 21270 17176 21284 17232
rect 21220 17172 21284 17176
rect 13492 17036 13556 17100
rect 3551 16892 3615 16896
rect 3551 16836 3555 16892
rect 3555 16836 3611 16892
rect 3611 16836 3615 16892
rect 3551 16832 3615 16836
rect 3631 16892 3695 16896
rect 3631 16836 3635 16892
rect 3635 16836 3691 16892
rect 3691 16836 3695 16892
rect 3631 16832 3695 16836
rect 3711 16892 3775 16896
rect 3711 16836 3715 16892
rect 3715 16836 3771 16892
rect 3771 16836 3775 16892
rect 3711 16832 3775 16836
rect 3791 16892 3855 16896
rect 3791 16836 3795 16892
rect 3795 16836 3851 16892
rect 3851 16836 3855 16892
rect 3791 16832 3855 16836
rect 8749 16892 8813 16896
rect 8749 16836 8753 16892
rect 8753 16836 8809 16892
rect 8809 16836 8813 16892
rect 8749 16832 8813 16836
rect 8829 16892 8893 16896
rect 8829 16836 8833 16892
rect 8833 16836 8889 16892
rect 8889 16836 8893 16892
rect 8829 16832 8893 16836
rect 8909 16892 8973 16896
rect 8909 16836 8913 16892
rect 8913 16836 8969 16892
rect 8969 16836 8973 16892
rect 8909 16832 8973 16836
rect 8989 16892 9053 16896
rect 8989 16836 8993 16892
rect 8993 16836 9049 16892
rect 9049 16836 9053 16892
rect 8989 16832 9053 16836
rect 13947 16892 14011 16896
rect 13947 16836 13951 16892
rect 13951 16836 14007 16892
rect 14007 16836 14011 16892
rect 13947 16832 14011 16836
rect 14027 16892 14091 16896
rect 14027 16836 14031 16892
rect 14031 16836 14087 16892
rect 14087 16836 14091 16892
rect 14027 16832 14091 16836
rect 14107 16892 14171 16896
rect 14107 16836 14111 16892
rect 14111 16836 14167 16892
rect 14167 16836 14171 16892
rect 14107 16832 14171 16836
rect 14187 16892 14251 16896
rect 14187 16836 14191 16892
rect 14191 16836 14247 16892
rect 14247 16836 14251 16892
rect 14187 16832 14251 16836
rect 796 16764 860 16828
rect 1900 16764 1964 16828
rect 2268 16824 2332 16828
rect 2268 16768 2318 16824
rect 2318 16768 2332 16824
rect 2268 16764 2332 16768
rect 4108 16628 4172 16692
rect 19145 16892 19209 16896
rect 19145 16836 19149 16892
rect 19149 16836 19205 16892
rect 19205 16836 19209 16892
rect 19145 16832 19209 16836
rect 19225 16892 19289 16896
rect 19225 16836 19229 16892
rect 19229 16836 19285 16892
rect 19285 16836 19289 16892
rect 19225 16832 19289 16836
rect 19305 16892 19369 16896
rect 19305 16836 19309 16892
rect 19309 16836 19365 16892
rect 19365 16836 19369 16892
rect 19305 16832 19369 16836
rect 19385 16892 19449 16896
rect 19385 16836 19389 16892
rect 19389 16836 19445 16892
rect 19445 16836 19449 16892
rect 19385 16832 19449 16836
rect 8156 16628 8220 16692
rect 10548 16688 10612 16692
rect 10548 16632 10562 16688
rect 10562 16632 10612 16688
rect 10548 16628 10612 16632
rect 10916 16628 10980 16692
rect 14596 16628 14660 16692
rect 3372 16492 3436 16556
rect 6868 16492 6932 16556
rect 10180 16492 10244 16556
rect 14780 16492 14844 16556
rect 6150 16348 6214 16352
rect 6150 16292 6154 16348
rect 6154 16292 6210 16348
rect 6210 16292 6214 16348
rect 6150 16288 6214 16292
rect 6230 16348 6294 16352
rect 6230 16292 6234 16348
rect 6234 16292 6290 16348
rect 6290 16292 6294 16348
rect 6230 16288 6294 16292
rect 6310 16348 6374 16352
rect 6310 16292 6314 16348
rect 6314 16292 6370 16348
rect 6370 16292 6374 16348
rect 6310 16288 6374 16292
rect 6390 16348 6454 16352
rect 6390 16292 6394 16348
rect 6394 16292 6450 16348
rect 6450 16292 6454 16348
rect 6390 16288 6454 16292
rect 11348 16348 11412 16352
rect 11348 16292 11352 16348
rect 11352 16292 11408 16348
rect 11408 16292 11412 16348
rect 11348 16288 11412 16292
rect 11428 16348 11492 16352
rect 11428 16292 11432 16348
rect 11432 16292 11488 16348
rect 11488 16292 11492 16348
rect 11428 16288 11492 16292
rect 11508 16348 11572 16352
rect 11508 16292 11512 16348
rect 11512 16292 11568 16348
rect 11568 16292 11572 16348
rect 11508 16288 11572 16292
rect 11588 16348 11652 16352
rect 11588 16292 11592 16348
rect 11592 16292 11648 16348
rect 11648 16292 11652 16348
rect 11588 16288 11652 16292
rect 16546 16348 16610 16352
rect 16546 16292 16550 16348
rect 16550 16292 16606 16348
rect 16606 16292 16610 16348
rect 16546 16288 16610 16292
rect 16626 16348 16690 16352
rect 16626 16292 16630 16348
rect 16630 16292 16686 16348
rect 16686 16292 16690 16348
rect 16626 16288 16690 16292
rect 16706 16348 16770 16352
rect 16706 16292 16710 16348
rect 16710 16292 16766 16348
rect 16766 16292 16770 16348
rect 16706 16288 16770 16292
rect 16786 16348 16850 16352
rect 16786 16292 16790 16348
rect 16790 16292 16846 16348
rect 16846 16292 16850 16348
rect 16786 16288 16850 16292
rect 21744 16348 21808 16352
rect 21744 16292 21748 16348
rect 21748 16292 21804 16348
rect 21804 16292 21808 16348
rect 21744 16288 21808 16292
rect 21824 16348 21888 16352
rect 21824 16292 21828 16348
rect 21828 16292 21884 16348
rect 21884 16292 21888 16348
rect 21824 16288 21888 16292
rect 21904 16348 21968 16352
rect 21904 16292 21908 16348
rect 21908 16292 21964 16348
rect 21964 16292 21968 16348
rect 21904 16288 21968 16292
rect 21984 16348 22048 16352
rect 21984 16292 21988 16348
rect 21988 16292 22044 16348
rect 22044 16292 22048 16348
rect 21984 16288 22048 16292
rect 10916 16220 10980 16284
rect 244 16084 308 16148
rect 1716 16084 1780 16148
rect 5396 16084 5460 16148
rect 11836 16084 11900 16148
rect 4844 15872 4908 15876
rect 4844 15816 4894 15872
rect 4894 15816 4908 15872
rect 4844 15812 4908 15816
rect 3551 15804 3615 15808
rect 3551 15748 3555 15804
rect 3555 15748 3611 15804
rect 3611 15748 3615 15804
rect 3551 15744 3615 15748
rect 3631 15804 3695 15808
rect 3631 15748 3635 15804
rect 3635 15748 3691 15804
rect 3691 15748 3695 15804
rect 3631 15744 3695 15748
rect 3711 15804 3775 15808
rect 3711 15748 3715 15804
rect 3715 15748 3771 15804
rect 3771 15748 3775 15804
rect 3711 15744 3775 15748
rect 3791 15804 3855 15808
rect 3791 15748 3795 15804
rect 3795 15748 3851 15804
rect 3851 15748 3855 15804
rect 3791 15744 3855 15748
rect 4108 15676 4172 15740
rect 7788 15948 7852 16012
rect 19012 15948 19076 16012
rect 13676 15812 13740 15876
rect 8749 15804 8813 15808
rect 8749 15748 8753 15804
rect 8753 15748 8809 15804
rect 8809 15748 8813 15804
rect 8749 15744 8813 15748
rect 8829 15804 8893 15808
rect 8829 15748 8833 15804
rect 8833 15748 8889 15804
rect 8889 15748 8893 15804
rect 8829 15744 8893 15748
rect 8909 15804 8973 15808
rect 8909 15748 8913 15804
rect 8913 15748 8969 15804
rect 8969 15748 8973 15804
rect 8909 15744 8973 15748
rect 8989 15804 9053 15808
rect 8989 15748 8993 15804
rect 8993 15748 9049 15804
rect 9049 15748 9053 15804
rect 8989 15744 9053 15748
rect 13947 15804 14011 15808
rect 13947 15748 13951 15804
rect 13951 15748 14007 15804
rect 14007 15748 14011 15804
rect 13947 15744 14011 15748
rect 14027 15804 14091 15808
rect 14027 15748 14031 15804
rect 14031 15748 14087 15804
rect 14087 15748 14091 15804
rect 14027 15744 14091 15748
rect 14107 15804 14171 15808
rect 14107 15748 14111 15804
rect 14111 15748 14167 15804
rect 14167 15748 14171 15804
rect 14107 15744 14171 15748
rect 14187 15804 14251 15808
rect 14187 15748 14191 15804
rect 14191 15748 14247 15804
rect 14247 15748 14251 15804
rect 14187 15744 14251 15748
rect 19145 15804 19209 15808
rect 19145 15748 19149 15804
rect 19149 15748 19205 15804
rect 19205 15748 19209 15804
rect 19145 15744 19209 15748
rect 19225 15804 19289 15808
rect 19225 15748 19229 15804
rect 19229 15748 19285 15804
rect 19285 15748 19289 15804
rect 19225 15744 19289 15748
rect 19305 15804 19369 15808
rect 19305 15748 19309 15804
rect 19309 15748 19365 15804
rect 19365 15748 19369 15804
rect 19305 15744 19369 15748
rect 19385 15804 19449 15808
rect 19385 15748 19389 15804
rect 19389 15748 19445 15804
rect 19445 15748 19449 15804
rect 19385 15744 19449 15748
rect 6684 15676 6748 15740
rect 4476 15600 4540 15604
rect 4476 15544 4526 15600
rect 4526 15544 4540 15600
rect 4476 15540 4540 15544
rect 7052 15540 7116 15604
rect 10180 15540 10244 15604
rect 16252 15600 16316 15604
rect 16252 15544 16302 15600
rect 16302 15544 16316 15600
rect 16252 15540 16316 15544
rect 1900 15404 1964 15468
rect 5764 15404 5828 15468
rect 796 15132 860 15196
rect 428 14996 492 15060
rect 18092 15268 18156 15332
rect 6150 15260 6214 15264
rect 6150 15204 6154 15260
rect 6154 15204 6210 15260
rect 6210 15204 6214 15260
rect 6150 15200 6214 15204
rect 6230 15260 6294 15264
rect 6230 15204 6234 15260
rect 6234 15204 6290 15260
rect 6290 15204 6294 15260
rect 6230 15200 6294 15204
rect 6310 15260 6374 15264
rect 6310 15204 6314 15260
rect 6314 15204 6370 15260
rect 6370 15204 6374 15260
rect 6310 15200 6374 15204
rect 6390 15260 6454 15264
rect 6390 15204 6394 15260
rect 6394 15204 6450 15260
rect 6450 15204 6454 15260
rect 6390 15200 6454 15204
rect 11348 15260 11412 15264
rect 11348 15204 11352 15260
rect 11352 15204 11408 15260
rect 11408 15204 11412 15260
rect 11348 15200 11412 15204
rect 11428 15260 11492 15264
rect 11428 15204 11432 15260
rect 11432 15204 11488 15260
rect 11488 15204 11492 15260
rect 11428 15200 11492 15204
rect 11508 15260 11572 15264
rect 11508 15204 11512 15260
rect 11512 15204 11568 15260
rect 11568 15204 11572 15260
rect 11508 15200 11572 15204
rect 11588 15260 11652 15264
rect 11588 15204 11592 15260
rect 11592 15204 11648 15260
rect 11648 15204 11652 15260
rect 11588 15200 11652 15204
rect 16546 15260 16610 15264
rect 16546 15204 16550 15260
rect 16550 15204 16606 15260
rect 16606 15204 16610 15260
rect 16546 15200 16610 15204
rect 16626 15260 16690 15264
rect 16626 15204 16630 15260
rect 16630 15204 16686 15260
rect 16686 15204 16690 15260
rect 16626 15200 16690 15204
rect 16706 15260 16770 15264
rect 16706 15204 16710 15260
rect 16710 15204 16766 15260
rect 16766 15204 16770 15260
rect 16706 15200 16770 15204
rect 16786 15260 16850 15264
rect 16786 15204 16790 15260
rect 16790 15204 16846 15260
rect 16846 15204 16850 15260
rect 16786 15200 16850 15204
rect 21744 15260 21808 15264
rect 21744 15204 21748 15260
rect 21748 15204 21804 15260
rect 21804 15204 21808 15260
rect 21744 15200 21808 15204
rect 21824 15260 21888 15264
rect 21824 15204 21828 15260
rect 21828 15204 21884 15260
rect 21884 15204 21888 15260
rect 21824 15200 21888 15204
rect 21904 15260 21968 15264
rect 21904 15204 21908 15260
rect 21908 15204 21964 15260
rect 21964 15204 21968 15260
rect 21904 15200 21968 15204
rect 21984 15260 22048 15264
rect 21984 15204 21988 15260
rect 21988 15204 22044 15260
rect 22044 15204 22048 15260
rect 21984 15200 22048 15204
rect 5028 15192 5092 15196
rect 5028 15136 5078 15192
rect 5078 15136 5092 15192
rect 5028 15132 5092 15136
rect 8340 15192 8404 15196
rect 8340 15136 8390 15192
rect 8390 15136 8404 15192
rect 8340 15132 8404 15136
rect 13124 15132 13188 15196
rect 15332 15132 15396 15196
rect 2636 15056 2700 15060
rect 2636 15000 2650 15056
rect 2650 15000 2700 15056
rect 2636 14996 2700 15000
rect 3372 14996 3436 15060
rect 6868 14860 6932 14924
rect 9628 14860 9692 14924
rect 12940 14860 13004 14924
rect 18460 14860 18524 14924
rect 20300 14860 20364 14924
rect 3551 14716 3615 14720
rect 3551 14660 3555 14716
rect 3555 14660 3611 14716
rect 3611 14660 3615 14716
rect 3551 14656 3615 14660
rect 3631 14716 3695 14720
rect 3631 14660 3635 14716
rect 3635 14660 3691 14716
rect 3691 14660 3695 14716
rect 3631 14656 3695 14660
rect 3711 14716 3775 14720
rect 3711 14660 3715 14716
rect 3715 14660 3771 14716
rect 3771 14660 3775 14716
rect 3711 14656 3775 14660
rect 3791 14716 3855 14720
rect 3791 14660 3795 14716
rect 3795 14660 3851 14716
rect 3851 14660 3855 14716
rect 3791 14656 3855 14660
rect 3372 14588 3436 14652
rect 4660 14588 4724 14652
rect 8749 14716 8813 14720
rect 8749 14660 8753 14716
rect 8753 14660 8809 14716
rect 8809 14660 8813 14716
rect 8749 14656 8813 14660
rect 8829 14716 8893 14720
rect 8829 14660 8833 14716
rect 8833 14660 8889 14716
rect 8889 14660 8893 14716
rect 8829 14656 8893 14660
rect 8909 14716 8973 14720
rect 8909 14660 8913 14716
rect 8913 14660 8969 14716
rect 8969 14660 8973 14716
rect 8909 14656 8973 14660
rect 8989 14716 9053 14720
rect 8989 14660 8993 14716
rect 8993 14660 9049 14716
rect 9049 14660 9053 14716
rect 8989 14656 9053 14660
rect 13947 14716 14011 14720
rect 13947 14660 13951 14716
rect 13951 14660 14007 14716
rect 14007 14660 14011 14716
rect 13947 14656 14011 14660
rect 14027 14716 14091 14720
rect 14027 14660 14031 14716
rect 14031 14660 14087 14716
rect 14087 14660 14091 14716
rect 14027 14656 14091 14660
rect 14107 14716 14171 14720
rect 14107 14660 14111 14716
rect 14111 14660 14167 14716
rect 14167 14660 14171 14716
rect 14107 14656 14171 14660
rect 14187 14716 14251 14720
rect 14187 14660 14191 14716
rect 14191 14660 14247 14716
rect 14247 14660 14251 14716
rect 14187 14656 14251 14660
rect 19145 14716 19209 14720
rect 19145 14660 19149 14716
rect 19149 14660 19205 14716
rect 19205 14660 19209 14716
rect 19145 14656 19209 14660
rect 19225 14716 19289 14720
rect 19225 14660 19229 14716
rect 19229 14660 19285 14716
rect 19285 14660 19289 14716
rect 19225 14656 19289 14660
rect 19305 14716 19369 14720
rect 19305 14660 19309 14716
rect 19309 14660 19365 14716
rect 19365 14660 19369 14716
rect 19305 14656 19369 14660
rect 19385 14716 19449 14720
rect 19385 14660 19389 14716
rect 19389 14660 19445 14716
rect 19445 14660 19449 14716
rect 19385 14656 19449 14660
rect 12204 14316 12268 14380
rect 3924 14240 3988 14244
rect 3924 14184 3938 14240
rect 3938 14184 3988 14240
rect 3924 14180 3988 14184
rect 6150 14172 6214 14176
rect 6150 14116 6154 14172
rect 6154 14116 6210 14172
rect 6210 14116 6214 14172
rect 6150 14112 6214 14116
rect 6230 14172 6294 14176
rect 6230 14116 6234 14172
rect 6234 14116 6290 14172
rect 6290 14116 6294 14172
rect 6230 14112 6294 14116
rect 6310 14172 6374 14176
rect 6310 14116 6314 14172
rect 6314 14116 6370 14172
rect 6370 14116 6374 14172
rect 6310 14112 6374 14116
rect 6390 14172 6454 14176
rect 6390 14116 6394 14172
rect 6394 14116 6450 14172
rect 6450 14116 6454 14172
rect 6390 14112 6454 14116
rect 11348 14172 11412 14176
rect 11348 14116 11352 14172
rect 11352 14116 11408 14172
rect 11408 14116 11412 14172
rect 11348 14112 11412 14116
rect 11428 14172 11492 14176
rect 11428 14116 11432 14172
rect 11432 14116 11488 14172
rect 11488 14116 11492 14172
rect 11428 14112 11492 14116
rect 11508 14172 11572 14176
rect 11508 14116 11512 14172
rect 11512 14116 11568 14172
rect 11568 14116 11572 14172
rect 11508 14112 11572 14116
rect 11588 14172 11652 14176
rect 11588 14116 11592 14172
rect 11592 14116 11648 14172
rect 11648 14116 11652 14172
rect 11588 14112 11652 14116
rect 16546 14172 16610 14176
rect 16546 14116 16550 14172
rect 16550 14116 16606 14172
rect 16606 14116 16610 14172
rect 16546 14112 16610 14116
rect 16626 14172 16690 14176
rect 16626 14116 16630 14172
rect 16630 14116 16686 14172
rect 16686 14116 16690 14172
rect 16626 14112 16690 14116
rect 16706 14172 16770 14176
rect 16706 14116 16710 14172
rect 16710 14116 16766 14172
rect 16766 14116 16770 14172
rect 16706 14112 16770 14116
rect 16786 14172 16850 14176
rect 16786 14116 16790 14172
rect 16790 14116 16846 14172
rect 16846 14116 16850 14172
rect 16786 14112 16850 14116
rect 21744 14172 21808 14176
rect 21744 14116 21748 14172
rect 21748 14116 21804 14172
rect 21804 14116 21808 14172
rect 21744 14112 21808 14116
rect 21824 14172 21888 14176
rect 21824 14116 21828 14172
rect 21828 14116 21884 14172
rect 21884 14116 21888 14172
rect 21824 14112 21888 14116
rect 21904 14172 21968 14176
rect 21904 14116 21908 14172
rect 21908 14116 21964 14172
rect 21964 14116 21968 14172
rect 21904 14112 21968 14116
rect 21984 14172 22048 14176
rect 21984 14116 21988 14172
rect 21988 14116 22044 14172
rect 22044 14116 22048 14172
rect 21984 14112 22048 14116
rect 5948 14044 6012 14108
rect 13308 14044 13372 14108
rect 17356 13908 17420 13972
rect 18828 13908 18892 13972
rect 244 13772 308 13836
rect 5580 13772 5644 13836
rect 3004 13636 3068 13700
rect 5028 13636 5092 13700
rect 7236 13636 7300 13700
rect 12572 13696 12636 13700
rect 12572 13640 12586 13696
rect 12586 13640 12636 13696
rect 12572 13636 12636 13640
rect 3551 13628 3615 13632
rect 3551 13572 3555 13628
rect 3555 13572 3611 13628
rect 3611 13572 3615 13628
rect 3551 13568 3615 13572
rect 3631 13628 3695 13632
rect 3631 13572 3635 13628
rect 3635 13572 3691 13628
rect 3691 13572 3695 13628
rect 3631 13568 3695 13572
rect 3711 13628 3775 13632
rect 3711 13572 3715 13628
rect 3715 13572 3771 13628
rect 3771 13572 3775 13628
rect 3711 13568 3775 13572
rect 3791 13628 3855 13632
rect 3791 13572 3795 13628
rect 3795 13572 3851 13628
rect 3851 13572 3855 13628
rect 3791 13568 3855 13572
rect 8749 13628 8813 13632
rect 8749 13572 8753 13628
rect 8753 13572 8809 13628
rect 8809 13572 8813 13628
rect 8749 13568 8813 13572
rect 8829 13628 8893 13632
rect 8829 13572 8833 13628
rect 8833 13572 8889 13628
rect 8889 13572 8893 13628
rect 8829 13568 8893 13572
rect 8909 13628 8973 13632
rect 8909 13572 8913 13628
rect 8913 13572 8969 13628
rect 8969 13572 8973 13628
rect 8909 13568 8973 13572
rect 8989 13628 9053 13632
rect 8989 13572 8993 13628
rect 8993 13572 9049 13628
rect 9049 13572 9053 13628
rect 8989 13568 9053 13572
rect 13947 13628 14011 13632
rect 13947 13572 13951 13628
rect 13951 13572 14007 13628
rect 14007 13572 14011 13628
rect 13947 13568 14011 13572
rect 14027 13628 14091 13632
rect 14027 13572 14031 13628
rect 14031 13572 14087 13628
rect 14087 13572 14091 13628
rect 14027 13568 14091 13572
rect 14107 13628 14171 13632
rect 14107 13572 14111 13628
rect 14111 13572 14167 13628
rect 14167 13572 14171 13628
rect 14107 13568 14171 13572
rect 14187 13628 14251 13632
rect 14187 13572 14191 13628
rect 14191 13572 14247 13628
rect 14247 13572 14251 13628
rect 14187 13568 14251 13572
rect 2820 13500 2884 13564
rect 9444 13500 9508 13564
rect 17908 13696 17972 13700
rect 17908 13640 17958 13696
rect 17958 13640 17972 13696
rect 17908 13636 17972 13640
rect 19145 13628 19209 13632
rect 19145 13572 19149 13628
rect 19149 13572 19205 13628
rect 19205 13572 19209 13628
rect 19145 13568 19209 13572
rect 19225 13628 19289 13632
rect 19225 13572 19229 13628
rect 19229 13572 19285 13628
rect 19285 13572 19289 13628
rect 19225 13568 19289 13572
rect 19305 13628 19369 13632
rect 19305 13572 19309 13628
rect 19309 13572 19365 13628
rect 19365 13572 19369 13628
rect 19305 13568 19369 13572
rect 19385 13628 19449 13632
rect 19385 13572 19389 13628
rect 19389 13572 19445 13628
rect 19445 13572 19449 13628
rect 19385 13568 19449 13572
rect 14596 13500 14660 13564
rect 1164 13228 1228 13292
rect 3924 13228 3988 13292
rect 4844 13228 4908 13292
rect 5948 13228 6012 13292
rect 6150 13084 6214 13088
rect 6150 13028 6154 13084
rect 6154 13028 6210 13084
rect 6210 13028 6214 13084
rect 6150 13024 6214 13028
rect 6230 13084 6294 13088
rect 6230 13028 6234 13084
rect 6234 13028 6290 13084
rect 6290 13028 6294 13084
rect 6230 13024 6294 13028
rect 6310 13084 6374 13088
rect 6310 13028 6314 13084
rect 6314 13028 6370 13084
rect 6370 13028 6374 13084
rect 6310 13024 6374 13028
rect 6390 13084 6454 13088
rect 6390 13028 6394 13084
rect 6394 13028 6450 13084
rect 6450 13028 6454 13084
rect 6390 13024 6454 13028
rect 428 12956 492 13020
rect 1348 12956 1412 13020
rect 2084 12956 2148 13020
rect 7236 12820 7300 12884
rect 9444 13228 9508 13292
rect 19932 13228 19996 13292
rect 18828 13092 18892 13156
rect 11348 13084 11412 13088
rect 11348 13028 11352 13084
rect 11352 13028 11408 13084
rect 11408 13028 11412 13084
rect 11348 13024 11412 13028
rect 11428 13084 11492 13088
rect 11428 13028 11432 13084
rect 11432 13028 11488 13084
rect 11488 13028 11492 13084
rect 11428 13024 11492 13028
rect 11508 13084 11572 13088
rect 11508 13028 11512 13084
rect 11512 13028 11568 13084
rect 11568 13028 11572 13084
rect 11508 13024 11572 13028
rect 11588 13084 11652 13088
rect 11588 13028 11592 13084
rect 11592 13028 11648 13084
rect 11648 13028 11652 13084
rect 11588 13024 11652 13028
rect 16546 13084 16610 13088
rect 16546 13028 16550 13084
rect 16550 13028 16606 13084
rect 16606 13028 16610 13084
rect 16546 13024 16610 13028
rect 16626 13084 16690 13088
rect 16626 13028 16630 13084
rect 16630 13028 16686 13084
rect 16686 13028 16690 13084
rect 16626 13024 16690 13028
rect 16706 13084 16770 13088
rect 16706 13028 16710 13084
rect 16710 13028 16766 13084
rect 16766 13028 16770 13084
rect 16706 13024 16770 13028
rect 16786 13084 16850 13088
rect 16786 13028 16790 13084
rect 16790 13028 16846 13084
rect 16846 13028 16850 13084
rect 16786 13024 16850 13028
rect 21744 13084 21808 13088
rect 21744 13028 21748 13084
rect 21748 13028 21804 13084
rect 21804 13028 21808 13084
rect 21744 13024 21808 13028
rect 21824 13084 21888 13088
rect 21824 13028 21828 13084
rect 21828 13028 21884 13084
rect 21884 13028 21888 13084
rect 21824 13024 21888 13028
rect 21904 13084 21968 13088
rect 21904 13028 21908 13084
rect 21908 13028 21964 13084
rect 21964 13028 21968 13084
rect 21904 13024 21968 13028
rect 21984 13084 22048 13088
rect 21984 13028 21988 13084
rect 21988 13028 22044 13084
rect 22044 13028 22048 13084
rect 21984 13024 22048 13028
rect 7052 12548 7116 12612
rect 7604 12608 7668 12612
rect 7604 12552 7654 12608
rect 7654 12552 7668 12608
rect 7604 12548 7668 12552
rect 12020 12548 12084 12612
rect 3551 12540 3615 12544
rect 3551 12484 3555 12540
rect 3555 12484 3611 12540
rect 3611 12484 3615 12540
rect 3551 12480 3615 12484
rect 3631 12540 3695 12544
rect 3631 12484 3635 12540
rect 3635 12484 3691 12540
rect 3691 12484 3695 12540
rect 3631 12480 3695 12484
rect 3711 12540 3775 12544
rect 3711 12484 3715 12540
rect 3715 12484 3771 12540
rect 3771 12484 3775 12540
rect 3711 12480 3775 12484
rect 3791 12540 3855 12544
rect 3791 12484 3795 12540
rect 3795 12484 3851 12540
rect 3851 12484 3855 12540
rect 3791 12480 3855 12484
rect 8749 12540 8813 12544
rect 8749 12484 8753 12540
rect 8753 12484 8809 12540
rect 8809 12484 8813 12540
rect 8749 12480 8813 12484
rect 8829 12540 8893 12544
rect 8829 12484 8833 12540
rect 8833 12484 8889 12540
rect 8889 12484 8893 12540
rect 8829 12480 8893 12484
rect 8909 12540 8973 12544
rect 8909 12484 8913 12540
rect 8913 12484 8969 12540
rect 8969 12484 8973 12540
rect 8909 12480 8973 12484
rect 8989 12540 9053 12544
rect 8989 12484 8993 12540
rect 8993 12484 9049 12540
rect 9049 12484 9053 12540
rect 8989 12480 9053 12484
rect 13947 12540 14011 12544
rect 13947 12484 13951 12540
rect 13951 12484 14007 12540
rect 14007 12484 14011 12540
rect 13947 12480 14011 12484
rect 14027 12540 14091 12544
rect 14027 12484 14031 12540
rect 14031 12484 14087 12540
rect 14087 12484 14091 12540
rect 14027 12480 14091 12484
rect 14107 12540 14171 12544
rect 14107 12484 14111 12540
rect 14111 12484 14167 12540
rect 14167 12484 14171 12540
rect 14107 12480 14171 12484
rect 14187 12540 14251 12544
rect 14187 12484 14191 12540
rect 14191 12484 14247 12540
rect 14247 12484 14251 12540
rect 14187 12480 14251 12484
rect 19145 12540 19209 12544
rect 19145 12484 19149 12540
rect 19149 12484 19205 12540
rect 19205 12484 19209 12540
rect 19145 12480 19209 12484
rect 19225 12540 19289 12544
rect 19225 12484 19229 12540
rect 19229 12484 19285 12540
rect 19285 12484 19289 12540
rect 19225 12480 19289 12484
rect 19305 12540 19369 12544
rect 19305 12484 19309 12540
rect 19309 12484 19365 12540
rect 19365 12484 19369 12540
rect 19305 12480 19369 12484
rect 19385 12540 19449 12544
rect 19385 12484 19389 12540
rect 19389 12484 19445 12540
rect 19445 12484 19449 12540
rect 19385 12480 19449 12484
rect 7788 12412 7852 12476
rect 11100 12412 11164 12476
rect 19748 12412 19812 12476
rect 4660 12276 4724 12340
rect 19012 12336 19076 12340
rect 19012 12280 19062 12336
rect 19062 12280 19076 12336
rect 19012 12276 19076 12280
rect 11100 12200 11164 12204
rect 11100 12144 11114 12200
rect 11114 12144 11164 12200
rect 11100 12140 11164 12144
rect 11836 12140 11900 12204
rect 1532 11792 1596 11796
rect 1532 11736 1582 11792
rect 1582 11736 1596 11792
rect 1532 11732 1596 11736
rect 1900 11732 1964 11796
rect 3188 11868 3252 11932
rect 3924 11868 3988 11932
rect 4108 11928 4172 11932
rect 4108 11872 4158 11928
rect 4158 11872 4172 11928
rect 4108 11868 4172 11872
rect 5580 12004 5644 12068
rect 17172 12004 17236 12068
rect 6150 11996 6214 12000
rect 6150 11940 6154 11996
rect 6154 11940 6210 11996
rect 6210 11940 6214 11996
rect 6150 11936 6214 11940
rect 6230 11996 6294 12000
rect 6230 11940 6234 11996
rect 6234 11940 6290 11996
rect 6290 11940 6294 11996
rect 6230 11936 6294 11940
rect 6310 11996 6374 12000
rect 6310 11940 6314 11996
rect 6314 11940 6370 11996
rect 6370 11940 6374 11996
rect 6310 11936 6374 11940
rect 6390 11996 6454 12000
rect 6390 11940 6394 11996
rect 6394 11940 6450 11996
rect 6450 11940 6454 11996
rect 6390 11936 6454 11940
rect 11348 11996 11412 12000
rect 11348 11940 11352 11996
rect 11352 11940 11408 11996
rect 11408 11940 11412 11996
rect 11348 11936 11412 11940
rect 11428 11996 11492 12000
rect 11428 11940 11432 11996
rect 11432 11940 11488 11996
rect 11488 11940 11492 11996
rect 11428 11936 11492 11940
rect 11508 11996 11572 12000
rect 11508 11940 11512 11996
rect 11512 11940 11568 11996
rect 11568 11940 11572 11996
rect 11508 11936 11572 11940
rect 11588 11996 11652 12000
rect 11588 11940 11592 11996
rect 11592 11940 11648 11996
rect 11648 11940 11652 11996
rect 11588 11936 11652 11940
rect 16546 11996 16610 12000
rect 16546 11940 16550 11996
rect 16550 11940 16606 11996
rect 16606 11940 16610 11996
rect 16546 11936 16610 11940
rect 16626 11996 16690 12000
rect 16626 11940 16630 11996
rect 16630 11940 16686 11996
rect 16686 11940 16690 11996
rect 16626 11936 16690 11940
rect 16706 11996 16770 12000
rect 16706 11940 16710 11996
rect 16710 11940 16766 11996
rect 16766 11940 16770 11996
rect 16706 11936 16770 11940
rect 16786 11996 16850 12000
rect 16786 11940 16790 11996
rect 16790 11940 16846 11996
rect 16846 11940 16850 11996
rect 16786 11936 16850 11940
rect 21744 11996 21808 12000
rect 21744 11940 21748 11996
rect 21748 11940 21804 11996
rect 21804 11940 21808 11996
rect 21744 11936 21808 11940
rect 21824 11996 21888 12000
rect 21824 11940 21828 11996
rect 21828 11940 21884 11996
rect 21884 11940 21888 11996
rect 21824 11936 21888 11940
rect 21904 11996 21968 12000
rect 21904 11940 21908 11996
rect 21908 11940 21964 11996
rect 21964 11940 21968 11996
rect 21904 11936 21968 11940
rect 21984 11996 22048 12000
rect 21984 11940 21988 11996
rect 21988 11940 22044 11996
rect 22044 11940 22048 11996
rect 21984 11936 22048 11940
rect 10180 11732 10244 11796
rect 10364 11732 10428 11796
rect 16988 11868 17052 11932
rect 2084 11596 2148 11660
rect 5212 11460 5276 11524
rect 3551 11452 3615 11456
rect 3551 11396 3555 11452
rect 3555 11396 3611 11452
rect 3611 11396 3615 11452
rect 3551 11392 3615 11396
rect 3631 11452 3695 11456
rect 3631 11396 3635 11452
rect 3635 11396 3691 11452
rect 3691 11396 3695 11452
rect 3631 11392 3695 11396
rect 3711 11452 3775 11456
rect 3711 11396 3715 11452
rect 3715 11396 3771 11452
rect 3771 11396 3775 11452
rect 3711 11392 3775 11396
rect 3791 11452 3855 11456
rect 3791 11396 3795 11452
rect 3795 11396 3851 11452
rect 3851 11396 3855 11452
rect 3791 11392 3855 11396
rect 8749 11452 8813 11456
rect 8749 11396 8753 11452
rect 8753 11396 8809 11452
rect 8809 11396 8813 11452
rect 8749 11392 8813 11396
rect 8829 11452 8893 11456
rect 8829 11396 8833 11452
rect 8833 11396 8889 11452
rect 8889 11396 8893 11452
rect 8829 11392 8893 11396
rect 8909 11452 8973 11456
rect 8909 11396 8913 11452
rect 8913 11396 8969 11452
rect 8969 11396 8973 11452
rect 8909 11392 8973 11396
rect 8989 11452 9053 11456
rect 8989 11396 8993 11452
rect 8993 11396 9049 11452
rect 9049 11396 9053 11452
rect 8989 11392 9053 11396
rect 13947 11452 14011 11456
rect 13947 11396 13951 11452
rect 13951 11396 14007 11452
rect 14007 11396 14011 11452
rect 13947 11392 14011 11396
rect 14027 11452 14091 11456
rect 14027 11396 14031 11452
rect 14031 11396 14087 11452
rect 14087 11396 14091 11452
rect 14027 11392 14091 11396
rect 14107 11452 14171 11456
rect 14107 11396 14111 11452
rect 14111 11396 14167 11452
rect 14167 11396 14171 11452
rect 14107 11392 14171 11396
rect 14187 11452 14251 11456
rect 14187 11396 14191 11452
rect 14191 11396 14247 11452
rect 14247 11396 14251 11452
rect 14187 11392 14251 11396
rect 19145 11452 19209 11456
rect 19145 11396 19149 11452
rect 19149 11396 19205 11452
rect 19205 11396 19209 11452
rect 19145 11392 19209 11396
rect 19225 11452 19289 11456
rect 19225 11396 19229 11452
rect 19229 11396 19285 11452
rect 19285 11396 19289 11452
rect 19225 11392 19289 11396
rect 19305 11452 19369 11456
rect 19305 11396 19309 11452
rect 19309 11396 19365 11452
rect 19365 11396 19369 11452
rect 19305 11392 19369 11396
rect 19385 11452 19449 11456
rect 19385 11396 19389 11452
rect 19389 11396 19445 11452
rect 19445 11396 19449 11452
rect 19385 11392 19449 11396
rect 4108 11324 4172 11388
rect 2820 11188 2884 11252
rect 16068 11324 16132 11388
rect 2268 11112 2332 11116
rect 2268 11056 2282 11112
rect 2282 11056 2332 11112
rect 2268 11052 2332 11056
rect 3188 10780 3252 10844
rect 4476 10916 4540 10980
rect 5396 10916 5460 10980
rect 5396 10780 5460 10844
rect 6868 10916 6932 10980
rect 10916 10976 10980 10980
rect 10916 10920 10966 10976
rect 10966 10920 10980 10976
rect 10916 10916 10980 10920
rect 16252 10916 16316 10980
rect 6150 10908 6214 10912
rect 6150 10852 6154 10908
rect 6154 10852 6210 10908
rect 6210 10852 6214 10908
rect 6150 10848 6214 10852
rect 6230 10908 6294 10912
rect 6230 10852 6234 10908
rect 6234 10852 6290 10908
rect 6290 10852 6294 10908
rect 6230 10848 6294 10852
rect 6310 10908 6374 10912
rect 6310 10852 6314 10908
rect 6314 10852 6370 10908
rect 6370 10852 6374 10908
rect 6310 10848 6374 10852
rect 6390 10908 6454 10912
rect 6390 10852 6394 10908
rect 6394 10852 6450 10908
rect 6450 10852 6454 10908
rect 6390 10848 6454 10852
rect 11348 10908 11412 10912
rect 11348 10852 11352 10908
rect 11352 10852 11408 10908
rect 11408 10852 11412 10908
rect 11348 10848 11412 10852
rect 11428 10908 11492 10912
rect 11428 10852 11432 10908
rect 11432 10852 11488 10908
rect 11488 10852 11492 10908
rect 11428 10848 11492 10852
rect 11508 10908 11572 10912
rect 11508 10852 11512 10908
rect 11512 10852 11568 10908
rect 11568 10852 11572 10908
rect 11508 10848 11572 10852
rect 11588 10908 11652 10912
rect 11588 10852 11592 10908
rect 11592 10852 11648 10908
rect 11648 10852 11652 10908
rect 11588 10848 11652 10852
rect 16546 10908 16610 10912
rect 16546 10852 16550 10908
rect 16550 10852 16606 10908
rect 16606 10852 16610 10908
rect 16546 10848 16610 10852
rect 16626 10908 16690 10912
rect 16626 10852 16630 10908
rect 16630 10852 16686 10908
rect 16686 10852 16690 10908
rect 16626 10848 16690 10852
rect 16706 10908 16770 10912
rect 16706 10852 16710 10908
rect 16710 10852 16766 10908
rect 16766 10852 16770 10908
rect 16706 10848 16770 10852
rect 16786 10908 16850 10912
rect 16786 10852 16790 10908
rect 16790 10852 16846 10908
rect 16846 10852 16850 10908
rect 16786 10848 16850 10852
rect 21744 10908 21808 10912
rect 21744 10852 21748 10908
rect 21748 10852 21804 10908
rect 21804 10852 21808 10908
rect 21744 10848 21808 10852
rect 21824 10908 21888 10912
rect 21824 10852 21828 10908
rect 21828 10852 21884 10908
rect 21884 10852 21888 10908
rect 21824 10848 21888 10852
rect 21904 10908 21968 10912
rect 21904 10852 21908 10908
rect 21908 10852 21964 10908
rect 21964 10852 21968 10908
rect 21904 10848 21968 10852
rect 21984 10908 22048 10912
rect 21984 10852 21988 10908
rect 21988 10852 22044 10908
rect 22044 10852 22048 10908
rect 21984 10848 22048 10852
rect 8156 10780 8220 10844
rect 3004 10508 3068 10572
rect 10732 10568 10796 10572
rect 10732 10512 10782 10568
rect 10782 10512 10796 10568
rect 10732 10508 10796 10512
rect 13308 10508 13372 10572
rect 20300 10508 20364 10572
rect 12204 10372 12268 10436
rect 3551 10364 3615 10368
rect 3551 10308 3555 10364
rect 3555 10308 3611 10364
rect 3611 10308 3615 10364
rect 3551 10304 3615 10308
rect 3631 10364 3695 10368
rect 3631 10308 3635 10364
rect 3635 10308 3691 10364
rect 3691 10308 3695 10364
rect 3631 10304 3695 10308
rect 3711 10364 3775 10368
rect 3711 10308 3715 10364
rect 3715 10308 3771 10364
rect 3771 10308 3775 10364
rect 3711 10304 3775 10308
rect 3791 10364 3855 10368
rect 3791 10308 3795 10364
rect 3795 10308 3851 10364
rect 3851 10308 3855 10364
rect 3791 10304 3855 10308
rect 8749 10364 8813 10368
rect 8749 10308 8753 10364
rect 8753 10308 8809 10364
rect 8809 10308 8813 10364
rect 8749 10304 8813 10308
rect 8829 10364 8893 10368
rect 8829 10308 8833 10364
rect 8833 10308 8889 10364
rect 8889 10308 8893 10364
rect 8829 10304 8893 10308
rect 8909 10364 8973 10368
rect 8909 10308 8913 10364
rect 8913 10308 8969 10364
rect 8969 10308 8973 10364
rect 8909 10304 8973 10308
rect 8989 10364 9053 10368
rect 8989 10308 8993 10364
rect 8993 10308 9049 10364
rect 9049 10308 9053 10364
rect 8989 10304 9053 10308
rect 13947 10364 14011 10368
rect 13947 10308 13951 10364
rect 13951 10308 14007 10364
rect 14007 10308 14011 10364
rect 13947 10304 14011 10308
rect 14027 10364 14091 10368
rect 14027 10308 14031 10364
rect 14031 10308 14087 10364
rect 14087 10308 14091 10364
rect 14027 10304 14091 10308
rect 14107 10364 14171 10368
rect 14107 10308 14111 10364
rect 14111 10308 14167 10364
rect 14167 10308 14171 10364
rect 14107 10304 14171 10308
rect 14187 10364 14251 10368
rect 14187 10308 14191 10364
rect 14191 10308 14247 10364
rect 14247 10308 14251 10364
rect 14187 10304 14251 10308
rect 19145 10364 19209 10368
rect 19145 10308 19149 10364
rect 19149 10308 19205 10364
rect 19205 10308 19209 10364
rect 19145 10304 19209 10308
rect 19225 10364 19289 10368
rect 19225 10308 19229 10364
rect 19229 10308 19285 10364
rect 19285 10308 19289 10364
rect 19225 10304 19289 10308
rect 19305 10364 19369 10368
rect 19305 10308 19309 10364
rect 19309 10308 19365 10364
rect 19365 10308 19369 10364
rect 19305 10304 19369 10308
rect 19385 10364 19449 10368
rect 19385 10308 19389 10364
rect 19389 10308 19445 10364
rect 19445 10308 19449 10364
rect 19385 10304 19449 10308
rect 5396 10236 5460 10300
rect 5028 9888 5092 9892
rect 5028 9832 5078 9888
rect 5078 9832 5092 9888
rect 5028 9828 5092 9832
rect 6150 9820 6214 9824
rect 6150 9764 6154 9820
rect 6154 9764 6210 9820
rect 6210 9764 6214 9820
rect 6150 9760 6214 9764
rect 6230 9820 6294 9824
rect 6230 9764 6234 9820
rect 6234 9764 6290 9820
rect 6290 9764 6294 9820
rect 6230 9760 6294 9764
rect 6310 9820 6374 9824
rect 6310 9764 6314 9820
rect 6314 9764 6370 9820
rect 6370 9764 6374 9820
rect 6310 9760 6374 9764
rect 6390 9820 6454 9824
rect 6390 9764 6394 9820
rect 6394 9764 6450 9820
rect 6450 9764 6454 9820
rect 6390 9760 6454 9764
rect 11348 9820 11412 9824
rect 11348 9764 11352 9820
rect 11352 9764 11408 9820
rect 11408 9764 11412 9820
rect 11348 9760 11412 9764
rect 11428 9820 11492 9824
rect 11428 9764 11432 9820
rect 11432 9764 11488 9820
rect 11488 9764 11492 9820
rect 11428 9760 11492 9764
rect 11508 9820 11572 9824
rect 11508 9764 11512 9820
rect 11512 9764 11568 9820
rect 11568 9764 11572 9820
rect 11508 9760 11572 9764
rect 11588 9820 11652 9824
rect 11588 9764 11592 9820
rect 11592 9764 11648 9820
rect 11648 9764 11652 9820
rect 11588 9760 11652 9764
rect 13492 9964 13556 10028
rect 13676 9964 13740 10028
rect 8340 9692 8404 9756
rect 16546 9820 16610 9824
rect 16546 9764 16550 9820
rect 16550 9764 16606 9820
rect 16606 9764 16610 9820
rect 16546 9760 16610 9764
rect 16626 9820 16690 9824
rect 16626 9764 16630 9820
rect 16630 9764 16686 9820
rect 16686 9764 16690 9820
rect 16626 9760 16690 9764
rect 16706 9820 16770 9824
rect 16706 9764 16710 9820
rect 16710 9764 16766 9820
rect 16766 9764 16770 9820
rect 16706 9760 16770 9764
rect 16786 9820 16850 9824
rect 16786 9764 16790 9820
rect 16790 9764 16846 9820
rect 16846 9764 16850 9820
rect 16786 9760 16850 9764
rect 21744 9820 21808 9824
rect 21744 9764 21748 9820
rect 21748 9764 21804 9820
rect 21804 9764 21808 9820
rect 21744 9760 21808 9764
rect 21824 9820 21888 9824
rect 21824 9764 21828 9820
rect 21828 9764 21884 9820
rect 21884 9764 21888 9820
rect 21824 9760 21888 9764
rect 21904 9820 21968 9824
rect 21904 9764 21908 9820
rect 21908 9764 21964 9820
rect 21964 9764 21968 9820
rect 21904 9760 21968 9764
rect 21984 9820 22048 9824
rect 21984 9764 21988 9820
rect 21988 9764 22044 9820
rect 22044 9764 22048 9820
rect 21984 9760 22048 9764
rect 14780 9692 14844 9756
rect 19932 9692 19996 9756
rect 16988 9556 17052 9620
rect 19012 9556 19076 9620
rect 17172 9420 17236 9484
rect 2636 9284 2700 9348
rect 20484 9420 20548 9484
rect 3551 9276 3615 9280
rect 3551 9220 3555 9276
rect 3555 9220 3611 9276
rect 3611 9220 3615 9276
rect 3551 9216 3615 9220
rect 3631 9276 3695 9280
rect 3631 9220 3635 9276
rect 3635 9220 3691 9276
rect 3691 9220 3695 9276
rect 3631 9216 3695 9220
rect 3711 9276 3775 9280
rect 3711 9220 3715 9276
rect 3715 9220 3771 9276
rect 3771 9220 3775 9276
rect 3711 9216 3775 9220
rect 3791 9276 3855 9280
rect 3791 9220 3795 9276
rect 3795 9220 3851 9276
rect 3851 9220 3855 9276
rect 3791 9216 3855 9220
rect 8749 9276 8813 9280
rect 8749 9220 8753 9276
rect 8753 9220 8809 9276
rect 8809 9220 8813 9276
rect 8749 9216 8813 9220
rect 8829 9276 8893 9280
rect 8829 9220 8833 9276
rect 8833 9220 8889 9276
rect 8889 9220 8893 9276
rect 8829 9216 8893 9220
rect 8909 9276 8973 9280
rect 8909 9220 8913 9276
rect 8913 9220 8969 9276
rect 8969 9220 8973 9276
rect 8909 9216 8973 9220
rect 8989 9276 9053 9280
rect 8989 9220 8993 9276
rect 8993 9220 9049 9276
rect 9049 9220 9053 9276
rect 8989 9216 9053 9220
rect 13947 9276 14011 9280
rect 13947 9220 13951 9276
rect 13951 9220 14007 9276
rect 14007 9220 14011 9276
rect 13947 9216 14011 9220
rect 14027 9276 14091 9280
rect 14027 9220 14031 9276
rect 14031 9220 14087 9276
rect 14087 9220 14091 9276
rect 14027 9216 14091 9220
rect 14107 9276 14171 9280
rect 14107 9220 14111 9276
rect 14111 9220 14167 9276
rect 14167 9220 14171 9276
rect 14107 9216 14171 9220
rect 14187 9276 14251 9280
rect 14187 9220 14191 9276
rect 14191 9220 14247 9276
rect 14247 9220 14251 9276
rect 14187 9216 14251 9220
rect 19145 9276 19209 9280
rect 19145 9220 19149 9276
rect 19149 9220 19205 9276
rect 19205 9220 19209 9276
rect 19145 9216 19209 9220
rect 19225 9276 19289 9280
rect 19225 9220 19229 9276
rect 19229 9220 19285 9276
rect 19285 9220 19289 9276
rect 19225 9216 19289 9220
rect 19305 9276 19369 9280
rect 19305 9220 19309 9276
rect 19309 9220 19365 9276
rect 19365 9220 19369 9276
rect 19305 9216 19369 9220
rect 19385 9276 19449 9280
rect 19385 9220 19389 9276
rect 19389 9220 19445 9276
rect 19445 9220 19449 9276
rect 19385 9216 19449 9220
rect 4292 9148 4356 9212
rect 5764 9012 5828 9076
rect 16252 9012 16316 9076
rect 2452 8740 2516 8804
rect 2268 8604 2332 8668
rect 12204 8740 12268 8804
rect 12940 8740 13004 8804
rect 6150 8732 6214 8736
rect 6150 8676 6154 8732
rect 6154 8676 6210 8732
rect 6210 8676 6214 8732
rect 6150 8672 6214 8676
rect 6230 8732 6294 8736
rect 6230 8676 6234 8732
rect 6234 8676 6290 8732
rect 6290 8676 6294 8732
rect 6230 8672 6294 8676
rect 6310 8732 6374 8736
rect 6310 8676 6314 8732
rect 6314 8676 6370 8732
rect 6370 8676 6374 8732
rect 6310 8672 6374 8676
rect 6390 8732 6454 8736
rect 6390 8676 6394 8732
rect 6394 8676 6450 8732
rect 6450 8676 6454 8732
rect 6390 8672 6454 8676
rect 11348 8732 11412 8736
rect 11348 8676 11352 8732
rect 11352 8676 11408 8732
rect 11408 8676 11412 8732
rect 11348 8672 11412 8676
rect 11428 8732 11492 8736
rect 11428 8676 11432 8732
rect 11432 8676 11488 8732
rect 11488 8676 11492 8732
rect 11428 8672 11492 8676
rect 11508 8732 11572 8736
rect 11508 8676 11512 8732
rect 11512 8676 11568 8732
rect 11568 8676 11572 8732
rect 11508 8672 11572 8676
rect 11588 8732 11652 8736
rect 11588 8676 11592 8732
rect 11592 8676 11648 8732
rect 11648 8676 11652 8732
rect 11588 8672 11652 8676
rect 3372 8604 3436 8668
rect 4476 8604 4540 8668
rect 6868 8604 6932 8668
rect 16546 8732 16610 8736
rect 16546 8676 16550 8732
rect 16550 8676 16606 8732
rect 16606 8676 16610 8732
rect 16546 8672 16610 8676
rect 16626 8732 16690 8736
rect 16626 8676 16630 8732
rect 16630 8676 16686 8732
rect 16686 8676 16690 8732
rect 16626 8672 16690 8676
rect 16706 8732 16770 8736
rect 16706 8676 16710 8732
rect 16710 8676 16766 8732
rect 16766 8676 16770 8732
rect 16706 8672 16770 8676
rect 16786 8732 16850 8736
rect 16786 8676 16790 8732
rect 16790 8676 16846 8732
rect 16846 8676 16850 8732
rect 16786 8672 16850 8676
rect 21744 8732 21808 8736
rect 21744 8676 21748 8732
rect 21748 8676 21804 8732
rect 21804 8676 21808 8732
rect 21744 8672 21808 8676
rect 21824 8732 21888 8736
rect 21824 8676 21828 8732
rect 21828 8676 21884 8732
rect 21884 8676 21888 8732
rect 21824 8672 21888 8676
rect 21904 8732 21968 8736
rect 21904 8676 21908 8732
rect 21908 8676 21964 8732
rect 21964 8676 21968 8732
rect 21904 8672 21968 8676
rect 21984 8732 22048 8736
rect 21984 8676 21988 8732
rect 21988 8676 22044 8732
rect 22044 8676 22048 8732
rect 21984 8672 22048 8676
rect 5028 8468 5092 8532
rect 9628 8468 9692 8532
rect 3188 8332 3252 8396
rect 3372 8332 3436 8396
rect 8340 8332 8404 8396
rect 9444 8332 9508 8396
rect 12940 8332 13004 8396
rect 13124 8332 13188 8396
rect 17540 8332 17604 8396
rect 2452 8196 2516 8260
rect 3551 8188 3615 8192
rect 3551 8132 3555 8188
rect 3555 8132 3611 8188
rect 3611 8132 3615 8188
rect 3551 8128 3615 8132
rect 3631 8188 3695 8192
rect 3631 8132 3635 8188
rect 3635 8132 3691 8188
rect 3691 8132 3695 8188
rect 3631 8128 3695 8132
rect 3711 8188 3775 8192
rect 3711 8132 3715 8188
rect 3715 8132 3771 8188
rect 3771 8132 3775 8188
rect 3711 8128 3775 8132
rect 3791 8188 3855 8192
rect 3791 8132 3795 8188
rect 3795 8132 3851 8188
rect 3851 8132 3855 8188
rect 3791 8128 3855 8132
rect 5212 8196 5276 8260
rect 8749 8188 8813 8192
rect 8749 8132 8753 8188
rect 8753 8132 8809 8188
rect 8809 8132 8813 8188
rect 8749 8128 8813 8132
rect 8829 8188 8893 8192
rect 8829 8132 8833 8188
rect 8833 8132 8889 8188
rect 8889 8132 8893 8188
rect 8829 8128 8893 8132
rect 8909 8188 8973 8192
rect 8909 8132 8913 8188
rect 8913 8132 8969 8188
rect 8969 8132 8973 8188
rect 8909 8128 8973 8132
rect 8989 8188 9053 8192
rect 8989 8132 8993 8188
rect 8993 8132 9049 8188
rect 9049 8132 9053 8188
rect 8989 8128 9053 8132
rect 10180 7924 10244 7988
rect 12204 7924 12268 7988
rect 3188 7848 3252 7852
rect 3188 7792 3238 7848
rect 3238 7792 3252 7848
rect 3188 7788 3252 7792
rect 13947 8188 14011 8192
rect 13947 8132 13951 8188
rect 13951 8132 14007 8188
rect 14007 8132 14011 8188
rect 13947 8128 14011 8132
rect 14027 8188 14091 8192
rect 14027 8132 14031 8188
rect 14031 8132 14087 8188
rect 14087 8132 14091 8188
rect 14027 8128 14091 8132
rect 14107 8188 14171 8192
rect 14107 8132 14111 8188
rect 14111 8132 14167 8188
rect 14167 8132 14171 8188
rect 14107 8128 14171 8132
rect 14187 8188 14251 8192
rect 14187 8132 14191 8188
rect 14191 8132 14247 8188
rect 14247 8132 14251 8188
rect 14187 8128 14251 8132
rect 19145 8188 19209 8192
rect 19145 8132 19149 8188
rect 19149 8132 19205 8188
rect 19205 8132 19209 8188
rect 19145 8128 19209 8132
rect 19225 8188 19289 8192
rect 19225 8132 19229 8188
rect 19229 8132 19285 8188
rect 19285 8132 19289 8188
rect 19225 8128 19289 8132
rect 19305 8188 19369 8192
rect 19305 8132 19309 8188
rect 19309 8132 19365 8188
rect 19365 8132 19369 8188
rect 19305 8128 19369 8132
rect 19385 8188 19449 8192
rect 19385 8132 19389 8188
rect 19389 8132 19445 8188
rect 19445 8132 19449 8188
rect 19385 8128 19449 8132
rect 2084 7516 2148 7580
rect 18828 7712 18892 7716
rect 18828 7656 18842 7712
rect 18842 7656 18892 7712
rect 18828 7652 18892 7656
rect 6150 7644 6214 7648
rect 6150 7588 6154 7644
rect 6154 7588 6210 7644
rect 6210 7588 6214 7644
rect 6150 7584 6214 7588
rect 6230 7644 6294 7648
rect 6230 7588 6234 7644
rect 6234 7588 6290 7644
rect 6290 7588 6294 7644
rect 6230 7584 6294 7588
rect 6310 7644 6374 7648
rect 6310 7588 6314 7644
rect 6314 7588 6370 7644
rect 6370 7588 6374 7644
rect 6310 7584 6374 7588
rect 6390 7644 6454 7648
rect 6390 7588 6394 7644
rect 6394 7588 6450 7644
rect 6450 7588 6454 7644
rect 6390 7584 6454 7588
rect 11348 7644 11412 7648
rect 11348 7588 11352 7644
rect 11352 7588 11408 7644
rect 11408 7588 11412 7644
rect 11348 7584 11412 7588
rect 11428 7644 11492 7648
rect 11428 7588 11432 7644
rect 11432 7588 11488 7644
rect 11488 7588 11492 7644
rect 11428 7584 11492 7588
rect 11508 7644 11572 7648
rect 11508 7588 11512 7644
rect 11512 7588 11568 7644
rect 11568 7588 11572 7644
rect 11508 7584 11572 7588
rect 11588 7644 11652 7648
rect 11588 7588 11592 7644
rect 11592 7588 11648 7644
rect 11648 7588 11652 7644
rect 11588 7584 11652 7588
rect 16546 7644 16610 7648
rect 16546 7588 16550 7644
rect 16550 7588 16606 7644
rect 16606 7588 16610 7644
rect 16546 7584 16610 7588
rect 16626 7644 16690 7648
rect 16626 7588 16630 7644
rect 16630 7588 16686 7644
rect 16686 7588 16690 7644
rect 16626 7584 16690 7588
rect 16706 7644 16770 7648
rect 16706 7588 16710 7644
rect 16710 7588 16766 7644
rect 16766 7588 16770 7644
rect 16706 7584 16770 7588
rect 16786 7644 16850 7648
rect 16786 7588 16790 7644
rect 16790 7588 16846 7644
rect 16846 7588 16850 7644
rect 16786 7584 16850 7588
rect 21744 7644 21808 7648
rect 21744 7588 21748 7644
rect 21748 7588 21804 7644
rect 21804 7588 21808 7644
rect 21744 7584 21808 7588
rect 21824 7644 21888 7648
rect 21824 7588 21828 7644
rect 21828 7588 21884 7644
rect 21884 7588 21888 7644
rect 21824 7584 21888 7588
rect 21904 7644 21968 7648
rect 21904 7588 21908 7644
rect 21908 7588 21964 7644
rect 21964 7588 21968 7644
rect 21904 7584 21968 7588
rect 21984 7644 22048 7648
rect 21984 7588 21988 7644
rect 21988 7588 22044 7644
rect 22044 7588 22048 7644
rect 21984 7584 22048 7588
rect 4476 7516 4540 7580
rect 5580 7516 5644 7580
rect 5764 7516 5828 7580
rect 13308 7516 13372 7580
rect 1900 7244 1964 7308
rect 11100 7244 11164 7308
rect 2268 7168 2332 7172
rect 2268 7112 2282 7168
rect 2282 7112 2332 7168
rect 2268 7108 2332 7112
rect 3551 7100 3615 7104
rect 3551 7044 3555 7100
rect 3555 7044 3611 7100
rect 3611 7044 3615 7100
rect 3551 7040 3615 7044
rect 3631 7100 3695 7104
rect 3631 7044 3635 7100
rect 3635 7044 3691 7100
rect 3691 7044 3695 7100
rect 3631 7040 3695 7044
rect 3711 7100 3775 7104
rect 3711 7044 3715 7100
rect 3715 7044 3771 7100
rect 3771 7044 3775 7100
rect 3711 7040 3775 7044
rect 3791 7100 3855 7104
rect 3791 7044 3795 7100
rect 3795 7044 3851 7100
rect 3851 7044 3855 7100
rect 3791 7040 3855 7044
rect 8749 7100 8813 7104
rect 8749 7044 8753 7100
rect 8753 7044 8809 7100
rect 8809 7044 8813 7100
rect 8749 7040 8813 7044
rect 8829 7100 8893 7104
rect 8829 7044 8833 7100
rect 8833 7044 8889 7100
rect 8889 7044 8893 7100
rect 8829 7040 8893 7044
rect 8909 7100 8973 7104
rect 8909 7044 8913 7100
rect 8913 7044 8969 7100
rect 8969 7044 8973 7100
rect 8909 7040 8973 7044
rect 8989 7100 9053 7104
rect 8989 7044 8993 7100
rect 8993 7044 9049 7100
rect 9049 7044 9053 7100
rect 8989 7040 9053 7044
rect 13947 7100 14011 7104
rect 13947 7044 13951 7100
rect 13951 7044 14007 7100
rect 14007 7044 14011 7100
rect 13947 7040 14011 7044
rect 14027 7100 14091 7104
rect 14027 7044 14031 7100
rect 14031 7044 14087 7100
rect 14087 7044 14091 7100
rect 14027 7040 14091 7044
rect 14107 7100 14171 7104
rect 14107 7044 14111 7100
rect 14111 7044 14167 7100
rect 14167 7044 14171 7100
rect 14107 7040 14171 7044
rect 14187 7100 14251 7104
rect 14187 7044 14191 7100
rect 14191 7044 14247 7100
rect 14247 7044 14251 7100
rect 14187 7040 14251 7044
rect 4292 6972 4356 7036
rect 4660 6972 4724 7036
rect 5212 6836 5276 6900
rect 7052 6972 7116 7036
rect 19145 7100 19209 7104
rect 19145 7044 19149 7100
rect 19149 7044 19205 7100
rect 19205 7044 19209 7100
rect 19145 7040 19209 7044
rect 19225 7100 19289 7104
rect 19225 7044 19229 7100
rect 19229 7044 19285 7100
rect 19285 7044 19289 7100
rect 19225 7040 19289 7044
rect 19305 7100 19369 7104
rect 19305 7044 19309 7100
rect 19309 7044 19365 7100
rect 19365 7044 19369 7100
rect 19305 7040 19369 7044
rect 19385 7100 19449 7104
rect 19385 7044 19389 7100
rect 19389 7044 19445 7100
rect 19445 7044 19449 7100
rect 19385 7040 19449 7044
rect 5764 6836 5828 6900
rect 7604 6836 7668 6900
rect 12756 6836 12820 6900
rect 14412 6836 14476 6900
rect 2820 6700 2884 6764
rect 3004 6700 3068 6764
rect 3924 6700 3988 6764
rect 2636 6564 2700 6628
rect 4476 6564 4540 6628
rect 10364 6564 10428 6628
rect 6150 6556 6214 6560
rect 6150 6500 6154 6556
rect 6154 6500 6210 6556
rect 6210 6500 6214 6556
rect 6150 6496 6214 6500
rect 6230 6556 6294 6560
rect 6230 6500 6234 6556
rect 6234 6500 6290 6556
rect 6290 6500 6294 6556
rect 6230 6496 6294 6500
rect 6310 6556 6374 6560
rect 6310 6500 6314 6556
rect 6314 6500 6370 6556
rect 6370 6500 6374 6556
rect 6310 6496 6374 6500
rect 6390 6556 6454 6560
rect 6390 6500 6394 6556
rect 6394 6500 6450 6556
rect 6450 6500 6454 6556
rect 6390 6496 6454 6500
rect 11348 6556 11412 6560
rect 11348 6500 11352 6556
rect 11352 6500 11408 6556
rect 11408 6500 11412 6556
rect 11348 6496 11412 6500
rect 11428 6556 11492 6560
rect 11428 6500 11432 6556
rect 11432 6500 11488 6556
rect 11488 6500 11492 6556
rect 11428 6496 11492 6500
rect 11508 6556 11572 6560
rect 11508 6500 11512 6556
rect 11512 6500 11568 6556
rect 11568 6500 11572 6556
rect 11508 6496 11572 6500
rect 11588 6556 11652 6560
rect 11588 6500 11592 6556
rect 11592 6500 11648 6556
rect 11648 6500 11652 6556
rect 11588 6496 11652 6500
rect 5396 6292 5460 6356
rect 16546 6556 16610 6560
rect 16546 6500 16550 6556
rect 16550 6500 16606 6556
rect 16606 6500 16610 6556
rect 16546 6496 16610 6500
rect 16626 6556 16690 6560
rect 16626 6500 16630 6556
rect 16630 6500 16686 6556
rect 16686 6500 16690 6556
rect 16626 6496 16690 6500
rect 16706 6556 16770 6560
rect 16706 6500 16710 6556
rect 16710 6500 16766 6556
rect 16766 6500 16770 6556
rect 16706 6496 16770 6500
rect 16786 6556 16850 6560
rect 16786 6500 16790 6556
rect 16790 6500 16846 6556
rect 16846 6500 16850 6556
rect 16786 6496 16850 6500
rect 21744 6556 21808 6560
rect 21744 6500 21748 6556
rect 21748 6500 21804 6556
rect 21804 6500 21808 6556
rect 21744 6496 21808 6500
rect 21824 6556 21888 6560
rect 21824 6500 21828 6556
rect 21828 6500 21884 6556
rect 21884 6500 21888 6556
rect 21824 6496 21888 6500
rect 21904 6556 21968 6560
rect 21904 6500 21908 6556
rect 21908 6500 21964 6556
rect 21964 6500 21968 6556
rect 21904 6496 21968 6500
rect 21984 6556 22048 6560
rect 21984 6500 21988 6556
rect 21988 6500 22044 6556
rect 22044 6500 22048 6556
rect 21984 6496 22048 6500
rect 15148 6292 15212 6356
rect 2820 6020 2884 6084
rect 10180 6156 10244 6220
rect 18092 6156 18156 6220
rect 3551 6012 3615 6016
rect 3551 5956 3555 6012
rect 3555 5956 3611 6012
rect 3611 5956 3615 6012
rect 3551 5952 3615 5956
rect 3631 6012 3695 6016
rect 3631 5956 3635 6012
rect 3635 5956 3691 6012
rect 3691 5956 3695 6012
rect 3631 5952 3695 5956
rect 3711 6012 3775 6016
rect 3711 5956 3715 6012
rect 3715 5956 3771 6012
rect 3771 5956 3775 6012
rect 3711 5952 3775 5956
rect 3791 6012 3855 6016
rect 3791 5956 3795 6012
rect 3795 5956 3851 6012
rect 3851 5956 3855 6012
rect 3791 5952 3855 5956
rect 8749 6012 8813 6016
rect 8749 5956 8753 6012
rect 8753 5956 8809 6012
rect 8809 5956 8813 6012
rect 8749 5952 8813 5956
rect 8829 6012 8893 6016
rect 8829 5956 8833 6012
rect 8833 5956 8889 6012
rect 8889 5956 8893 6012
rect 8829 5952 8893 5956
rect 8909 6012 8973 6016
rect 8909 5956 8913 6012
rect 8913 5956 8969 6012
rect 8969 5956 8973 6012
rect 8909 5952 8973 5956
rect 8989 6012 9053 6016
rect 8989 5956 8993 6012
rect 8993 5956 9049 6012
rect 9049 5956 9053 6012
rect 8989 5952 9053 5956
rect 13947 6012 14011 6016
rect 13947 5956 13951 6012
rect 13951 5956 14007 6012
rect 14007 5956 14011 6012
rect 13947 5952 14011 5956
rect 14027 6012 14091 6016
rect 14027 5956 14031 6012
rect 14031 5956 14087 6012
rect 14087 5956 14091 6012
rect 14027 5952 14091 5956
rect 14107 6012 14171 6016
rect 14107 5956 14111 6012
rect 14111 5956 14167 6012
rect 14167 5956 14171 6012
rect 14107 5952 14171 5956
rect 14187 6012 14251 6016
rect 14187 5956 14191 6012
rect 14191 5956 14247 6012
rect 14247 5956 14251 6012
rect 14187 5952 14251 5956
rect 19145 6012 19209 6016
rect 19145 5956 19149 6012
rect 19149 5956 19205 6012
rect 19205 5956 19209 6012
rect 19145 5952 19209 5956
rect 19225 6012 19289 6016
rect 19225 5956 19229 6012
rect 19229 5956 19285 6012
rect 19285 5956 19289 6012
rect 19225 5952 19289 5956
rect 19305 6012 19369 6016
rect 19305 5956 19309 6012
rect 19309 5956 19365 6012
rect 19365 5956 19369 6012
rect 19305 5952 19369 5956
rect 19385 6012 19449 6016
rect 19385 5956 19389 6012
rect 19389 5956 19445 6012
rect 19445 5956 19449 6012
rect 19385 5952 19449 5956
rect 4476 5748 4540 5812
rect 9628 5612 9692 5676
rect 19012 5612 19076 5676
rect 18460 5536 18524 5540
rect 18460 5480 18474 5536
rect 18474 5480 18524 5536
rect 18460 5476 18524 5480
rect 6150 5468 6214 5472
rect 6150 5412 6154 5468
rect 6154 5412 6210 5468
rect 6210 5412 6214 5468
rect 6150 5408 6214 5412
rect 6230 5468 6294 5472
rect 6230 5412 6234 5468
rect 6234 5412 6290 5468
rect 6290 5412 6294 5468
rect 6230 5408 6294 5412
rect 6310 5468 6374 5472
rect 6310 5412 6314 5468
rect 6314 5412 6370 5468
rect 6370 5412 6374 5468
rect 6310 5408 6374 5412
rect 6390 5468 6454 5472
rect 6390 5412 6394 5468
rect 6394 5412 6450 5468
rect 6450 5412 6454 5468
rect 6390 5408 6454 5412
rect 11348 5468 11412 5472
rect 11348 5412 11352 5468
rect 11352 5412 11408 5468
rect 11408 5412 11412 5468
rect 11348 5408 11412 5412
rect 11428 5468 11492 5472
rect 11428 5412 11432 5468
rect 11432 5412 11488 5468
rect 11488 5412 11492 5468
rect 11428 5408 11492 5412
rect 11508 5468 11572 5472
rect 11508 5412 11512 5468
rect 11512 5412 11568 5468
rect 11568 5412 11572 5468
rect 11508 5408 11572 5412
rect 11588 5468 11652 5472
rect 11588 5412 11592 5468
rect 11592 5412 11648 5468
rect 11648 5412 11652 5468
rect 11588 5408 11652 5412
rect 16546 5468 16610 5472
rect 16546 5412 16550 5468
rect 16550 5412 16606 5468
rect 16606 5412 16610 5468
rect 16546 5408 16610 5412
rect 16626 5468 16690 5472
rect 16626 5412 16630 5468
rect 16630 5412 16686 5468
rect 16686 5412 16690 5468
rect 16626 5408 16690 5412
rect 16706 5468 16770 5472
rect 16706 5412 16710 5468
rect 16710 5412 16766 5468
rect 16766 5412 16770 5468
rect 16706 5408 16770 5412
rect 16786 5468 16850 5472
rect 16786 5412 16790 5468
rect 16790 5412 16846 5468
rect 16846 5412 16850 5468
rect 16786 5408 16850 5412
rect 3372 5340 3436 5404
rect 17724 5340 17788 5404
rect 21744 5468 21808 5472
rect 21744 5412 21748 5468
rect 21748 5412 21804 5468
rect 21804 5412 21808 5468
rect 21744 5408 21808 5412
rect 21824 5468 21888 5472
rect 21824 5412 21828 5468
rect 21828 5412 21884 5468
rect 21884 5412 21888 5468
rect 21824 5408 21888 5412
rect 21904 5468 21968 5472
rect 21904 5412 21908 5468
rect 21908 5412 21964 5468
rect 21964 5412 21968 5468
rect 21904 5408 21968 5412
rect 21984 5468 22048 5472
rect 21984 5412 21988 5468
rect 21988 5412 22044 5468
rect 22044 5412 22048 5468
rect 21984 5408 22048 5412
rect 5028 5068 5092 5132
rect 5212 5068 5276 5132
rect 3551 4924 3615 4928
rect 3551 4868 3555 4924
rect 3555 4868 3611 4924
rect 3611 4868 3615 4924
rect 3551 4864 3615 4868
rect 3631 4924 3695 4928
rect 3631 4868 3635 4924
rect 3635 4868 3691 4924
rect 3691 4868 3695 4924
rect 3631 4864 3695 4868
rect 3711 4924 3775 4928
rect 3711 4868 3715 4924
rect 3715 4868 3771 4924
rect 3771 4868 3775 4924
rect 3711 4864 3775 4868
rect 3791 4924 3855 4928
rect 3791 4868 3795 4924
rect 3795 4868 3851 4924
rect 3851 4868 3855 4924
rect 3791 4864 3855 4868
rect 8749 4924 8813 4928
rect 8749 4868 8753 4924
rect 8753 4868 8809 4924
rect 8809 4868 8813 4924
rect 8749 4864 8813 4868
rect 8829 4924 8893 4928
rect 8829 4868 8833 4924
rect 8833 4868 8889 4924
rect 8889 4868 8893 4924
rect 8829 4864 8893 4868
rect 8909 4924 8973 4928
rect 8909 4868 8913 4924
rect 8913 4868 8969 4924
rect 8969 4868 8973 4924
rect 8909 4864 8973 4868
rect 8989 4924 9053 4928
rect 8989 4868 8993 4924
rect 8993 4868 9049 4924
rect 9049 4868 9053 4924
rect 8989 4864 9053 4868
rect 13947 4924 14011 4928
rect 13947 4868 13951 4924
rect 13951 4868 14007 4924
rect 14007 4868 14011 4924
rect 13947 4864 14011 4868
rect 14027 4924 14091 4928
rect 14027 4868 14031 4924
rect 14031 4868 14087 4924
rect 14087 4868 14091 4924
rect 14027 4864 14091 4868
rect 14107 4924 14171 4928
rect 14107 4868 14111 4924
rect 14111 4868 14167 4924
rect 14167 4868 14171 4924
rect 14107 4864 14171 4868
rect 14187 4924 14251 4928
rect 14187 4868 14191 4924
rect 14191 4868 14247 4924
rect 14247 4868 14251 4924
rect 14187 4864 14251 4868
rect 19145 4924 19209 4928
rect 19145 4868 19149 4924
rect 19149 4868 19205 4924
rect 19205 4868 19209 4924
rect 19145 4864 19209 4868
rect 19225 4924 19289 4928
rect 19225 4868 19229 4924
rect 19229 4868 19285 4924
rect 19285 4868 19289 4924
rect 19225 4864 19289 4868
rect 19305 4924 19369 4928
rect 19305 4868 19309 4924
rect 19309 4868 19365 4924
rect 19365 4868 19369 4924
rect 19305 4864 19369 4868
rect 19385 4924 19449 4928
rect 19385 4868 19389 4924
rect 19389 4868 19445 4924
rect 19445 4868 19449 4924
rect 19385 4864 19449 4868
rect 2452 4524 2516 4588
rect 4108 4524 4172 4588
rect 4292 4584 4356 4588
rect 4292 4528 4342 4584
rect 4342 4528 4356 4584
rect 4292 4524 4356 4528
rect 4660 4388 4724 4452
rect 8156 4524 8220 4588
rect 12572 4524 12636 4588
rect 10548 4388 10612 4452
rect 18644 4388 18708 4452
rect 6150 4380 6214 4384
rect 6150 4324 6154 4380
rect 6154 4324 6210 4380
rect 6210 4324 6214 4380
rect 6150 4320 6214 4324
rect 6230 4380 6294 4384
rect 6230 4324 6234 4380
rect 6234 4324 6290 4380
rect 6290 4324 6294 4380
rect 6230 4320 6294 4324
rect 6310 4380 6374 4384
rect 6310 4324 6314 4380
rect 6314 4324 6370 4380
rect 6370 4324 6374 4380
rect 6310 4320 6374 4324
rect 6390 4380 6454 4384
rect 6390 4324 6394 4380
rect 6394 4324 6450 4380
rect 6450 4324 6454 4380
rect 6390 4320 6454 4324
rect 11348 4380 11412 4384
rect 11348 4324 11352 4380
rect 11352 4324 11408 4380
rect 11408 4324 11412 4380
rect 11348 4320 11412 4324
rect 11428 4380 11492 4384
rect 11428 4324 11432 4380
rect 11432 4324 11488 4380
rect 11488 4324 11492 4380
rect 11428 4320 11492 4324
rect 11508 4380 11572 4384
rect 11508 4324 11512 4380
rect 11512 4324 11568 4380
rect 11568 4324 11572 4380
rect 11508 4320 11572 4324
rect 11588 4380 11652 4384
rect 11588 4324 11592 4380
rect 11592 4324 11648 4380
rect 11648 4324 11652 4380
rect 11588 4320 11652 4324
rect 16546 4380 16610 4384
rect 16546 4324 16550 4380
rect 16550 4324 16606 4380
rect 16606 4324 16610 4380
rect 16546 4320 16610 4324
rect 16626 4380 16690 4384
rect 16626 4324 16630 4380
rect 16630 4324 16686 4380
rect 16686 4324 16690 4380
rect 16626 4320 16690 4324
rect 16706 4380 16770 4384
rect 16706 4324 16710 4380
rect 16710 4324 16766 4380
rect 16766 4324 16770 4380
rect 16706 4320 16770 4324
rect 16786 4380 16850 4384
rect 16786 4324 16790 4380
rect 16790 4324 16846 4380
rect 16846 4324 16850 4380
rect 16786 4320 16850 4324
rect 21744 4380 21808 4384
rect 21744 4324 21748 4380
rect 21748 4324 21804 4380
rect 21804 4324 21808 4380
rect 21744 4320 21808 4324
rect 21824 4380 21888 4384
rect 21824 4324 21828 4380
rect 21828 4324 21884 4380
rect 21884 4324 21888 4380
rect 21824 4320 21888 4324
rect 21904 4380 21968 4384
rect 21904 4324 21908 4380
rect 21908 4324 21964 4380
rect 21964 4324 21968 4380
rect 21904 4320 21968 4324
rect 21984 4380 22048 4384
rect 21984 4324 21988 4380
rect 21988 4324 22044 4380
rect 22044 4324 22048 4380
rect 21984 4320 22048 4324
rect 4108 4116 4172 4180
rect 14596 4252 14660 4316
rect 15700 4040 15764 4044
rect 15700 3984 15714 4040
rect 15714 3984 15764 4040
rect 15700 3980 15764 3984
rect 5580 3844 5644 3908
rect 18276 4040 18340 4044
rect 18276 3984 18290 4040
rect 18290 3984 18340 4040
rect 18276 3980 18340 3984
rect 20116 4040 20180 4044
rect 20116 3984 20130 4040
rect 20130 3984 20180 4040
rect 3551 3836 3615 3840
rect 3551 3780 3555 3836
rect 3555 3780 3611 3836
rect 3611 3780 3615 3836
rect 3551 3776 3615 3780
rect 3631 3836 3695 3840
rect 3631 3780 3635 3836
rect 3635 3780 3691 3836
rect 3691 3780 3695 3836
rect 3631 3776 3695 3780
rect 3711 3836 3775 3840
rect 3711 3780 3715 3836
rect 3715 3780 3771 3836
rect 3771 3780 3775 3836
rect 3711 3776 3775 3780
rect 3791 3836 3855 3840
rect 3791 3780 3795 3836
rect 3795 3780 3851 3836
rect 3851 3780 3855 3836
rect 3791 3776 3855 3780
rect 8749 3836 8813 3840
rect 8749 3780 8753 3836
rect 8753 3780 8809 3836
rect 8809 3780 8813 3836
rect 8749 3776 8813 3780
rect 8829 3836 8893 3840
rect 8829 3780 8833 3836
rect 8833 3780 8889 3836
rect 8889 3780 8893 3836
rect 8829 3776 8893 3780
rect 8909 3836 8973 3840
rect 8909 3780 8913 3836
rect 8913 3780 8969 3836
rect 8969 3780 8973 3836
rect 8909 3776 8973 3780
rect 8989 3836 9053 3840
rect 8989 3780 8993 3836
rect 8993 3780 9049 3836
rect 9049 3780 9053 3836
rect 8989 3776 9053 3780
rect 13947 3836 14011 3840
rect 13947 3780 13951 3836
rect 13951 3780 14007 3836
rect 14007 3780 14011 3836
rect 13947 3776 14011 3780
rect 14027 3836 14091 3840
rect 14027 3780 14031 3836
rect 14031 3780 14087 3836
rect 14087 3780 14091 3836
rect 14027 3776 14091 3780
rect 14107 3836 14171 3840
rect 14107 3780 14111 3836
rect 14111 3780 14167 3836
rect 14167 3780 14171 3836
rect 14107 3776 14171 3780
rect 14187 3836 14251 3840
rect 14187 3780 14191 3836
rect 14191 3780 14247 3836
rect 14247 3780 14251 3836
rect 14187 3776 14251 3780
rect 19145 3836 19209 3840
rect 19145 3780 19149 3836
rect 19149 3780 19205 3836
rect 19205 3780 19209 3836
rect 19145 3776 19209 3780
rect 19225 3836 19289 3840
rect 19225 3780 19229 3836
rect 19229 3780 19285 3836
rect 19285 3780 19289 3836
rect 19225 3776 19289 3780
rect 19305 3836 19369 3840
rect 19305 3780 19309 3836
rect 19309 3780 19365 3836
rect 19365 3780 19369 3836
rect 19305 3776 19369 3780
rect 19385 3836 19449 3840
rect 19385 3780 19389 3836
rect 19389 3780 19445 3836
rect 19445 3780 19449 3836
rect 19385 3776 19449 3780
rect 20116 3980 20180 3984
rect 7972 3572 8036 3636
rect 15148 3572 15212 3636
rect 15516 3632 15580 3636
rect 15516 3576 15530 3632
rect 15530 3576 15580 3632
rect 15516 3572 15580 3576
rect 16252 3360 16316 3364
rect 16252 3304 16302 3360
rect 16302 3304 16316 3360
rect 16252 3300 16316 3304
rect 17724 3300 17788 3364
rect 18092 3360 18156 3364
rect 18092 3304 18106 3360
rect 18106 3304 18156 3360
rect 18092 3300 18156 3304
rect 18828 3300 18892 3364
rect 6150 3292 6214 3296
rect 6150 3236 6154 3292
rect 6154 3236 6210 3292
rect 6210 3236 6214 3292
rect 6150 3232 6214 3236
rect 6230 3292 6294 3296
rect 6230 3236 6234 3292
rect 6234 3236 6290 3292
rect 6290 3236 6294 3292
rect 6230 3232 6294 3236
rect 6310 3292 6374 3296
rect 6310 3236 6314 3292
rect 6314 3236 6370 3292
rect 6370 3236 6374 3292
rect 6310 3232 6374 3236
rect 6390 3292 6454 3296
rect 6390 3236 6394 3292
rect 6394 3236 6450 3292
rect 6450 3236 6454 3292
rect 6390 3232 6454 3236
rect 11348 3292 11412 3296
rect 11348 3236 11352 3292
rect 11352 3236 11408 3292
rect 11408 3236 11412 3292
rect 11348 3232 11412 3236
rect 11428 3292 11492 3296
rect 11428 3236 11432 3292
rect 11432 3236 11488 3292
rect 11488 3236 11492 3292
rect 11428 3232 11492 3236
rect 11508 3292 11572 3296
rect 11508 3236 11512 3292
rect 11512 3236 11568 3292
rect 11568 3236 11572 3292
rect 11508 3232 11572 3236
rect 11588 3292 11652 3296
rect 11588 3236 11592 3292
rect 11592 3236 11648 3292
rect 11648 3236 11652 3292
rect 11588 3232 11652 3236
rect 16546 3292 16610 3296
rect 16546 3236 16550 3292
rect 16550 3236 16606 3292
rect 16606 3236 16610 3292
rect 16546 3232 16610 3236
rect 16626 3292 16690 3296
rect 16626 3236 16630 3292
rect 16630 3236 16686 3292
rect 16686 3236 16690 3292
rect 16626 3232 16690 3236
rect 16706 3292 16770 3296
rect 16706 3236 16710 3292
rect 16710 3236 16766 3292
rect 16766 3236 16770 3292
rect 16706 3232 16770 3236
rect 16786 3292 16850 3296
rect 16786 3236 16790 3292
rect 16790 3236 16846 3292
rect 16846 3236 16850 3292
rect 16786 3232 16850 3236
rect 21744 3292 21808 3296
rect 21744 3236 21748 3292
rect 21748 3236 21804 3292
rect 21804 3236 21808 3292
rect 21744 3232 21808 3236
rect 21824 3292 21888 3296
rect 21824 3236 21828 3292
rect 21828 3236 21884 3292
rect 21884 3236 21888 3292
rect 21824 3232 21888 3236
rect 21904 3292 21968 3296
rect 21904 3236 21908 3292
rect 21908 3236 21964 3292
rect 21964 3236 21968 3292
rect 21904 3232 21968 3236
rect 21984 3292 22048 3296
rect 21984 3236 21988 3292
rect 21988 3236 22044 3292
rect 22044 3236 22048 3292
rect 21984 3232 22048 3236
rect 8340 3164 8404 3228
rect 8524 3164 8588 3228
rect 9812 3164 9876 3228
rect 19012 3164 19076 3228
rect 12020 3028 12084 3092
rect 5948 2756 6012 2820
rect 3551 2748 3615 2752
rect 3551 2692 3555 2748
rect 3555 2692 3611 2748
rect 3611 2692 3615 2748
rect 3551 2688 3615 2692
rect 3631 2748 3695 2752
rect 3631 2692 3635 2748
rect 3635 2692 3691 2748
rect 3691 2692 3695 2748
rect 3631 2688 3695 2692
rect 3711 2748 3775 2752
rect 3711 2692 3715 2748
rect 3715 2692 3771 2748
rect 3771 2692 3775 2748
rect 3711 2688 3775 2692
rect 3791 2748 3855 2752
rect 3791 2692 3795 2748
rect 3795 2692 3851 2748
rect 3851 2692 3855 2748
rect 3791 2688 3855 2692
rect 8156 2620 8220 2684
rect 2820 2544 2884 2548
rect 2820 2488 2870 2544
rect 2870 2488 2884 2544
rect 2820 2484 2884 2488
rect 7604 2484 7668 2548
rect 6868 2348 6932 2412
rect 796 2212 860 2276
rect 5212 2212 5276 2276
rect 5396 2272 5460 2276
rect 9260 2756 9324 2820
rect 8749 2748 8813 2752
rect 8749 2692 8753 2748
rect 8753 2692 8809 2748
rect 8809 2692 8813 2748
rect 8749 2688 8813 2692
rect 8829 2748 8893 2752
rect 8829 2692 8833 2748
rect 8833 2692 8889 2748
rect 8889 2692 8893 2748
rect 8829 2688 8893 2692
rect 8909 2748 8973 2752
rect 8909 2692 8913 2748
rect 8913 2692 8969 2748
rect 8969 2692 8973 2748
rect 8909 2688 8973 2692
rect 8989 2748 9053 2752
rect 8989 2692 8993 2748
rect 8993 2692 9049 2748
rect 9049 2692 9053 2748
rect 8989 2688 9053 2692
rect 13947 2748 14011 2752
rect 13947 2692 13951 2748
rect 13951 2692 14007 2748
rect 14007 2692 14011 2748
rect 13947 2688 14011 2692
rect 14027 2748 14091 2752
rect 14027 2692 14031 2748
rect 14031 2692 14087 2748
rect 14087 2692 14091 2748
rect 14027 2688 14091 2692
rect 14107 2748 14171 2752
rect 14107 2692 14111 2748
rect 14111 2692 14167 2748
rect 14167 2692 14171 2748
rect 14107 2688 14171 2692
rect 14187 2748 14251 2752
rect 14187 2692 14191 2748
rect 14191 2692 14247 2748
rect 14247 2692 14251 2748
rect 14187 2688 14251 2692
rect 19145 2748 19209 2752
rect 19145 2692 19149 2748
rect 19149 2692 19205 2748
rect 19205 2692 19209 2748
rect 19145 2688 19209 2692
rect 19225 2748 19289 2752
rect 19225 2692 19229 2748
rect 19229 2692 19285 2748
rect 19285 2692 19289 2748
rect 19225 2688 19289 2692
rect 19305 2748 19369 2752
rect 19305 2692 19309 2748
rect 19309 2692 19365 2748
rect 19365 2692 19369 2748
rect 19305 2688 19369 2692
rect 19385 2748 19449 2752
rect 19385 2692 19389 2748
rect 19389 2692 19445 2748
rect 19445 2692 19449 2748
rect 19385 2688 19449 2692
rect 17356 2620 17420 2684
rect 17908 2620 17972 2684
rect 17356 2484 17420 2548
rect 5396 2216 5446 2272
rect 5446 2216 5460 2272
rect 5396 2212 5460 2216
rect 21036 2272 21100 2276
rect 21036 2216 21050 2272
rect 21050 2216 21100 2272
rect 21036 2212 21100 2216
rect 21404 2272 21468 2276
rect 21404 2216 21418 2272
rect 21418 2216 21468 2272
rect 21404 2212 21468 2216
rect 6150 2204 6214 2208
rect 6150 2148 6154 2204
rect 6154 2148 6210 2204
rect 6210 2148 6214 2204
rect 6150 2144 6214 2148
rect 6230 2204 6294 2208
rect 6230 2148 6234 2204
rect 6234 2148 6290 2204
rect 6290 2148 6294 2204
rect 6230 2144 6294 2148
rect 6310 2204 6374 2208
rect 6310 2148 6314 2204
rect 6314 2148 6370 2204
rect 6370 2148 6374 2204
rect 6310 2144 6374 2148
rect 6390 2204 6454 2208
rect 6390 2148 6394 2204
rect 6394 2148 6450 2204
rect 6450 2148 6454 2204
rect 6390 2144 6454 2148
rect 11348 2204 11412 2208
rect 11348 2148 11352 2204
rect 11352 2148 11408 2204
rect 11408 2148 11412 2204
rect 11348 2144 11412 2148
rect 11428 2204 11492 2208
rect 11428 2148 11432 2204
rect 11432 2148 11488 2204
rect 11488 2148 11492 2204
rect 11428 2144 11492 2148
rect 11508 2204 11572 2208
rect 11508 2148 11512 2204
rect 11512 2148 11568 2204
rect 11568 2148 11572 2204
rect 11508 2144 11572 2148
rect 11588 2204 11652 2208
rect 11588 2148 11592 2204
rect 11592 2148 11648 2204
rect 11648 2148 11652 2204
rect 11588 2144 11652 2148
rect 16546 2204 16610 2208
rect 16546 2148 16550 2204
rect 16550 2148 16606 2204
rect 16606 2148 16610 2204
rect 16546 2144 16610 2148
rect 16626 2204 16690 2208
rect 16626 2148 16630 2204
rect 16630 2148 16686 2204
rect 16686 2148 16690 2204
rect 16626 2144 16690 2148
rect 16706 2204 16770 2208
rect 16706 2148 16710 2204
rect 16710 2148 16766 2204
rect 16766 2148 16770 2204
rect 16706 2144 16770 2148
rect 16786 2204 16850 2208
rect 16786 2148 16790 2204
rect 16790 2148 16846 2204
rect 16846 2148 16850 2204
rect 16786 2144 16850 2148
rect 21744 2204 21808 2208
rect 21744 2148 21748 2204
rect 21748 2148 21804 2204
rect 21804 2148 21808 2204
rect 21744 2144 21808 2148
rect 21824 2204 21888 2208
rect 21824 2148 21828 2204
rect 21828 2148 21884 2204
rect 21884 2148 21888 2204
rect 21824 2144 21888 2148
rect 21904 2204 21968 2208
rect 21904 2148 21908 2204
rect 21908 2148 21964 2204
rect 21964 2148 21968 2204
rect 21904 2144 21968 2148
rect 21984 2204 22048 2208
rect 21984 2148 21988 2204
rect 21988 2148 22044 2204
rect 22044 2148 22048 2204
rect 21984 2144 22048 2148
rect 980 1940 1044 2004
rect 612 1804 676 1868
rect 7420 1804 7484 1868
rect 18644 1804 18708 1868
rect 3551 1660 3615 1664
rect 3551 1604 3555 1660
rect 3555 1604 3611 1660
rect 3611 1604 3615 1660
rect 3551 1600 3615 1604
rect 3631 1660 3695 1664
rect 3631 1604 3635 1660
rect 3635 1604 3691 1660
rect 3691 1604 3695 1660
rect 3631 1600 3695 1604
rect 3711 1660 3775 1664
rect 3711 1604 3715 1660
rect 3715 1604 3771 1660
rect 3771 1604 3775 1660
rect 3711 1600 3775 1604
rect 3791 1660 3855 1664
rect 3791 1604 3795 1660
rect 3795 1604 3851 1660
rect 3851 1604 3855 1660
rect 3791 1600 3855 1604
rect 8749 1660 8813 1664
rect 8749 1604 8753 1660
rect 8753 1604 8809 1660
rect 8809 1604 8813 1660
rect 8749 1600 8813 1604
rect 8829 1660 8893 1664
rect 8829 1604 8833 1660
rect 8833 1604 8889 1660
rect 8889 1604 8893 1660
rect 8829 1600 8893 1604
rect 8909 1660 8973 1664
rect 8909 1604 8913 1660
rect 8913 1604 8969 1660
rect 8969 1604 8973 1660
rect 8909 1600 8973 1604
rect 8989 1660 9053 1664
rect 8989 1604 8993 1660
rect 8993 1604 9049 1660
rect 9049 1604 9053 1660
rect 8989 1600 9053 1604
rect 13947 1660 14011 1664
rect 13947 1604 13951 1660
rect 13951 1604 14007 1660
rect 14007 1604 14011 1660
rect 13947 1600 14011 1604
rect 14027 1660 14091 1664
rect 14027 1604 14031 1660
rect 14031 1604 14087 1660
rect 14087 1604 14091 1660
rect 14027 1600 14091 1604
rect 14107 1660 14171 1664
rect 14107 1604 14111 1660
rect 14111 1604 14167 1660
rect 14167 1604 14171 1660
rect 14107 1600 14171 1604
rect 14187 1660 14251 1664
rect 14187 1604 14191 1660
rect 14191 1604 14247 1660
rect 14247 1604 14251 1660
rect 14187 1600 14251 1604
rect 16988 1728 17052 1732
rect 16988 1672 17038 1728
rect 17038 1672 17052 1728
rect 16988 1668 17052 1672
rect 19145 1660 19209 1664
rect 19145 1604 19149 1660
rect 19149 1604 19205 1660
rect 19205 1604 19209 1660
rect 19145 1600 19209 1604
rect 19225 1660 19289 1664
rect 19225 1604 19229 1660
rect 19229 1604 19285 1660
rect 19285 1604 19289 1660
rect 19225 1600 19289 1604
rect 19305 1660 19369 1664
rect 19305 1604 19309 1660
rect 19309 1604 19365 1660
rect 19365 1604 19369 1660
rect 19305 1600 19369 1604
rect 19385 1660 19449 1664
rect 19385 1604 19389 1660
rect 19389 1604 19445 1660
rect 19445 1604 19449 1660
rect 19385 1600 19449 1604
rect 1164 1260 1228 1324
rect 4108 1260 4172 1324
rect 7236 1260 7300 1324
rect 9812 1320 9876 1324
rect 9812 1264 9862 1320
rect 9862 1264 9876 1320
rect 9812 1260 9876 1264
rect 19012 1124 19076 1188
rect 6150 1116 6214 1120
rect 6150 1060 6154 1116
rect 6154 1060 6210 1116
rect 6210 1060 6214 1116
rect 6150 1056 6214 1060
rect 6230 1116 6294 1120
rect 6230 1060 6234 1116
rect 6234 1060 6290 1116
rect 6290 1060 6294 1116
rect 6230 1056 6294 1060
rect 6310 1116 6374 1120
rect 6310 1060 6314 1116
rect 6314 1060 6370 1116
rect 6370 1060 6374 1116
rect 6310 1056 6374 1060
rect 6390 1116 6454 1120
rect 6390 1060 6394 1116
rect 6394 1060 6450 1116
rect 6450 1060 6454 1116
rect 6390 1056 6454 1060
rect 11348 1116 11412 1120
rect 11348 1060 11352 1116
rect 11352 1060 11408 1116
rect 11408 1060 11412 1116
rect 11348 1056 11412 1060
rect 11428 1116 11492 1120
rect 11428 1060 11432 1116
rect 11432 1060 11488 1116
rect 11488 1060 11492 1116
rect 11428 1056 11492 1060
rect 11508 1116 11572 1120
rect 11508 1060 11512 1116
rect 11512 1060 11568 1116
rect 11568 1060 11572 1116
rect 11508 1056 11572 1060
rect 11588 1116 11652 1120
rect 11588 1060 11592 1116
rect 11592 1060 11648 1116
rect 11648 1060 11652 1116
rect 11588 1056 11652 1060
rect 16546 1116 16610 1120
rect 16546 1060 16550 1116
rect 16550 1060 16606 1116
rect 16606 1060 16610 1116
rect 16546 1056 16610 1060
rect 16626 1116 16690 1120
rect 16626 1060 16630 1116
rect 16630 1060 16686 1116
rect 16686 1060 16690 1116
rect 16626 1056 16690 1060
rect 16706 1116 16770 1120
rect 16706 1060 16710 1116
rect 16710 1060 16766 1116
rect 16766 1060 16770 1116
rect 16706 1056 16770 1060
rect 16786 1116 16850 1120
rect 16786 1060 16790 1116
rect 16790 1060 16846 1116
rect 16846 1060 16850 1116
rect 16786 1056 16850 1060
rect 21744 1116 21808 1120
rect 21744 1060 21748 1116
rect 21748 1060 21804 1116
rect 21804 1060 21808 1116
rect 21744 1056 21808 1060
rect 21824 1116 21888 1120
rect 21824 1060 21828 1116
rect 21828 1060 21884 1116
rect 21884 1060 21888 1116
rect 21824 1056 21888 1060
rect 21904 1116 21968 1120
rect 21904 1060 21908 1116
rect 21908 1060 21964 1116
rect 21964 1060 21968 1116
rect 21904 1056 21968 1060
rect 21984 1116 22048 1120
rect 21984 1060 21988 1116
rect 21988 1060 22044 1116
rect 22044 1060 22048 1116
rect 21984 1056 22048 1060
rect 9628 852 9692 916
rect 19932 852 19996 916
rect 20668 852 20732 916
rect 18828 580 18892 644
rect 8524 36 8588 100
<< metal4 >>
rect 3543 43008 3863 43568
rect 3543 42944 3551 43008
rect 3615 42944 3631 43008
rect 3695 42944 3711 43008
rect 3775 42944 3791 43008
rect 3855 42944 3863 43008
rect 3543 41920 3863 42944
rect 6142 43552 6462 43568
rect 6142 43488 6150 43552
rect 6214 43488 6230 43552
rect 6294 43488 6310 43552
rect 6374 43488 6390 43552
rect 6454 43488 6462 43552
rect 5027 42940 5093 42941
rect 5027 42876 5028 42940
rect 5092 42876 5093 42940
rect 5027 42875 5093 42876
rect 3543 41856 3551 41920
rect 3615 41856 3631 41920
rect 3695 41856 3711 41920
rect 3775 41856 3791 41920
rect 3855 41856 3863 41920
rect 795 41716 861 41717
rect 795 41652 796 41716
rect 860 41652 861 41716
rect 795 41651 861 41652
rect 611 40628 677 40629
rect 611 40564 612 40628
rect 676 40564 677 40628
rect 611 40563 677 40564
rect 243 16148 309 16149
rect 243 16084 244 16148
rect 308 16084 309 16148
rect 243 16083 309 16084
rect 246 13837 306 16083
rect 427 15060 493 15061
rect 427 14996 428 15060
rect 492 14996 493 15060
rect 427 14995 493 14996
rect 243 13836 309 13837
rect 243 13772 244 13836
rect 308 13772 309 13836
rect 243 13771 309 13772
rect 430 13021 490 14995
rect 427 13020 493 13021
rect 427 12956 428 13020
rect 492 12956 493 13020
rect 427 12955 493 12956
rect 614 1869 674 40563
rect 798 16829 858 41651
rect 3543 40832 3863 41856
rect 4659 41580 4725 41581
rect 4659 41516 4660 41580
rect 4724 41516 4725 41580
rect 4659 41515 4725 41516
rect 3543 40768 3551 40832
rect 3615 40768 3631 40832
rect 3695 40768 3711 40832
rect 3775 40768 3791 40832
rect 3855 40768 3863 40832
rect 3543 39744 3863 40768
rect 3543 39680 3551 39744
rect 3615 39680 3631 39744
rect 3695 39680 3711 39744
rect 3775 39680 3791 39744
rect 3855 39680 3863 39744
rect 2267 38724 2333 38725
rect 2267 38660 2268 38724
rect 2332 38660 2333 38724
rect 2267 38659 2333 38660
rect 2270 36685 2330 38659
rect 3543 38656 3863 39680
rect 3543 38592 3551 38656
rect 3615 38592 3631 38656
rect 3695 38592 3711 38656
rect 3775 38592 3791 38656
rect 3855 38592 3863 38656
rect 3543 37568 3863 38592
rect 3543 37504 3551 37568
rect 3615 37504 3631 37568
rect 3695 37504 3711 37568
rect 3775 37504 3791 37568
rect 3855 37504 3863 37568
rect 2267 36684 2333 36685
rect 2267 36620 2268 36684
rect 2332 36620 2333 36684
rect 2267 36619 2333 36620
rect 1715 35324 1781 35325
rect 1715 35260 1716 35324
rect 1780 35260 1781 35324
rect 1715 35259 1781 35260
rect 979 34508 1045 34509
rect 979 34444 980 34508
rect 1044 34444 1045 34508
rect 979 34443 1045 34444
rect 795 16828 861 16829
rect 795 16764 796 16828
rect 860 16764 861 16828
rect 795 16763 861 16764
rect 795 15196 861 15197
rect 795 15132 796 15196
rect 860 15132 861 15196
rect 795 15131 861 15132
rect 798 2277 858 15131
rect 795 2276 861 2277
rect 795 2212 796 2276
rect 860 2212 861 2276
rect 795 2211 861 2212
rect 982 2005 1042 34443
rect 1531 33420 1597 33421
rect 1531 33356 1532 33420
rect 1596 33356 1597 33420
rect 1531 33355 1597 33356
rect 1534 31770 1594 33355
rect 1166 31710 1594 31770
rect 1166 19005 1226 31710
rect 1531 31244 1597 31245
rect 1531 31180 1532 31244
rect 1596 31180 1597 31244
rect 1531 31179 1597 31180
rect 1534 26893 1594 31179
rect 1531 26892 1597 26893
rect 1531 26828 1532 26892
rect 1596 26828 1597 26892
rect 1531 26827 1597 26828
rect 1347 26212 1413 26213
rect 1347 26148 1348 26212
rect 1412 26148 1413 26212
rect 1347 26147 1413 26148
rect 1163 19004 1229 19005
rect 1163 18940 1164 19004
rect 1228 18940 1229 19004
rect 1163 18939 1229 18940
rect 1350 18730 1410 26147
rect 1718 26077 1778 35259
rect 1899 32332 1965 32333
rect 1899 32268 1900 32332
rect 1964 32268 1965 32332
rect 1899 32267 1965 32268
rect 1902 27301 1962 32267
rect 2270 31925 2330 36619
rect 3543 36480 3863 37504
rect 3543 36416 3551 36480
rect 3615 36416 3631 36480
rect 3695 36416 3711 36480
rect 3775 36416 3791 36480
rect 3855 36416 3863 36480
rect 3543 35392 3863 36416
rect 3543 35328 3551 35392
rect 3615 35328 3631 35392
rect 3695 35328 3711 35392
rect 3775 35328 3791 35392
rect 3855 35328 3863 35392
rect 2451 35324 2517 35325
rect 2451 35260 2452 35324
rect 2516 35260 2517 35324
rect 2451 35259 2517 35260
rect 2267 31924 2333 31925
rect 2267 31860 2268 31924
rect 2332 31860 2333 31924
rect 2267 31859 2333 31860
rect 2083 31788 2149 31789
rect 2083 31724 2084 31788
rect 2148 31724 2149 31788
rect 2083 31723 2149 31724
rect 2086 30701 2146 31723
rect 2083 30700 2149 30701
rect 2083 30636 2084 30700
rect 2148 30636 2149 30700
rect 2083 30635 2149 30636
rect 2267 28524 2333 28525
rect 2267 28460 2268 28524
rect 2332 28460 2333 28524
rect 2267 28459 2333 28460
rect 1899 27300 1965 27301
rect 1899 27236 1900 27300
rect 1964 27236 1965 27300
rect 1899 27235 1965 27236
rect 2083 27164 2149 27165
rect 2083 27100 2084 27164
rect 2148 27100 2149 27164
rect 2083 27099 2149 27100
rect 1715 26076 1781 26077
rect 1715 26012 1716 26076
rect 1780 26012 1781 26076
rect 1715 26011 1781 26012
rect 1715 25804 1781 25805
rect 1715 25740 1716 25804
rect 1780 25740 1781 25804
rect 1715 25739 1781 25740
rect 1166 18670 1410 18730
rect 1166 13293 1226 18670
rect 1531 17644 1597 17645
rect 1531 17580 1532 17644
rect 1596 17580 1597 17644
rect 1531 17579 1597 17580
rect 1163 13292 1229 13293
rect 1163 13228 1164 13292
rect 1228 13228 1229 13292
rect 1163 13227 1229 13228
rect 1347 13020 1413 13021
rect 1347 12956 1348 13020
rect 1412 12956 1413 13020
rect 1347 12955 1413 12956
rect 1350 2790 1410 12955
rect 1534 11797 1594 17579
rect 1718 16149 1778 25739
rect 2086 21181 2146 27099
rect 2083 21180 2149 21181
rect 2083 21116 2084 21180
rect 2148 21116 2149 21180
rect 2083 21115 2149 21116
rect 2270 16962 2330 28459
rect 2454 26485 2514 35259
rect 3003 34644 3069 34645
rect 3003 34580 3004 34644
rect 3068 34580 3069 34644
rect 3003 34579 3069 34580
rect 3006 29205 3066 34579
rect 3543 34304 3863 35328
rect 3543 34240 3551 34304
rect 3615 34240 3631 34304
rect 3695 34240 3711 34304
rect 3775 34240 3791 34304
rect 3855 34240 3863 34304
rect 3187 33692 3253 33693
rect 3187 33628 3188 33692
rect 3252 33628 3253 33692
rect 3187 33627 3253 33628
rect 3190 32877 3250 33627
rect 3543 33216 3863 34240
rect 3923 33964 3989 33965
rect 3923 33900 3924 33964
rect 3988 33900 3989 33964
rect 3923 33899 3989 33900
rect 3543 33152 3551 33216
rect 3615 33152 3631 33216
rect 3695 33152 3711 33216
rect 3775 33152 3791 33216
rect 3855 33152 3863 33216
rect 3187 32876 3253 32877
rect 3187 32812 3188 32876
rect 3252 32812 3253 32876
rect 3187 32811 3253 32812
rect 3190 30293 3250 32811
rect 3543 32128 3863 33152
rect 3543 32064 3551 32128
rect 3615 32064 3631 32128
rect 3695 32064 3711 32128
rect 3775 32064 3791 32128
rect 3855 32064 3863 32128
rect 3543 31040 3863 32064
rect 3543 30976 3551 31040
rect 3615 30976 3631 31040
rect 3695 30976 3711 31040
rect 3775 30976 3791 31040
rect 3855 30976 3863 31040
rect 3187 30292 3253 30293
rect 3187 30228 3188 30292
rect 3252 30228 3253 30292
rect 3187 30227 3253 30228
rect 3543 29952 3863 30976
rect 3543 29888 3551 29952
rect 3615 29888 3631 29952
rect 3695 29888 3711 29952
rect 3775 29888 3791 29952
rect 3855 29888 3863 29952
rect 3371 29748 3437 29749
rect 3371 29684 3372 29748
rect 3436 29684 3437 29748
rect 3371 29683 3437 29684
rect 3003 29204 3069 29205
rect 3003 29140 3004 29204
rect 3068 29140 3069 29204
rect 3003 29139 3069 29140
rect 2635 28388 2701 28389
rect 2635 28324 2636 28388
rect 2700 28324 2701 28388
rect 2635 28323 2701 28324
rect 2451 26484 2517 26485
rect 2451 26420 2452 26484
rect 2516 26420 2517 26484
rect 2451 26419 2517 26420
rect 2638 22949 2698 28323
rect 2819 27436 2885 27437
rect 2819 27372 2820 27436
rect 2884 27372 2885 27436
rect 2819 27371 2885 27372
rect 2822 23493 2882 27371
rect 3187 27300 3253 27301
rect 3187 27236 3188 27300
rect 3252 27236 3253 27300
rect 3187 27235 3253 27236
rect 3003 25396 3069 25397
rect 3003 25332 3004 25396
rect 3068 25332 3069 25396
rect 3003 25331 3069 25332
rect 2819 23492 2885 23493
rect 2819 23428 2820 23492
rect 2884 23428 2885 23492
rect 2819 23427 2885 23428
rect 2635 22948 2701 22949
rect 2635 22884 2636 22948
rect 2700 22884 2701 22948
rect 2635 22883 2701 22884
rect 2638 20637 2698 22883
rect 2635 20636 2701 20637
rect 2635 20572 2636 20636
rect 2700 20572 2701 20636
rect 2635 20571 2701 20572
rect 2451 19820 2517 19821
rect 2451 19756 2452 19820
rect 2516 19756 2517 19820
rect 2451 19755 2517 19756
rect 2086 16902 2330 16962
rect 1899 16828 1965 16829
rect 1899 16764 1900 16828
rect 1964 16764 1965 16828
rect 1899 16763 1965 16764
rect 1715 16148 1781 16149
rect 1715 16084 1716 16148
rect 1780 16084 1781 16148
rect 1715 16083 1781 16084
rect 1902 15469 1962 16763
rect 1899 15468 1965 15469
rect 1899 15404 1900 15468
rect 1964 15404 1965 15468
rect 1899 15403 1965 15404
rect 2086 13021 2146 16902
rect 2267 16828 2333 16829
rect 2267 16764 2268 16828
rect 2332 16764 2333 16828
rect 2267 16763 2333 16764
rect 2083 13020 2149 13021
rect 2083 12956 2084 13020
rect 2148 12956 2149 13020
rect 2083 12955 2149 12956
rect 1531 11796 1597 11797
rect 1531 11732 1532 11796
rect 1596 11732 1597 11796
rect 1531 11731 1597 11732
rect 1899 11796 1965 11797
rect 1899 11732 1900 11796
rect 1964 11732 1965 11796
rect 1899 11731 1965 11732
rect 1902 7309 1962 11731
rect 2083 11660 2149 11661
rect 2083 11596 2084 11660
rect 2148 11596 2149 11660
rect 2083 11595 2149 11596
rect 2086 7581 2146 11595
rect 2270 11117 2330 16763
rect 2267 11116 2333 11117
rect 2267 11052 2268 11116
rect 2332 11052 2333 11116
rect 2267 11051 2333 11052
rect 2454 8805 2514 19755
rect 3006 19549 3066 25331
rect 3190 25261 3250 27235
rect 3374 26757 3434 29683
rect 3543 28864 3863 29888
rect 3543 28800 3551 28864
rect 3615 28800 3631 28864
rect 3695 28800 3711 28864
rect 3775 28800 3791 28864
rect 3855 28800 3863 28864
rect 3543 27776 3863 28800
rect 3543 27712 3551 27776
rect 3615 27712 3631 27776
rect 3695 27712 3711 27776
rect 3775 27712 3791 27776
rect 3855 27712 3863 27776
rect 3371 26756 3437 26757
rect 3371 26692 3372 26756
rect 3436 26692 3437 26756
rect 3371 26691 3437 26692
rect 3543 26688 3863 27712
rect 3926 27437 3986 33899
rect 4107 31924 4173 31925
rect 4107 31860 4108 31924
rect 4172 31860 4173 31924
rect 4107 31859 4173 31860
rect 4110 29885 4170 31859
rect 4291 31788 4357 31789
rect 4291 31724 4292 31788
rect 4356 31724 4357 31788
rect 4291 31723 4357 31724
rect 4107 29884 4173 29885
rect 4107 29820 4108 29884
rect 4172 29820 4173 29884
rect 4107 29819 4173 29820
rect 3923 27436 3989 27437
rect 3923 27372 3924 27436
rect 3988 27372 3989 27436
rect 3923 27371 3989 27372
rect 3923 27164 3989 27165
rect 3923 27100 3924 27164
rect 3988 27100 3989 27164
rect 3923 27099 3989 27100
rect 3543 26624 3551 26688
rect 3615 26624 3631 26688
rect 3695 26624 3711 26688
rect 3775 26624 3791 26688
rect 3855 26624 3863 26688
rect 3543 25600 3863 26624
rect 3543 25536 3551 25600
rect 3615 25536 3631 25600
rect 3695 25536 3711 25600
rect 3775 25536 3791 25600
rect 3855 25536 3863 25600
rect 3187 25260 3253 25261
rect 3187 25196 3188 25260
rect 3252 25196 3253 25260
rect 3187 25195 3253 25196
rect 3543 24512 3863 25536
rect 3543 24448 3551 24512
rect 3615 24448 3631 24512
rect 3695 24448 3711 24512
rect 3775 24448 3791 24512
rect 3855 24448 3863 24512
rect 3543 23424 3863 24448
rect 3543 23360 3551 23424
rect 3615 23360 3631 23424
rect 3695 23360 3711 23424
rect 3775 23360 3791 23424
rect 3855 23360 3863 23424
rect 3543 22336 3863 23360
rect 3543 22272 3551 22336
rect 3615 22272 3631 22336
rect 3695 22272 3711 22336
rect 3775 22272 3791 22336
rect 3855 22272 3863 22336
rect 3543 21248 3863 22272
rect 3543 21184 3551 21248
rect 3615 21184 3631 21248
rect 3695 21184 3711 21248
rect 3775 21184 3791 21248
rect 3855 21184 3863 21248
rect 3543 20160 3863 21184
rect 3926 20501 3986 27099
rect 3923 20500 3989 20501
rect 3923 20436 3924 20500
rect 3988 20436 3989 20500
rect 3923 20435 3989 20436
rect 3543 20096 3551 20160
rect 3615 20096 3631 20160
rect 3695 20096 3711 20160
rect 3775 20096 3791 20160
rect 3855 20096 3863 20160
rect 3003 19548 3069 19549
rect 3003 19484 3004 19548
rect 3068 19484 3069 19548
rect 3003 19483 3069 19484
rect 3006 19350 3066 19483
rect 2638 19290 3066 19350
rect 2638 17373 2698 19290
rect 3543 19072 3863 20096
rect 3543 19008 3551 19072
rect 3615 19008 3631 19072
rect 3695 19008 3711 19072
rect 3775 19008 3791 19072
rect 3855 19008 3863 19072
rect 3187 19004 3253 19005
rect 3187 18940 3188 19004
rect 3252 18940 3253 19004
rect 3187 18939 3253 18940
rect 2635 17372 2701 17373
rect 2635 17308 2636 17372
rect 2700 17308 2701 17372
rect 2635 17307 2701 17308
rect 2819 17372 2885 17373
rect 2819 17308 2820 17372
rect 2884 17308 2885 17372
rect 2819 17307 2885 17308
rect 2635 15060 2701 15061
rect 2635 14996 2636 15060
rect 2700 14996 2701 15060
rect 2635 14995 2701 14996
rect 2638 9349 2698 14995
rect 2822 13565 2882 17307
rect 3190 15058 3250 18939
rect 3543 17984 3863 19008
rect 3543 17920 3551 17984
rect 3615 17920 3631 17984
rect 3695 17920 3711 17984
rect 3775 17920 3791 17984
rect 3855 17920 3863 17984
rect 3371 17916 3437 17917
rect 3371 17852 3372 17916
rect 3436 17852 3437 17916
rect 3371 17851 3437 17852
rect 3374 16557 3434 17851
rect 3543 16896 3863 17920
rect 4110 17917 4170 29819
rect 4294 29610 4354 31723
rect 4662 31517 4722 41515
rect 5030 39949 5090 42875
rect 6142 42464 6462 43488
rect 8741 43008 9061 43568
rect 8741 42944 8749 43008
rect 8813 42944 8829 43008
rect 8893 42944 8909 43008
rect 8973 42944 8989 43008
rect 9053 42944 9061 43008
rect 6683 42532 6749 42533
rect 6683 42468 6684 42532
rect 6748 42468 6749 42532
rect 6683 42467 6749 42468
rect 6142 42400 6150 42464
rect 6214 42400 6230 42464
rect 6294 42400 6310 42464
rect 6374 42400 6390 42464
rect 6454 42400 6462 42464
rect 6142 41376 6462 42400
rect 6142 41312 6150 41376
rect 6214 41312 6230 41376
rect 6294 41312 6310 41376
rect 6374 41312 6390 41376
rect 6454 41312 6462 41376
rect 6142 40288 6462 41312
rect 6142 40224 6150 40288
rect 6214 40224 6230 40288
rect 6294 40224 6310 40288
rect 6374 40224 6390 40288
rect 6454 40224 6462 40288
rect 5395 40220 5461 40221
rect 5395 40156 5396 40220
rect 5460 40156 5461 40220
rect 5395 40155 5461 40156
rect 5027 39948 5093 39949
rect 5027 39884 5028 39948
rect 5092 39884 5093 39948
rect 5027 39883 5093 39884
rect 4843 37636 4909 37637
rect 4843 37572 4844 37636
rect 4908 37572 4909 37636
rect 4843 37571 4909 37572
rect 4846 33149 4906 37571
rect 5027 36548 5093 36549
rect 5027 36484 5028 36548
rect 5092 36484 5093 36548
rect 5027 36483 5093 36484
rect 5030 33285 5090 36483
rect 5398 35461 5458 40155
rect 6142 39200 6462 40224
rect 6142 39136 6150 39200
rect 6214 39136 6230 39200
rect 6294 39136 6310 39200
rect 6374 39136 6390 39200
rect 6454 39136 6462 39200
rect 6142 38112 6462 39136
rect 6142 38048 6150 38112
rect 6214 38048 6230 38112
rect 6294 38048 6310 38112
rect 6374 38048 6390 38112
rect 6454 38048 6462 38112
rect 6142 37024 6462 38048
rect 6142 36960 6150 37024
rect 6214 36960 6230 37024
rect 6294 36960 6310 37024
rect 6374 36960 6390 37024
rect 6454 36960 6462 37024
rect 6142 35936 6462 36960
rect 6686 36821 6746 42467
rect 8339 42260 8405 42261
rect 8339 42196 8340 42260
rect 8404 42196 8405 42260
rect 8339 42195 8405 42196
rect 7419 41580 7485 41581
rect 7419 41516 7420 41580
rect 7484 41516 7485 41580
rect 7419 41515 7485 41516
rect 6683 36820 6749 36821
rect 6683 36756 6684 36820
rect 6748 36756 6749 36820
rect 6683 36755 6749 36756
rect 6867 36820 6933 36821
rect 6867 36756 6868 36820
rect 6932 36756 6933 36820
rect 6867 36755 6933 36756
rect 6142 35872 6150 35936
rect 6214 35872 6230 35936
rect 6294 35872 6310 35936
rect 6374 35872 6390 35936
rect 6454 35872 6462 35936
rect 5763 35868 5829 35869
rect 5763 35804 5764 35868
rect 5828 35804 5829 35868
rect 5763 35803 5829 35804
rect 5395 35460 5461 35461
rect 5395 35396 5396 35460
rect 5460 35396 5461 35460
rect 5395 35395 5461 35396
rect 5027 33284 5093 33285
rect 5027 33220 5028 33284
rect 5092 33220 5093 33284
rect 5027 33219 5093 33220
rect 4843 33148 4909 33149
rect 4843 33084 4844 33148
rect 4908 33084 4909 33148
rect 4843 33083 4909 33084
rect 4659 31516 4725 31517
rect 4659 31452 4660 31516
rect 4724 31452 4725 31516
rect 4659 31451 4725 31452
rect 4294 29550 4722 29610
rect 4291 28660 4357 28661
rect 4291 28596 4292 28660
rect 4356 28596 4357 28660
rect 4291 28595 4357 28596
rect 4294 24445 4354 28595
rect 4475 27164 4541 27165
rect 4475 27100 4476 27164
rect 4540 27100 4541 27164
rect 4475 27099 4541 27100
rect 4478 25669 4538 27099
rect 4475 25668 4541 25669
rect 4475 25604 4476 25668
rect 4540 25604 4541 25668
rect 4475 25603 4541 25604
rect 4291 24444 4357 24445
rect 4291 24380 4292 24444
rect 4356 24380 4357 24444
rect 4291 24379 4357 24380
rect 4291 24172 4357 24173
rect 4291 24108 4292 24172
rect 4356 24108 4357 24172
rect 4291 24107 4357 24108
rect 4294 18733 4354 24107
rect 4662 23493 4722 29550
rect 5030 29341 5090 33219
rect 5579 31380 5645 31381
rect 5579 31316 5580 31380
rect 5644 31316 5645 31380
rect 5579 31315 5645 31316
rect 5211 30156 5277 30157
rect 5211 30092 5212 30156
rect 5276 30092 5277 30156
rect 5211 30091 5277 30092
rect 5027 29340 5093 29341
rect 5027 29276 5028 29340
rect 5092 29276 5093 29340
rect 5027 29275 5093 29276
rect 4843 29068 4909 29069
rect 4843 29004 4844 29068
rect 4908 29004 4909 29068
rect 4843 29003 4909 29004
rect 4659 23492 4725 23493
rect 4659 23428 4660 23492
rect 4724 23428 4725 23492
rect 4659 23427 4725 23428
rect 4662 22405 4722 23427
rect 4659 22404 4725 22405
rect 4659 22340 4660 22404
rect 4724 22340 4725 22404
rect 4659 22339 4725 22340
rect 4659 20092 4725 20093
rect 4659 20028 4660 20092
rect 4724 20028 4725 20092
rect 4659 20027 4725 20028
rect 4291 18732 4357 18733
rect 4291 18668 4292 18732
rect 4356 18668 4357 18732
rect 4291 18667 4357 18668
rect 4107 17916 4173 17917
rect 4107 17852 4108 17916
rect 4172 17852 4173 17916
rect 4107 17851 4173 17852
rect 3923 17372 3989 17373
rect 3923 17308 3924 17372
rect 3988 17308 3989 17372
rect 3923 17307 3989 17308
rect 3543 16832 3551 16896
rect 3615 16832 3631 16896
rect 3695 16832 3711 16896
rect 3775 16832 3791 16896
rect 3855 16832 3863 16896
rect 3371 16556 3437 16557
rect 3371 16492 3372 16556
rect 3436 16492 3437 16556
rect 3371 16491 3437 16492
rect 3543 15808 3863 16832
rect 3543 15744 3551 15808
rect 3615 15744 3631 15808
rect 3695 15744 3711 15808
rect 3775 15744 3791 15808
rect 3855 15744 3863 15808
rect 3371 15060 3437 15061
rect 3371 15058 3372 15060
rect 3190 14998 3372 15058
rect 3371 14996 3372 14998
rect 3436 14996 3437 15060
rect 3371 14995 3437 14996
rect 3543 14720 3863 15744
rect 3543 14656 3551 14720
rect 3615 14656 3631 14720
rect 3695 14656 3711 14720
rect 3775 14656 3791 14720
rect 3855 14656 3863 14720
rect 3371 14652 3437 14653
rect 3371 14588 3372 14652
rect 3436 14588 3437 14652
rect 3371 14587 3437 14588
rect 3003 13700 3069 13701
rect 3003 13636 3004 13700
rect 3068 13636 3069 13700
rect 3003 13635 3069 13636
rect 2819 13564 2885 13565
rect 2819 13500 2820 13564
rect 2884 13500 2885 13564
rect 2819 13499 2885 13500
rect 2819 11252 2885 11253
rect 2819 11188 2820 11252
rect 2884 11188 2885 11252
rect 2819 11187 2885 11188
rect 2635 9348 2701 9349
rect 2635 9284 2636 9348
rect 2700 9284 2701 9348
rect 2635 9283 2701 9284
rect 2451 8804 2517 8805
rect 2451 8740 2452 8804
rect 2516 8740 2517 8804
rect 2451 8739 2517 8740
rect 2267 8668 2333 8669
rect 2267 8604 2268 8668
rect 2332 8604 2333 8668
rect 2267 8603 2333 8604
rect 2083 7580 2149 7581
rect 2083 7516 2084 7580
rect 2148 7516 2149 7580
rect 2083 7515 2149 7516
rect 1899 7308 1965 7309
rect 1899 7244 1900 7308
rect 1964 7244 1965 7308
rect 1899 7243 1965 7244
rect 2270 7173 2330 8603
rect 2451 8260 2517 8261
rect 2451 8196 2452 8260
rect 2516 8196 2517 8260
rect 2451 8195 2517 8196
rect 2267 7172 2333 7173
rect 2267 7108 2268 7172
rect 2332 7108 2333 7172
rect 2267 7107 2333 7108
rect 2454 4589 2514 8195
rect 2638 6629 2698 9283
rect 2822 6765 2882 11187
rect 3006 10573 3066 13635
rect 3187 11932 3253 11933
rect 3187 11868 3188 11932
rect 3252 11868 3253 11932
rect 3187 11867 3253 11868
rect 3190 10845 3250 11867
rect 3187 10844 3253 10845
rect 3187 10780 3188 10844
rect 3252 10780 3253 10844
rect 3187 10779 3253 10780
rect 3003 10572 3069 10573
rect 3003 10508 3004 10572
rect 3068 10508 3069 10572
rect 3003 10507 3069 10508
rect 3006 6765 3066 10507
rect 3374 8669 3434 14587
rect 3543 13632 3863 14656
rect 3926 14245 3986 17307
rect 4110 16693 4170 17851
rect 4107 16692 4173 16693
rect 4107 16628 4108 16692
rect 4172 16628 4173 16692
rect 4107 16627 4173 16628
rect 4110 15741 4170 16627
rect 4107 15740 4173 15741
rect 4107 15676 4108 15740
rect 4172 15676 4173 15740
rect 4107 15675 4173 15676
rect 3923 14244 3989 14245
rect 3923 14180 3924 14244
rect 3988 14180 3989 14244
rect 3923 14179 3989 14180
rect 3543 13568 3551 13632
rect 3615 13568 3631 13632
rect 3695 13568 3711 13632
rect 3775 13568 3791 13632
rect 3855 13568 3863 13632
rect 3543 12544 3863 13568
rect 3923 13292 3989 13293
rect 3923 13228 3924 13292
rect 3988 13228 3989 13292
rect 3923 13227 3989 13228
rect 3543 12480 3551 12544
rect 3615 12480 3631 12544
rect 3695 12480 3711 12544
rect 3775 12480 3791 12544
rect 3855 12480 3863 12544
rect 3543 11456 3863 12480
rect 3926 11933 3986 13227
rect 4110 11933 4170 15675
rect 4475 15604 4541 15605
rect 4475 15540 4476 15604
rect 4540 15540 4541 15604
rect 4475 15539 4541 15540
rect 3923 11932 3989 11933
rect 3923 11868 3924 11932
rect 3988 11868 3989 11932
rect 3923 11867 3989 11868
rect 4107 11932 4173 11933
rect 4107 11868 4108 11932
rect 4172 11868 4173 11932
rect 4107 11867 4173 11868
rect 3543 11392 3551 11456
rect 3615 11392 3631 11456
rect 3695 11392 3711 11456
rect 3775 11392 3791 11456
rect 3855 11392 3863 11456
rect 3543 10368 3863 11392
rect 4107 11388 4173 11389
rect 4107 11324 4108 11388
rect 4172 11324 4173 11388
rect 4107 11323 4173 11324
rect 3543 10304 3551 10368
rect 3615 10304 3631 10368
rect 3695 10304 3711 10368
rect 3775 10304 3791 10368
rect 3855 10304 3863 10368
rect 3543 9280 3863 10304
rect 3543 9216 3551 9280
rect 3615 9216 3631 9280
rect 3695 9216 3711 9280
rect 3775 9216 3791 9280
rect 3855 9216 3863 9280
rect 3371 8668 3437 8669
rect 3371 8604 3372 8668
rect 3436 8604 3437 8668
rect 3371 8603 3437 8604
rect 3187 8396 3253 8397
rect 3187 8332 3188 8396
rect 3252 8332 3253 8396
rect 3187 8331 3253 8332
rect 3371 8396 3437 8397
rect 3371 8332 3372 8396
rect 3436 8332 3437 8396
rect 3371 8331 3437 8332
rect 3190 7853 3250 8331
rect 3187 7852 3253 7853
rect 3187 7788 3188 7852
rect 3252 7788 3253 7852
rect 3187 7787 3253 7788
rect 2819 6764 2885 6765
rect 2819 6700 2820 6764
rect 2884 6700 2885 6764
rect 2819 6699 2885 6700
rect 3003 6764 3069 6765
rect 3003 6700 3004 6764
rect 3068 6700 3069 6764
rect 3003 6699 3069 6700
rect 2635 6628 2701 6629
rect 2635 6564 2636 6628
rect 2700 6564 2701 6628
rect 2635 6563 2701 6564
rect 2819 6084 2885 6085
rect 2819 6020 2820 6084
rect 2884 6020 2885 6084
rect 2819 6019 2885 6020
rect 2451 4588 2517 4589
rect 2451 4524 2452 4588
rect 2516 4524 2517 4588
rect 2451 4523 2517 4524
rect 1166 2730 1410 2790
rect 979 2004 1045 2005
rect 979 1940 980 2004
rect 1044 1940 1045 2004
rect 979 1939 1045 1940
rect 611 1868 677 1869
rect 611 1804 612 1868
rect 676 1804 677 1868
rect 611 1803 677 1804
rect 1166 1325 1226 2730
rect 2822 2549 2882 6019
rect 3374 5405 3434 8331
rect 3543 8192 3863 9216
rect 4110 8530 4170 11323
rect 4478 10981 4538 15539
rect 4662 14653 4722 20027
rect 4846 17509 4906 29003
rect 5027 27708 5093 27709
rect 5027 27644 5028 27708
rect 5092 27644 5093 27708
rect 5027 27643 5093 27644
rect 5030 24037 5090 27643
rect 5214 24717 5274 30091
rect 5395 26212 5461 26213
rect 5395 26148 5396 26212
rect 5460 26148 5461 26212
rect 5395 26147 5461 26148
rect 5211 24716 5277 24717
rect 5211 24652 5212 24716
rect 5276 24652 5277 24716
rect 5211 24651 5277 24652
rect 5027 24036 5093 24037
rect 5027 23972 5028 24036
rect 5092 23972 5093 24036
rect 5027 23971 5093 23972
rect 5027 19548 5093 19549
rect 5027 19484 5028 19548
rect 5092 19484 5093 19548
rect 5027 19483 5093 19484
rect 4843 17508 4909 17509
rect 4843 17444 4844 17508
rect 4908 17444 4909 17508
rect 4843 17443 4909 17444
rect 4843 15876 4909 15877
rect 4843 15812 4844 15876
rect 4908 15812 4909 15876
rect 4843 15811 4909 15812
rect 4659 14652 4725 14653
rect 4659 14588 4660 14652
rect 4724 14588 4725 14652
rect 4659 14587 4725 14588
rect 4662 12341 4722 14587
rect 4846 13293 4906 15811
rect 5030 15197 5090 19483
rect 5214 19413 5274 24651
rect 5211 19412 5277 19413
rect 5211 19348 5212 19412
rect 5276 19348 5277 19412
rect 5211 19347 5277 19348
rect 5211 19004 5277 19005
rect 5211 18940 5212 19004
rect 5276 18940 5277 19004
rect 5211 18939 5277 18940
rect 5027 15196 5093 15197
rect 5027 15132 5028 15196
rect 5092 15132 5093 15196
rect 5027 15131 5093 15132
rect 5027 13700 5093 13701
rect 5027 13636 5028 13700
rect 5092 13636 5093 13700
rect 5027 13635 5093 13636
rect 4843 13292 4909 13293
rect 4843 13228 4844 13292
rect 4908 13228 4909 13292
rect 4843 13227 4909 13228
rect 4659 12340 4725 12341
rect 4659 12276 4660 12340
rect 4724 12276 4725 12340
rect 4659 12275 4725 12276
rect 4475 10980 4541 10981
rect 4475 10916 4476 10980
rect 4540 10916 4541 10980
rect 4475 10915 4541 10916
rect 5030 9893 5090 13635
rect 5214 11525 5274 18939
rect 5398 16149 5458 26147
rect 5395 16148 5461 16149
rect 5395 16084 5396 16148
rect 5460 16084 5461 16148
rect 5395 16083 5461 16084
rect 5582 16010 5642 31315
rect 5766 31109 5826 35803
rect 5947 34916 6013 34917
rect 5947 34852 5948 34916
rect 6012 34852 6013 34916
rect 5947 34851 6013 34852
rect 5763 31108 5829 31109
rect 5763 31044 5764 31108
rect 5828 31044 5829 31108
rect 5763 31043 5829 31044
rect 5950 30565 6010 34851
rect 6142 34848 6462 35872
rect 6142 34784 6150 34848
rect 6214 34784 6230 34848
rect 6294 34784 6310 34848
rect 6374 34784 6390 34848
rect 6454 34784 6462 34848
rect 6142 33760 6462 34784
rect 6683 34236 6749 34237
rect 6683 34172 6684 34236
rect 6748 34172 6749 34236
rect 6683 34171 6749 34172
rect 6142 33696 6150 33760
rect 6214 33696 6230 33760
rect 6294 33696 6310 33760
rect 6374 33696 6390 33760
rect 6454 33696 6462 33760
rect 6142 32672 6462 33696
rect 6142 32608 6150 32672
rect 6214 32608 6230 32672
rect 6294 32608 6310 32672
rect 6374 32608 6390 32672
rect 6454 32608 6462 32672
rect 6142 31584 6462 32608
rect 6142 31520 6150 31584
rect 6214 31520 6230 31584
rect 6294 31520 6310 31584
rect 6374 31520 6390 31584
rect 6454 31520 6462 31584
rect 5947 30564 6013 30565
rect 5947 30500 5948 30564
rect 6012 30500 6013 30564
rect 5947 30499 6013 30500
rect 6142 30496 6462 31520
rect 6142 30432 6150 30496
rect 6214 30432 6230 30496
rect 6294 30432 6310 30496
rect 6374 30432 6390 30496
rect 6454 30432 6462 30496
rect 6142 29408 6462 30432
rect 6142 29344 6150 29408
rect 6214 29344 6230 29408
rect 6294 29344 6310 29408
rect 6374 29344 6390 29408
rect 6454 29344 6462 29408
rect 5947 28796 6013 28797
rect 5947 28732 5948 28796
rect 6012 28732 6013 28796
rect 5947 28731 6013 28732
rect 5950 28389 6010 28731
rect 5947 28388 6013 28389
rect 5947 28324 5948 28388
rect 6012 28324 6013 28388
rect 5947 28323 6013 28324
rect 5763 25668 5829 25669
rect 5763 25604 5764 25668
rect 5828 25604 5829 25668
rect 5763 25603 5829 25604
rect 5766 20773 5826 25603
rect 5950 24309 6010 28323
rect 6142 28320 6462 29344
rect 6686 28661 6746 34171
rect 6870 32333 6930 36755
rect 7235 36684 7301 36685
rect 7235 36620 7236 36684
rect 7300 36620 7301 36684
rect 7235 36619 7301 36620
rect 6867 32332 6933 32333
rect 6867 32268 6868 32332
rect 6932 32268 6933 32332
rect 6867 32267 6933 32268
rect 7238 30565 7298 36619
rect 7235 30564 7301 30565
rect 7235 30500 7236 30564
rect 7300 30500 7301 30564
rect 7235 30499 7301 30500
rect 6683 28660 6749 28661
rect 6683 28596 6684 28660
rect 6748 28596 6749 28660
rect 6683 28595 6749 28596
rect 6142 28256 6150 28320
rect 6214 28256 6230 28320
rect 6294 28256 6310 28320
rect 6374 28256 6390 28320
rect 6454 28256 6462 28320
rect 6142 27232 6462 28256
rect 7235 27708 7301 27709
rect 7235 27644 7236 27708
rect 7300 27644 7301 27708
rect 7235 27643 7301 27644
rect 6142 27168 6150 27232
rect 6214 27168 6230 27232
rect 6294 27168 6310 27232
rect 6374 27168 6390 27232
rect 6454 27168 6462 27232
rect 6142 26144 6462 27168
rect 6683 26756 6749 26757
rect 6683 26692 6684 26756
rect 6748 26692 6749 26756
rect 6683 26691 6749 26692
rect 6142 26080 6150 26144
rect 6214 26080 6230 26144
rect 6294 26080 6310 26144
rect 6374 26080 6390 26144
rect 6454 26080 6462 26144
rect 6142 25056 6462 26080
rect 6142 24992 6150 25056
rect 6214 24992 6230 25056
rect 6294 24992 6310 25056
rect 6374 24992 6390 25056
rect 6454 24992 6462 25056
rect 5947 24308 6013 24309
rect 5947 24244 5948 24308
rect 6012 24244 6013 24308
rect 5947 24243 6013 24244
rect 6142 23968 6462 24992
rect 6142 23904 6150 23968
rect 6214 23904 6230 23968
rect 6294 23904 6310 23968
rect 6374 23904 6390 23968
rect 6454 23904 6462 23968
rect 6142 22880 6462 23904
rect 6142 22816 6150 22880
rect 6214 22816 6230 22880
rect 6294 22816 6310 22880
rect 6374 22816 6390 22880
rect 6454 22816 6462 22880
rect 6142 21792 6462 22816
rect 6142 21728 6150 21792
rect 6214 21728 6230 21792
rect 6294 21728 6310 21792
rect 6374 21728 6390 21792
rect 6454 21728 6462 21792
rect 5763 20772 5829 20773
rect 5763 20708 5764 20772
rect 5828 20708 5829 20772
rect 5763 20707 5829 20708
rect 6142 20704 6462 21728
rect 6142 20640 6150 20704
rect 6214 20640 6230 20704
rect 6294 20640 6310 20704
rect 6374 20640 6390 20704
rect 6454 20640 6462 20704
rect 6142 19616 6462 20640
rect 6142 19552 6150 19616
rect 6214 19552 6230 19616
rect 6294 19552 6310 19616
rect 6374 19552 6390 19616
rect 6454 19552 6462 19616
rect 5947 19140 6013 19141
rect 5947 19076 5948 19140
rect 6012 19076 6013 19140
rect 5947 19075 6013 19076
rect 5398 15950 5642 16010
rect 5211 11524 5277 11525
rect 5211 11460 5212 11524
rect 5276 11460 5277 11524
rect 5211 11459 5277 11460
rect 5027 9892 5093 9893
rect 5027 9828 5028 9892
rect 5092 9828 5093 9892
rect 5027 9827 5093 9828
rect 5030 9690 5090 9827
rect 4662 9630 5090 9690
rect 4291 9212 4357 9213
rect 4291 9148 4292 9212
rect 4356 9148 4357 9212
rect 4291 9147 4357 9148
rect 3543 8128 3551 8192
rect 3615 8128 3631 8192
rect 3695 8128 3711 8192
rect 3775 8128 3791 8192
rect 3855 8128 3863 8192
rect 3543 7104 3863 8128
rect 3543 7040 3551 7104
rect 3615 7040 3631 7104
rect 3695 7040 3711 7104
rect 3775 7040 3791 7104
rect 3855 7040 3863 7104
rect 3543 6016 3863 7040
rect 3926 8470 4170 8530
rect 3926 6765 3986 8470
rect 4294 7170 4354 9147
rect 4475 8668 4541 8669
rect 4475 8604 4476 8668
rect 4540 8604 4541 8668
rect 4475 8603 4541 8604
rect 4478 7581 4538 8603
rect 4475 7580 4541 7581
rect 4475 7516 4476 7580
rect 4540 7516 4541 7580
rect 4475 7515 4541 7516
rect 4110 7110 4354 7170
rect 3923 6764 3989 6765
rect 3923 6700 3924 6764
rect 3988 6700 3989 6764
rect 3923 6699 3989 6700
rect 3543 5952 3551 6016
rect 3615 5952 3631 6016
rect 3695 5952 3711 6016
rect 3775 5952 3791 6016
rect 3855 5952 3863 6016
rect 3371 5404 3437 5405
rect 3371 5340 3372 5404
rect 3436 5340 3437 5404
rect 3371 5339 3437 5340
rect 3543 4928 3863 5952
rect 3543 4864 3551 4928
rect 3615 4864 3631 4928
rect 3695 4864 3711 4928
rect 3775 4864 3791 4928
rect 3855 4864 3863 4928
rect 3543 3840 3863 4864
rect 4110 4589 4170 7110
rect 4662 7037 4722 9630
rect 5027 8532 5093 8533
rect 5027 8468 5028 8532
rect 5092 8468 5093 8532
rect 5027 8467 5093 8468
rect 4291 7036 4357 7037
rect 4291 6972 4292 7036
rect 4356 6972 4357 7036
rect 4291 6971 4357 6972
rect 4659 7036 4725 7037
rect 4659 6972 4660 7036
rect 4724 6972 4725 7036
rect 4659 6971 4725 6972
rect 4294 4589 4354 6971
rect 4475 6628 4541 6629
rect 4475 6564 4476 6628
rect 4540 6564 4541 6628
rect 4475 6563 4541 6564
rect 4478 5813 4538 6563
rect 4475 5812 4541 5813
rect 4475 5748 4476 5812
rect 4540 5748 4541 5812
rect 4475 5747 4541 5748
rect 4107 4588 4173 4589
rect 4107 4524 4108 4588
rect 4172 4524 4173 4588
rect 4107 4523 4173 4524
rect 4291 4588 4357 4589
rect 4291 4524 4292 4588
rect 4356 4524 4357 4588
rect 4291 4523 4357 4524
rect 4662 4453 4722 6971
rect 5030 5133 5090 8467
rect 5214 8261 5274 11459
rect 5398 10981 5458 15950
rect 5763 15468 5829 15469
rect 5763 15404 5764 15468
rect 5828 15404 5829 15468
rect 5763 15403 5829 15404
rect 5579 13836 5645 13837
rect 5579 13772 5580 13836
rect 5644 13772 5645 13836
rect 5579 13771 5645 13772
rect 5582 12069 5642 13771
rect 5579 12068 5645 12069
rect 5579 12004 5580 12068
rect 5644 12004 5645 12068
rect 5579 12003 5645 12004
rect 5395 10980 5461 10981
rect 5395 10916 5396 10980
rect 5460 10916 5461 10980
rect 5395 10915 5461 10916
rect 5395 10844 5461 10845
rect 5395 10780 5396 10844
rect 5460 10780 5461 10844
rect 5395 10779 5461 10780
rect 5398 10301 5458 10779
rect 5395 10300 5461 10301
rect 5395 10236 5396 10300
rect 5460 10236 5461 10300
rect 5395 10235 5461 10236
rect 5766 9690 5826 15403
rect 5950 14109 6010 19075
rect 6142 18528 6462 19552
rect 6142 18464 6150 18528
rect 6214 18464 6230 18528
rect 6294 18464 6310 18528
rect 6374 18464 6390 18528
rect 6454 18464 6462 18528
rect 6142 17440 6462 18464
rect 6686 18053 6746 26691
rect 7051 25668 7117 25669
rect 7051 25604 7052 25668
rect 7116 25604 7117 25668
rect 7051 25603 7117 25604
rect 6867 25532 6933 25533
rect 6867 25468 6868 25532
rect 6932 25468 6933 25532
rect 6867 25467 6933 25468
rect 6870 22269 6930 25467
rect 7054 23901 7114 25603
rect 7051 23900 7117 23901
rect 7051 23836 7052 23900
rect 7116 23836 7117 23900
rect 7051 23835 7117 23836
rect 6867 22268 6933 22269
rect 6867 22204 6868 22268
rect 6932 22204 6933 22268
rect 6867 22203 6933 22204
rect 6867 21452 6933 21453
rect 6867 21388 6868 21452
rect 6932 21388 6933 21452
rect 6867 21387 6933 21388
rect 6870 19350 6930 21387
rect 7054 20093 7114 23835
rect 7238 23221 7298 27643
rect 7235 23220 7301 23221
rect 7235 23156 7236 23220
rect 7300 23156 7301 23220
rect 7235 23155 7301 23156
rect 7051 20092 7117 20093
rect 7051 20028 7052 20092
rect 7116 20028 7117 20092
rect 7051 20027 7117 20028
rect 6870 19290 7298 19350
rect 7051 18596 7117 18597
rect 7051 18532 7052 18596
rect 7116 18532 7117 18596
rect 7051 18531 7117 18532
rect 6683 18052 6749 18053
rect 6683 17988 6684 18052
rect 6748 17988 6749 18052
rect 6683 17987 6749 17988
rect 6142 17376 6150 17440
rect 6214 17376 6230 17440
rect 6294 17376 6310 17440
rect 6374 17376 6390 17440
rect 6454 17376 6462 17440
rect 6142 16352 6462 17376
rect 6867 16556 6933 16557
rect 6867 16492 6868 16556
rect 6932 16492 6933 16556
rect 6867 16491 6933 16492
rect 6142 16288 6150 16352
rect 6214 16288 6230 16352
rect 6294 16288 6310 16352
rect 6374 16288 6390 16352
rect 6454 16288 6462 16352
rect 6142 15264 6462 16288
rect 6683 15740 6749 15741
rect 6683 15676 6684 15740
rect 6748 15676 6749 15740
rect 6683 15675 6749 15676
rect 6142 15200 6150 15264
rect 6214 15200 6230 15264
rect 6294 15200 6310 15264
rect 6374 15200 6390 15264
rect 6454 15200 6462 15264
rect 6142 14176 6462 15200
rect 6142 14112 6150 14176
rect 6214 14112 6230 14176
rect 6294 14112 6310 14176
rect 6374 14112 6390 14176
rect 6454 14112 6462 14176
rect 5947 14108 6013 14109
rect 5947 14044 5948 14108
rect 6012 14044 6013 14108
rect 5947 14043 6013 14044
rect 5947 13292 6013 13293
rect 5947 13228 5948 13292
rect 6012 13228 6013 13292
rect 5947 13227 6013 13228
rect 5398 9630 5826 9690
rect 5211 8260 5277 8261
rect 5211 8196 5212 8260
rect 5276 8196 5277 8260
rect 5211 8195 5277 8196
rect 5398 7034 5458 9630
rect 5763 9076 5829 9077
rect 5763 9012 5764 9076
rect 5828 9012 5829 9076
rect 5763 9011 5829 9012
rect 5766 7581 5826 9011
rect 5579 7580 5645 7581
rect 5579 7516 5580 7580
rect 5644 7516 5645 7580
rect 5579 7515 5645 7516
rect 5763 7580 5829 7581
rect 5763 7516 5764 7580
rect 5828 7516 5829 7580
rect 5763 7515 5829 7516
rect 5214 6974 5458 7034
rect 5214 6901 5274 6974
rect 5211 6900 5277 6901
rect 5211 6836 5212 6900
rect 5276 6836 5277 6900
rect 5211 6835 5277 6836
rect 5395 6356 5461 6357
rect 5395 6292 5396 6356
rect 5460 6292 5461 6356
rect 5395 6291 5461 6292
rect 5027 5132 5093 5133
rect 5027 5068 5028 5132
rect 5092 5068 5093 5132
rect 5027 5067 5093 5068
rect 5211 5132 5277 5133
rect 5211 5068 5212 5132
rect 5276 5068 5277 5132
rect 5211 5067 5277 5068
rect 4659 4452 4725 4453
rect 4659 4388 4660 4452
rect 4724 4388 4725 4452
rect 4659 4387 4725 4388
rect 4107 4180 4173 4181
rect 4107 4116 4108 4180
rect 4172 4116 4173 4180
rect 4107 4115 4173 4116
rect 3543 3776 3551 3840
rect 3615 3776 3631 3840
rect 3695 3776 3711 3840
rect 3775 3776 3791 3840
rect 3855 3776 3863 3840
rect 3543 2752 3863 3776
rect 3543 2688 3551 2752
rect 3615 2688 3631 2752
rect 3695 2688 3711 2752
rect 3775 2688 3791 2752
rect 3855 2688 3863 2752
rect 2819 2548 2885 2549
rect 2819 2484 2820 2548
rect 2884 2484 2885 2548
rect 2819 2483 2885 2484
rect 3543 1664 3863 2688
rect 3543 1600 3551 1664
rect 3615 1600 3631 1664
rect 3695 1600 3711 1664
rect 3775 1600 3791 1664
rect 3855 1600 3863 1664
rect 1163 1324 1229 1325
rect 1163 1260 1164 1324
rect 1228 1260 1229 1324
rect 1163 1259 1229 1260
rect 3543 1040 3863 1600
rect 4110 1325 4170 4115
rect 5214 2277 5274 5067
rect 5398 2277 5458 6291
rect 5582 3909 5642 7515
rect 5766 6901 5826 7515
rect 5763 6900 5829 6901
rect 5763 6836 5764 6900
rect 5828 6836 5829 6900
rect 5763 6835 5829 6836
rect 5579 3908 5645 3909
rect 5579 3844 5580 3908
rect 5644 3844 5645 3908
rect 5579 3843 5645 3844
rect 5950 2821 6010 13227
rect 6142 13088 6462 14112
rect 6142 13024 6150 13088
rect 6214 13024 6230 13088
rect 6294 13024 6310 13088
rect 6374 13024 6390 13088
rect 6454 13024 6462 13088
rect 6142 12000 6462 13024
rect 6686 13018 6746 15675
rect 6870 14925 6930 16491
rect 7054 15605 7114 18531
rect 7238 18461 7298 19290
rect 7235 18460 7301 18461
rect 7235 18396 7236 18460
rect 7300 18396 7301 18460
rect 7235 18395 7301 18396
rect 7051 15604 7117 15605
rect 7051 15540 7052 15604
rect 7116 15540 7117 15604
rect 7051 15539 7117 15540
rect 6867 14924 6933 14925
rect 6867 14860 6868 14924
rect 6932 14860 6933 14924
rect 6867 14859 6933 14860
rect 7238 13701 7298 18395
rect 7235 13700 7301 13701
rect 7235 13636 7236 13700
rect 7300 13636 7301 13700
rect 7235 13635 7301 13636
rect 6686 12958 6930 13018
rect 6142 11936 6150 12000
rect 6214 11936 6230 12000
rect 6294 11936 6310 12000
rect 6374 11936 6390 12000
rect 6454 11936 6462 12000
rect 6142 10912 6462 11936
rect 6870 10981 6930 12958
rect 7235 12884 7301 12885
rect 7235 12820 7236 12884
rect 7300 12820 7301 12884
rect 7235 12819 7301 12820
rect 7051 12612 7117 12613
rect 7051 12548 7052 12612
rect 7116 12548 7117 12612
rect 7051 12547 7117 12548
rect 6867 10980 6933 10981
rect 6867 10916 6868 10980
rect 6932 10916 6933 10980
rect 6867 10915 6933 10916
rect 6142 10848 6150 10912
rect 6214 10848 6230 10912
rect 6294 10848 6310 10912
rect 6374 10848 6390 10912
rect 6454 10848 6462 10912
rect 6142 9824 6462 10848
rect 6142 9760 6150 9824
rect 6214 9760 6230 9824
rect 6294 9760 6310 9824
rect 6374 9760 6390 9824
rect 6454 9760 6462 9824
rect 6142 8736 6462 9760
rect 6142 8672 6150 8736
rect 6214 8672 6230 8736
rect 6294 8672 6310 8736
rect 6374 8672 6390 8736
rect 6454 8672 6462 8736
rect 6142 7648 6462 8672
rect 6867 8668 6933 8669
rect 6867 8604 6868 8668
rect 6932 8604 6933 8668
rect 6867 8603 6933 8604
rect 6142 7584 6150 7648
rect 6214 7584 6230 7648
rect 6294 7584 6310 7648
rect 6374 7584 6390 7648
rect 6454 7584 6462 7648
rect 6142 6560 6462 7584
rect 6142 6496 6150 6560
rect 6214 6496 6230 6560
rect 6294 6496 6310 6560
rect 6374 6496 6390 6560
rect 6454 6496 6462 6560
rect 6142 5472 6462 6496
rect 6142 5408 6150 5472
rect 6214 5408 6230 5472
rect 6294 5408 6310 5472
rect 6374 5408 6390 5472
rect 6454 5408 6462 5472
rect 6142 4384 6462 5408
rect 6142 4320 6150 4384
rect 6214 4320 6230 4384
rect 6294 4320 6310 4384
rect 6374 4320 6390 4384
rect 6454 4320 6462 4384
rect 6142 3296 6462 4320
rect 6142 3232 6150 3296
rect 6214 3232 6230 3296
rect 6294 3232 6310 3296
rect 6374 3232 6390 3296
rect 6454 3232 6462 3296
rect 5947 2820 6013 2821
rect 5947 2756 5948 2820
rect 6012 2756 6013 2820
rect 5947 2755 6013 2756
rect 5211 2276 5277 2277
rect 5211 2212 5212 2276
rect 5276 2212 5277 2276
rect 5211 2211 5277 2212
rect 5395 2276 5461 2277
rect 5395 2212 5396 2276
rect 5460 2212 5461 2276
rect 5395 2211 5461 2212
rect 6142 2208 6462 3232
rect 6870 2413 6930 8603
rect 7054 7037 7114 12547
rect 7051 7036 7117 7037
rect 7051 6972 7052 7036
rect 7116 6972 7117 7036
rect 7051 6971 7117 6972
rect 6867 2412 6933 2413
rect 6867 2348 6868 2412
rect 6932 2348 6933 2412
rect 6867 2347 6933 2348
rect 6142 2144 6150 2208
rect 6214 2144 6230 2208
rect 6294 2144 6310 2208
rect 6374 2144 6390 2208
rect 6454 2144 6462 2208
rect 4107 1324 4173 1325
rect 4107 1260 4108 1324
rect 4172 1260 4173 1324
rect 4107 1259 4173 1260
rect 6142 1120 6462 2144
rect 7238 1325 7298 12819
rect 7422 1869 7482 41515
rect 8155 38452 8221 38453
rect 8155 38388 8156 38452
rect 8220 38388 8221 38452
rect 8155 38387 8221 38388
rect 7971 37364 8037 37365
rect 7971 37300 7972 37364
rect 8036 37300 8037 37364
rect 7971 37299 8037 37300
rect 7787 37092 7853 37093
rect 7787 37028 7788 37092
rect 7852 37028 7853 37092
rect 7787 37027 7853 37028
rect 7603 36004 7669 36005
rect 7603 35940 7604 36004
rect 7668 35940 7669 36004
rect 7603 35939 7669 35940
rect 7606 24445 7666 35939
rect 7790 31245 7850 37027
rect 7787 31244 7853 31245
rect 7787 31180 7788 31244
rect 7852 31180 7853 31244
rect 7787 31179 7853 31180
rect 7787 27708 7853 27709
rect 7787 27644 7788 27708
rect 7852 27644 7853 27708
rect 7787 27643 7853 27644
rect 7790 25941 7850 27643
rect 7787 25940 7853 25941
rect 7787 25876 7788 25940
rect 7852 25876 7853 25940
rect 7787 25875 7853 25876
rect 7603 24444 7669 24445
rect 7603 24380 7604 24444
rect 7668 24380 7669 24444
rect 7603 24379 7669 24380
rect 7603 24308 7669 24309
rect 7603 24244 7604 24308
rect 7668 24244 7669 24308
rect 7603 24243 7669 24244
rect 7606 19685 7666 24243
rect 7787 22948 7853 22949
rect 7787 22884 7788 22948
rect 7852 22884 7853 22948
rect 7787 22883 7853 22884
rect 7790 22405 7850 22883
rect 7787 22404 7853 22405
rect 7787 22340 7788 22404
rect 7852 22340 7853 22404
rect 7787 22339 7853 22340
rect 7603 19684 7669 19685
rect 7603 19620 7604 19684
rect 7668 19620 7669 19684
rect 7603 19619 7669 19620
rect 7603 17508 7669 17509
rect 7603 17444 7604 17508
rect 7668 17444 7669 17508
rect 7603 17443 7669 17444
rect 7606 12613 7666 17443
rect 7790 16013 7850 22339
rect 7787 16012 7853 16013
rect 7787 15948 7788 16012
rect 7852 15948 7853 16012
rect 7787 15947 7853 15948
rect 7603 12612 7669 12613
rect 7603 12548 7604 12612
rect 7668 12548 7669 12612
rect 7603 12547 7669 12548
rect 7790 12477 7850 15947
rect 7787 12476 7853 12477
rect 7787 12412 7788 12476
rect 7852 12412 7853 12476
rect 7787 12411 7853 12412
rect 7603 6900 7669 6901
rect 7603 6836 7604 6900
rect 7668 6836 7669 6900
rect 7603 6835 7669 6836
rect 7606 2549 7666 6835
rect 7974 3637 8034 37299
rect 8158 31789 8218 38387
rect 8342 35869 8402 42195
rect 8741 41920 9061 42944
rect 11340 43552 11660 43568
rect 11340 43488 11348 43552
rect 11412 43488 11428 43552
rect 11492 43488 11508 43552
rect 11572 43488 11588 43552
rect 11652 43488 11660 43552
rect 11340 42464 11660 43488
rect 11835 43212 11901 43213
rect 11835 43148 11836 43212
rect 11900 43148 11901 43212
rect 11835 43147 11901 43148
rect 11340 42400 11348 42464
rect 11412 42400 11428 42464
rect 11492 42400 11508 42464
rect 11572 42400 11588 42464
rect 11652 42400 11660 42464
rect 9259 42396 9325 42397
rect 9259 42332 9260 42396
rect 9324 42332 9325 42396
rect 9259 42331 9325 42332
rect 9443 42396 9509 42397
rect 9443 42332 9444 42396
rect 9508 42332 9509 42396
rect 9443 42331 9509 42332
rect 8741 41856 8749 41920
rect 8813 41856 8829 41920
rect 8893 41856 8909 41920
rect 8973 41856 8989 41920
rect 9053 41856 9061 41920
rect 8741 40832 9061 41856
rect 8741 40768 8749 40832
rect 8813 40768 8829 40832
rect 8893 40768 8909 40832
rect 8973 40768 8989 40832
rect 9053 40768 9061 40832
rect 8741 39744 9061 40768
rect 8741 39680 8749 39744
rect 8813 39680 8829 39744
rect 8893 39680 8909 39744
rect 8973 39680 8989 39744
rect 9053 39680 9061 39744
rect 8741 38656 9061 39680
rect 8741 38592 8749 38656
rect 8813 38592 8829 38656
rect 8893 38592 8909 38656
rect 8973 38592 8989 38656
rect 9053 38592 9061 38656
rect 8741 37568 9061 38592
rect 8741 37504 8749 37568
rect 8813 37504 8829 37568
rect 8893 37504 8909 37568
rect 8973 37504 8989 37568
rect 9053 37504 9061 37568
rect 8523 37228 8589 37229
rect 8523 37164 8524 37228
rect 8588 37164 8589 37228
rect 8523 37163 8589 37164
rect 8339 35868 8405 35869
rect 8339 35804 8340 35868
rect 8404 35804 8405 35868
rect 8339 35803 8405 35804
rect 8339 33012 8405 33013
rect 8339 32948 8340 33012
rect 8404 32948 8405 33012
rect 8339 32947 8405 32948
rect 8155 31788 8221 31789
rect 8155 31724 8156 31788
rect 8220 31724 8221 31788
rect 8155 31723 8221 31724
rect 8155 28388 8221 28389
rect 8155 28324 8156 28388
rect 8220 28324 8221 28388
rect 8155 28323 8221 28324
rect 8158 18325 8218 28323
rect 8342 20093 8402 32947
rect 8526 31381 8586 37163
rect 8741 36480 9061 37504
rect 8741 36416 8749 36480
rect 8813 36416 8829 36480
rect 8893 36416 8909 36480
rect 8973 36416 8989 36480
rect 9053 36416 9061 36480
rect 8741 35392 9061 36416
rect 8741 35328 8749 35392
rect 8813 35328 8829 35392
rect 8893 35328 8909 35392
rect 8973 35328 8989 35392
rect 9053 35328 9061 35392
rect 8741 34304 9061 35328
rect 8741 34240 8749 34304
rect 8813 34240 8829 34304
rect 8893 34240 8909 34304
rect 8973 34240 8989 34304
rect 9053 34240 9061 34304
rect 8741 33216 9061 34240
rect 8741 33152 8749 33216
rect 8813 33152 8829 33216
rect 8893 33152 8909 33216
rect 8973 33152 8989 33216
rect 9053 33152 9061 33216
rect 8741 32128 9061 33152
rect 8741 32064 8749 32128
rect 8813 32064 8829 32128
rect 8893 32064 8909 32128
rect 8973 32064 8989 32128
rect 9053 32064 9061 32128
rect 8523 31380 8589 31381
rect 8523 31316 8524 31380
rect 8588 31316 8589 31380
rect 8523 31315 8589 31316
rect 8741 31040 9061 32064
rect 8741 30976 8749 31040
rect 8813 30976 8829 31040
rect 8893 30976 8909 31040
rect 8973 30976 8989 31040
rect 9053 30976 9061 31040
rect 8741 29952 9061 30976
rect 8741 29888 8749 29952
rect 8813 29888 8829 29952
rect 8893 29888 8909 29952
rect 8973 29888 8989 29952
rect 9053 29888 9061 29952
rect 8741 28864 9061 29888
rect 8741 28800 8749 28864
rect 8813 28800 8829 28864
rect 8893 28800 8909 28864
rect 8973 28800 8989 28864
rect 9053 28800 9061 28864
rect 8523 28796 8589 28797
rect 8523 28732 8524 28796
rect 8588 28732 8589 28796
rect 8523 28731 8589 28732
rect 8526 27165 8586 28731
rect 8741 27776 9061 28800
rect 8741 27712 8749 27776
rect 8813 27712 8829 27776
rect 8893 27712 8909 27776
rect 8973 27712 8989 27776
rect 9053 27712 9061 27776
rect 8523 27164 8589 27165
rect 8523 27100 8524 27164
rect 8588 27100 8589 27164
rect 8523 27099 8589 27100
rect 8523 27028 8589 27029
rect 8523 26964 8524 27028
rect 8588 26964 8589 27028
rect 8523 26963 8589 26964
rect 8526 23493 8586 26963
rect 8741 26688 9061 27712
rect 8741 26624 8749 26688
rect 8813 26624 8829 26688
rect 8893 26624 8909 26688
rect 8973 26624 8989 26688
rect 9053 26624 9061 26688
rect 8741 25600 9061 26624
rect 8741 25536 8749 25600
rect 8813 25536 8829 25600
rect 8893 25536 8909 25600
rect 8973 25536 8989 25600
rect 9053 25536 9061 25600
rect 8741 24512 9061 25536
rect 8741 24448 8749 24512
rect 8813 24448 8829 24512
rect 8893 24448 8909 24512
rect 8973 24448 8989 24512
rect 9053 24448 9061 24512
rect 8523 23492 8589 23493
rect 8523 23428 8524 23492
rect 8588 23428 8589 23492
rect 8523 23427 8589 23428
rect 8339 20092 8405 20093
rect 8339 20028 8340 20092
rect 8404 20028 8405 20092
rect 8339 20027 8405 20028
rect 8526 19821 8586 23427
rect 8741 23424 9061 24448
rect 8741 23360 8749 23424
rect 8813 23360 8829 23424
rect 8893 23360 8909 23424
rect 8973 23360 8989 23424
rect 9053 23360 9061 23424
rect 8741 22336 9061 23360
rect 8741 22272 8749 22336
rect 8813 22272 8829 22336
rect 8893 22272 8909 22336
rect 8973 22272 8989 22336
rect 9053 22272 9061 22336
rect 8741 21248 9061 22272
rect 8741 21184 8749 21248
rect 8813 21184 8829 21248
rect 8893 21184 8909 21248
rect 8973 21184 8989 21248
rect 9053 21184 9061 21248
rect 8741 20160 9061 21184
rect 8741 20096 8749 20160
rect 8813 20096 8829 20160
rect 8893 20096 8909 20160
rect 8973 20096 8989 20160
rect 9053 20096 9061 20160
rect 8523 19820 8589 19821
rect 8523 19756 8524 19820
rect 8588 19756 8589 19820
rect 8523 19755 8589 19756
rect 8741 19072 9061 20096
rect 8741 19008 8749 19072
rect 8813 19008 8829 19072
rect 8893 19008 8909 19072
rect 8973 19008 8989 19072
rect 9053 19008 9061 19072
rect 8155 18324 8221 18325
rect 8155 18260 8156 18324
rect 8220 18260 8221 18324
rect 8155 18259 8221 18260
rect 8741 17984 9061 19008
rect 8741 17920 8749 17984
rect 8813 17920 8829 17984
rect 8893 17920 8909 17984
rect 8973 17920 8989 17984
rect 9053 17920 9061 17984
rect 8741 16896 9061 17920
rect 8741 16832 8749 16896
rect 8813 16832 8829 16896
rect 8893 16832 8909 16896
rect 8973 16832 8989 16896
rect 9053 16832 9061 16896
rect 8155 16692 8221 16693
rect 8155 16628 8156 16692
rect 8220 16628 8221 16692
rect 8155 16627 8221 16628
rect 8158 10845 8218 16627
rect 8741 15808 9061 16832
rect 8741 15744 8749 15808
rect 8813 15744 8829 15808
rect 8893 15744 8909 15808
rect 8973 15744 8989 15808
rect 9053 15744 9061 15808
rect 8339 15196 8405 15197
rect 8339 15132 8340 15196
rect 8404 15132 8405 15196
rect 8339 15131 8405 15132
rect 8155 10844 8221 10845
rect 8155 10780 8156 10844
rect 8220 10780 8221 10844
rect 8155 10779 8221 10780
rect 8342 9757 8402 15131
rect 8741 14720 9061 15744
rect 8741 14656 8749 14720
rect 8813 14656 8829 14720
rect 8893 14656 8909 14720
rect 8973 14656 8989 14720
rect 9053 14656 9061 14720
rect 8741 13632 9061 14656
rect 8741 13568 8749 13632
rect 8813 13568 8829 13632
rect 8893 13568 8909 13632
rect 8973 13568 8989 13632
rect 9053 13568 9061 13632
rect 8741 12544 9061 13568
rect 8741 12480 8749 12544
rect 8813 12480 8829 12544
rect 8893 12480 8909 12544
rect 8973 12480 8989 12544
rect 9053 12480 9061 12544
rect 8741 11456 9061 12480
rect 8741 11392 8749 11456
rect 8813 11392 8829 11456
rect 8893 11392 8909 11456
rect 8973 11392 8989 11456
rect 9053 11392 9061 11456
rect 8741 10368 9061 11392
rect 8741 10304 8749 10368
rect 8813 10304 8829 10368
rect 8893 10304 8909 10368
rect 8973 10304 8989 10368
rect 9053 10304 9061 10368
rect 8339 9756 8405 9757
rect 8339 9692 8340 9756
rect 8404 9692 8405 9756
rect 8339 9691 8405 9692
rect 8741 9280 9061 10304
rect 8741 9216 8749 9280
rect 8813 9216 8829 9280
rect 8893 9216 8909 9280
rect 8973 9216 8989 9280
rect 9053 9216 9061 9280
rect 8339 8396 8405 8397
rect 8339 8332 8340 8396
rect 8404 8332 8405 8396
rect 8339 8331 8405 8332
rect 8155 4588 8221 4589
rect 8155 4524 8156 4588
rect 8220 4524 8221 4588
rect 8155 4523 8221 4524
rect 7971 3636 8037 3637
rect 7971 3572 7972 3636
rect 8036 3572 8037 3636
rect 7971 3571 8037 3572
rect 8158 2685 8218 4523
rect 8342 3229 8402 8331
rect 8741 8192 9061 9216
rect 8741 8128 8749 8192
rect 8813 8128 8829 8192
rect 8893 8128 8909 8192
rect 8973 8128 8989 8192
rect 9053 8128 9061 8192
rect 8741 7104 9061 8128
rect 8741 7040 8749 7104
rect 8813 7040 8829 7104
rect 8893 7040 8909 7104
rect 8973 7040 8989 7104
rect 9053 7040 9061 7104
rect 8741 6016 9061 7040
rect 8741 5952 8749 6016
rect 8813 5952 8829 6016
rect 8893 5952 8909 6016
rect 8973 5952 8989 6016
rect 9053 5952 9061 6016
rect 8741 4928 9061 5952
rect 8741 4864 8749 4928
rect 8813 4864 8829 4928
rect 8893 4864 8909 4928
rect 8973 4864 8989 4928
rect 9053 4864 9061 4928
rect 8741 3840 9061 4864
rect 8741 3776 8749 3840
rect 8813 3776 8829 3840
rect 8893 3776 8909 3840
rect 8973 3776 8989 3840
rect 9053 3776 9061 3840
rect 8339 3228 8405 3229
rect 8339 3164 8340 3228
rect 8404 3164 8405 3228
rect 8339 3163 8405 3164
rect 8523 3228 8589 3229
rect 8523 3164 8524 3228
rect 8588 3164 8589 3228
rect 8523 3163 8589 3164
rect 8155 2684 8221 2685
rect 8155 2620 8156 2684
rect 8220 2620 8221 2684
rect 8155 2619 8221 2620
rect 7603 2548 7669 2549
rect 7603 2484 7604 2548
rect 7668 2484 7669 2548
rect 7603 2483 7669 2484
rect 7419 1868 7485 1869
rect 7419 1804 7420 1868
rect 7484 1804 7485 1868
rect 7419 1803 7485 1804
rect 7235 1324 7301 1325
rect 7235 1260 7236 1324
rect 7300 1260 7301 1324
rect 7235 1259 7301 1260
rect 6142 1056 6150 1120
rect 6214 1056 6230 1120
rect 6294 1056 6310 1120
rect 6374 1056 6390 1120
rect 6454 1056 6462 1120
rect 6142 1040 6462 1056
rect 8526 101 8586 3163
rect 8741 2752 9061 3776
rect 9262 2821 9322 42331
rect 9446 35461 9506 42331
rect 10179 41988 10245 41989
rect 10179 41924 10180 41988
rect 10244 41924 10245 41988
rect 10179 41923 10245 41924
rect 9811 37772 9877 37773
rect 9811 37708 9812 37772
rect 9876 37708 9877 37772
rect 9811 37707 9877 37708
rect 9443 35460 9509 35461
rect 9443 35396 9444 35460
rect 9508 35396 9509 35460
rect 9443 35395 9509 35396
rect 9627 32196 9693 32197
rect 9627 32132 9628 32196
rect 9692 32132 9693 32196
rect 9627 32131 9693 32132
rect 9630 31770 9690 32131
rect 9446 31710 9690 31770
rect 9446 29477 9506 31710
rect 9627 30836 9693 30837
rect 9627 30772 9628 30836
rect 9692 30772 9693 30836
rect 9627 30771 9693 30772
rect 9443 29476 9509 29477
rect 9443 29412 9444 29476
rect 9508 29412 9509 29476
rect 9443 29411 9509 29412
rect 9443 27164 9509 27165
rect 9443 27100 9444 27164
rect 9508 27100 9509 27164
rect 9443 27099 9509 27100
rect 9446 20637 9506 27099
rect 9630 24173 9690 30771
rect 9814 30429 9874 37707
rect 9995 36004 10061 36005
rect 9995 35940 9996 36004
rect 10060 35940 10061 36004
rect 9995 35939 10061 35940
rect 9998 32197 10058 35939
rect 9995 32196 10061 32197
rect 9995 32132 9996 32196
rect 10060 32132 10061 32196
rect 9995 32131 10061 32132
rect 9811 30428 9877 30429
rect 9811 30364 9812 30428
rect 9876 30364 9877 30428
rect 9811 30363 9877 30364
rect 10182 28661 10242 41923
rect 11340 41376 11660 42400
rect 11340 41312 11348 41376
rect 11412 41312 11428 41376
rect 11492 41312 11508 41376
rect 11572 41312 11588 41376
rect 11652 41312 11660 41376
rect 11838 41430 11898 43147
rect 13939 43008 14259 43568
rect 13939 42944 13947 43008
rect 14011 42944 14027 43008
rect 14091 42944 14107 43008
rect 14171 42944 14187 43008
rect 14251 42944 14259 43008
rect 13123 42940 13189 42941
rect 13123 42876 13124 42940
rect 13188 42876 13189 42940
rect 13123 42875 13189 42876
rect 11838 41370 12082 41430
rect 11340 40288 11660 41312
rect 11340 40224 11348 40288
rect 11412 40224 11428 40288
rect 11492 40224 11508 40288
rect 11572 40224 11588 40288
rect 11652 40224 11660 40288
rect 11340 39200 11660 40224
rect 11340 39136 11348 39200
rect 11412 39136 11428 39200
rect 11492 39136 11508 39200
rect 11572 39136 11588 39200
rect 11652 39136 11660 39200
rect 11340 38112 11660 39136
rect 11340 38048 11348 38112
rect 11412 38048 11428 38112
rect 11492 38048 11508 38112
rect 11572 38048 11588 38112
rect 11652 38048 11660 38112
rect 11340 37024 11660 38048
rect 11340 36960 11348 37024
rect 11412 36960 11428 37024
rect 11492 36960 11508 37024
rect 11572 36960 11588 37024
rect 11652 36960 11660 37024
rect 10731 36004 10797 36005
rect 10731 35940 10732 36004
rect 10796 35940 10797 36004
rect 10731 35939 10797 35940
rect 10363 32060 10429 32061
rect 10363 31996 10364 32060
rect 10428 31996 10429 32060
rect 10363 31995 10429 31996
rect 10179 28660 10245 28661
rect 10179 28596 10180 28660
rect 10244 28596 10245 28660
rect 10179 28595 10245 28596
rect 10179 26348 10245 26349
rect 10179 26284 10180 26348
rect 10244 26284 10245 26348
rect 10179 26283 10245 26284
rect 9811 24852 9877 24853
rect 9811 24788 9812 24852
rect 9876 24788 9877 24852
rect 9811 24787 9877 24788
rect 9627 24172 9693 24173
rect 9627 24108 9628 24172
rect 9692 24108 9693 24172
rect 9627 24107 9693 24108
rect 9814 21181 9874 24787
rect 10182 22405 10242 26283
rect 10179 22404 10245 22405
rect 10179 22340 10180 22404
rect 10244 22340 10245 22404
rect 10179 22339 10245 22340
rect 9811 21180 9877 21181
rect 9811 21116 9812 21180
rect 9876 21116 9877 21180
rect 9811 21115 9877 21116
rect 9443 20636 9509 20637
rect 9443 20572 9444 20636
rect 9508 20572 9509 20636
rect 9443 20571 9509 20572
rect 9814 19350 9874 21115
rect 9446 19290 9874 19350
rect 9446 17917 9506 19290
rect 9443 17916 9509 17917
rect 9443 17852 9444 17916
rect 9508 17852 9509 17916
rect 9443 17851 9509 17852
rect 9446 13565 9506 17851
rect 10182 16557 10242 22339
rect 10366 20637 10426 31995
rect 10547 29068 10613 29069
rect 10547 29004 10548 29068
rect 10612 29004 10613 29068
rect 10547 29003 10613 29004
rect 10550 27165 10610 29003
rect 10547 27164 10613 27165
rect 10547 27100 10548 27164
rect 10612 27100 10613 27164
rect 10547 27099 10613 27100
rect 10547 23900 10613 23901
rect 10547 23836 10548 23900
rect 10612 23836 10613 23900
rect 10547 23835 10613 23836
rect 10550 21453 10610 23835
rect 10547 21452 10613 21453
rect 10547 21388 10548 21452
rect 10612 21388 10613 21452
rect 10547 21387 10613 21388
rect 10363 20636 10429 20637
rect 10363 20572 10364 20636
rect 10428 20572 10429 20636
rect 10363 20571 10429 20572
rect 10547 18596 10613 18597
rect 10547 18532 10548 18596
rect 10612 18532 10613 18596
rect 10547 18531 10613 18532
rect 10550 17098 10610 18531
rect 10734 17509 10794 35939
rect 11340 35936 11660 36960
rect 11340 35872 11348 35936
rect 11412 35872 11428 35936
rect 11492 35872 11508 35936
rect 11572 35872 11588 35936
rect 11652 35872 11660 35936
rect 11099 35868 11165 35869
rect 11099 35804 11100 35868
rect 11164 35804 11165 35868
rect 11099 35803 11165 35804
rect 10915 34644 10981 34645
rect 10915 34580 10916 34644
rect 10980 34580 10981 34644
rect 10915 34579 10981 34580
rect 10918 30157 10978 34579
rect 10915 30156 10981 30157
rect 10915 30092 10916 30156
rect 10980 30092 10981 30156
rect 10915 30091 10981 30092
rect 11102 29341 11162 35803
rect 11340 34848 11660 35872
rect 11340 34784 11348 34848
rect 11412 34784 11428 34848
rect 11492 34784 11508 34848
rect 11572 34784 11588 34848
rect 11652 34784 11660 34848
rect 11340 33760 11660 34784
rect 11835 34644 11901 34645
rect 11835 34580 11836 34644
rect 11900 34580 11901 34644
rect 11835 34579 11901 34580
rect 11340 33696 11348 33760
rect 11412 33696 11428 33760
rect 11492 33696 11508 33760
rect 11572 33696 11588 33760
rect 11652 33696 11660 33760
rect 11340 32672 11660 33696
rect 11340 32608 11348 32672
rect 11412 32608 11428 32672
rect 11492 32608 11508 32672
rect 11572 32608 11588 32672
rect 11652 32608 11660 32672
rect 11340 31584 11660 32608
rect 11340 31520 11348 31584
rect 11412 31520 11428 31584
rect 11492 31520 11508 31584
rect 11572 31520 11588 31584
rect 11652 31520 11660 31584
rect 11340 30496 11660 31520
rect 11340 30432 11348 30496
rect 11412 30432 11428 30496
rect 11492 30432 11508 30496
rect 11572 30432 11588 30496
rect 11652 30432 11660 30496
rect 11340 29408 11660 30432
rect 11340 29344 11348 29408
rect 11412 29344 11428 29408
rect 11492 29344 11508 29408
rect 11572 29344 11588 29408
rect 11652 29344 11660 29408
rect 11099 29340 11165 29341
rect 11099 29276 11100 29340
rect 11164 29276 11165 29340
rect 11099 29275 11165 29276
rect 11340 28320 11660 29344
rect 11340 28256 11348 28320
rect 11412 28256 11428 28320
rect 11492 28256 11508 28320
rect 11572 28256 11588 28320
rect 11652 28256 11660 28320
rect 11340 27232 11660 28256
rect 11340 27168 11348 27232
rect 11412 27168 11428 27232
rect 11492 27168 11508 27232
rect 11572 27168 11588 27232
rect 11652 27168 11660 27232
rect 11340 26144 11660 27168
rect 11340 26080 11348 26144
rect 11412 26080 11428 26144
rect 11492 26080 11508 26144
rect 11572 26080 11588 26144
rect 11652 26080 11660 26144
rect 11340 25056 11660 26080
rect 11340 24992 11348 25056
rect 11412 24992 11428 25056
rect 11492 24992 11508 25056
rect 11572 24992 11588 25056
rect 11652 24992 11660 25056
rect 11340 23968 11660 24992
rect 11340 23904 11348 23968
rect 11412 23904 11428 23968
rect 11492 23904 11508 23968
rect 11572 23904 11588 23968
rect 11652 23904 11660 23968
rect 11099 23628 11165 23629
rect 11099 23564 11100 23628
rect 11164 23564 11165 23628
rect 11099 23563 11165 23564
rect 11102 22677 11162 23563
rect 11340 22880 11660 23904
rect 11340 22816 11348 22880
rect 11412 22816 11428 22880
rect 11492 22816 11508 22880
rect 11572 22816 11588 22880
rect 11652 22816 11660 22880
rect 11099 22676 11165 22677
rect 11099 22612 11100 22676
rect 11164 22612 11165 22676
rect 11099 22611 11165 22612
rect 10915 22268 10981 22269
rect 10915 22204 10916 22268
rect 10980 22204 10981 22268
rect 10915 22203 10981 22204
rect 10731 17508 10797 17509
rect 10731 17444 10732 17508
rect 10796 17444 10797 17508
rect 10731 17443 10797 17444
rect 10550 17038 10794 17098
rect 10547 16692 10613 16693
rect 10547 16628 10548 16692
rect 10612 16628 10613 16692
rect 10547 16627 10613 16628
rect 10179 16556 10245 16557
rect 10179 16492 10180 16556
rect 10244 16492 10245 16556
rect 10179 16491 10245 16492
rect 10182 15605 10242 16491
rect 10179 15604 10245 15605
rect 10179 15540 10180 15604
rect 10244 15540 10245 15604
rect 10179 15539 10245 15540
rect 9627 14924 9693 14925
rect 9627 14860 9628 14924
rect 9692 14860 9693 14924
rect 9627 14859 9693 14860
rect 9443 13564 9509 13565
rect 9443 13500 9444 13564
rect 9508 13500 9509 13564
rect 9443 13499 9509 13500
rect 9443 13292 9509 13293
rect 9443 13228 9444 13292
rect 9508 13228 9509 13292
rect 9443 13227 9509 13228
rect 9446 8397 9506 13227
rect 9630 8533 9690 14859
rect 10179 11796 10245 11797
rect 10179 11732 10180 11796
rect 10244 11732 10245 11796
rect 10179 11731 10245 11732
rect 10363 11796 10429 11797
rect 10363 11732 10364 11796
rect 10428 11732 10429 11796
rect 10363 11731 10429 11732
rect 9627 8532 9693 8533
rect 9627 8468 9628 8532
rect 9692 8468 9693 8532
rect 9627 8467 9693 8468
rect 9443 8396 9509 8397
rect 9443 8332 9444 8396
rect 9508 8332 9509 8396
rect 9443 8331 9509 8332
rect 10182 7989 10242 11731
rect 10179 7988 10245 7989
rect 10179 7924 10180 7988
rect 10244 7924 10245 7988
rect 10179 7923 10245 7924
rect 10182 6221 10242 7923
rect 10366 6629 10426 11731
rect 10363 6628 10429 6629
rect 10363 6564 10364 6628
rect 10428 6564 10429 6628
rect 10363 6563 10429 6564
rect 10179 6220 10245 6221
rect 10179 6156 10180 6220
rect 10244 6156 10245 6220
rect 10179 6155 10245 6156
rect 9627 5676 9693 5677
rect 9627 5612 9628 5676
rect 9692 5612 9693 5676
rect 9627 5611 9693 5612
rect 9259 2820 9325 2821
rect 9259 2756 9260 2820
rect 9324 2756 9325 2820
rect 9259 2755 9325 2756
rect 8741 2688 8749 2752
rect 8813 2688 8829 2752
rect 8893 2688 8909 2752
rect 8973 2688 8989 2752
rect 9053 2688 9061 2752
rect 8741 1664 9061 2688
rect 8741 1600 8749 1664
rect 8813 1600 8829 1664
rect 8893 1600 8909 1664
rect 8973 1600 8989 1664
rect 9053 1600 9061 1664
rect 8741 1040 9061 1600
rect 9630 917 9690 5611
rect 10550 4453 10610 16627
rect 10734 10573 10794 17038
rect 10918 16693 10978 22203
rect 11099 22132 11165 22133
rect 11099 22068 11100 22132
rect 11164 22068 11165 22132
rect 11099 22067 11165 22068
rect 10915 16692 10981 16693
rect 10915 16628 10916 16692
rect 10980 16628 10981 16692
rect 10915 16627 10981 16628
rect 10915 16284 10981 16285
rect 10915 16220 10916 16284
rect 10980 16220 10981 16284
rect 10915 16219 10981 16220
rect 10918 10981 10978 16219
rect 11102 12477 11162 22067
rect 11340 21792 11660 22816
rect 11838 21997 11898 34579
rect 12022 33149 12082 41370
rect 12571 38452 12637 38453
rect 12571 38388 12572 38452
rect 12636 38388 12637 38452
rect 12571 38387 12637 38388
rect 12019 33148 12085 33149
rect 12019 33084 12020 33148
rect 12084 33084 12085 33148
rect 12019 33083 12085 33084
rect 12203 30564 12269 30565
rect 12203 30500 12204 30564
rect 12268 30500 12269 30564
rect 12203 30499 12269 30500
rect 12206 24853 12266 30499
rect 12387 26756 12453 26757
rect 12387 26692 12388 26756
rect 12452 26692 12453 26756
rect 12387 26691 12453 26692
rect 12019 24852 12085 24853
rect 12019 24788 12020 24852
rect 12084 24788 12085 24852
rect 12019 24787 12085 24788
rect 12203 24852 12269 24853
rect 12203 24788 12204 24852
rect 12268 24788 12269 24852
rect 12203 24787 12269 24788
rect 11835 21996 11901 21997
rect 11835 21932 11836 21996
rect 11900 21932 11901 21996
rect 11835 21931 11901 21932
rect 11340 21728 11348 21792
rect 11412 21728 11428 21792
rect 11492 21728 11508 21792
rect 11572 21728 11588 21792
rect 11652 21728 11660 21792
rect 11340 20704 11660 21728
rect 11340 20640 11348 20704
rect 11412 20640 11428 20704
rect 11492 20640 11508 20704
rect 11572 20640 11588 20704
rect 11652 20640 11660 20704
rect 11340 19616 11660 20640
rect 11340 19552 11348 19616
rect 11412 19552 11428 19616
rect 11492 19552 11508 19616
rect 11572 19552 11588 19616
rect 11652 19552 11660 19616
rect 11340 18528 11660 19552
rect 11340 18464 11348 18528
rect 11412 18464 11428 18528
rect 11492 18464 11508 18528
rect 11572 18464 11588 18528
rect 11652 18464 11660 18528
rect 11340 17440 11660 18464
rect 11340 17376 11348 17440
rect 11412 17376 11428 17440
rect 11492 17376 11508 17440
rect 11572 17376 11588 17440
rect 11652 17376 11660 17440
rect 11340 16352 11660 17376
rect 11340 16288 11348 16352
rect 11412 16288 11428 16352
rect 11492 16288 11508 16352
rect 11572 16288 11588 16352
rect 11652 16288 11660 16352
rect 11340 15264 11660 16288
rect 11835 16148 11901 16149
rect 11835 16084 11836 16148
rect 11900 16084 11901 16148
rect 11835 16083 11901 16084
rect 11340 15200 11348 15264
rect 11412 15200 11428 15264
rect 11492 15200 11508 15264
rect 11572 15200 11588 15264
rect 11652 15200 11660 15264
rect 11340 14176 11660 15200
rect 11340 14112 11348 14176
rect 11412 14112 11428 14176
rect 11492 14112 11508 14176
rect 11572 14112 11588 14176
rect 11652 14112 11660 14176
rect 11340 13088 11660 14112
rect 11340 13024 11348 13088
rect 11412 13024 11428 13088
rect 11492 13024 11508 13088
rect 11572 13024 11588 13088
rect 11652 13024 11660 13088
rect 11099 12476 11165 12477
rect 11099 12412 11100 12476
rect 11164 12412 11165 12476
rect 11099 12411 11165 12412
rect 11099 12204 11165 12205
rect 11099 12140 11100 12204
rect 11164 12140 11165 12204
rect 11099 12139 11165 12140
rect 10915 10980 10981 10981
rect 10915 10916 10916 10980
rect 10980 10916 10981 10980
rect 10915 10915 10981 10916
rect 10731 10572 10797 10573
rect 10731 10508 10732 10572
rect 10796 10508 10797 10572
rect 10731 10507 10797 10508
rect 11102 7309 11162 12139
rect 11340 12000 11660 13024
rect 11838 12205 11898 16083
rect 12022 12746 12082 24787
rect 12390 22130 12450 26691
rect 12206 22070 12450 22130
rect 12206 21725 12266 22070
rect 12203 21724 12269 21725
rect 12203 21660 12204 21724
rect 12268 21660 12269 21724
rect 12203 21659 12269 21660
rect 12203 21452 12269 21453
rect 12203 21388 12204 21452
rect 12268 21388 12269 21452
rect 12203 21387 12269 21388
rect 12206 14381 12266 21387
rect 12574 20773 12634 38387
rect 12755 33556 12821 33557
rect 12755 33492 12756 33556
rect 12820 33492 12821 33556
rect 12755 33491 12821 33492
rect 12571 20772 12637 20773
rect 12571 20708 12572 20772
rect 12636 20708 12637 20772
rect 12571 20707 12637 20708
rect 12203 14380 12269 14381
rect 12203 14316 12204 14380
rect 12268 14316 12269 14380
rect 12203 14315 12269 14316
rect 12571 13700 12637 13701
rect 12571 13636 12572 13700
rect 12636 13636 12637 13700
rect 12571 13635 12637 13636
rect 12022 12686 12266 12746
rect 12019 12612 12085 12613
rect 12019 12548 12020 12612
rect 12084 12548 12085 12612
rect 12019 12547 12085 12548
rect 11835 12204 11901 12205
rect 11835 12140 11836 12204
rect 11900 12140 11901 12204
rect 11835 12139 11901 12140
rect 11340 11936 11348 12000
rect 11412 11936 11428 12000
rect 11492 11936 11508 12000
rect 11572 11936 11588 12000
rect 11652 11936 11660 12000
rect 11340 10912 11660 11936
rect 11340 10848 11348 10912
rect 11412 10848 11428 10912
rect 11492 10848 11508 10912
rect 11572 10848 11588 10912
rect 11652 10848 11660 10912
rect 11340 9824 11660 10848
rect 11340 9760 11348 9824
rect 11412 9760 11428 9824
rect 11492 9760 11508 9824
rect 11572 9760 11588 9824
rect 11652 9760 11660 9824
rect 11340 8736 11660 9760
rect 11340 8672 11348 8736
rect 11412 8672 11428 8736
rect 11492 8672 11508 8736
rect 11572 8672 11588 8736
rect 11652 8672 11660 8736
rect 11340 7648 11660 8672
rect 11340 7584 11348 7648
rect 11412 7584 11428 7648
rect 11492 7584 11508 7648
rect 11572 7584 11588 7648
rect 11652 7584 11660 7648
rect 11099 7308 11165 7309
rect 11099 7244 11100 7308
rect 11164 7244 11165 7308
rect 11099 7243 11165 7244
rect 11340 6560 11660 7584
rect 11340 6496 11348 6560
rect 11412 6496 11428 6560
rect 11492 6496 11508 6560
rect 11572 6496 11588 6560
rect 11652 6496 11660 6560
rect 11340 5472 11660 6496
rect 11340 5408 11348 5472
rect 11412 5408 11428 5472
rect 11492 5408 11508 5472
rect 11572 5408 11588 5472
rect 11652 5408 11660 5472
rect 10547 4452 10613 4453
rect 10547 4388 10548 4452
rect 10612 4388 10613 4452
rect 10547 4387 10613 4388
rect 11340 4384 11660 5408
rect 11340 4320 11348 4384
rect 11412 4320 11428 4384
rect 11492 4320 11508 4384
rect 11572 4320 11588 4384
rect 11652 4320 11660 4384
rect 11340 3296 11660 4320
rect 11340 3232 11348 3296
rect 11412 3232 11428 3296
rect 11492 3232 11508 3296
rect 11572 3232 11588 3296
rect 11652 3232 11660 3296
rect 9811 3228 9877 3229
rect 9811 3164 9812 3228
rect 9876 3164 9877 3228
rect 9811 3163 9877 3164
rect 9814 1325 9874 3163
rect 11340 2208 11660 3232
rect 12022 3093 12082 12547
rect 12206 10437 12266 12686
rect 12203 10436 12269 10437
rect 12203 10372 12204 10436
rect 12268 10372 12269 10436
rect 12203 10371 12269 10372
rect 12203 8804 12269 8805
rect 12203 8740 12204 8804
rect 12268 8740 12269 8804
rect 12203 8739 12269 8740
rect 12206 7989 12266 8739
rect 12203 7988 12269 7989
rect 12203 7924 12204 7988
rect 12268 7924 12269 7988
rect 12203 7923 12269 7924
rect 12574 4589 12634 13635
rect 12758 6901 12818 33491
rect 13126 31770 13186 42875
rect 13939 41920 14259 42944
rect 13939 41856 13947 41920
rect 14011 41856 14027 41920
rect 14091 41856 14107 41920
rect 14171 41856 14187 41920
rect 14251 41856 14259 41920
rect 13939 40832 14259 41856
rect 16538 43552 16858 43568
rect 16538 43488 16546 43552
rect 16610 43488 16626 43552
rect 16690 43488 16706 43552
rect 16770 43488 16786 43552
rect 16850 43488 16858 43552
rect 16538 42464 16858 43488
rect 19137 43008 19457 43568
rect 19137 42944 19145 43008
rect 19209 42944 19225 43008
rect 19289 42944 19305 43008
rect 19369 42944 19385 43008
rect 19449 42944 19457 43008
rect 17907 42940 17973 42941
rect 17907 42876 17908 42940
rect 17972 42876 17973 42940
rect 17907 42875 17973 42876
rect 16538 42400 16546 42464
rect 16610 42400 16626 42464
rect 16690 42400 16706 42464
rect 16770 42400 16786 42464
rect 16850 42400 16858 42464
rect 15147 41716 15213 41717
rect 15147 41652 15148 41716
rect 15212 41652 15213 41716
rect 15147 41651 15213 41652
rect 16067 41716 16133 41717
rect 16067 41652 16068 41716
rect 16132 41652 16133 41716
rect 16067 41651 16133 41652
rect 13939 40768 13947 40832
rect 14011 40768 14027 40832
rect 14091 40768 14107 40832
rect 14171 40768 14187 40832
rect 14251 40768 14259 40832
rect 13939 39744 14259 40768
rect 13939 39680 13947 39744
rect 14011 39680 14027 39744
rect 14091 39680 14107 39744
rect 14171 39680 14187 39744
rect 14251 39680 14259 39744
rect 13939 38656 14259 39680
rect 13939 38592 13947 38656
rect 14011 38592 14027 38656
rect 14091 38592 14107 38656
rect 14171 38592 14187 38656
rect 14251 38592 14259 38656
rect 13939 37568 14259 38592
rect 13939 37504 13947 37568
rect 14011 37504 14027 37568
rect 14091 37504 14107 37568
rect 14171 37504 14187 37568
rect 14251 37504 14259 37568
rect 13939 36480 14259 37504
rect 14411 37228 14477 37229
rect 14411 37164 14412 37228
rect 14476 37164 14477 37228
rect 14411 37163 14477 37164
rect 13939 36416 13947 36480
rect 14011 36416 14027 36480
rect 14091 36416 14107 36480
rect 14171 36416 14187 36480
rect 14251 36416 14259 36480
rect 13939 35392 14259 36416
rect 13939 35328 13947 35392
rect 14011 35328 14027 35392
rect 14091 35328 14107 35392
rect 14171 35328 14187 35392
rect 14251 35328 14259 35392
rect 13939 34304 14259 35328
rect 13939 34240 13947 34304
rect 14011 34240 14027 34304
rect 14091 34240 14107 34304
rect 14171 34240 14187 34304
rect 14251 34240 14259 34304
rect 13939 33216 14259 34240
rect 13939 33152 13947 33216
rect 14011 33152 14027 33216
rect 14091 33152 14107 33216
rect 14171 33152 14187 33216
rect 14251 33152 14259 33216
rect 13939 32128 14259 33152
rect 13939 32064 13947 32128
rect 14011 32064 14027 32128
rect 14091 32064 14107 32128
rect 14171 32064 14187 32128
rect 14251 32064 14259 32128
rect 13675 31924 13741 31925
rect 13675 31860 13676 31924
rect 13740 31860 13741 31924
rect 13675 31859 13741 31860
rect 12942 31710 13186 31770
rect 12942 22405 13002 31710
rect 13307 30700 13373 30701
rect 13307 30636 13308 30700
rect 13372 30636 13373 30700
rect 13307 30635 13373 30636
rect 13123 28524 13189 28525
rect 13123 28460 13124 28524
rect 13188 28460 13189 28524
rect 13123 28459 13189 28460
rect 13126 22949 13186 28459
rect 13310 25261 13370 30635
rect 13491 28796 13557 28797
rect 13491 28732 13492 28796
rect 13556 28732 13557 28796
rect 13491 28731 13557 28732
rect 13307 25260 13373 25261
rect 13307 25196 13308 25260
rect 13372 25196 13373 25260
rect 13307 25195 13373 25196
rect 13494 23221 13554 28731
rect 13491 23220 13557 23221
rect 13491 23156 13492 23220
rect 13556 23156 13557 23220
rect 13491 23155 13557 23156
rect 13123 22948 13189 22949
rect 13123 22884 13124 22948
rect 13188 22884 13189 22948
rect 13123 22883 13189 22884
rect 13123 22812 13189 22813
rect 13123 22748 13124 22812
rect 13188 22748 13189 22812
rect 13123 22747 13189 22748
rect 12939 22404 13005 22405
rect 12939 22340 12940 22404
rect 13004 22340 13005 22404
rect 12939 22339 13005 22340
rect 13126 20773 13186 22747
rect 13678 22110 13738 31859
rect 13310 22050 13738 22110
rect 13939 31040 14259 32064
rect 13939 30976 13947 31040
rect 14011 30976 14027 31040
rect 14091 30976 14107 31040
rect 14171 30976 14187 31040
rect 14251 30976 14259 31040
rect 13939 29952 14259 30976
rect 13939 29888 13947 29952
rect 14011 29888 14027 29952
rect 14091 29888 14107 29952
rect 14171 29888 14187 29952
rect 14251 29888 14259 29952
rect 13939 28864 14259 29888
rect 13939 28800 13947 28864
rect 14011 28800 14027 28864
rect 14091 28800 14107 28864
rect 14171 28800 14187 28864
rect 14251 28800 14259 28864
rect 13939 27776 14259 28800
rect 13939 27712 13947 27776
rect 14011 27712 14027 27776
rect 14091 27712 14107 27776
rect 14171 27712 14187 27776
rect 14251 27712 14259 27776
rect 13939 26688 14259 27712
rect 13939 26624 13947 26688
rect 14011 26624 14027 26688
rect 14091 26624 14107 26688
rect 14171 26624 14187 26688
rect 14251 26624 14259 26688
rect 13939 25600 14259 26624
rect 13939 25536 13947 25600
rect 14011 25536 14027 25600
rect 14091 25536 14107 25600
rect 14171 25536 14187 25600
rect 14251 25536 14259 25600
rect 13939 24512 14259 25536
rect 13939 24448 13947 24512
rect 14011 24448 14027 24512
rect 14091 24448 14107 24512
rect 14171 24448 14187 24512
rect 14251 24448 14259 24512
rect 13939 23424 14259 24448
rect 13939 23360 13947 23424
rect 14011 23360 14027 23424
rect 14091 23360 14107 23424
rect 14171 23360 14187 23424
rect 14251 23360 14259 23424
rect 13939 22336 14259 23360
rect 13939 22272 13947 22336
rect 14011 22272 14027 22336
rect 14091 22272 14107 22336
rect 14171 22272 14187 22336
rect 14251 22272 14259 22336
rect 13123 20772 13189 20773
rect 13123 20708 13124 20772
rect 13188 20708 13189 20772
rect 13123 20707 13189 20708
rect 12939 20500 13005 20501
rect 12939 20436 12940 20500
rect 13004 20436 13005 20500
rect 12939 20435 13005 20436
rect 12942 17781 13002 20435
rect 12939 17780 13005 17781
rect 12939 17716 12940 17780
rect 13004 17716 13005 17780
rect 12939 17715 13005 17716
rect 12942 14925 13002 17715
rect 13123 15196 13189 15197
rect 13123 15132 13124 15196
rect 13188 15132 13189 15196
rect 13123 15131 13189 15132
rect 12939 14924 13005 14925
rect 12939 14860 12940 14924
rect 13004 14860 13005 14924
rect 12939 14859 13005 14860
rect 12939 8804 13005 8805
rect 12939 8740 12940 8804
rect 13004 8740 13005 8804
rect 12939 8739 13005 8740
rect 12942 8397 13002 8739
rect 13126 8397 13186 15131
rect 13310 14109 13370 22050
rect 13939 21248 14259 22272
rect 13939 21184 13947 21248
rect 14011 21184 14027 21248
rect 14091 21184 14107 21248
rect 14171 21184 14187 21248
rect 14251 21184 14259 21248
rect 13675 20908 13741 20909
rect 13675 20844 13676 20908
rect 13740 20844 13741 20908
rect 13675 20843 13741 20844
rect 13678 17373 13738 20843
rect 13939 20160 14259 21184
rect 13939 20096 13947 20160
rect 14011 20096 14027 20160
rect 14091 20096 14107 20160
rect 14171 20096 14187 20160
rect 14251 20096 14259 20160
rect 13939 19072 14259 20096
rect 14414 19821 14474 37163
rect 14779 36684 14845 36685
rect 14779 36620 14780 36684
rect 14844 36620 14845 36684
rect 14779 36619 14845 36620
rect 14782 32741 14842 36619
rect 15150 33149 15210 41651
rect 15331 41444 15397 41445
rect 15331 41380 15332 41444
rect 15396 41380 15397 41444
rect 15331 41379 15397 41380
rect 15334 38725 15394 41379
rect 15331 38724 15397 38725
rect 15331 38660 15332 38724
rect 15396 38660 15397 38724
rect 15331 38659 15397 38660
rect 15515 36276 15581 36277
rect 15515 36212 15516 36276
rect 15580 36212 15581 36276
rect 15515 36211 15581 36212
rect 15331 35596 15397 35597
rect 15331 35532 15332 35596
rect 15396 35532 15397 35596
rect 15331 35531 15397 35532
rect 15147 33148 15213 33149
rect 15147 33084 15148 33148
rect 15212 33084 15213 33148
rect 15147 33083 15213 33084
rect 14779 32740 14845 32741
rect 14779 32676 14780 32740
rect 14844 32676 14845 32740
rect 14779 32675 14845 32676
rect 14782 30973 14842 32675
rect 15334 31789 15394 35531
rect 14963 31788 15029 31789
rect 14963 31724 14964 31788
rect 15028 31724 15029 31788
rect 14963 31723 15029 31724
rect 15331 31788 15397 31789
rect 15331 31724 15332 31788
rect 15396 31724 15397 31788
rect 15331 31723 15397 31724
rect 14966 31378 15026 31723
rect 14966 31318 15394 31378
rect 15147 31108 15213 31109
rect 15147 31044 15148 31108
rect 15212 31044 15213 31108
rect 15147 31043 15213 31044
rect 14779 30972 14845 30973
rect 14779 30908 14780 30972
rect 14844 30908 14845 30972
rect 14779 30907 14845 30908
rect 14595 28660 14661 28661
rect 14595 28596 14596 28660
rect 14660 28596 14661 28660
rect 14595 28595 14661 28596
rect 14411 19820 14477 19821
rect 14411 19756 14412 19820
rect 14476 19756 14477 19820
rect 14411 19755 14477 19756
rect 13939 19008 13947 19072
rect 14011 19008 14027 19072
rect 14091 19008 14107 19072
rect 14171 19008 14187 19072
rect 14251 19008 14259 19072
rect 13939 17984 14259 19008
rect 13939 17920 13947 17984
rect 14011 17920 14027 17984
rect 14091 17920 14107 17984
rect 14171 17920 14187 17984
rect 14251 17920 14259 17984
rect 13675 17372 13741 17373
rect 13675 17308 13676 17372
rect 13740 17308 13741 17372
rect 13675 17307 13741 17308
rect 13491 17100 13557 17101
rect 13491 17036 13492 17100
rect 13556 17036 13557 17100
rect 13491 17035 13557 17036
rect 13307 14108 13373 14109
rect 13307 14044 13308 14108
rect 13372 14044 13373 14108
rect 13307 14043 13373 14044
rect 13307 10572 13373 10573
rect 13307 10508 13308 10572
rect 13372 10508 13373 10572
rect 13307 10507 13373 10508
rect 12939 8396 13005 8397
rect 12939 8332 12940 8396
rect 13004 8332 13005 8396
rect 12939 8331 13005 8332
rect 13123 8396 13189 8397
rect 13123 8332 13124 8396
rect 13188 8332 13189 8396
rect 13123 8331 13189 8332
rect 13310 7581 13370 10507
rect 13494 10029 13554 17035
rect 13939 16896 14259 17920
rect 14411 17508 14477 17509
rect 14411 17444 14412 17508
rect 14476 17444 14477 17508
rect 14411 17443 14477 17444
rect 13939 16832 13947 16896
rect 14011 16832 14027 16896
rect 14091 16832 14107 16896
rect 14171 16832 14187 16896
rect 14251 16832 14259 16896
rect 13675 15876 13741 15877
rect 13675 15812 13676 15876
rect 13740 15812 13741 15876
rect 13675 15811 13741 15812
rect 13678 10029 13738 15811
rect 13939 15808 14259 16832
rect 13939 15744 13947 15808
rect 14011 15744 14027 15808
rect 14091 15744 14107 15808
rect 14171 15744 14187 15808
rect 14251 15744 14259 15808
rect 13939 14720 14259 15744
rect 13939 14656 13947 14720
rect 14011 14656 14027 14720
rect 14091 14656 14107 14720
rect 14171 14656 14187 14720
rect 14251 14656 14259 14720
rect 13939 13632 14259 14656
rect 13939 13568 13947 13632
rect 14011 13568 14027 13632
rect 14091 13568 14107 13632
rect 14171 13568 14187 13632
rect 14251 13568 14259 13632
rect 13939 12544 14259 13568
rect 13939 12480 13947 12544
rect 14011 12480 14027 12544
rect 14091 12480 14107 12544
rect 14171 12480 14187 12544
rect 14251 12480 14259 12544
rect 13939 11456 14259 12480
rect 13939 11392 13947 11456
rect 14011 11392 14027 11456
rect 14091 11392 14107 11456
rect 14171 11392 14187 11456
rect 14251 11392 14259 11456
rect 13939 10368 14259 11392
rect 13939 10304 13947 10368
rect 14011 10304 14027 10368
rect 14091 10304 14107 10368
rect 14171 10304 14187 10368
rect 14251 10304 14259 10368
rect 13491 10028 13557 10029
rect 13491 9964 13492 10028
rect 13556 9964 13557 10028
rect 13491 9963 13557 9964
rect 13675 10028 13741 10029
rect 13675 9964 13676 10028
rect 13740 9964 13741 10028
rect 13675 9963 13741 9964
rect 13939 9280 14259 10304
rect 13939 9216 13947 9280
rect 14011 9216 14027 9280
rect 14091 9216 14107 9280
rect 14171 9216 14187 9280
rect 14251 9216 14259 9280
rect 13939 8192 14259 9216
rect 13939 8128 13947 8192
rect 14011 8128 14027 8192
rect 14091 8128 14107 8192
rect 14171 8128 14187 8192
rect 14251 8128 14259 8192
rect 13307 7580 13373 7581
rect 13307 7516 13308 7580
rect 13372 7516 13373 7580
rect 13307 7515 13373 7516
rect 13939 7104 14259 8128
rect 13939 7040 13947 7104
rect 14011 7040 14027 7104
rect 14091 7040 14107 7104
rect 14171 7040 14187 7104
rect 14251 7040 14259 7104
rect 12755 6900 12821 6901
rect 12755 6836 12756 6900
rect 12820 6836 12821 6900
rect 12755 6835 12821 6836
rect 13939 6016 14259 7040
rect 14414 6901 14474 17443
rect 14598 16693 14658 28595
rect 14963 27980 15029 27981
rect 14963 27916 14964 27980
rect 15028 27916 15029 27980
rect 14963 27915 15029 27916
rect 14966 24717 15026 27915
rect 14779 24716 14845 24717
rect 14779 24652 14780 24716
rect 14844 24652 14845 24716
rect 14779 24651 14845 24652
rect 14963 24716 15029 24717
rect 14963 24652 14964 24716
rect 15028 24652 15029 24716
rect 14963 24651 15029 24652
rect 14782 22269 14842 24651
rect 14963 24580 15029 24581
rect 14963 24516 14964 24580
rect 15028 24516 15029 24580
rect 14963 24515 15029 24516
rect 14779 22268 14845 22269
rect 14779 22204 14780 22268
rect 14844 22204 14845 22268
rect 14779 22203 14845 22204
rect 14966 17645 15026 24515
rect 15150 24037 15210 31043
rect 15147 24036 15213 24037
rect 15147 23972 15148 24036
rect 15212 23972 15213 24036
rect 15147 23971 15213 23972
rect 15334 22110 15394 31318
rect 15518 24989 15578 36211
rect 15883 33828 15949 33829
rect 15883 33764 15884 33828
rect 15948 33764 15949 33828
rect 15883 33763 15949 33764
rect 15699 32876 15765 32877
rect 15699 32812 15700 32876
rect 15764 32812 15765 32876
rect 15699 32811 15765 32812
rect 15515 24988 15581 24989
rect 15515 24924 15516 24988
rect 15580 24924 15581 24988
rect 15515 24923 15581 24924
rect 15334 22050 15578 22110
rect 15147 20772 15213 20773
rect 15147 20708 15148 20772
rect 15212 20708 15213 20772
rect 15147 20707 15213 20708
rect 14963 17644 15029 17645
rect 14963 17580 14964 17644
rect 15028 17580 15029 17644
rect 14963 17579 15029 17580
rect 15150 17509 15210 20707
rect 15331 20500 15397 20501
rect 15331 20436 15332 20500
rect 15396 20436 15397 20500
rect 15331 20435 15397 20436
rect 15147 17508 15213 17509
rect 15147 17444 15148 17508
rect 15212 17444 15213 17508
rect 15147 17443 15213 17444
rect 14595 16692 14661 16693
rect 14595 16628 14596 16692
rect 14660 16628 14661 16692
rect 14595 16627 14661 16628
rect 14779 16556 14845 16557
rect 14779 16492 14780 16556
rect 14844 16492 14845 16556
rect 14779 16491 14845 16492
rect 14595 13564 14661 13565
rect 14595 13500 14596 13564
rect 14660 13500 14661 13564
rect 14595 13499 14661 13500
rect 14411 6900 14477 6901
rect 14411 6836 14412 6900
rect 14476 6836 14477 6900
rect 14411 6835 14477 6836
rect 13939 5952 13947 6016
rect 14011 5952 14027 6016
rect 14091 5952 14107 6016
rect 14171 5952 14187 6016
rect 14251 5952 14259 6016
rect 13939 4928 14259 5952
rect 13939 4864 13947 4928
rect 14011 4864 14027 4928
rect 14091 4864 14107 4928
rect 14171 4864 14187 4928
rect 14251 4864 14259 4928
rect 12571 4588 12637 4589
rect 12571 4524 12572 4588
rect 12636 4524 12637 4588
rect 12571 4523 12637 4524
rect 13939 3840 14259 4864
rect 14598 4317 14658 13499
rect 14782 9757 14842 16491
rect 15334 15197 15394 20435
rect 15331 15196 15397 15197
rect 15331 15132 15332 15196
rect 15396 15132 15397 15196
rect 15331 15131 15397 15132
rect 14779 9756 14845 9757
rect 14779 9692 14780 9756
rect 14844 9692 14845 9756
rect 14779 9691 14845 9692
rect 15147 6356 15213 6357
rect 15147 6292 15148 6356
rect 15212 6292 15213 6356
rect 15147 6291 15213 6292
rect 14595 4316 14661 4317
rect 14595 4252 14596 4316
rect 14660 4252 14661 4316
rect 14595 4251 14661 4252
rect 13939 3776 13947 3840
rect 14011 3776 14027 3840
rect 14091 3776 14107 3840
rect 14171 3776 14187 3840
rect 14251 3776 14259 3840
rect 12019 3092 12085 3093
rect 12019 3028 12020 3092
rect 12084 3028 12085 3092
rect 12019 3027 12085 3028
rect 11340 2144 11348 2208
rect 11412 2144 11428 2208
rect 11492 2144 11508 2208
rect 11572 2144 11588 2208
rect 11652 2144 11660 2208
rect 9811 1324 9877 1325
rect 9811 1260 9812 1324
rect 9876 1260 9877 1324
rect 9811 1259 9877 1260
rect 11340 1120 11660 2144
rect 11340 1056 11348 1120
rect 11412 1056 11428 1120
rect 11492 1056 11508 1120
rect 11572 1056 11588 1120
rect 11652 1056 11660 1120
rect 11340 1040 11660 1056
rect 13939 2752 14259 3776
rect 15150 3637 15210 6291
rect 15518 3637 15578 22050
rect 15702 4045 15762 32811
rect 15886 30021 15946 33763
rect 15883 30020 15949 30021
rect 15883 29956 15884 30020
rect 15948 29956 15949 30020
rect 15883 29955 15949 29956
rect 16070 29069 16130 41651
rect 16538 41376 16858 42400
rect 17723 42124 17789 42125
rect 17723 42060 17724 42124
rect 17788 42060 17789 42124
rect 17723 42059 17789 42060
rect 17355 41580 17421 41581
rect 17355 41516 17356 41580
rect 17420 41516 17421 41580
rect 17355 41515 17421 41516
rect 16538 41312 16546 41376
rect 16610 41312 16626 41376
rect 16690 41312 16706 41376
rect 16770 41312 16786 41376
rect 16850 41312 16858 41376
rect 16538 40288 16858 41312
rect 16538 40224 16546 40288
rect 16610 40224 16626 40288
rect 16690 40224 16706 40288
rect 16770 40224 16786 40288
rect 16850 40224 16858 40288
rect 16538 39200 16858 40224
rect 16538 39136 16546 39200
rect 16610 39136 16626 39200
rect 16690 39136 16706 39200
rect 16770 39136 16786 39200
rect 16850 39136 16858 39200
rect 16538 38112 16858 39136
rect 16538 38048 16546 38112
rect 16610 38048 16626 38112
rect 16690 38048 16706 38112
rect 16770 38048 16786 38112
rect 16850 38048 16858 38112
rect 16538 37024 16858 38048
rect 16538 36960 16546 37024
rect 16610 36960 16626 37024
rect 16690 36960 16706 37024
rect 16770 36960 16786 37024
rect 16850 36960 16858 37024
rect 16538 35936 16858 36960
rect 16538 35872 16546 35936
rect 16610 35872 16626 35936
rect 16690 35872 16706 35936
rect 16770 35872 16786 35936
rect 16850 35872 16858 35936
rect 16538 34848 16858 35872
rect 16538 34784 16546 34848
rect 16610 34784 16626 34848
rect 16690 34784 16706 34848
rect 16770 34784 16786 34848
rect 16850 34784 16858 34848
rect 16538 33760 16858 34784
rect 16538 33696 16546 33760
rect 16610 33696 16626 33760
rect 16690 33696 16706 33760
rect 16770 33696 16786 33760
rect 16850 33696 16858 33760
rect 16538 32672 16858 33696
rect 16538 32608 16546 32672
rect 16610 32608 16626 32672
rect 16690 32608 16706 32672
rect 16770 32608 16786 32672
rect 16850 32608 16858 32672
rect 16538 31584 16858 32608
rect 16538 31520 16546 31584
rect 16610 31520 16626 31584
rect 16690 31520 16706 31584
rect 16770 31520 16786 31584
rect 16850 31520 16858 31584
rect 16538 30496 16858 31520
rect 16538 30432 16546 30496
rect 16610 30432 16626 30496
rect 16690 30432 16706 30496
rect 16770 30432 16786 30496
rect 16850 30432 16858 30496
rect 16538 29408 16858 30432
rect 16538 29344 16546 29408
rect 16610 29344 16626 29408
rect 16690 29344 16706 29408
rect 16770 29344 16786 29408
rect 16850 29344 16858 29408
rect 16067 29068 16133 29069
rect 16067 29004 16068 29068
rect 16132 29004 16133 29068
rect 16067 29003 16133 29004
rect 16538 28320 16858 29344
rect 17171 29068 17237 29069
rect 17171 29004 17172 29068
rect 17236 29004 17237 29068
rect 17171 29003 17237 29004
rect 16538 28256 16546 28320
rect 16610 28256 16626 28320
rect 16690 28256 16706 28320
rect 16770 28256 16786 28320
rect 16850 28256 16858 28320
rect 16067 27708 16133 27709
rect 16067 27644 16068 27708
rect 16132 27644 16133 27708
rect 16067 27643 16133 27644
rect 15883 21180 15949 21181
rect 15883 21116 15884 21180
rect 15948 21116 15949 21180
rect 15883 21115 15949 21116
rect 15886 17781 15946 21115
rect 16070 20773 16130 27643
rect 16538 27232 16858 28256
rect 16538 27168 16546 27232
rect 16610 27168 16626 27232
rect 16690 27168 16706 27232
rect 16770 27168 16786 27232
rect 16850 27168 16858 27232
rect 16538 26144 16858 27168
rect 16538 26080 16546 26144
rect 16610 26080 16626 26144
rect 16690 26080 16706 26144
rect 16770 26080 16786 26144
rect 16850 26080 16858 26144
rect 16538 25056 16858 26080
rect 16538 24992 16546 25056
rect 16610 24992 16626 25056
rect 16690 24992 16706 25056
rect 16770 24992 16786 25056
rect 16850 24992 16858 25056
rect 16538 23968 16858 24992
rect 16987 24716 17053 24717
rect 16987 24652 16988 24716
rect 17052 24652 17053 24716
rect 16987 24651 17053 24652
rect 16538 23904 16546 23968
rect 16610 23904 16626 23968
rect 16690 23904 16706 23968
rect 16770 23904 16786 23968
rect 16850 23904 16858 23968
rect 16251 23492 16317 23493
rect 16251 23428 16252 23492
rect 16316 23428 16317 23492
rect 16251 23427 16317 23428
rect 16067 20772 16133 20773
rect 16067 20708 16068 20772
rect 16132 20708 16133 20772
rect 16067 20707 16133 20708
rect 16067 20364 16133 20365
rect 16067 20300 16068 20364
rect 16132 20300 16133 20364
rect 16067 20299 16133 20300
rect 16070 18869 16130 20299
rect 16067 18868 16133 18869
rect 16067 18804 16068 18868
rect 16132 18804 16133 18868
rect 16067 18803 16133 18804
rect 15883 17780 15949 17781
rect 15883 17716 15884 17780
rect 15948 17716 15949 17780
rect 15883 17715 15949 17716
rect 16070 11389 16130 18803
rect 16254 18053 16314 23427
rect 16538 22880 16858 23904
rect 16538 22816 16546 22880
rect 16610 22816 16626 22880
rect 16690 22816 16706 22880
rect 16770 22816 16786 22880
rect 16850 22816 16858 22880
rect 16538 21792 16858 22816
rect 16538 21728 16546 21792
rect 16610 21728 16626 21792
rect 16690 21728 16706 21792
rect 16770 21728 16786 21792
rect 16850 21728 16858 21792
rect 16538 20704 16858 21728
rect 16538 20640 16546 20704
rect 16610 20640 16626 20704
rect 16690 20640 16706 20704
rect 16770 20640 16786 20704
rect 16850 20640 16858 20704
rect 16538 19616 16858 20640
rect 16538 19552 16546 19616
rect 16610 19552 16626 19616
rect 16690 19552 16706 19616
rect 16770 19552 16786 19616
rect 16850 19552 16858 19616
rect 16538 18528 16858 19552
rect 16538 18464 16546 18528
rect 16610 18464 16626 18528
rect 16690 18464 16706 18528
rect 16770 18464 16786 18528
rect 16850 18464 16858 18528
rect 16251 18052 16317 18053
rect 16251 17988 16252 18052
rect 16316 17988 16317 18052
rect 16251 17987 16317 17988
rect 16538 17440 16858 18464
rect 16990 18189 17050 24651
rect 16987 18188 17053 18189
rect 16987 18124 16988 18188
rect 17052 18124 17053 18188
rect 16987 18123 17053 18124
rect 16987 18052 17053 18053
rect 16987 17988 16988 18052
rect 17052 17988 17053 18052
rect 16987 17987 17053 17988
rect 16538 17376 16546 17440
rect 16610 17376 16626 17440
rect 16690 17376 16706 17440
rect 16770 17376 16786 17440
rect 16850 17376 16858 17440
rect 16538 16352 16858 17376
rect 16538 16288 16546 16352
rect 16610 16288 16626 16352
rect 16690 16288 16706 16352
rect 16770 16288 16786 16352
rect 16850 16288 16858 16352
rect 16251 15604 16317 15605
rect 16251 15540 16252 15604
rect 16316 15540 16317 15604
rect 16251 15539 16317 15540
rect 16067 11388 16133 11389
rect 16067 11324 16068 11388
rect 16132 11324 16133 11388
rect 16067 11323 16133 11324
rect 16254 10981 16314 15539
rect 16538 15264 16858 16288
rect 16538 15200 16546 15264
rect 16610 15200 16626 15264
rect 16690 15200 16706 15264
rect 16770 15200 16786 15264
rect 16850 15200 16858 15264
rect 16538 14176 16858 15200
rect 16538 14112 16546 14176
rect 16610 14112 16626 14176
rect 16690 14112 16706 14176
rect 16770 14112 16786 14176
rect 16850 14112 16858 14176
rect 16538 13088 16858 14112
rect 16538 13024 16546 13088
rect 16610 13024 16626 13088
rect 16690 13024 16706 13088
rect 16770 13024 16786 13088
rect 16850 13024 16858 13088
rect 16538 12000 16858 13024
rect 16538 11936 16546 12000
rect 16610 11936 16626 12000
rect 16690 11936 16706 12000
rect 16770 11936 16786 12000
rect 16850 11936 16858 12000
rect 16251 10980 16317 10981
rect 16251 10916 16252 10980
rect 16316 10916 16317 10980
rect 16251 10915 16317 10916
rect 16538 10912 16858 11936
rect 16990 11933 17050 17987
rect 17174 12069 17234 29003
rect 17358 28933 17418 41515
rect 17726 40901 17786 42059
rect 17723 40900 17789 40901
rect 17723 40836 17724 40900
rect 17788 40836 17789 40900
rect 17723 40835 17789 40836
rect 17910 40629 17970 42875
rect 19137 41920 19457 42944
rect 21736 43552 22056 43568
rect 21736 43488 21744 43552
rect 21808 43488 21824 43552
rect 21888 43488 21904 43552
rect 21968 43488 21984 43552
rect 22048 43488 22056 43552
rect 21736 42464 22056 43488
rect 21736 42400 21744 42464
rect 21808 42400 21824 42464
rect 21888 42400 21904 42464
rect 21968 42400 21984 42464
rect 22048 42400 22056 42464
rect 19747 42396 19813 42397
rect 19747 42332 19748 42396
rect 19812 42332 19813 42396
rect 19747 42331 19813 42332
rect 19137 41856 19145 41920
rect 19209 41856 19225 41920
rect 19289 41856 19305 41920
rect 19369 41856 19385 41920
rect 19449 41856 19457 41920
rect 18091 41852 18157 41853
rect 18091 41788 18092 41852
rect 18156 41788 18157 41852
rect 18091 41787 18157 41788
rect 17907 40628 17973 40629
rect 17907 40564 17908 40628
rect 17972 40564 17973 40628
rect 17907 40563 17973 40564
rect 18094 38997 18154 41787
rect 18275 41308 18341 41309
rect 18275 41244 18276 41308
rect 18340 41244 18341 41308
rect 18275 41243 18341 41244
rect 18091 38996 18157 38997
rect 18091 38932 18092 38996
rect 18156 38932 18157 38996
rect 18091 38931 18157 38932
rect 18278 38725 18338 41243
rect 19137 40832 19457 41856
rect 19137 40768 19145 40832
rect 19209 40768 19225 40832
rect 19289 40768 19305 40832
rect 19369 40768 19385 40832
rect 19449 40768 19457 40832
rect 19011 40084 19077 40085
rect 19011 40020 19012 40084
rect 19076 40020 19077 40084
rect 19011 40019 19077 40020
rect 18275 38724 18341 38725
rect 18275 38660 18276 38724
rect 18340 38660 18341 38724
rect 18275 38659 18341 38660
rect 17723 36276 17789 36277
rect 17723 36212 17724 36276
rect 17788 36212 17789 36276
rect 17723 36211 17789 36212
rect 17355 28932 17421 28933
rect 17355 28868 17356 28932
rect 17420 28868 17421 28932
rect 17355 28867 17421 28868
rect 17539 27844 17605 27845
rect 17539 27780 17540 27844
rect 17604 27780 17605 27844
rect 17539 27779 17605 27780
rect 17355 24172 17421 24173
rect 17355 24108 17356 24172
rect 17420 24108 17421 24172
rect 17355 24107 17421 24108
rect 17358 17370 17418 24107
rect 17542 18050 17602 27779
rect 17726 19413 17786 36211
rect 18091 34100 18157 34101
rect 18091 34036 18092 34100
rect 18156 34036 18157 34100
rect 18091 34035 18157 34036
rect 17907 33692 17973 33693
rect 17907 33628 17908 33692
rect 17972 33628 17973 33692
rect 17907 33627 17973 33628
rect 17723 19412 17789 19413
rect 17723 19348 17724 19412
rect 17788 19348 17789 19412
rect 17723 19347 17789 19348
rect 17542 17990 17786 18050
rect 17358 17310 17602 17370
rect 17355 13972 17421 13973
rect 17355 13908 17356 13972
rect 17420 13908 17421 13972
rect 17355 13907 17421 13908
rect 17171 12068 17237 12069
rect 17171 12004 17172 12068
rect 17236 12004 17237 12068
rect 17171 12003 17237 12004
rect 16987 11932 17053 11933
rect 16987 11868 16988 11932
rect 17052 11868 17053 11932
rect 16987 11867 17053 11868
rect 16538 10848 16546 10912
rect 16610 10848 16626 10912
rect 16690 10848 16706 10912
rect 16770 10848 16786 10912
rect 16850 10848 16858 10912
rect 16538 9824 16858 10848
rect 16538 9760 16546 9824
rect 16610 9760 16626 9824
rect 16690 9760 16706 9824
rect 16770 9760 16786 9824
rect 16850 9760 16858 9824
rect 16251 9076 16317 9077
rect 16251 9012 16252 9076
rect 16316 9012 16317 9076
rect 16251 9011 16317 9012
rect 15699 4044 15765 4045
rect 15699 3980 15700 4044
rect 15764 3980 15765 4044
rect 15699 3979 15765 3980
rect 15147 3636 15213 3637
rect 15147 3572 15148 3636
rect 15212 3572 15213 3636
rect 15147 3571 15213 3572
rect 15515 3636 15581 3637
rect 15515 3572 15516 3636
rect 15580 3572 15581 3636
rect 15515 3571 15581 3572
rect 16254 3365 16314 9011
rect 16538 8736 16858 9760
rect 16987 9620 17053 9621
rect 16987 9556 16988 9620
rect 17052 9556 17053 9620
rect 16987 9555 17053 9556
rect 16538 8672 16546 8736
rect 16610 8672 16626 8736
rect 16690 8672 16706 8736
rect 16770 8672 16786 8736
rect 16850 8672 16858 8736
rect 16538 7648 16858 8672
rect 16538 7584 16546 7648
rect 16610 7584 16626 7648
rect 16690 7584 16706 7648
rect 16770 7584 16786 7648
rect 16850 7584 16858 7648
rect 16538 6560 16858 7584
rect 16538 6496 16546 6560
rect 16610 6496 16626 6560
rect 16690 6496 16706 6560
rect 16770 6496 16786 6560
rect 16850 6496 16858 6560
rect 16538 5472 16858 6496
rect 16538 5408 16546 5472
rect 16610 5408 16626 5472
rect 16690 5408 16706 5472
rect 16770 5408 16786 5472
rect 16850 5408 16858 5472
rect 16538 4384 16858 5408
rect 16538 4320 16546 4384
rect 16610 4320 16626 4384
rect 16690 4320 16706 4384
rect 16770 4320 16786 4384
rect 16850 4320 16858 4384
rect 16251 3364 16317 3365
rect 16251 3300 16252 3364
rect 16316 3300 16317 3364
rect 16251 3299 16317 3300
rect 13939 2688 13947 2752
rect 14011 2688 14027 2752
rect 14091 2688 14107 2752
rect 14171 2688 14187 2752
rect 14251 2688 14259 2752
rect 13939 1664 14259 2688
rect 13939 1600 13947 1664
rect 14011 1600 14027 1664
rect 14091 1600 14107 1664
rect 14171 1600 14187 1664
rect 14251 1600 14259 1664
rect 13939 1040 14259 1600
rect 16538 3296 16858 4320
rect 16538 3232 16546 3296
rect 16610 3232 16626 3296
rect 16690 3232 16706 3296
rect 16770 3232 16786 3296
rect 16850 3232 16858 3296
rect 16538 2208 16858 3232
rect 16538 2144 16546 2208
rect 16610 2144 16626 2208
rect 16690 2144 16706 2208
rect 16770 2144 16786 2208
rect 16850 2144 16858 2208
rect 16538 1120 16858 2144
rect 16990 1733 17050 9555
rect 17171 9484 17237 9485
rect 17171 9420 17172 9484
rect 17236 9420 17237 9484
rect 17171 9419 17237 9420
rect 17174 2410 17234 9419
rect 17358 2685 17418 13907
rect 17542 8397 17602 17310
rect 17726 12450 17786 17990
rect 17910 13701 17970 33627
rect 18094 26213 18154 34035
rect 18827 29068 18893 29069
rect 18827 29004 18828 29068
rect 18892 29004 18893 29068
rect 18827 29003 18893 29004
rect 18091 26212 18157 26213
rect 18091 26148 18092 26212
rect 18156 26148 18157 26212
rect 18091 26147 18157 26148
rect 18275 25396 18341 25397
rect 18275 25332 18276 25396
rect 18340 25332 18341 25396
rect 18275 25331 18341 25332
rect 18091 18732 18157 18733
rect 18091 18668 18092 18732
rect 18156 18668 18157 18732
rect 18091 18667 18157 18668
rect 18094 15333 18154 18667
rect 18091 15332 18157 15333
rect 18091 15268 18092 15332
rect 18156 15268 18157 15332
rect 18091 15267 18157 15268
rect 17907 13700 17973 13701
rect 17907 13636 17908 13700
rect 17972 13636 17973 13700
rect 17907 13635 17973 13636
rect 17726 12390 17970 12450
rect 17539 8396 17605 8397
rect 17539 8332 17540 8396
rect 17604 8332 17605 8396
rect 17539 8331 17605 8332
rect 17723 5404 17789 5405
rect 17723 5340 17724 5404
rect 17788 5340 17789 5404
rect 17723 5339 17789 5340
rect 17726 3365 17786 5339
rect 17723 3364 17789 3365
rect 17723 3300 17724 3364
rect 17788 3300 17789 3364
rect 17723 3299 17789 3300
rect 17910 2685 17970 12390
rect 18091 6220 18157 6221
rect 18091 6156 18092 6220
rect 18156 6156 18157 6220
rect 18091 6155 18157 6156
rect 18094 3365 18154 6155
rect 18278 4045 18338 25331
rect 18643 24852 18709 24853
rect 18643 24788 18644 24852
rect 18708 24788 18709 24852
rect 18643 24787 18709 24788
rect 18646 19277 18706 24787
rect 18643 19276 18709 19277
rect 18643 19212 18644 19276
rect 18708 19212 18709 19276
rect 18643 19211 18709 19212
rect 18459 14924 18525 14925
rect 18459 14860 18460 14924
rect 18524 14860 18525 14924
rect 18459 14859 18525 14860
rect 18462 5541 18522 14859
rect 18830 13973 18890 29003
rect 19014 20909 19074 40019
rect 19137 39744 19457 40768
rect 19750 40493 19810 42331
rect 20483 42260 20549 42261
rect 20483 42196 20484 42260
rect 20548 42196 20549 42260
rect 20483 42195 20549 42196
rect 19931 40764 19997 40765
rect 19931 40700 19932 40764
rect 19996 40700 19997 40764
rect 19931 40699 19997 40700
rect 19747 40492 19813 40493
rect 19747 40428 19748 40492
rect 19812 40428 19813 40492
rect 19747 40427 19813 40428
rect 19563 40084 19629 40085
rect 19563 40020 19564 40084
rect 19628 40020 19629 40084
rect 19563 40019 19629 40020
rect 19137 39680 19145 39744
rect 19209 39680 19225 39744
rect 19289 39680 19305 39744
rect 19369 39680 19385 39744
rect 19449 39680 19457 39744
rect 19137 38656 19457 39680
rect 19137 38592 19145 38656
rect 19209 38592 19225 38656
rect 19289 38592 19305 38656
rect 19369 38592 19385 38656
rect 19449 38592 19457 38656
rect 19137 37568 19457 38592
rect 19137 37504 19145 37568
rect 19209 37504 19225 37568
rect 19289 37504 19305 37568
rect 19369 37504 19385 37568
rect 19449 37504 19457 37568
rect 19137 36480 19457 37504
rect 19137 36416 19145 36480
rect 19209 36416 19225 36480
rect 19289 36416 19305 36480
rect 19369 36416 19385 36480
rect 19449 36416 19457 36480
rect 19137 35392 19457 36416
rect 19137 35328 19145 35392
rect 19209 35328 19225 35392
rect 19289 35328 19305 35392
rect 19369 35328 19385 35392
rect 19449 35328 19457 35392
rect 19137 34304 19457 35328
rect 19137 34240 19145 34304
rect 19209 34240 19225 34304
rect 19289 34240 19305 34304
rect 19369 34240 19385 34304
rect 19449 34240 19457 34304
rect 19137 33216 19457 34240
rect 19137 33152 19145 33216
rect 19209 33152 19225 33216
rect 19289 33152 19305 33216
rect 19369 33152 19385 33216
rect 19449 33152 19457 33216
rect 19137 32128 19457 33152
rect 19137 32064 19145 32128
rect 19209 32064 19225 32128
rect 19289 32064 19305 32128
rect 19369 32064 19385 32128
rect 19449 32064 19457 32128
rect 19137 31040 19457 32064
rect 19137 30976 19145 31040
rect 19209 30976 19225 31040
rect 19289 30976 19305 31040
rect 19369 30976 19385 31040
rect 19449 30976 19457 31040
rect 19137 29952 19457 30976
rect 19137 29888 19145 29952
rect 19209 29888 19225 29952
rect 19289 29888 19305 29952
rect 19369 29888 19385 29952
rect 19449 29888 19457 29952
rect 19137 28864 19457 29888
rect 19137 28800 19145 28864
rect 19209 28800 19225 28864
rect 19289 28800 19305 28864
rect 19369 28800 19385 28864
rect 19449 28800 19457 28864
rect 19137 27776 19457 28800
rect 19137 27712 19145 27776
rect 19209 27712 19225 27776
rect 19289 27712 19305 27776
rect 19369 27712 19385 27776
rect 19449 27712 19457 27776
rect 19137 26688 19457 27712
rect 19137 26624 19145 26688
rect 19209 26624 19225 26688
rect 19289 26624 19305 26688
rect 19369 26624 19385 26688
rect 19449 26624 19457 26688
rect 19137 25600 19457 26624
rect 19137 25536 19145 25600
rect 19209 25536 19225 25600
rect 19289 25536 19305 25600
rect 19369 25536 19385 25600
rect 19449 25536 19457 25600
rect 19137 24512 19457 25536
rect 19137 24448 19145 24512
rect 19209 24448 19225 24512
rect 19289 24448 19305 24512
rect 19369 24448 19385 24512
rect 19449 24448 19457 24512
rect 19137 23424 19457 24448
rect 19137 23360 19145 23424
rect 19209 23360 19225 23424
rect 19289 23360 19305 23424
rect 19369 23360 19385 23424
rect 19449 23360 19457 23424
rect 19137 22336 19457 23360
rect 19566 22541 19626 40019
rect 19934 39949 19994 40699
rect 19931 39948 19997 39949
rect 19931 39884 19932 39948
rect 19996 39884 19997 39948
rect 19931 39883 19997 39884
rect 20115 38724 20181 38725
rect 20115 38660 20116 38724
rect 20180 38660 20181 38724
rect 20115 38659 20181 38660
rect 20118 31770 20178 38659
rect 20299 32876 20365 32877
rect 20299 32812 20300 32876
rect 20364 32812 20365 32876
rect 20299 32811 20365 32812
rect 19750 31710 20178 31770
rect 19563 22540 19629 22541
rect 19563 22476 19564 22540
rect 19628 22476 19629 22540
rect 19563 22475 19629 22476
rect 19137 22272 19145 22336
rect 19209 22272 19225 22336
rect 19289 22272 19305 22336
rect 19369 22272 19385 22336
rect 19449 22272 19457 22336
rect 19137 21248 19457 22272
rect 19750 22110 19810 31710
rect 19137 21184 19145 21248
rect 19209 21184 19225 21248
rect 19289 21184 19305 21248
rect 19369 21184 19385 21248
rect 19449 21184 19457 21248
rect 19011 20908 19077 20909
rect 19011 20844 19012 20908
rect 19076 20844 19077 20908
rect 19011 20843 19077 20844
rect 19137 20160 19457 21184
rect 19137 20096 19145 20160
rect 19209 20096 19225 20160
rect 19289 20096 19305 20160
rect 19369 20096 19385 20160
rect 19449 20096 19457 20160
rect 19137 19072 19457 20096
rect 19566 22050 19810 22110
rect 19931 22132 19997 22133
rect 19931 22068 19932 22132
rect 19996 22068 19997 22132
rect 20302 22110 20362 32811
rect 19931 22067 19997 22068
rect 19566 19821 19626 22050
rect 19747 20908 19813 20909
rect 19747 20844 19748 20908
rect 19812 20844 19813 20908
rect 19747 20843 19813 20844
rect 19563 19820 19629 19821
rect 19563 19756 19564 19820
rect 19628 19756 19629 19820
rect 19563 19755 19629 19756
rect 19137 19008 19145 19072
rect 19209 19008 19225 19072
rect 19289 19008 19305 19072
rect 19369 19008 19385 19072
rect 19449 19008 19457 19072
rect 19137 17984 19457 19008
rect 19137 17920 19145 17984
rect 19209 17920 19225 17984
rect 19289 17920 19305 17984
rect 19369 17920 19385 17984
rect 19449 17920 19457 17984
rect 19137 16896 19457 17920
rect 19137 16832 19145 16896
rect 19209 16832 19225 16896
rect 19289 16832 19305 16896
rect 19369 16832 19385 16896
rect 19449 16832 19457 16896
rect 19011 16012 19077 16013
rect 19011 15948 19012 16012
rect 19076 15948 19077 16012
rect 19011 15947 19077 15948
rect 18827 13972 18893 13973
rect 18827 13908 18828 13972
rect 18892 13908 18893 13972
rect 18827 13907 18893 13908
rect 18827 13156 18893 13157
rect 18827 13092 18828 13156
rect 18892 13092 18893 13156
rect 18827 13091 18893 13092
rect 18830 7717 18890 13091
rect 19014 12341 19074 15947
rect 19137 15808 19457 16832
rect 19137 15744 19145 15808
rect 19209 15744 19225 15808
rect 19289 15744 19305 15808
rect 19369 15744 19385 15808
rect 19449 15744 19457 15808
rect 19137 14720 19457 15744
rect 19137 14656 19145 14720
rect 19209 14656 19225 14720
rect 19289 14656 19305 14720
rect 19369 14656 19385 14720
rect 19449 14656 19457 14720
rect 19137 13632 19457 14656
rect 19137 13568 19145 13632
rect 19209 13568 19225 13632
rect 19289 13568 19305 13632
rect 19369 13568 19385 13632
rect 19449 13568 19457 13632
rect 19137 12544 19457 13568
rect 19137 12480 19145 12544
rect 19209 12480 19225 12544
rect 19289 12480 19305 12544
rect 19369 12480 19385 12544
rect 19449 12480 19457 12544
rect 19011 12340 19077 12341
rect 19011 12276 19012 12340
rect 19076 12276 19077 12340
rect 19011 12275 19077 12276
rect 19137 11456 19457 12480
rect 19750 12477 19810 20843
rect 19934 13293 19994 22067
rect 20118 22050 20362 22110
rect 19931 13292 19997 13293
rect 19931 13228 19932 13292
rect 19996 13228 19997 13292
rect 19931 13227 19997 13228
rect 19747 12476 19813 12477
rect 19747 12412 19748 12476
rect 19812 12412 19813 12476
rect 19747 12411 19813 12412
rect 19137 11392 19145 11456
rect 19209 11392 19225 11456
rect 19289 11392 19305 11456
rect 19369 11392 19385 11456
rect 19449 11392 19457 11456
rect 19137 10368 19457 11392
rect 19137 10304 19145 10368
rect 19209 10304 19225 10368
rect 19289 10304 19305 10368
rect 19369 10304 19385 10368
rect 19449 10304 19457 10368
rect 19011 9620 19077 9621
rect 19011 9556 19012 9620
rect 19076 9556 19077 9620
rect 19011 9555 19077 9556
rect 18827 7716 18893 7717
rect 18827 7652 18828 7716
rect 18892 7652 18893 7716
rect 18827 7651 18893 7652
rect 19014 5677 19074 9555
rect 19137 9280 19457 10304
rect 19931 9756 19997 9757
rect 19931 9692 19932 9756
rect 19996 9692 19997 9756
rect 19931 9691 19997 9692
rect 19137 9216 19145 9280
rect 19209 9216 19225 9280
rect 19289 9216 19305 9280
rect 19369 9216 19385 9280
rect 19449 9216 19457 9280
rect 19137 8192 19457 9216
rect 19137 8128 19145 8192
rect 19209 8128 19225 8192
rect 19289 8128 19305 8192
rect 19369 8128 19385 8192
rect 19449 8128 19457 8192
rect 19137 7104 19457 8128
rect 19137 7040 19145 7104
rect 19209 7040 19225 7104
rect 19289 7040 19305 7104
rect 19369 7040 19385 7104
rect 19449 7040 19457 7104
rect 19137 6016 19457 7040
rect 19137 5952 19145 6016
rect 19209 5952 19225 6016
rect 19289 5952 19305 6016
rect 19369 5952 19385 6016
rect 19449 5952 19457 6016
rect 19011 5676 19077 5677
rect 19011 5612 19012 5676
rect 19076 5612 19077 5676
rect 19011 5611 19077 5612
rect 18459 5540 18525 5541
rect 18459 5476 18460 5540
rect 18524 5476 18525 5540
rect 18459 5475 18525 5476
rect 19137 4928 19457 5952
rect 19137 4864 19145 4928
rect 19209 4864 19225 4928
rect 19289 4864 19305 4928
rect 19369 4864 19385 4928
rect 19449 4864 19457 4928
rect 18643 4452 18709 4453
rect 18643 4388 18644 4452
rect 18708 4388 18709 4452
rect 18643 4387 18709 4388
rect 18275 4044 18341 4045
rect 18275 3980 18276 4044
rect 18340 3980 18341 4044
rect 18275 3979 18341 3980
rect 18091 3364 18157 3365
rect 18091 3300 18092 3364
rect 18156 3300 18157 3364
rect 18091 3299 18157 3300
rect 17355 2684 17421 2685
rect 17355 2620 17356 2684
rect 17420 2620 17421 2684
rect 17355 2619 17421 2620
rect 17907 2684 17973 2685
rect 17907 2620 17908 2684
rect 17972 2620 17973 2684
rect 17907 2619 17973 2620
rect 17355 2548 17421 2549
rect 17355 2484 17356 2548
rect 17420 2484 17421 2548
rect 17355 2483 17421 2484
rect 17358 2410 17418 2483
rect 17174 2350 17418 2410
rect 18646 1869 18706 4387
rect 19137 3840 19457 4864
rect 19137 3776 19145 3840
rect 19209 3776 19225 3840
rect 19289 3776 19305 3840
rect 19369 3776 19385 3840
rect 19449 3776 19457 3840
rect 18827 3364 18893 3365
rect 18827 3300 18828 3364
rect 18892 3300 18893 3364
rect 18827 3299 18893 3300
rect 18643 1868 18709 1869
rect 18643 1804 18644 1868
rect 18708 1804 18709 1868
rect 18643 1803 18709 1804
rect 16987 1732 17053 1733
rect 16987 1668 16988 1732
rect 17052 1668 17053 1732
rect 16987 1667 17053 1668
rect 16538 1056 16546 1120
rect 16610 1056 16626 1120
rect 16690 1056 16706 1120
rect 16770 1056 16786 1120
rect 16850 1056 16858 1120
rect 16538 1040 16858 1056
rect 9627 916 9693 917
rect 9627 852 9628 916
rect 9692 852 9693 916
rect 9627 851 9693 852
rect 18830 645 18890 3299
rect 19011 3228 19077 3229
rect 19011 3164 19012 3228
rect 19076 3164 19077 3228
rect 19011 3163 19077 3164
rect 19014 1189 19074 3163
rect 19137 2752 19457 3776
rect 19137 2688 19145 2752
rect 19209 2688 19225 2752
rect 19289 2688 19305 2752
rect 19369 2688 19385 2752
rect 19449 2688 19457 2752
rect 19137 1664 19457 2688
rect 19137 1600 19145 1664
rect 19209 1600 19225 1664
rect 19289 1600 19305 1664
rect 19369 1600 19385 1664
rect 19449 1600 19457 1664
rect 19011 1188 19077 1189
rect 19011 1124 19012 1188
rect 19076 1124 19077 1188
rect 19011 1123 19077 1124
rect 19137 1040 19457 1600
rect 19934 917 19994 9691
rect 20118 4045 20178 22050
rect 20299 14924 20365 14925
rect 20299 14860 20300 14924
rect 20364 14860 20365 14924
rect 20299 14859 20365 14860
rect 20302 10573 20362 14859
rect 20299 10572 20365 10573
rect 20299 10508 20300 10572
rect 20364 10508 20365 10572
rect 20299 10507 20365 10508
rect 20486 9485 20546 42195
rect 21736 41376 22056 42400
rect 21736 41312 21744 41376
rect 21808 41312 21824 41376
rect 21888 41312 21904 41376
rect 21968 41312 21984 41376
rect 22048 41312 22056 41376
rect 21736 40288 22056 41312
rect 21736 40224 21744 40288
rect 21808 40224 21824 40288
rect 21888 40224 21904 40288
rect 21968 40224 21984 40288
rect 22048 40224 22056 40288
rect 21736 39200 22056 40224
rect 21736 39136 21744 39200
rect 21808 39136 21824 39200
rect 21888 39136 21904 39200
rect 21968 39136 21984 39200
rect 22048 39136 22056 39200
rect 21736 38112 22056 39136
rect 21736 38048 21744 38112
rect 21808 38048 21824 38112
rect 21888 38048 21904 38112
rect 21968 38048 21984 38112
rect 22048 38048 22056 38112
rect 21736 37024 22056 38048
rect 21736 36960 21744 37024
rect 21808 36960 21824 37024
rect 21888 36960 21904 37024
rect 21968 36960 21984 37024
rect 22048 36960 22056 37024
rect 21736 35936 22056 36960
rect 21736 35872 21744 35936
rect 21808 35872 21824 35936
rect 21888 35872 21904 35936
rect 21968 35872 21984 35936
rect 22048 35872 22056 35936
rect 21736 34848 22056 35872
rect 21736 34784 21744 34848
rect 21808 34784 21824 34848
rect 21888 34784 21904 34848
rect 21968 34784 21984 34848
rect 22048 34784 22056 34848
rect 21035 34508 21101 34509
rect 21035 34444 21036 34508
rect 21100 34444 21101 34508
rect 21035 34443 21101 34444
rect 20851 30428 20917 30429
rect 20851 30364 20852 30428
rect 20916 30364 20917 30428
rect 20851 30363 20917 30364
rect 20667 30156 20733 30157
rect 20667 30092 20668 30156
rect 20732 30092 20733 30156
rect 20667 30091 20733 30092
rect 20483 9484 20549 9485
rect 20483 9420 20484 9484
rect 20548 9420 20549 9484
rect 20483 9419 20549 9420
rect 20115 4044 20181 4045
rect 20115 3980 20116 4044
rect 20180 3980 20181 4044
rect 20115 3979 20181 3980
rect 20670 917 20730 30091
rect 20854 19413 20914 30363
rect 20851 19412 20917 19413
rect 20851 19348 20852 19412
rect 20916 19348 20917 19412
rect 20851 19347 20917 19348
rect 21038 2277 21098 34443
rect 21736 33760 22056 34784
rect 21736 33696 21744 33760
rect 21808 33696 21824 33760
rect 21888 33696 21904 33760
rect 21968 33696 21984 33760
rect 22048 33696 22056 33760
rect 21736 32672 22056 33696
rect 21736 32608 21744 32672
rect 21808 32608 21824 32672
rect 21888 32608 21904 32672
rect 21968 32608 21984 32672
rect 22048 32608 22056 32672
rect 21736 31584 22056 32608
rect 21736 31520 21744 31584
rect 21808 31520 21824 31584
rect 21888 31520 21904 31584
rect 21968 31520 21984 31584
rect 22048 31520 22056 31584
rect 21736 30496 22056 31520
rect 21736 30432 21744 30496
rect 21808 30432 21824 30496
rect 21888 30432 21904 30496
rect 21968 30432 21984 30496
rect 22048 30432 22056 30496
rect 21736 29408 22056 30432
rect 21736 29344 21744 29408
rect 21808 29344 21824 29408
rect 21888 29344 21904 29408
rect 21968 29344 21984 29408
rect 22048 29344 22056 29408
rect 21736 28320 22056 29344
rect 21736 28256 21744 28320
rect 21808 28256 21824 28320
rect 21888 28256 21904 28320
rect 21968 28256 21984 28320
rect 22048 28256 22056 28320
rect 21736 27232 22056 28256
rect 21736 27168 21744 27232
rect 21808 27168 21824 27232
rect 21888 27168 21904 27232
rect 21968 27168 21984 27232
rect 22048 27168 22056 27232
rect 21736 26144 22056 27168
rect 21736 26080 21744 26144
rect 21808 26080 21824 26144
rect 21888 26080 21904 26144
rect 21968 26080 21984 26144
rect 22048 26080 22056 26144
rect 21736 25056 22056 26080
rect 21736 24992 21744 25056
rect 21808 24992 21824 25056
rect 21888 24992 21904 25056
rect 21968 24992 21984 25056
rect 22048 24992 22056 25056
rect 21736 23968 22056 24992
rect 21736 23904 21744 23968
rect 21808 23904 21824 23968
rect 21888 23904 21904 23968
rect 21968 23904 21984 23968
rect 22048 23904 22056 23968
rect 21403 23492 21469 23493
rect 21403 23428 21404 23492
rect 21468 23428 21469 23492
rect 21403 23427 21469 23428
rect 21219 23356 21285 23357
rect 21219 23292 21220 23356
rect 21284 23292 21285 23356
rect 21219 23291 21285 23292
rect 21222 17237 21282 23291
rect 21219 17236 21285 17237
rect 21219 17172 21220 17236
rect 21284 17172 21285 17236
rect 21219 17171 21285 17172
rect 21406 2277 21466 23427
rect 21736 22880 22056 23904
rect 21736 22816 21744 22880
rect 21808 22816 21824 22880
rect 21888 22816 21904 22880
rect 21968 22816 21984 22880
rect 22048 22816 22056 22880
rect 21736 21792 22056 22816
rect 21736 21728 21744 21792
rect 21808 21728 21824 21792
rect 21888 21728 21904 21792
rect 21968 21728 21984 21792
rect 22048 21728 22056 21792
rect 21736 20704 22056 21728
rect 21736 20640 21744 20704
rect 21808 20640 21824 20704
rect 21888 20640 21904 20704
rect 21968 20640 21984 20704
rect 22048 20640 22056 20704
rect 21736 19616 22056 20640
rect 21736 19552 21744 19616
rect 21808 19552 21824 19616
rect 21888 19552 21904 19616
rect 21968 19552 21984 19616
rect 22048 19552 22056 19616
rect 21736 18528 22056 19552
rect 21736 18464 21744 18528
rect 21808 18464 21824 18528
rect 21888 18464 21904 18528
rect 21968 18464 21984 18528
rect 22048 18464 22056 18528
rect 21736 17440 22056 18464
rect 21736 17376 21744 17440
rect 21808 17376 21824 17440
rect 21888 17376 21904 17440
rect 21968 17376 21984 17440
rect 22048 17376 22056 17440
rect 21736 16352 22056 17376
rect 21736 16288 21744 16352
rect 21808 16288 21824 16352
rect 21888 16288 21904 16352
rect 21968 16288 21984 16352
rect 22048 16288 22056 16352
rect 21736 15264 22056 16288
rect 21736 15200 21744 15264
rect 21808 15200 21824 15264
rect 21888 15200 21904 15264
rect 21968 15200 21984 15264
rect 22048 15200 22056 15264
rect 21736 14176 22056 15200
rect 21736 14112 21744 14176
rect 21808 14112 21824 14176
rect 21888 14112 21904 14176
rect 21968 14112 21984 14176
rect 22048 14112 22056 14176
rect 21736 13088 22056 14112
rect 21736 13024 21744 13088
rect 21808 13024 21824 13088
rect 21888 13024 21904 13088
rect 21968 13024 21984 13088
rect 22048 13024 22056 13088
rect 21736 12000 22056 13024
rect 21736 11936 21744 12000
rect 21808 11936 21824 12000
rect 21888 11936 21904 12000
rect 21968 11936 21984 12000
rect 22048 11936 22056 12000
rect 21736 10912 22056 11936
rect 21736 10848 21744 10912
rect 21808 10848 21824 10912
rect 21888 10848 21904 10912
rect 21968 10848 21984 10912
rect 22048 10848 22056 10912
rect 21736 9824 22056 10848
rect 21736 9760 21744 9824
rect 21808 9760 21824 9824
rect 21888 9760 21904 9824
rect 21968 9760 21984 9824
rect 22048 9760 22056 9824
rect 21736 8736 22056 9760
rect 21736 8672 21744 8736
rect 21808 8672 21824 8736
rect 21888 8672 21904 8736
rect 21968 8672 21984 8736
rect 22048 8672 22056 8736
rect 21736 7648 22056 8672
rect 21736 7584 21744 7648
rect 21808 7584 21824 7648
rect 21888 7584 21904 7648
rect 21968 7584 21984 7648
rect 22048 7584 22056 7648
rect 21736 6560 22056 7584
rect 21736 6496 21744 6560
rect 21808 6496 21824 6560
rect 21888 6496 21904 6560
rect 21968 6496 21984 6560
rect 22048 6496 22056 6560
rect 21736 5472 22056 6496
rect 21736 5408 21744 5472
rect 21808 5408 21824 5472
rect 21888 5408 21904 5472
rect 21968 5408 21984 5472
rect 22048 5408 22056 5472
rect 21736 4384 22056 5408
rect 21736 4320 21744 4384
rect 21808 4320 21824 4384
rect 21888 4320 21904 4384
rect 21968 4320 21984 4384
rect 22048 4320 22056 4384
rect 21736 3296 22056 4320
rect 21736 3232 21744 3296
rect 21808 3232 21824 3296
rect 21888 3232 21904 3296
rect 21968 3232 21984 3296
rect 22048 3232 22056 3296
rect 21035 2276 21101 2277
rect 21035 2212 21036 2276
rect 21100 2212 21101 2276
rect 21035 2211 21101 2212
rect 21403 2276 21469 2277
rect 21403 2212 21404 2276
rect 21468 2212 21469 2276
rect 21403 2211 21469 2212
rect 21736 2208 22056 3232
rect 21736 2144 21744 2208
rect 21808 2144 21824 2208
rect 21888 2144 21904 2208
rect 21968 2144 21984 2208
rect 22048 2144 22056 2208
rect 21736 1120 22056 2144
rect 21736 1056 21744 1120
rect 21808 1056 21824 1120
rect 21888 1056 21904 1120
rect 21968 1056 21984 1120
rect 22048 1056 22056 1120
rect 21736 1040 22056 1056
rect 19931 916 19997 917
rect 19931 852 19932 916
rect 19996 852 19997 916
rect 19931 851 19997 852
rect 20667 916 20733 917
rect 20667 852 20668 916
rect 20732 852 20733 916
rect 20667 851 20733 852
rect 18827 644 18893 645
rect 18827 580 18828 644
rect 18892 580 18893 644
rect 18827 579 18893 580
rect 8523 100 8589 101
rect 8523 36 8524 100
rect 8588 36 8589 100
rect 8523 35 8589 36
use sky130_fd_sc_hd__clkbuf_1  _000_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 21344 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _001_
timestamp 1688980957
transform 1 0 20976 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _002_
timestamp 1688980957
transform 1 0 20700 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _003_
timestamp 1688980957
transform 1 0 20608 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _004_
timestamp 1688980957
transform 1 0 20792 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _005_
timestamp 1688980957
transform 1 0 20792 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _006_
timestamp 1688980957
transform 1 0 20976 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _007_
timestamp 1688980957
transform 1 0 21344 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _008_
timestamp 1688980957
transform 1 0 20976 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _009_
timestamp 1688980957
transform 1 0 20792 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _010_
timestamp 1688980957
transform 1 0 18952 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _011_
timestamp 1688980957
transform 1 0 19688 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _012_
timestamp 1688980957
transform 1 0 20792 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _013_
timestamp 1688980957
transform 1 0 20516 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _014_
timestamp 1688980957
transform 1 0 20792 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _015_
timestamp 1688980957
transform 1 0 19504 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _016_
timestamp 1688980957
transform 1 0 20792 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _017_
timestamp 1688980957
transform 1 0 20056 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _018_
timestamp 1688980957
transform 1 0 20792 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _019_
timestamp 1688980957
transform 1 0 20792 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _020_
timestamp 1688980957
transform 1 0 20792 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _021_
timestamp 1688980957
transform 1 0 20516 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _022_
timestamp 1688980957
transform 1 0 20792 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _023_
timestamp 1688980957
transform 1 0 20516 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _024_
timestamp 1688980957
transform 1 0 20792 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _025_
timestamp 1688980957
transform 1 0 20056 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _026_
timestamp 1688980957
transform 1 0 20792 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _027_
timestamp 1688980957
transform 1 0 19964 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _028_
timestamp 1688980957
transform 1 0 19504 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _029_
timestamp 1688980957
transform 1 0 20240 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _030_
timestamp 1688980957
transform 1 0 20516 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _031_
timestamp 1688980957
transform 1 0 18584 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _032_
timestamp 1688980957
transform 1 0 16100 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _033_
timestamp 1688980957
transform 1 0 18952 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _034_
timestamp 1688980957
transform 1 0 18216 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _035_
timestamp 1688980957
transform 1 0 20240 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _036_
timestamp 1688980957
transform 1 0 20792 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _037_
timestamp 1688980957
transform 1 0 18676 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _038_
timestamp 1688980957
transform 1 0 17940 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _039_
timestamp 1688980957
transform 1 0 17756 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _040_
timestamp 1688980957
transform 1 0 17664 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _041_
timestamp 1688980957
transform 1 0 19412 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _042_
timestamp 1688980957
transform 1 0 18032 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _043_
timestamp 1688980957
transform 1 0 19228 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _044_
timestamp 1688980957
transform 1 0 17756 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _045_
timestamp 1688980957
transform 1 0 19136 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _046_
timestamp 1688980957
transform 1 0 18032 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _047_
timestamp 1688980957
transform 1 0 17480 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _048_
timestamp 1688980957
transform 1 0 19964 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _049_
timestamp 1688980957
transform 1 0 18308 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _050_
timestamp 1688980957
transform 1 0 18584 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _051_
timestamp 1688980957
transform 1 0 19412 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _052_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 17204 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _053_
timestamp 1688980957
transform 1 0 1748 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _054_
timestamp 1688980957
transform 1 0 3404 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _055_
timestamp 1688980957
transform 1 0 3956 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _056_
timestamp 1688980957
transform 1 0 1748 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _057_
timestamp 1688980957
transform 1 0 2484 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _058_
timestamp 1688980957
transform 1 0 3128 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _059_
timestamp 1688980957
transform 1 0 3772 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _060_
timestamp 1688980957
transform 1 0 10304 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _061_
timestamp 1688980957
transform 1 0 2760 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _062_
timestamp 1688980957
transform 1 0 3036 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _063_
timestamp 1688980957
transform 1 0 5152 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _064_
timestamp 1688980957
transform 1 0 4324 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _065_
timestamp 1688980957
transform 1 0 4600 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _066_
timestamp 1688980957
transform 1 0 4048 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _067_
timestamp 1688980957
transform 1 0 4876 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _068_
timestamp 1688980957
transform 1 0 5428 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _069_
timestamp 1688980957
transform 1 0 5428 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _070_
timestamp 1688980957
transform 1 0 5980 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _071_
timestamp 1688980957
transform 1 0 6164 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _072_
timestamp 1688980957
transform 1 0 5704 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _073_
timestamp 1688980957
transform 1 0 5428 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _074_
timestamp 1688980957
transform 1 0 5704 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _075_
timestamp 1688980957
transform 1 0 5980 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _076_
timestamp 1688980957
transform 1 0 7268 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _077_
timestamp 1688980957
transform 1 0 5980 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _078_
timestamp 1688980957
transform 1 0 8372 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _079_
timestamp 1688980957
transform 1 0 7452 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _080_
timestamp 1688980957
transform 1 0 7728 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _081_
timestamp 1688980957
transform 1 0 8556 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _082_
timestamp 1688980957
transform 1 0 9752 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _083_
timestamp 1688980957
transform 1 0 9200 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _084_
timestamp 1688980957
transform 1 0 9476 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _085_
timestamp 1688980957
transform 1 0 10580 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _086_
timestamp 1688980957
transform 1 0 8924 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _087_
timestamp 1688980957
transform 1 0 11040 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _088_
timestamp 1688980957
transform 1 0 10028 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _089_
timestamp 1688980957
transform 1 0 9200 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _090_
timestamp 1688980957
transform 1 0 9844 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _091_
timestamp 1688980957
transform 1 0 13616 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _092_
timestamp 1688980957
transform 1 0 12328 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _093_
timestamp 1688980957
transform 1 0 10488 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _094_
timestamp 1688980957
transform 1 0 4692 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _095_
timestamp 1688980957
transform 1 0 11684 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _096_
timestamp 1688980957
transform 1 0 12604 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _097_
timestamp 1688980957
transform 1 0 7084 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _098_
timestamp 1688980957
transform 1 0 12052 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _099_
timestamp 1688980957
transform 1 0 12880 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _100_
timestamp 1688980957
transform 1 0 9292 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _101_
timestamp 1688980957
transform 1 0 10488 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _102_
timestamp 1688980957
transform 1 0 8464 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _103_
timestamp 1688980957
transform 1 0 9936 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _104_
timestamp 1688980957
transform 1 0 11500 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _105_
timestamp 1688980957
transform 1 0 10212 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _106_
timestamp 1688980957
transform 1 0 10764 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _107_
timestamp 1688980957
transform 1 0 11408 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _108_
timestamp 1688980957
transform 1 0 13340 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _109_
timestamp 1688980957
transform 1 0 18308 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _110_
timestamp 1688980957
transform 1 0 14904 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _111_
timestamp 1688980957
transform 1 0 15180 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _112_
timestamp 1688980957
transform 1 0 16100 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _113_
timestamp 1688980957
transform 1 0 14904 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _114_
timestamp 1688980957
transform 1 0 16468 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _115_
timestamp 1688980957
transform 1 0 15180 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _116_
timestamp 1688980957
transform 1 0 15456 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _117_
timestamp 1688980957
transform 1 0 17756 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _118_
timestamp 1688980957
transform 1 0 17020 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _119_
timestamp 1688980957
transform 1 0 17296 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _120_
timestamp 1688980957
transform 1 0 16744 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _121_
timestamp 1688980957
transform 1 0 8924 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _122_
timestamp 1688980957
transform 1 0 15180 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _123_
timestamp 1688980957
transform 1 0 18032 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _124_
timestamp 1688980957
transform 1 0 5704 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _125_
timestamp 1688980957
transform 1 0 7912 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _126_
timestamp 1688980957
transform 1 0 5244 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _127_
timestamp 1688980957
transform 1 0 11592 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _128_
timestamp 1688980957
transform 1 0 10672 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _129_
timestamp 1688980957
transform 1 0 5704 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _130_
timestamp 1688980957
transform 1 0 4968 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _131_
timestamp 1688980957
transform 1 0 8096 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _132_
timestamp 1688980957
transform 1 0 10948 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _133_
timestamp 1688980957
transform 1 0 1380 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _134_
timestamp 1688980957
transform 1 0 8924 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _135_
timestamp 1688980957
transform 1 0 13708 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _136_
timestamp 1688980957
transform 1 0 3772 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _137_
timestamp 1688980957
transform 1 0 1472 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _138_
timestamp 1688980957
transform 1 0 3956 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _139_
timestamp 1688980957
transform 1 0 8556 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _140_
timestamp 1688980957
transform 1 0 10672 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _141_
timestamp 1688980957
transform 1 0 3864 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _142_
timestamp 1688980957
transform 1 0 5152 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _143_
timestamp 1688980957
transform 1 0 8372 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _144_
timestamp 1688980957
transform 1 0 15732 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _145_
timestamp 1688980957
transform 1 0 4232 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _146_
timestamp 1688980957
transform 1 0 1380 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _147_
timestamp 1688980957
transform 1 0 14076 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _148_
timestamp 1688980957
transform 1 0 14076 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _149_
timestamp 1688980957
transform 1 0 4600 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _150_
timestamp 1688980957
transform 1 0 6900 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _151_
timestamp 1688980957
transform 1 0 5704 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _152_
timestamp 1688980957
transform 1 0 11500 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _153_
timestamp 1688980957
transform 1 0 2852 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _154_
timestamp 1688980957
transform 1 0 3404 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _155_
timestamp 1688980957
transform 1 0 14812 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _156_
timestamp 1688980957
transform 1 0 3404 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _157_
timestamp 1688980957
transform 1 0 6900 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _158_
timestamp 1688980957
transform 1 0 8924 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _159_
timestamp 1688980957
transform 1 0 2024 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _160_
timestamp 1688980957
transform 1 0 6440 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _161_
timestamp 1688980957
transform 1 0 8924 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _162_
timestamp 1688980957
transform 1 0 1380 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _163_
timestamp 1688980957
transform 1 0 3772 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _164_
timestamp 1688980957
transform 1 0 11040 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _165_
timestamp 1688980957
transform 1 0 3772 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _166_
timestamp 1688980957
transform 1 0 8372 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _167_
timestamp 1688980957
transform 1 0 2024 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _168_
timestamp 1688980957
transform 1 0 10764 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _169_
timestamp 1688980957
transform 1 0 5796 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _170_
timestamp 1688980957
transform 1 0 5980 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _171_
timestamp 1688980957
transform 1 0 15456 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4784 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1688980957
transform 1 0 9936 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1688980957
transform 1 0 9660 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_4
timestamp 1688980957
transform 1 0 13248 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_5
timestamp 1688980957
transform 1 0 11224 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_6
timestamp 1688980957
transform 1 0 12512 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_7
timestamp 1688980957
transform 1 0 12880 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_8
timestamp 1688980957
transform 1 0 14260 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_9
timestamp 1688980957
transform 1 0 9568 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_10
timestamp 1688980957
transform 1 0 9200 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_11
timestamp 1688980957
transform 1 0 6440 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_12
timestamp 1688980957
transform 1 0 8556 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_13
timestamp 1688980957
transform 1 0 8188 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_14
timestamp 1688980957
transform 1 0 6808 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_15
timestamp 1688980957
transform 1 0 13156 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_16
timestamp 1688980957
transform 1 0 19688 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_17
timestamp 1688980957
transform 1 0 21160 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_18
timestamp 1688980957
transform 1 0 15640 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_19
timestamp 1688980957
transform 1 0 11132 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_20
timestamp 1688980957
transform 1 0 5244 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_21
timestamp 1688980957
transform 1 0 9660 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_22
timestamp 1688980957
transform 1 0 1564 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_23
timestamp 1688980957
transform 1 0 7728 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_24
timestamp 1688980957
transform 1 0 6716 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_25
timestamp 1688980957
transform 1 0 5612 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_26
timestamp 1688980957
transform 1 0 10764 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_27
timestamp 1688980957
transform 1 0 5796 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_28
timestamp 1688980957
transform 1 0 12236 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_29
timestamp 1688980957
transform 1 0 19504 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_30
timestamp 1688980957
transform 1 0 7084 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_31
timestamp 1688980957
transform 1 0 2852 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_32
timestamp 1688980957
transform 1 0 7728 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_33
timestamp 1688980957
transform 1 0 5336 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_34
timestamp 1688980957
transform 1 0 5612 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_35
timestamp 1688980957
transform 1 0 1564 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_36
timestamp 1688980957
transform 1 0 2116 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_37
timestamp 1688980957
transform 1 0 3036 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__diode_2  ANTENNA_38
timestamp 1688980957
transform 1 0 6900 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_0._0_
timestamp 1688980957
transform 1 0 19320 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_1._0_
timestamp 1688980957
transform 1 0 19964 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_2._0_
timestamp 1688980957
transform 1 0 19412 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_3._0_
timestamp 1688980957
transform 1 0 19964 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_4._0_
timestamp 1688980957
transform 1 0 20700 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_5._0_
timestamp 1688980957
transform 1 0 19780 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_6._0_
timestamp 1688980957
transform 1 0 19228 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_7._0_
timestamp 1688980957
transform 1 0 19872 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_8._0_
timestamp 1688980957
transform 1 0 18492 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_9._0_
timestamp 1688980957
transform 1 0 18676 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_10._0_
timestamp 1688980957
transform 1 0 19228 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_11._0_
timestamp 1688980957
transform 1 0 18860 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_12._0_
timestamp 1688980957
transform 1 0 19136 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_13._0_
timestamp 1688980957
transform 1 0 19228 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_14._0_
timestamp 1688980957
transform 1 0 19964 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_15._0_
timestamp 1688980957
transform 1 0 18860 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_16._0_
timestamp 1688980957
transform 1 0 20424 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_17._0_
timestamp 1688980957
transform 1 0 18400 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_18._0_
timestamp 1688980957
transform 1 0 19872 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_19._0_
timestamp 1688980957
transform 1 0 18768 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_20._0_
timestamp 1688980957
transform 1 0 19964 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_21._0_
timestamp 1688980957
transform 1 0 20516 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_22._0_
timestamp 1688980957
transform 1 0 20240 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_23._0_
timestamp 1688980957
transform 1 0 18584 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_24._0_
timestamp 1688980957
transform 1 0 19872 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_25._0_
timestamp 1688980957
transform 1 0 17848 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_26._0_
timestamp 1688980957
transform 1 0 19688 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_27._0_
timestamp 1688980957
transform 1 0 18032 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_28._0_
timestamp 1688980957
transform 1 0 19780 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_29._0_
timestamp 1688980957
transform 1 0 18860 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_30._0_
timestamp 1688980957
transform 1 0 19688 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_inbuf_31._0_
timestamp 1688980957
transform 1 0 18308 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_0._0_
timestamp 1688980957
transform 1 0 20056 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_1._0_
timestamp 1688980957
transform 1 0 20332 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_2._0_
timestamp 1688980957
transform 1 0 20424 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_3._0_
timestamp 1688980957
transform 1 0 20424 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_4._0_
timestamp 1688980957
transform 1 0 20332 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_5._0_
timestamp 1688980957
transform 1 0 20056 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_6._0_
timestamp 1688980957
transform 1 0 20332 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_7._0_
timestamp 1688980957
transform 1 0 20240 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_8._0_
timestamp 1688980957
transform 1 0 19596 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_9._0_
timestamp 1688980957
transform 1 0 19228 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_10._0_
timestamp 1688980957
transform 1 0 19964 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_11._0_
timestamp 1688980957
transform 1 0 19964 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_12._0_
timestamp 1688980957
transform 1 0 19964 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_13._0_
timestamp 1688980957
transform 1 0 20240 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_14._0_
timestamp 1688980957
transform 1 0 19412 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_15._0_
timestamp 1688980957
transform 1 0 20148 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_16._0_
timestamp 1688980957
transform 1 0 19688 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_17._0_
timestamp 1688980957
transform 1 0 19780 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_18._0_
timestamp 1688980957
transform 1 0 20884 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_19._0_
timestamp 1688980957
transform 1 0 19688 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_20._0_
timestamp 1688980957
transform 1 0 20240 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_21._0_
timestamp 1688980957
transform 1 0 20516 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_22._0_
timestamp 1688980957
transform 1 0 20240 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_23._0_
timestamp 1688980957
transform 1 0 19688 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_24._0_
timestamp 1688980957
transform 1 0 19964 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_25._0_
timestamp 1688980957
transform 1 0 18768 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_26._0_
timestamp 1688980957
transform 1 0 20332 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_27._0_
timestamp 1688980957
transform 1 0 19136 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_28._0_
timestamp 1688980957
transform 1 0 20516 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_29._0_
timestamp 1688980957
transform 1 0 20240 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_30._0_
timestamp 1688980957
transform 1 0 17204 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  data_outbuf_31._0_
timestamp 1688980957
transform 1 0 19412 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_9 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1932 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_29
timestamp 1688980957
transform 1 0 3772 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_57 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 6348 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_62
timestamp 1688980957
transform 1 0 6808 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_0_101
timestamp 1688980957
transform 1 0 10396 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_110 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 11224 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_139
timestamp 1688980957
transform 1 0 13892 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_175
timestamp 1688980957
transform 1 0 17204 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_221
timestamp 1688980957
transform 1 0 21436 0 1 1088
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_21
timestamp 1688980957
transform 1 0 3036 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_55
timestamp 1688980957
transform 1 0 6164 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_1_57
timestamp 1688980957
transform 1 0 6348 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_125
timestamp 1688980957
transform 1 0 12604 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_130
timestamp 1688980957
transform 1 0 13064 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_167
timestamp 1688980957
transform 1 0 16468 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_1_221
timestamp 1688980957
transform 1 0 21436 0 -1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_3
timestamp 1688980957
transform 1 0 1380 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_7
timestamp 1688980957
transform 1 0 1748 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_21
timestamp 1688980957
transform 1 0 3036 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_38
timestamp 1688980957
transform 1 0 4600 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_45
timestamp 1688980957
transform 1 0 5244 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_50
timestamp 1688980957
transform 1 0 5704 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_61
timestamp 1688980957
transform 1 0 6716 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_2_85
timestamp 1688980957
transform 1 0 8924 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_90
timestamp 1688980957
transform 1 0 9384 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_94
timestamp 1688980957
transform 1 0 9752 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_108
timestamp 1688980957
transform 1 0 11040 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_118
timestamp 1688980957
transform 1 0 11960 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_122
timestamp 1688980957
transform 1 0 12328 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_126
timestamp 1688980957
transform 1 0 12696 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_130
timestamp 1688980957
transform 1 0 13064 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_134
timestamp 1688980957
transform 1 0 13432 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_139
timestamp 1688980957
transform 1 0 13892 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_141
timestamp 1688980957
transform 1 0 14076 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_148
timestamp 1688980957
transform 1 0 14720 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_153
timestamp 1688980957
transform 1 0 15180 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_173
timestamp 1688980957
transform 1 0 17020 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_190
timestamp 1688980957
transform 1 0 18584 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_2_221
timestamp 1688980957
transform 1 0 21436 0 1 2176
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_3
timestamp 1688980957
transform 1 0 1380 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_48 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5520 0 -1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_57
timestamp 1688980957
transform 1 0 6348 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_96
timestamp 1688980957
transform 1 0 9936 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_100
timestamp 1688980957
transform 1 0 10304 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_105
timestamp 1688980957
transform 1 0 10764 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_3_116 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 11776 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_3_128
timestamp 1688980957
transform 1 0 12880 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_133
timestamp 1688980957
transform 1 0 13340 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_156
timestamp 1688980957
transform 1 0 15456 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_166
timestamp 1688980957
transform 1 0 16376 0 -1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_3
timestamp 1688980957
transform 1 0 1380 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_20
timestamp 1688980957
transform 1 0 2944 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_53 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5980 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_4_65 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 7084 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_72
timestamp 1688980957
transform 1 0 7728 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_76
timestamp 1688980957
transform 1 0 8096 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_91
timestamp 1688980957
transform 1 0 9476 0 1 3264
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_98
timestamp 1688980957
transform 1 0 10120 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_110
timestamp 1688980957
transform 1 0 11224 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_122
timestamp 1688980957
transform 1 0 12328 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_131
timestamp 1688980957
transform 1 0 13156 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_136
timestamp 1688980957
transform 1 0 13616 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_159
timestamp 1688980957
transform 1 0 15732 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_194
timestamp 1688980957
transform 1 0 18952 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_4_221
timestamp 1688980957
transform 1 0 21436 0 1 3264
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_3
timestamp 1688980957
transform 1 0 1380 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_5_53
timestamp 1688980957
transform 1 0 5980 0 -1 4352
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_57
timestamp 1688980957
transform 1 0 6348 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_69
timestamp 1688980957
transform 1 0 7452 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_81
timestamp 1688980957
transform 1 0 8556 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_93
timestamp 1688980957
transform 1 0 9660 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_5_105
timestamp 1688980957
transform 1 0 10764 0 -1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_111
timestamp 1688980957
transform 1 0 11316 0 -1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_113
timestamp 1688980957
transform 1 0 11500 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_125
timestamp 1688980957
transform 1 0 12604 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_137
timestamp 1688980957
transform 1 0 13708 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_141
timestamp 1688980957
transform 1 0 14076 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_148
timestamp 1688980957
transform 1 0 14720 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_5_169
timestamp 1688980957
transform 1 0 16652 0 -1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_177
timestamp 1688980957
transform 1 0 17388 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_200
timestamp 1688980957
transform 1 0 19504 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_6
timestamp 1688980957
transform 1 0 1656 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_29
timestamp 1688980957
transform 1 0 3772 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_60
timestamp 1688980957
transform 1 0 6624 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_72
timestamp 1688980957
transform 1 0 7728 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_85
timestamp 1688980957
transform 1 0 8924 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_97
timestamp 1688980957
transform 1 0 10028 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_109
timestamp 1688980957
transform 1 0 11132 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_121
timestamp 1688980957
transform 1 0 12236 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_6_133
timestamp 1688980957
transform 1 0 13340 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_139
timestamp 1688980957
transform 1 0 13892 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_141
timestamp 1688980957
transform 1 0 14076 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_6_161
timestamp 1688980957
transform 1 0 15916 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_203
timestamp 1688980957
transform 1 0 19780 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_221
timestamp 1688980957
transform 1 0 21436 0 1 4352
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_7_9
timestamp 1688980957
transform 1 0 1932 0 -1 5440
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_57
timestamp 1688980957
transform 1 0 6348 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_69
timestamp 1688980957
transform 1 0 7452 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_81
timestamp 1688980957
transform 1 0 8556 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_93
timestamp 1688980957
transform 1 0 9660 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_7_105
timestamp 1688980957
transform 1 0 10764 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_111
timestamp 1688980957
transform 1 0 11316 0 -1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_113
timestamp 1688980957
transform 1 0 11500 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_7_125
timestamp 1688980957
transform 1 0 12604 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_222
timestamp 1688980957
transform 1 0 21528 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_3
timestamp 1688980957
transform 1 0 1380 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_8_77
timestamp 1688980957
transform 1 0 8188 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_83
timestamp 1688980957
transform 1 0 8740 0 1 5440
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_85
timestamp 1688980957
transform 1 0 8924 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_8_97
timestamp 1688980957
transform 1 0 10028 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_104
timestamp 1688980957
transform 1 0 10672 0 1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_116
timestamp 1688980957
transform 1 0 11776 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_128
timestamp 1688980957
transform 1 0 12880 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_8_136
timestamp 1688980957
transform 1 0 13616 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_141
timestamp 1688980957
transform 1 0 14076 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_191
timestamp 1688980957
transform 1 0 18676 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_218
timestamp 1688980957
transform 1 0 21160 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_3
timestamp 1688980957
transform 1 0 1380 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_19
timestamp 1688980957
transform 1 0 2852 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_23
timestamp 1688980957
transform 1 0 3220 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_28
timestamp 1688980957
transform 1 0 3680 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_75
timestamp 1688980957
transform 1 0 8004 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_87
timestamp 1688980957
transform 1 0 9108 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_9_110
timestamp 1688980957
transform 1 0 11224 0 -1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_113
timestamp 1688980957
transform 1 0 11500 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_117
timestamp 1688980957
transform 1 0 11868 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_9_129
timestamp 1688980957
transform 1 0 12972 0 -1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_137
timestamp 1688980957
transform 1 0 13708 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_162
timestamp 1688980957
transform 1 0 16008 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_182
timestamp 1688980957
transform 1 0 17848 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_9
timestamp 1688980957
transform 1 0 1932 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_10_85
timestamp 1688980957
transform 1 0 8924 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_91
timestamp 1688980957
transform 1 0 9476 0 1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_122
timestamp 1688980957
transform 1 0 12328 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_134
timestamp 1688980957
transform 1 0 13432 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_10_159
timestamp 1688980957
transform 1 0 15732 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_167
timestamp 1688980957
transform 1 0 16468 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_197
timestamp 1688980957
transform 1 0 19228 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_221
timestamp 1688980957
transform 1 0 21436 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_3
timestamp 1688980957
transform 1 0 1380 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_55
timestamp 1688980957
transform 1 0 6164 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_69
timestamp 1688980957
transform 1 0 7452 0 -1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_128
timestamp 1688980957
transform 1 0 12880 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_11_140
timestamp 1688980957
transform 1 0 13984 0 -1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_154
timestamp 1688980957
transform 1 0 15272 0 -1 7616
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_188
timestamp 1688980957
transform 1 0 18400 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_221
timestamp 1688980957
transform 1 0 21436 0 -1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_9
timestamp 1688980957
transform 1 0 1932 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_29
timestamp 1688980957
transform 1 0 3772 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_48
timestamp 1688980957
transform 1 0 5520 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_82
timestamp 1688980957
transform 1 0 8648 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_88
timestamp 1688980957
transform 1 0 9200 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_107
timestamp 1688980957
transform 1 0 10948 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_12_130
timestamp 1688980957
transform 1 0 13064 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_136
timestamp 1688980957
transform 1 0 13616 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_156
timestamp 1688980957
transform 1 0 15456 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_197
timestamp 1688980957
transform 1 0 19228 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_12_218
timestamp 1688980957
transform 1 0 21160 0 1 7616
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_13_9
timestamp 1688980957
transform 1 0 1932 0 -1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_55
timestamp 1688980957
transform 1 0 6164 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_57
timestamp 1688980957
transform 1 0 6348 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_73
timestamp 1688980957
transform 1 0 7820 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_13_111
timestamp 1688980957
transform 1 0 11316 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_13_158
timestamp 1688980957
transform 1 0 15640 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_166
timestamp 1688980957
transform 1 0 16376 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_13_188
timestamp 1688980957
transform 1 0 18400 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_9
timestamp 1688980957
transform 1 0 1932 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_26
timestamp 1688980957
transform 1 0 3496 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_47
timestamp 1688980957
transform 1 0 5428 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_82
timestamp 1688980957
transform 1 0 8648 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_85
timestamp 1688980957
transform 1 0 8924 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_14_101
timestamp 1688980957
transform 1 0 10396 0 1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_14_133
timestamp 1688980957
transform 1 0 13340 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_139
timestamp 1688980957
transform 1 0 13892 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_195
timestamp 1688980957
transform 1 0 19044 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_14_197
timestamp 1688980957
transform 1 0 19228 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_9
timestamp 1688980957
transform 1 0 1932 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_13
timestamp 1688980957
transform 1 0 2300 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_15_66
timestamp 1688980957
transform 1 0 7176 0 -1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_15_107
timestamp 1688980957
transform 1 0 10948 0 -1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_111
timestamp 1688980957
transform 1 0 11316 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_113
timestamp 1688980957
transform 1 0 11500 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_15_140
timestamp 1688980957
transform 1 0 13984 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_146
timestamp 1688980957
transform 1 0 14536 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_15_165
timestamp 1688980957
transform 1 0 16284 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_15_169
timestamp 1688980957
transform 1 0 16652 0 -1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_177
timestamp 1688980957
transform 1 0 17388 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_15_222
timestamp 1688980957
transform 1 0 21528 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_3
timestamp 1688980957
transform 1 0 1380 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_41
timestamp 1688980957
transform 1 0 4876 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_58
timestamp 1688980957
transform 1 0 6440 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_85
timestamp 1688980957
transform 1 0 8924 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_89
timestamp 1688980957
transform 1 0 9292 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_16_105
timestamp 1688980957
transform 1 0 10764 0 1 9792
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_16_113
timestamp 1688980957
transform 1 0 11500 0 1 9792
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_16_136
timestamp 1688980957
transform 1 0 13616 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_16_141
timestamp 1688980957
transform 1 0 14076 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_16_177
timestamp 1688980957
transform 1 0 17388 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_16_212
timestamp 1688980957
transform 1 0 20608 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_3
timestamp 1688980957
transform 1 0 1380 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_11
timestamp 1688980957
transform 1 0 2116 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_34
timestamp 1688980957
transform 1 0 4232 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_57
timestamp 1688980957
transform 1 0 6348 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_61
timestamp 1688980957
transform 1 0 6716 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_65
timestamp 1688980957
transform 1 0 7084 0 -1 10880
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_17_113
timestamp 1688980957
transform 1 0 11500 0 -1 10880
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_161
timestamp 1688980957
transform 1 0 15916 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_167
timestamp 1688980957
transform 1 0 16468 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_169
timestamp 1688980957
transform 1 0 16652 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_17_175
timestamp 1688980957
transform 1 0 17204 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_17_191
timestamp 1688980957
transform 1 0 18676 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_17_215
timestamp 1688980957
transform 1 0 20884 0 -1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_3
timestamp 1688980957
transform 1 0 1380 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_11
timestamp 1688980957
transform 1 0 2116 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_18_29
timestamp 1688980957
transform 1 0 3772 0 1 10880
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_39
timestamp 1688980957
transform 1 0 4692 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_68
timestamp 1688980957
transform 1 0 7360 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_18_130
timestamp 1688980957
transform 1 0 13064 0 1 10880
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_138
timestamp 1688980957
transform 1 0 13800 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_18_156
timestamp 1688980957
transform 1 0 15456 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_18_172
timestamp 1688980957
transform 1 0 16928 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_194
timestamp 1688980957
transform 1 0 18952 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_197
timestamp 1688980957
transform 1 0 19228 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_18_221
timestamp 1688980957
transform 1 0 21436 0 1 10880
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_21
timestamp 1688980957
transform 1 0 3036 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_54
timestamp 1688980957
transform 1 0 6072 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_66
timestamp 1688980957
transform 1 0 7176 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_89
timestamp 1688980957
transform 1 0 9292 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_19_113
timestamp 1688980957
transform 1 0 11500 0 -1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_19_121
timestamp 1688980957
transform 1 0 12236 0 -1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_19_144
timestamp 1688980957
transform 1 0 14352 0 -1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_148
timestamp 1688980957
transform 1 0 14720 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_167
timestamp 1688980957
transform 1 0 16468 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_19_169
timestamp 1688980957
transform 1 0 16652 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_19_191
timestamp 1688980957
transform 1 0 18676 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_9
timestamp 1688980957
transform 1 0 1932 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_32
timestamp 1688980957
transform 1 0 4048 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_85
timestamp 1688980957
transform 1 0 8924 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_93
timestamp 1688980957
transform 1 0 9660 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_116
timestamp 1688980957
transform 1 0 11776 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_124
timestamp 1688980957
transform 1 0 12512 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_20_141
timestamp 1688980957
transform 1 0 14076 0 1 11968
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_149
timestamp 1688980957
transform 1 0 14812 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_166
timestamp 1688980957
transform 1 0 16376 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_20_170
timestamp 1688980957
transform 1 0 16744 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_20_192
timestamp 1688980957
transform 1 0 18768 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_20_197
timestamp 1688980957
transform 1 0 19228 0 1 11968
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_3
timestamp 1688980957
transform 1 0 1380 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_11
timestamp 1688980957
transform 1 0 2116 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_34
timestamp 1688980957
transform 1 0 4232 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_38
timestamp 1688980957
transform 1 0 4600 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_21_54
timestamp 1688980957
transform 1 0 6072 0 -1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_57
timestamp 1688980957
transform 1 0 6348 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_76
timestamp 1688980957
transform 1 0 8096 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_0_21_113
timestamp 1688980957
transform 1 0 11500 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_21_164
timestamp 1688980957
transform 1 0 16192 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_21_169
timestamp 1688980957
transform 1 0 16652 0 -1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_177
timestamp 1688980957
transform 1 0 17388 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_21_184
timestamp 1688980957
transform 1 0 18032 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_21_209
timestamp 1688980957
transform 1 0 20332 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_3
timestamp 1688980957
transform 1 0 1380 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_11
timestamp 1688980957
transform 1 0 2116 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_27
timestamp 1688980957
transform 1 0 3588 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_50
timestamp 1688980957
transform 1 0 5704 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_22_88
timestamp 1688980957
transform 1 0 9200 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_22_130
timestamp 1688980957
transform 1 0 13064 0 1 13056
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_138
timestamp 1688980957
transform 1 0 13800 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_162
timestamp 1688980957
transform 1 0 16008 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_178
timestamp 1688980957
transform 1 0 17480 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_22_200
timestamp 1688980957
transform 1 0 19504 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_22_216
timestamp 1688980957
transform 1 0 20976 0 1 13056
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_12
timestamp 1688980957
transform 1 0 2208 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_18
timestamp 1688980957
transform 1 0 2760 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_21
timestamp 1688980957
transform 1 0 3036 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_23_38
timestamp 1688980957
transform 1 0 4600 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_57
timestamp 1688980957
transform 1 0 6348 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_77
timestamp 1688980957
transform 1 0 8188 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_83
timestamp 1688980957
transform 1 0 8740 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_23_111
timestamp 1688980957
transform 1 0 11316 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_23_113
timestamp 1688980957
transform 1 0 11500 0 -1 14144
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_23_132
timestamp 1688980957
transform 1 0 13248 0 -1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_23_144
timestamp 1688980957
transform 1 0 14352 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_23_184
timestamp 1688980957
transform 1 0 18032 0 -1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_192
timestamp 1688980957
transform 1 0 18768 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_197
timestamp 1688980957
transform 1 0 19228 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_23_215
timestamp 1688980957
transform 1 0 20884 0 -1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_3
timestamp 1688980957
transform 1 0 1380 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_11
timestamp 1688980957
transform 1 0 2116 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_29
timestamp 1688980957
transform 1 0 3772 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_33
timestamp 1688980957
transform 1 0 4140 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_24_79
timestamp 1688980957
transform 1 0 8372 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_24_83
timestamp 1688980957
transform 1 0 8740 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_85
timestamp 1688980957
transform 1 0 8924 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_93
timestamp 1688980957
transform 1 0 9660 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_137
timestamp 1688980957
transform 1 0 13708 0 1 14144
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_162
timestamp 1688980957
transform 1 0 16008 0 1 14144
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_24_174
timestamp 1688980957
transform 1 0 17112 0 1 14144
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_24_186
timestamp 1688980957
transform 1 0 18216 0 1 14144
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_24_194
timestamp 1688980957
transform 1 0 18952 0 1 14144
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_24_197
timestamp 1688980957
transform 1 0 19228 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_3
timestamp 1688980957
transform 1 0 1380 0 -1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_78
timestamp 1688980957
transform 1 0 8280 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_25_113
timestamp 1688980957
transform 1 0 11500 0 -1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_25_134
timestamp 1688980957
transform 1 0 13432 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_25_158
timestamp 1688980957
transform 1 0 15640 0 -1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_25_166
timestamp 1688980957
transform 1 0 16376 0 -1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_25_169
timestamp 1688980957
transform 1 0 16652 0 -1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_196
timestamp 1688980957
transform 1 0 19136 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_200
timestamp 1688980957
transform 1 0 19504 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_25_204
timestamp 1688980957
transform 1 0 19872 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_211
timestamp 1688980957
transform 1 0 20516 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_25_218
timestamp 1688980957
transform 1 0 21160 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_18
timestamp 1688980957
transform 1 0 2760 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_56
timestamp 1688980957
transform 1 0 6256 0 1 15232
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_26_76
timestamp 1688980957
transform 1 0 8096 0 1 15232
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_26_85
timestamp 1688980957
transform 1 0 8924 0 1 15232
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_103
timestamp 1688980957
transform 1 0 10580 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_26_115
timestamp 1688980957
transform 1 0 11684 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_26_144
timestamp 1688980957
transform 1 0 14352 0 1 15232
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_26_161
timestamp 1688980957
transform 1 0 15916 0 1 15232
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_26_213
timestamp 1688980957
transform 1 0 20700 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_9
timestamp 1688980957
transform 1 0 1932 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_39
timestamp 1688980957
transform 1 0 4692 0 -1 16320
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_27_57
timestamp 1688980957
transform 1 0 6348 0 -1 16320
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_69
timestamp 1688980957
transform 1 0 7452 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_74
timestamp 1688980957
transform 1 0 7912 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27_113
timestamp 1688980957
transform 1 0 11500 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_165
timestamp 1688980957
transform 1 0 16284 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_184
timestamp 1688980957
transform 1 0 18032 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_27_190
timestamp 1688980957
transform 1 0 18584 0 -1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_27_198
timestamp 1688980957
transform 1 0 19320 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_28_3
timestamp 1688980957
transform 1 0 1380 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_7
timestamp 1688980957
transform 1 0 1748 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_23
timestamp 1688980957
transform 1 0 3220 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_41
timestamp 1688980957
transform 1 0 4876 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_63
timestamp 1688980957
transform 1 0 6900 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_67
timestamp 1688980957
transform 1 0 7268 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_121
timestamp 1688980957
transform 1 0 12236 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_138
timestamp 1688980957
transform 1 0 13800 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_28_144
timestamp 1688980957
transform 1 0 14352 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_28_186
timestamp 1688980957
transform 1 0 18216 0 1 16320
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_28_194
timestamp 1688980957
transform 1 0 18952 0 1 16320
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_28_197
timestamp 1688980957
transform 1 0 19228 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_3
timestamp 1688980957
transform 1 0 1380 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_8
timestamp 1688980957
transform 1 0 1840 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_29_53
timestamp 1688980957
transform 1 0 5980 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_29_57
timestamp 1688980957
transform 1 0 6348 0 -1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_63
timestamp 1688980957
transform 1 0 6900 0 -1 17408
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_29_82
timestamp 1688980957
transform 1 0 8648 0 -1 17408
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_29_94
timestamp 1688980957
transform 1 0 9752 0 -1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_111
timestamp 1688980957
transform 1 0 11316 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_29_116
timestamp 1688980957
transform 1 0 11776 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_29_141
timestamp 1688980957
transform 1 0 14076 0 -1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_152
timestamp 1688980957
transform 1 0 15088 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_29_193
timestamp 1688980957
transform 1 0 18860 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_30_29
timestamp 1688980957
transform 1 0 3772 0 1 17408
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_37
timestamp 1688980957
transform 1 0 4508 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_41
timestamp 1688980957
transform 1 0 4876 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_45
timestamp 1688980957
transform 1 0 5244 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_48
timestamp 1688980957
transform 1 0 5520 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_65
timestamp 1688980957
transform 1 0 7084 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_30_100
timestamp 1688980957
transform 1 0 10304 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_30_119
timestamp 1688980957
transform 1 0 12052 0 1 17408
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_195
timestamp 1688980957
transform 1 0 19044 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_200
timestamp 1688980957
transform 1 0 19504 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_208
timestamp 1688980957
transform 1 0 20240 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_30_213
timestamp 1688980957
transform 1 0 20700 0 1 17408
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_30_218
timestamp 1688980957
transform 1 0 21160 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_13
timestamp 1688980957
transform 1 0 2300 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_50
timestamp 1688980957
transform 1 0 5704 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_57
timestamp 1688980957
transform 1 0 6348 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_61
timestamp 1688980957
transform 1 0 6716 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_95
timestamp 1688980957
transform 1 0 9844 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_113
timestamp 1688980957
transform 1 0 11500 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_31_134
timestamp 1688980957
transform 1 0 13432 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_138
timestamp 1688980957
transform 1 0 13800 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_31_154
timestamp 1688980957
transform 1 0 15272 0 -1 18496
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_162
timestamp 1688980957
transform 1 0 16008 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_166
timestamp 1688980957
transform 1 0 16376 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_31_184
timestamp 1688980957
transform 1 0 18032 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_31_190
timestamp 1688980957
transform 1 0 18584 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_207
timestamp 1688980957
transform 1 0 20148 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_31_215
timestamp 1688980957
transform 1 0 20884 0 -1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_88
timestamp 1688980957
transform 1 0 9200 0 1 18496
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_32_105
timestamp 1688980957
transform 1 0 10764 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_129
timestamp 1688980957
transform 1 0 12972 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_32_136
timestamp 1688980957
transform 1 0 13616 0 1 18496
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_141
timestamp 1688980957
transform 1 0 14076 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_32_153
timestamp 1688980957
transform 1 0 15180 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_32_157
timestamp 1688980957
transform 1 0 15548 0 1 18496
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_32_184
timestamp 1688980957
transform 1 0 18032 0 1 18496
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_3
timestamp 1688980957
transform 1 0 1380 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_33_22
timestamp 1688980957
transform 1 0 3128 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_57
timestamp 1688980957
transform 1 0 6348 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_65
timestamp 1688980957
transform 1 0 7084 0 -1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_33_84
timestamp 1688980957
transform 1 0 8832 0 -1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_33_96
timestamp 1688980957
transform 1 0 9936 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_113
timestamp 1688980957
transform 1 0 11500 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_121
timestamp 1688980957
transform 1 0 12236 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_166
timestamp 1688980957
transform 1 0 16376 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_33_184
timestamp 1688980957
transform 1 0 18032 0 -1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_33_215
timestamp 1688980957
transform 1 0 20884 0 -1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_11
timestamp 1688980957
transform 1 0 2116 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_34_32
timestamp 1688980957
transform 1 0 4048 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_36
timestamp 1688980957
transform 1 0 4416 0 1 19584
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_34_70
timestamp 1688980957
transform 1 0 7544 0 1 19584
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_82
timestamp 1688980957
transform 1 0 8648 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_85
timestamp 1688980957
transform 1 0 8924 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_93
timestamp 1688980957
transform 1 0 9660 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_116
timestamp 1688980957
transform 1 0 11776 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_124
timestamp 1688980957
transform 1 0 12512 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_34_180
timestamp 1688980957
transform 1 0 17664 0 1 19584
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_188
timestamp 1688980957
transform 1 0 18400 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_34_213
timestamp 1688980957
transform 1 0 20700 0 1 19584
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_34_218
timestamp 1688980957
transform 1 0 21160 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_6
timestamp 1688980957
transform 1 0 1656 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_35_51
timestamp 1688980957
transform 1 0 5796 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_55
timestamp 1688980957
transform 1 0 6164 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_57
timestamp 1688980957
transform 1 0 6348 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_35_61
timestamp 1688980957
transform 1 0 6716 0 -1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_67
timestamp 1688980957
transform 1 0 7268 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_35_86
timestamp 1688980957
transform 1 0 9016 0 -1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_35_94
timestamp 1688980957
transform 1 0 9752 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_128
timestamp 1688980957
transform 1 0 12880 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_35_166
timestamp 1688980957
transform 1 0 16376 0 -1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_169
timestamp 1688980957
transform 1 0 16652 0 -1 20672
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_35_185
timestamp 1688980957
transform 1 0 18124 0 -1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_35_215
timestamp 1688980957
transform 1 0 20884 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_47
timestamp 1688980957
transform 1 0 5428 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_51
timestamp 1688980957
transform 1 0 5796 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_71
timestamp 1688980957
transform 1 0 7636 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_83
timestamp 1688980957
transform 1 0 8740 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_100
timestamp 1688980957
transform 1 0 10304 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_108
timestamp 1688980957
transform 1 0 11040 0 1 20672
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_125
timestamp 1688980957
transform 1 0 12604 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_137
timestamp 1688980957
transform 1 0 13708 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_156
timestamp 1688980957
transform 1 0 15456 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_36_166
timestamp 1688980957
transform 1 0 16376 0 1 20672
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_36_184
timestamp 1688980957
transform 1 0 18032 0 1 20672
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_36_197
timestamp 1688980957
transform 1 0 19228 0 1 20672
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_36_205
timestamp 1688980957
transform 1 0 19964 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_36_221
timestamp 1688980957
transform 1 0 21436 0 1 20672
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_3
timestamp 1688980957
transform 1 0 1380 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_37_49
timestamp 1688980957
transform 1 0 5612 0 -1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_53
timestamp 1688980957
transform 1 0 5980 0 -1 21760
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_57
timestamp 1688980957
transform 1 0 6348 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_69
timestamp 1688980957
transform 1 0 7452 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_37_106
timestamp 1688980957
transform 1 0 10856 0 -1 21760
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_131
timestamp 1688980957
transform 1 0 13156 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_143
timestamp 1688980957
transform 1 0 14260 0 -1 21760
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_37_155
timestamp 1688980957
transform 1 0 15364 0 -1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_37_167
timestamp 1688980957
transform 1 0 16468 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_37_190
timestamp 1688980957
transform 1 0 18584 0 -1 21760
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_37_198
timestamp 1688980957
transform 1 0 19320 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_26
timestamp 1688980957
transform 1 0 3496 0 1 21760
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_29
timestamp 1688980957
transform 1 0 3772 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_38_77
timestamp 1688980957
transform 1 0 8188 0 1 21760
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_83
timestamp 1688980957
transform 1 0 8740 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_85
timestamp 1688980957
transform 1 0 8924 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_102
timestamp 1688980957
transform 1 0 10488 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_38_118
timestamp 1688980957
transform 1 0 11960 0 1 21760
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_38_141
timestamp 1688980957
transform 1 0 14076 0 1 21760
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_153
timestamp 1688980957
transform 1 0 15180 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_191
timestamp 1688980957
transform 1 0 18676 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_38_197
timestamp 1688980957
transform 1 0 19228 0 1 21760
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_3
timestamp 1688980957
transform 1 0 1380 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_40
timestamp 1688980957
transform 1 0 4784 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_52
timestamp 1688980957
transform 1 0 5888 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_39_57
timestamp 1688980957
transform 1 0 6348 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_61
timestamp 1688980957
transform 1 0 6716 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_90
timestamp 1688980957
transform 1 0 9384 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_111
timestamp 1688980957
transform 1 0 11316 0 -1 22848
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_113
timestamp 1688980957
transform 1 0 11500 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_125
timestamp 1688980957
transform 1 0 12604 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_149
timestamp 1688980957
transform 1 0 14812 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_39_165
timestamp 1688980957
transform 1 0 16284 0 -1 22848
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_39_169
timestamp 1688980957
transform 1 0 16652 0 -1 22848
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_39_181
timestamp 1688980957
transform 1 0 17756 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_39_213
timestamp 1688980957
transform 1 0 20700 0 -1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_27
timestamp 1688980957
transform 1 0 3588 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_44
timestamp 1688980957
transform 1 0 5152 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_85
timestamp 1688980957
transform 1 0 8924 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_138
timestamp 1688980957
transform 1 0 13800 0 1 22848
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_40_141
timestamp 1688980957
transform 1 0 14076 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_40_150
timestamp 1688980957
transform 1 0 14904 0 1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_40_154
timestamp 1688980957
transform 1 0 15272 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_40_176
timestamp 1688980957
transform 1 0 17296 0 1 22848
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_184
timestamp 1688980957
transform 1 0 18032 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_40_190
timestamp 1688980957
transform 1 0 18584 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40_215
timestamp 1688980957
transform 1 0 20884 0 1 22848
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_28
timestamp 1688980957
transform 1 0 3680 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_40
timestamp 1688980957
transform 1 0 4784 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_57
timestamp 1688980957
transform 1 0 6348 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_61
timestamp 1688980957
transform 1 0 6716 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_65
timestamp 1688980957
transform 1 0 7084 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41_71
timestamp 1688980957
transform 1 0 7636 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_41_93
timestamp 1688980957
transform 1 0 9660 0 -1 23936
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_41_113
timestamp 1688980957
transform 1 0 11500 0 -1 23936
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_125
timestamp 1688980957
transform 1 0 12604 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_41_164
timestamp 1688980957
transform 1 0 16192 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_41_184
timestamp 1688980957
transform 1 0 18032 0 -1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_41_192
timestamp 1688980957
transform 1 0 18768 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_21
timestamp 1688980957
transform 1 0 3036 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_27
timestamp 1688980957
transform 1 0 3588 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_29
timestamp 1688980957
transform 1 0 3772 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_37
timestamp 1688980957
transform 1 0 4508 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_60
timestamp 1688980957
transform 1 0 6624 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_81
timestamp 1688980957
transform 1 0 8556 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_42_85
timestamp 1688980957
transform 1 0 8924 0 1 23936
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_93
timestamp 1688980957
transform 1 0 9660 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_42_116
timestamp 1688980957
transform 1 0 11776 0 1 23936
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_42_122
timestamp 1688980957
transform 1 0 12328 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_138
timestamp 1688980957
transform 1 0 13800 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_42_151
timestamp 1688980957
transform 1 0 14996 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_42_176
timestamp 1688980957
transform 1 0 17296 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_194
timestamp 1688980957
transform 1 0 18952 0 1 23936
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_42_217
timestamp 1688980957
transform 1 0 21068 0 1 23936
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_24
timestamp 1688980957
transform 1 0 3312 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_51
timestamp 1688980957
transform 1 0 5796 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_55
timestamp 1688980957
transform 1 0 6164 0 -1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_43_57
timestamp 1688980957
transform 1 0 6348 0 -1 25024
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_69
timestamp 1688980957
transform 1 0 7452 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_43_107
timestamp 1688980957
transform 1 0 10948 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_111
timestamp 1688980957
transform 1 0 11316 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_43_128
timestamp 1688980957
transform 1 0 12880 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_149
timestamp 1688980957
transform 1 0 14812 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_166
timestamp 1688980957
transform 1 0 16376 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_43_169
timestamp 1688980957
transform 1 0 16652 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_43_175
timestamp 1688980957
transform 1 0 17204 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_43_199
timestamp 1688980957
transform 1 0 19412 0 -1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_32
timestamp 1688980957
transform 1 0 4048 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_71
timestamp 1688980957
transform 1 0 7636 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_44_78
timestamp 1688980957
transform 1 0 8280 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_0_44_106
timestamp 1688980957
transform 1 0 10856 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_110
timestamp 1688980957
transform 1 0 11224 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_129
timestamp 1688980957
transform 1 0 12972 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_137
timestamp 1688980957
transform 1 0 13708 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_44_144
timestamp 1688980957
transform 1 0 14352 0 1 25024
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_44_185
timestamp 1688980957
transform 1 0 18124 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_194
timestamp 1688980957
transform 1 0 18952 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_44_197
timestamp 1688980957
transform 1 0 19228 0 1 25024
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_209
timestamp 1688980957
transform 1 0 20332 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_44_216
timestamp 1688980957
transform 1 0 20976 0 1 25024
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_39
timestamp 1688980957
transform 1 0 4692 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_51
timestamp 1688980957
transform 1 0 5796 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_55
timestamp 1688980957
transform 1 0 6164 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_45_108
timestamp 1688980957
transform 1 0 11040 0 -1 26112
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_143
timestamp 1688980957
transform 1 0 14260 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_155
timestamp 1688980957
transform 1 0 15364 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_163
timestamp 1688980957
transform 1 0 16100 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_167
timestamp 1688980957
transform 1 0 16468 0 -1 26112
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_45_169
timestamp 1688980957
transform 1 0 16652 0 -1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_45_212
timestamp 1688980957
transform 1 0 20608 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_27
timestamp 1688980957
transform 1 0 3588 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_44
timestamp 1688980957
transform 1 0 5152 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_67
timestamp 1688980957
transform 1 0 7268 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_92
timestamp 1688980957
transform 1 0 9568 0 1 26112
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_46_127
timestamp 1688980957
transform 1 0 12788 0 1 26112
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_139
timestamp 1688980957
transform 1 0 13892 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_180
timestamp 1688980957
transform 1 0 17664 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_46_186
timestamp 1688980957
transform 1 0 18216 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_46_190
timestamp 1688980957
transform 1 0 18584 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_46_203
timestamp 1688980957
transform 1 0 19780 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_46_212
timestamp 1688980957
transform 1 0 20608 0 1 26112
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_47_37
timestamp 1688980957
transform 1 0 4508 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_96
timestamp 1688980957
transform 1 0 9936 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_47_131
timestamp 1688980957
transform 1 0 13156 0 -1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_47_167
timestamp 1688980957
transform 1 0 16468 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_47_187
timestamp 1688980957
transform 1 0 18308 0 -1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_47_195
timestamp 1688980957
transform 1 0 19044 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_3
timestamp 1688980957
transform 1 0 1380 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_26
timestamp 1688980957
transform 1 0 3496 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_32
timestamp 1688980957
transform 1 0 4048 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_64
timestamp 1688980957
transform 1 0 6992 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_85
timestamp 1688980957
transform 1 0 8924 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_48_93
timestamp 1688980957
transform 1 0 9660 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_48_129
timestamp 1688980957
transform 1 0 12972 0 1 27200
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_48_137
timestamp 1688980957
transform 1 0 13708 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_48_156
timestamp 1688980957
transform 1 0 15456 0 1 27200
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_48_183
timestamp 1688980957
transform 1 0 17940 0 1 27200
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_48_195
timestamp 1688980957
transform 1 0 19044 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_213
timestamp 1688980957
transform 1 0 20700 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_48_221
timestamp 1688980957
transform 1 0 21436 0 1 27200
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_10
timestamp 1688980957
transform 1 0 2024 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_47
timestamp 1688980957
transform 1 0 5428 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_55
timestamp 1688980957
transform 1 0 6164 0 -1 28288
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_49_57
timestamp 1688980957
transform 1 0 6348 0 -1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_69
timestamp 1688980957
transform 1 0 7452 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_101
timestamp 1688980957
transform 1 0 10396 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49_109
timestamp 1688980957
transform 1 0 11132 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_113
timestamp 1688980957
transform 1 0 11500 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_129
timestamp 1688980957
transform 1 0 12972 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_49_137
timestamp 1688980957
transform 1 0 13708 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_49_155
timestamp 1688980957
transform 1 0 15364 0 -1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_163
timestamp 1688980957
transform 1 0 16100 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_167
timestamp 1688980957
transform 1 0 16468 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_49_169
timestamp 1688980957
transform 1 0 16652 0 -1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_49_208
timestamp 1688980957
transform 1 0 20240 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_10
timestamp 1688980957
transform 1 0 2024 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_27
timestamp 1688980957
transform 1 0 3588 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_29
timestamp 1688980957
transform 1 0 3772 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_50_55
timestamp 1688980957
transform 1 0 6164 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_50_63
timestamp 1688980957
transform 1 0 6900 0 1 28288
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_80
timestamp 1688980957
transform 1 0 8464 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_50_85
timestamp 1688980957
transform 1 0 8924 0 1 28288
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_50_108
timestamp 1688980957
transform 1 0 11040 0 1 28288
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_50_127
timestamp 1688980957
transform 1 0 12788 0 1 28288
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_50_139
timestamp 1688980957
transform 1 0 13892 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_3
timestamp 1688980957
transform 1 0 1380 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_51_38
timestamp 1688980957
transform 1 0 4600 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_51_57
timestamp 1688980957
transform 1 0 6348 0 -1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_51_65
timestamp 1688980957
transform 1 0 7084 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_107
timestamp 1688980957
transform 1 0 10948 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_111
timestamp 1688980957
transform 1 0 11316 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_51_128
timestamp 1688980957
transform 1 0 12880 0 -1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_185
timestamp 1688980957
transform 1 0 18124 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_51_202
timestamp 1688980957
transform 1 0 19688 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_51_208
timestamp 1688980957
transform 1 0 20240 0 -1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_51_216
timestamp 1688980957
transform 1 0 20976 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_7
timestamp 1688980957
transform 1 0 1748 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_26
timestamp 1688980957
transform 1 0 3496 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52_29
timestamp 1688980957
transform 1 0 3772 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_33
timestamp 1688980957
transform 1 0 4140 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_62
timestamp 1688980957
transform 1 0 6808 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_68
timestamp 1688980957
transform 1 0 7360 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_52_85
timestamp 1688980957
transform 1 0 8924 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_93
timestamp 1688980957
transform 1 0 9660 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_52_130
timestamp 1688980957
transform 1 0 13064 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_138
timestamp 1688980957
transform 1 0 13800 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_52_165
timestamp 1688980957
transform 1 0 16284 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_52_178
timestamp 1688980957
transform 1 0 17480 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_52_182
timestamp 1688980957
transform 1 0 17848 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_52_186
timestamp 1688980957
transform 1 0 18216 0 1 29376
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_52_194
timestamp 1688980957
transform 1 0 18952 0 1 29376
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_52_197
timestamp 1688980957
transform 1 0 19228 0 1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_53_39
timestamp 1688980957
transform 1 0 4692 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_53_72
timestamp 1688980957
transform 1 0 7728 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_80
timestamp 1688980957
transform 1 0 8464 0 -1 30464
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_53_96
timestamp 1688980957
transform 1 0 9936 0 -1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_53_108
timestamp 1688980957
transform 1 0 11040 0 -1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_53_164
timestamp 1688980957
transform 1 0 16192 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_53_184
timestamp 1688980957
transform 1 0 18032 0 -1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_53_192
timestamp 1688980957
transform 1 0 18768 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_53_215
timestamp 1688980957
transform 1 0 20884 0 -1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_50
timestamp 1688980957
transform 1 0 5704 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_54_70
timestamp 1688980957
transform 1 0 7544 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_54_81
timestamp 1688980957
transform 1 0 8556 0 1 30464
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_85
timestamp 1688980957
transform 1 0 8924 0 1 30464
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_54_97
timestamp 1688980957
transform 1 0 10028 0 1 30464
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_54_109
timestamp 1688980957
transform 1 0 11132 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_119
timestamp 1688980957
transform 1 0 12052 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_54_129
timestamp 1688980957
transform 1 0 12972 0 1 30464
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_54_137
timestamp 1688980957
transform 1 0 13708 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_54_156
timestamp 1688980957
transform 1 0 15456 0 1 30464
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_180
timestamp 1688980957
transform 1 0 17664 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_184
timestamp 1688980957
transform 1 0 18032 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_54_192
timestamp 1688980957
transform 1 0 18768 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_54_213
timestamp 1688980957
transform 1 0 20700 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_18
timestamp 1688980957
transform 1 0 2760 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_40
timestamp 1688980957
transform 1 0 4784 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_60
timestamp 1688980957
transform 1 0 6624 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_66
timestamp 1688980957
transform 1 0 7176 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_55_88
timestamp 1688980957
transform 1 0 9200 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_0_55_109
timestamp 1688980957
transform 1 0 11132 0 -1 31552
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_55_131
timestamp 1688980957
transform 1 0 13156 0 -1 31552
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_55_143
timestamp 1688980957
transform 1 0 14260 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_55_160
timestamp 1688980957
transform 1 0 15824 0 -1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_55_200
timestamp 1688980957
transform 1 0 19504 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_55_207
timestamp 1688980957
transform 1 0 20148 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_55_212
timestamp 1688980957
transform 1 0 20608 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_55_217
timestamp 1688980957
transform 1 0 21068 0 -1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_6
timestamp 1688980957
transform 1 0 1656 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_56_35
timestamp 1688980957
transform 1 0 4324 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_56_40
timestamp 1688980957
transform 1 0 4784 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_63
timestamp 1688980957
transform 1 0 6900 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_56_85
timestamp 1688980957
transform 1 0 8924 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_93
timestamp 1688980957
transform 1 0 9660 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_56_115
timestamp 1688980957
transform 1 0 11684 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_121
timestamp 1688980957
transform 1 0 12236 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_56_177
timestamp 1688980957
transform 1 0 17388 0 1 31552
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_56_194
timestamp 1688980957
transform 1 0 18952 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_200
timestamp 1688980957
transform 1 0 19504 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_204
timestamp 1688980957
transform 1 0 19872 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_56_211
timestamp 1688980957
transform 1 0 20516 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_56_215
timestamp 1688980957
transform 1 0 20884 0 1 31552
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57_3
timestamp 1688980957
transform 1 0 1380 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57_26
timestamp 1688980957
transform 1 0 3496 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_57_49
timestamp 1688980957
transform 1 0 5612 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_55
timestamp 1688980957
transform 1 0 6164 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_57_60
timestamp 1688980957
transform 1 0 6624 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  FILLER_0_57_82
timestamp 1688980957
transform 1 0 8648 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57_103
timestamp 1688980957
transform 1 0 10580 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_111
timestamp 1688980957
transform 1 0 11316 0 -1 32640
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_57_113
timestamp 1688980957
transform 1 0 11500 0 -1 32640
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_155
timestamp 1688980957
transform 1 0 15364 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_57_159
timestamp 1688980957
transform 1 0 15732 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_167
timestamp 1688980957
transform 1 0 16468 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_57_169
timestamp 1688980957
transform 1 0 16652 0 -1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_57_186
timestamp 1688980957
transform 1 0 18216 0 -1 32640
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_57_200
timestamp 1688980957
transform 1 0 19504 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_58_7
timestamp 1688980957
transform 1 0 1748 0 1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_44
timestamp 1688980957
transform 1 0 5152 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_85
timestamp 1688980957
transform 1 0 8924 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58_119
timestamp 1688980957
transform 1 0 12052 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_58_123
timestamp 1688980957
transform 1 0 12420 0 1 32640
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_58_141
timestamp 1688980957
transform 1 0 14076 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_58_145
timestamp 1688980957
transform 1 0 14444 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_59_15
timestamp 1688980957
transform 1 0 2484 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_59_35
timestamp 1688980957
transform 1 0 4324 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_59_53
timestamp 1688980957
transform 1 0 5980 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_59_57
timestamp 1688980957
transform 1 0 6348 0 -1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_65
timestamp 1688980957
transform 1 0 7084 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_59_81
timestamp 1688980957
transform 1 0 8556 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_85
timestamp 1688980957
transform 1 0 8924 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_59_101
timestamp 1688980957
transform 1 0 10396 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_59_107
timestamp 1688980957
transform 1 0 10948 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_111
timestamp 1688980957
transform 1 0 11316 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_128
timestamp 1688980957
transform 1 0 12880 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_59_162
timestamp 1688980957
transform 1 0 16008 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_172
timestamp 1688980957
transform 1 0 16928 0 -1 33728
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_59_179
timestamp 1688980957
transform 1 0 17572 0 -1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_59_191
timestamp 1688980957
transform 1 0 18676 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_195
timestamp 1688980957
transform 1 0 19044 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_59_199
timestamp 1688980957
transform 1 0 19412 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_59_208
timestamp 1688980957
transform 1 0 20240 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_59_221
timestamp 1688980957
transform 1 0 21436 0 -1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_60_3
timestamp 1688980957
transform 1 0 1380 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_60_26
timestamp 1688980957
transform 1 0 3496 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_60_35
timestamp 1688980957
transform 1 0 4324 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_60_76
timestamp 1688980957
transform 1 0 8096 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_60_85
timestamp 1688980957
transform 1 0 8924 0 1 33728
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_60_119
timestamp 1688980957
transform 1 0 12052 0 1 33728
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_60_131
timestamp 1688980957
transform 1 0 13156 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_139
timestamp 1688980957
transform 1 0 13892 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_60_141
timestamp 1688980957
transform 1 0 14076 0 1 33728
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_149
timestamp 1688980957
transform 1 0 14812 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_181
timestamp 1688980957
transform 1 0 17756 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_195
timestamp 1688980957
transform 1 0 19044 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_60_200
timestamp 1688980957
transform 1 0 19504 0 1 33728
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_208
timestamp 1688980957
transform 1 0 20240 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_60_215
timestamp 1688980957
transform 1 0 20884 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_61_3
timestamp 1688980957
transform 1 0 1380 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_7
timestamp 1688980957
transform 1 0 1748 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_61_60
timestamp 1688980957
transform 1 0 6624 0 -1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_61_68
timestamp 1688980957
transform 1 0 7360 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_61_108
timestamp 1688980957
transform 1 0 11040 0 -1 34816
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_61_113
timestamp 1688980957
transform 1 0 11500 0 -1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_61_125
timestamp 1688980957
transform 1 0 12604 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_61_159
timestamp 1688980957
transform 1 0 15732 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_164
timestamp 1688980957
transform 1 0 16192 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_61_169
timestamp 1688980957
transform 1 0 16652 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_61_173
timestamp 1688980957
transform 1 0 17020 0 -1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_61_190
timestamp 1688980957
transform 1 0 18584 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_61_196
timestamp 1688980957
transform 1 0 19136 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_9
timestamp 1688980957
transform 1 0 1932 0 1 34816
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_62_71
timestamp 1688980957
transform 1 0 7636 0 1 34816
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_83
timestamp 1688980957
transform 1 0 8740 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_62_103
timestamp 1688980957
transform 1 0 10580 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_62_111
timestamp 1688980957
transform 1 0 11316 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_62_135
timestamp 1688980957
transform 1 0 13524 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_62_139
timestamp 1688980957
transform 1 0 13892 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_62_141
timestamp 1688980957
transform 1 0 14076 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_62_183
timestamp 1688980957
transform 1 0 17940 0 1 34816
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_62_191
timestamp 1688980957
transform 1 0 18676 0 1 34816
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_3
timestamp 1688980957
transform 1 0 1380 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_40
timestamp 1688980957
transform 1 0 4784 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_63
timestamp 1688980957
transform 1 0 6900 0 -1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_100
timestamp 1688980957
transform 1 0 10304 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_63_113
timestamp 1688980957
transform 1 0 11500 0 -1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_134
timestamp 1688980957
transform 1 0 13432 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_63_146
timestamp 1688980957
transform 1 0 14536 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_0_63_157
timestamp 1688980957
transform 1 0 15548 0 -1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_63_165
timestamp 1688980957
transform 1 0 16284 0 -1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_63_176
timestamp 1688980957
transform 1 0 17296 0 -1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_63_210
timestamp 1688980957
transform 1 0 20424 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_63_217
timestamp 1688980957
transform 1 0 21068 0 -1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_9
timestamp 1688980957
transform 1 0 1932 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_27
timestamp 1688980957
transform 1 0 3588 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_64_29
timestamp 1688980957
transform 1 0 3772 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_64_34
timestamp 1688980957
transform 1 0 4232 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_42
timestamp 1688980957
transform 1 0 4968 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_64_47
timestamp 1688980957
transform 1 0 5428 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_64_67
timestamp 1688980957
transform 1 0 7268 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_100
timestamp 1688980957
transform 1 0 10304 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_64_105
timestamp 1688980957
transform 1 0 10764 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_109
timestamp 1688980957
transform 1 0 11132 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_125
timestamp 1688980957
transform 1 0 12604 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_64_137
timestamp 1688980957
transform 1 0 13708 0 1 35904
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_64_144
timestamp 1688980957
transform 1 0 14352 0 1 35904
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_64_156
timestamp 1688980957
transform 1 0 15456 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_160
timestamp 1688980957
transform 1 0 15824 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_64_164
timestamp 1688980957
transform 1 0 16192 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_64_186
timestamp 1688980957
transform 1 0 18216 0 1 35904
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_64_194
timestamp 1688980957
transform 1 0 18952 0 1 35904
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_209
timestamp 1688980957
transform 1 0 20332 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_64_213
timestamp 1688980957
transform 1 0 20700 0 1 35904
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_65_3
timestamp 1688980957
transform 1 0 1380 0 -1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_65_15
timestamp 1688980957
transform 1 0 2484 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_65_47
timestamp 1688980957
transform 1 0 5428 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_65_51
timestamp 1688980957
transform 1 0 5796 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_65_63
timestamp 1688980957
transform 1 0 6900 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_65_117
timestamp 1688980957
transform 1 0 11868 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_65_125
timestamp 1688980957
transform 1 0 12604 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_65_152
timestamp 1688980957
transform 1 0 15088 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_163
timestamp 1688980957
transform 1 0 16100 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_167
timestamp 1688980957
transform 1 0 16468 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_65_192
timestamp 1688980957
transform 1 0 18768 0 -1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_65_202
timestamp 1688980957
transform 1 0 19688 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_65_207
timestamp 1688980957
transform 1 0 20148 0 -1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_65_218
timestamp 1688980957
transform 1 0 21160 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_3
timestamp 1688980957
transform 1 0 1380 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_66_19
timestamp 1688980957
transform 1 0 2852 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_27
timestamp 1688980957
transform 1 0 3588 0 1 36992
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_66_71
timestamp 1688980957
transform 1 0 7636 0 1 36992
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_83
timestamp 1688980957
transform 1 0 8740 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_66_85
timestamp 1688980957
transform 1 0 8924 0 1 36992
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_66_95
timestamp 1688980957
transform 1 0 9844 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_66_119
timestamp 1688980957
transform 1 0 12052 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_0_66_137
timestamp 1688980957
transform 1 0 13708 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_66_141
timestamp 1688980957
transform 1 0 14076 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66_168
timestamp 1688980957
transform 1 0 16560 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_174
timestamp 1688980957
transform 1 0 17112 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_66_178
timestamp 1688980957
transform 1 0 17480 0 1 36992
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_66_186
timestamp 1688980957
transform 1 0 18216 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_195
timestamp 1688980957
transform 1 0 19044 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_66_197
timestamp 1688980957
transform 1 0 19228 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_66_201
timestamp 1688980957
transform 1 0 19596 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_67_30
timestamp 1688980957
transform 1 0 3864 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_34
timestamp 1688980957
transform 1 0 4232 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_57
timestamp 1688980957
transform 1 0 6348 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_67_61
timestamp 1688980957
transform 1 0 6716 0 -1 38080
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_81
timestamp 1688980957
transform 1 0 8556 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_67_108
timestamp 1688980957
transform 1 0 11040 0 -1 38080
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_113
timestamp 1688980957
transform 1 0 11500 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_67_125
timestamp 1688980957
transform 1 0 12604 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_67_144
timestamp 1688980957
transform 1 0 14352 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_67_161
timestamp 1688980957
transform 1 0 15916 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_167
timestamp 1688980957
transform 1 0 16468 0 -1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_67_169
timestamp 1688980957
transform 1 0 16652 0 -1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_67_181
timestamp 1688980957
transform 1 0 17756 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_189
timestamp 1688980957
transform 1 0 18492 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_67_193
timestamp 1688980957
transform 1 0 18860 0 -1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_67_201
timestamp 1688980957
transform 1 0 19596 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_67_207
timestamp 1688980957
transform 1 0 20148 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_67_217
timestamp 1688980957
transform 1 0 21068 0 -1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_68_3
timestamp 1688980957
transform 1 0 1380 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_21
timestamp 1688980957
transform 1 0 3036 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_29
timestamp 1688980957
transform 1 0 3772 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_45
timestamp 1688980957
transform 1 0 5244 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_68_76
timestamp 1688980957
transform 1 0 8096 0 1 38080
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_85
timestamp 1688980957
transform 1 0 8924 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_97
timestamp 1688980957
transform 1 0 10028 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_109
timestamp 1688980957
transform 1 0 11132 0 1 38080
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_121
timestamp 1688980957
transform 1 0 12236 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_68_133
timestamp 1688980957
transform 1 0 13340 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_139
timestamp 1688980957
transform 1 0 13892 0 1 38080
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_68_141
timestamp 1688980957
transform 1 0 14076 0 1 38080
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_68_153
timestamp 1688980957
transform 1 0 15180 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_68_161
timestamp 1688980957
transform 1 0 15916 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_68_166
timestamp 1688980957
transform 1 0 16376 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_68_174
timestamp 1688980957
transform 1 0 17112 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_68_179
timestamp 1688980957
transform 1 0 17572 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_0_68_185
timestamp 1688980957
transform 1 0 18124 0 1 38080
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_68_193
timestamp 1688980957
transform 1 0 18860 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_0_68_197
timestamp 1688980957
transform 1 0 19228 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_68_201
timestamp 1688980957
transform 1 0 19596 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_68_217
timestamp 1688980957
transform 1 0 21068 0 1 38080
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_69_24
timestamp 1688980957
transform 1 0 3312 0 -1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_28
timestamp 1688980957
transform 1 0 3680 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_69_44
timestamp 1688980957
transform 1 0 5152 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_52
timestamp 1688980957
transform 1 0 5888 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_72
timestamp 1688980957
transform 1 0 7728 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_84
timestamp 1688980957
transform 1 0 8832 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_96
timestamp 1688980957
transform 1 0 9936 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_69_108
timestamp 1688980957
transform 1 0 11040 0 -1 39168
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_113
timestamp 1688980957
transform 1 0 11500 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_125
timestamp 1688980957
transform 1 0 12604 0 -1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_137
timestamp 1688980957
transform 1 0 13708 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_69_149
timestamp 1688980957
transform 1 0 14812 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_157
timestamp 1688980957
transform 1 0 15548 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_69_161
timestamp 1688980957
transform 1 0 15916 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_167
timestamp 1688980957
transform 1 0 16468 0 -1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_69_169
timestamp 1688980957
transform 1 0 16652 0 -1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_69_181
timestamp 1688980957
transform 1 0 17756 0 -1 39168
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_69_189
timestamp 1688980957
transform 1 0 18492 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_69_195
timestamp 1688980957
transform 1 0 19044 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_201
timestamp 1688980957
transform 1 0 19596 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_69_205
timestamp 1688980957
transform 1 0 19964 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_69_209
timestamp 1688980957
transform 1 0 20332 0 -1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_3
timestamp 1688980957
transform 1 0 1380 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_70_25
timestamp 1688980957
transform 1 0 3404 0 1 39168
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_35
timestamp 1688980957
transform 1 0 4324 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_70_47
timestamp 1688980957
transform 1 0 5428 0 1 39168
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_58
timestamp 1688980957
transform 1 0 6440 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_70
timestamp 1688980957
transform 1 0 7544 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_70_82
timestamp 1688980957
transform 1 0 8648 0 1 39168
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_85
timestamp 1688980957
transform 1 0 8924 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_97
timestamp 1688980957
transform 1 0 10028 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_109
timestamp 1688980957
transform 1 0 11132 0 1 39168
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_121
timestamp 1688980957
transform 1 0 12236 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_70_133
timestamp 1688980957
transform 1 0 13340 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_139
timestamp 1688980957
transform 1 0 13892 0 1 39168
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_141
timestamp 1688980957
transform 1 0 14076 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_70_153
timestamp 1688980957
transform 1 0 15180 0 1 39168
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_70_164
timestamp 1688980957
transform 1 0 16192 0 1 39168
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_176
timestamp 1688980957
transform 1 0 17296 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_70_183
timestamp 1688980957
transform 1 0 17940 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_70_187
timestamp 1688980957
transform 1 0 18308 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_70_212
timestamp 1688980957
transform 1 0 20608 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_70_217
timestamp 1688980957
transform 1 0 21068 0 1 39168
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_71_3
timestamp 1688980957
transform 1 0 1380 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_71_19
timestamp 1688980957
transform 1 0 2852 0 -1 40256
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_27
timestamp 1688980957
transform 1 0 3588 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_39
timestamp 1688980957
transform 1 0 4692 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_71_51
timestamp 1688980957
transform 1 0 5796 0 -1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_55
timestamp 1688980957
transform 1 0 6164 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_57
timestamp 1688980957
transform 1 0 6348 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_69
timestamp 1688980957
transform 1 0 7452 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_81
timestamp 1688980957
transform 1 0 8556 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_93
timestamp 1688980957
transform 1 0 9660 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_71_105
timestamp 1688980957
transform 1 0 10764 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_111
timestamp 1688980957
transform 1 0 11316 0 -1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_113
timestamp 1688980957
transform 1 0 11500 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_125
timestamp 1688980957
transform 1 0 12604 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_137
timestamp 1688980957
transform 1 0 13708 0 -1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_71_149
timestamp 1688980957
transform 1 0 14812 0 -1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_71_161
timestamp 1688980957
transform 1 0 15916 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_71_166
timestamp 1688980957
transform 1 0 16376 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_71_169
timestamp 1688980957
transform 1 0 16652 0 -1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_177
timestamp 1688980957
transform 1 0 17388 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_71_202
timestamp 1688980957
transform 1 0 19688 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_71_206
timestamp 1688980957
transform 1 0 20056 0 -1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_72_21
timestamp 1688980957
transform 1 0 3036 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_27
timestamp 1688980957
transform 1 0 3588 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_29
timestamp 1688980957
transform 1 0 3772 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_72_41
timestamp 1688980957
transform 1 0 4876 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_0_72_50
timestamp 1688980957
transform 1 0 5704 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_72_58
timestamp 1688980957
transform 1 0 6440 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_72_63
timestamp 1688980957
transform 1 0 6900 0 1 40256
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_68
timestamp 1688980957
transform 1 0 7360 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_72_80
timestamp 1688980957
transform 1 0 8464 0 1 40256
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_85
timestamp 1688980957
transform 1 0 8924 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_97
timestamp 1688980957
transform 1 0 10028 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_109
timestamp 1688980957
transform 1 0 11132 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_121
timestamp 1688980957
transform 1 0 12236 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_72_133
timestamp 1688980957
transform 1 0 13340 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_72_139
timestamp 1688980957
transform 1 0 13892 0 1 40256
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_141
timestamp 1688980957
transform 1 0 14076 0 1 40256
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_72_153
timestamp 1688980957
transform 1 0 15180 0 1 40256
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_72_165
timestamp 1688980957
transform 1 0 16284 0 1 40256
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_72_173
timestamp 1688980957
transform 1 0 17020 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_72_197
timestamp 1688980957
transform 1 0 19228 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_72_217
timestamp 1688980957
transform 1 0 21068 0 1 40256
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_73_21
timestamp 1688980957
transform 1 0 3036 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_73_29
timestamp 1688980957
transform 1 0 3772 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_73_34
timestamp 1688980957
transform 1 0 4232 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_0_73_42
timestamp 1688980957
transform 1 0 4968 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_73_60
timestamp 1688980957
transform 1 0 6624 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_73_70
timestamp 1688980957
transform 1 0 7544 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_73_74
timestamp 1688980957
transform 1 0 7912 0 -1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_82
timestamp 1688980957
transform 1 0 8648 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_94
timestamp 1688980957
transform 1 0 9752 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_73_106
timestamp 1688980957
transform 1 0 10856 0 -1 41344
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_113
timestamp 1688980957
transform 1 0 11500 0 -1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_73_125
timestamp 1688980957
transform 1 0 12604 0 -1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_73_137
timestamp 1688980957
transform 1 0 13708 0 -1 41344
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_73_145
timestamp 1688980957
transform 1 0 14444 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_73_159
timestamp 1688980957
transform 1 0 15732 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_164
timestamp 1688980957
transform 1 0 16192 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_73_178
timestamp 1688980957
transform 1 0 17480 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_73_189
timestamp 1688980957
transform 1 0 18492 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_73_217
timestamp 1688980957
transform 1 0 21068 0 -1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_74_15
timestamp 1688980957
transform 1 0 2484 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_21
timestamp 1688980957
transform 1 0 3036 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_74_56
timestamp 1688980957
transform 1 0 6256 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_74_60
timestamp 1688980957
transform 1 0 6624 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_65
timestamp 1688980957
transform 1 0 7084 0 1 41344
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_97
timestamp 1688980957
transform 1 0 10028 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_109
timestamp 1688980957
transform 1 0 11132 0 1 41344
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_74_121
timestamp 1688980957
transform 1 0 12236 0 1 41344
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_74_133
timestamp 1688980957
transform 1 0 13340 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_139
timestamp 1688980957
transform 1 0 13892 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_74_141
timestamp 1688980957
transform 1 0 14076 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_74_194
timestamp 1688980957
transform 1 0 18952 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_74_200
timestamp 1688980957
transform 1 0 19504 0 1 41344
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_74_204
timestamp 1688980957
transform 1 0 19872 0 1 41344
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_3
timestamp 1688980957
transform 1 0 1380 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_28
timestamp 1688980957
transform 1 0 3680 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_75_45
timestamp 1688980957
transform 1 0 5244 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_75_61
timestamp 1688980957
transform 1 0 6716 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_75_73
timestamp 1688980957
transform 1 0 7820 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_75_79
timestamp 1688980957
transform 1 0 8372 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_75_83
timestamp 1688980957
transform 1 0 8740 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_75_94
timestamp 1688980957
transform 1 0 9752 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_75_98
timestamp 1688980957
transform 1 0 10120 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_75_106
timestamp 1688980957
transform 1 0 10856 0 -1 42432
box -38 -48 590 592
use sky130_ef_sc_hd__decap_12  FILLER_0_75_113
timestamp 1688980957
transform 1 0 11500 0 -1 42432
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_75_125
timestamp 1688980957
transform 1 0 12604 0 -1 42432
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_75_133
timestamp 1688980957
transform 1 0 13340 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_75_139
timestamp 1688980957
transform 1 0 13892 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_75_167
timestamp 1688980957
transform 1 0 16468 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_75_179
timestamp 1688980957
transform 1 0 17572 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_75_197
timestamp 1688980957
transform 1 0 19228 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_75_221
timestamp 1688980957
transform 1 0 21436 0 -1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_76_3
timestamp 1688980957
transform 1 0 1380 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_29
timestamp 1688980957
transform 1 0 3772 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_88
timestamp 1688980957
transform 1 0 9200 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_99
timestamp 1688980957
transform 1 0 10212 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_112
timestamp 1688980957
transform 1 0 11408 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_116
timestamp 1688980957
transform 1 0 11776 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_76_123
timestamp 1688980957
transform 1 0 12420 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_134
timestamp 1688980957
transform 1 0 13432 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_139
timestamp 1688980957
transform 1 0 13892 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_151
timestamp 1688980957
transform 1 0 14996 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_76_172
timestamp 1688980957
transform 1 0 16928 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_76_194
timestamp 1688980957
transform 1 0 18952 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_76_221
timestamp 1688980957
transform 1 0 21436 0 1 42432
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_0_77_3
timestamp 1688980957
transform 1 0 1380 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_0_77_26
timestamp 1688980957
transform 1 0 3496 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_55
timestamp 1688980957
transform 1 0 6164 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_57
timestamp 1688980957
transform 1 0 6348 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_77_103
timestamp 1688980957
transform 1 0 10580 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_77_113
timestamp 1688980957
transform 1 0 11500 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_77_125
timestamp 1688980957
transform 1 0 12604 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  FILLER_0_77_131
timestamp 1688980957
transform 1 0 13156 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_167
timestamp 1688980957
transform 1 0 16468 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_77_195
timestamp 1688980957
transform 1 0 19044 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_77_221
timestamp 1688980957
transform 1 0 21436 0 -1 43520
box -38 -48 222 592
use sky130_fd_sc_hd__clkbuf_2  input1 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1472 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input2
timestamp 1688980957
transform 1 0 1748 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input3
timestamp 1688980957
transform 1 0 1932 0 -1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input4 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1380 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input5
timestamp 1688980957
transform 1 0 1380 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input6
timestamp 1688980957
transform 1 0 2852 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input7
timestamp 1688980957
transform 1 0 2576 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input8 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 1380 0 1 21760
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input9
timestamp 1688980957
transform 1 0 2300 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input10
timestamp 1688980957
transform 1 0 3312 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input11
timestamp 1688980957
transform 1 0 3036 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input12
timestamp 1688980957
transform 1 0 2760 0 -1 23936
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input13
timestamp 1688980957
transform 1 0 2852 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input14
timestamp 1688980957
transform 1 0 3772 0 1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input15
timestamp 1688980957
transform 1 0 3772 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input16
timestamp 1688980957
transform 1 0 1380 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input17
timestamp 1688980957
transform 1 0 1380 0 1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input18
timestamp 1688980957
transform 1 0 3220 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input19
timestamp 1688980957
transform 1 0 3772 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input20
timestamp 1688980957
transform 1 0 1380 0 1 20672
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input21
timestamp 1688980957
transform 1 0 1380 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input22
timestamp 1688980957
transform 1 0 1380 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input23
timestamp 1688980957
transform 1 0 6348 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input24
timestamp 1688980957
transform 1 0 2944 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input25
timestamp 1688980957
transform 1 0 1380 0 -1 27200
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input26
timestamp 1688980957
transform 1 0 5244 0 1 28288
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input27
timestamp 1688980957
transform 1 0 1380 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input28
timestamp 1688980957
transform 1 0 3036 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input29
timestamp 1688980957
transform 1 0 4232 0 1 29376
box -38 -48 958 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input30
timestamp 1688980957
transform 1 0 2760 0 1 30464
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input31
timestamp 1688980957
transform 1 0 1380 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input32
timestamp 1688980957
transform 1 0 1380 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input33
timestamp 1688980957
transform 1 0 1380 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input34
timestamp 1688980957
transform 1 0 1748 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input35
timestamp 1688980957
transform 1 0 1748 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input36
timestamp 1688980957
transform 1 0 2944 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input37
timestamp 1688980957
transform 1 0 3220 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input38
timestamp 1688980957
transform 1 0 3772 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input39
timestamp 1688980957
transform 1 0 1380 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input40
timestamp 1688980957
transform 1 0 1380 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input41
timestamp 1688980957
transform 1 0 1380 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input42
timestamp 1688980957
transform 1 0 1380 0 1 25024
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  input43
timestamp 1688980957
transform 1 0 3772 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input44
timestamp 1688980957
transform 1 0 1380 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input45
timestamp 1688980957
transform 1 0 2300 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input46
timestamp 1688980957
transform 1 0 2760 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input47
timestamp 1688980957
transform 1 0 3036 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input48
timestamp 1688980957
transform 1 0 3312 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__buf_4  input49 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 4232 0 -1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input50 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3680 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input51
timestamp 1688980957
transform 1 0 4324 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input52
timestamp 1688980957
transform 1 0 4232 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input53
timestamp 1688980957
transform 1 0 1380 0 -1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input54
timestamp 1688980957
transform 1 0 1380 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input55
timestamp 1688980957
transform 1 0 3036 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input56
timestamp 1688980957
transform 1 0 6348 0 -1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input57
timestamp 1688980957
transform 1 0 1380 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input58
timestamp 1688980957
transform 1 0 1748 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input59
timestamp 1688980957
transform 1 0 2852 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input60
timestamp 1688980957
transform 1 0 3772 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input61
timestamp 1688980957
transform 1 0 6348 0 -1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input62
timestamp 1688980957
transform 1 0 1380 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input63
timestamp 1688980957
transform 1 0 1932 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input64
timestamp 1688980957
transform 1 0 2300 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input65
timestamp 1688980957
transform 1 0 3128 0 1 38080
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input66
timestamp 1688980957
transform 1 0 1380 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input67
timestamp 1688980957
transform 1 0 1932 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input68
timestamp 1688980957
transform 1 0 2484 0 1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input69
timestamp 1688980957
transform 1 0 3036 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input70
timestamp 1688980957
transform 1 0 3772 0 1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input71
timestamp 1688980957
transform 1 0 1380 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input72
timestamp 1688980957
transform 1 0 1932 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input73
timestamp 1688980957
transform 1 0 2484 0 -1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input74
timestamp 1688980957
transform 1 0 2944 0 -1 32640
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input75
timestamp 1688980957
transform 1 0 1932 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input76
timestamp 1688980957
transform 1 0 1380 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input77
timestamp 1688980957
transform 1 0 2944 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input78
timestamp 1688980957
transform 1 0 3772 0 1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__buf_4  input79
timestamp 1688980957
transform 1 0 1380 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  input80
timestamp 1688980957
transform 1 0 3772 0 1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__buf_8  input81 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 19228 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  input82
timestamp 1688980957
transform 1 0 18308 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input83
timestamp 1688980957
transform 1 0 14352 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input84
timestamp 1688980957
transform 1 0 13800 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input85
timestamp 1688980957
transform 1 0 16284 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input86
timestamp 1688980957
transform 1 0 16008 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input87
timestamp 1688980957
transform 1 0 15732 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input88
timestamp 1688980957
transform 1 0 16836 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input89
timestamp 1688980957
transform 1 0 13708 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input90
timestamp 1688980957
transform 1 0 21344 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input91
timestamp 1688980957
transform 1 0 21344 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_8  input92
timestamp 1688980957
transform 1 0 16652 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_16  input93 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 17296 0 1 1088
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_16  input94
timestamp 1688980957
transform 1 0 17756 0 -1 2176
box -38 -48 1878 592
use sky130_fd_sc_hd__buf_8  input95
timestamp 1688980957
transform 1 0 17204 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  input96
timestamp 1688980957
transform 1 0 15456 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  input97
timestamp 1688980957
transform 1 0 19228 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  input98
timestamp 1688980957
transform 1 0 20332 0 1 1088
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  input99
timestamp 1688980957
transform 1 0 19596 0 -1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_8  input100
timestamp 1688980957
transform 1 0 20332 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  input101
timestamp 1688980957
transform 1 0 2208 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input102
timestamp 1688980957
transform 1 0 3220 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input103
timestamp 1688980957
transform 1 0 2576 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input104
timestamp 1688980957
transform 1 0 3588 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input105
timestamp 1688980957
transform 1 0 5244 0 -1 2176
box -38 -48 958 592
use sky130_fd_sc_hd__buf_2  input106
timestamp 1688980957
transform 1 0 5152 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input107
timestamp 1688980957
transform 1 0 5428 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input108
timestamp 1688980957
transform 1 0 4416 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input109
timestamp 1688980957
transform 1 0 5980 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input110
timestamp 1688980957
transform 1 0 6348 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input111
timestamp 1688980957
transform 1 0 4784 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input112
timestamp 1688980957
transform 1 0 6532 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input113
timestamp 1688980957
transform 1 0 2944 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input114
timestamp 1688980957
transform 1 0 4140 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input115
timestamp 1688980957
transform 1 0 4324 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input116
timestamp 1688980957
transform 1 0 3312 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input117
timestamp 1688980957
transform 1 0 4508 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input118
timestamp 1688980957
transform 1 0 4968 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input119
timestamp 1688980957
transform 1 0 4876 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input120
timestamp 1688980957
transform 1 0 4048 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input121
timestamp 1688980957
transform 1 0 6440 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input122
timestamp 1688980957
transform 1 0 8188 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input123
timestamp 1688980957
transform 1 0 8280 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input124
timestamp 1688980957
transform 1 0 8740 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input125
timestamp 1688980957
transform 1 0 8556 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input126
timestamp 1688980957
transform 1 0 9016 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input127
timestamp 1688980957
transform 1 0 8004 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input128
timestamp 1688980957
transform 1 0 5520 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__dlymetal6s2s_1  input129
timestamp 1688980957
transform 1 0 7084 0 1 1088
box -38 -48 958 592
use sky130_fd_sc_hd__clkbuf_2  input130
timestamp 1688980957
transform 1 0 5888 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input131
timestamp 1688980957
transform 1 0 7452 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input132
timestamp 1688980957
transform 1 0 6808 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input133
timestamp 1688980957
transform 1 0 7820 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input134
timestamp 1688980957
transform 1 0 7360 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input135
timestamp 1688980957
transform 1 0 7636 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input136
timestamp 1688980957
transform 1 0 7912 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input137
timestamp 1688980957
transform 1 0 18860 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input138
timestamp 1688980957
transform 1 0 18308 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input139
timestamp 1688980957
transform 1 0 18216 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input140
timestamp 1688980957
transform 1 0 18860 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input141
timestamp 1688980957
transform 1 0 13524 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input142
timestamp 1688980957
transform 1 0 14076 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input143
timestamp 1688980957
transform 1 0 14904 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input144
timestamp 1688980957
transform 1 0 16008 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input145
timestamp 1688980957
transform 1 0 19228 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input146
timestamp 1688980957
transform 1 0 19228 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input147
timestamp 1688980957
transform 1 0 14444 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input148
timestamp 1688980957
transform 1 0 12788 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input149
timestamp 1688980957
transform 1 0 18124 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input150
timestamp 1688980957
transform 1 0 18400 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input151
timestamp 1688980957
transform 1 0 18952 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input152
timestamp 1688980957
transform 1 0 18676 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input153
timestamp 1688980957
transform 1 0 9844 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input154
timestamp 1688980957
transform 1 0 9292 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  input155
timestamp 1688980957
transform 1 0 9660 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  input156
timestamp 1688980957
transform 1 0 10212 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input157
timestamp 1688980957
transform 1 0 10304 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input158
timestamp 1688980957
transform 1 0 10580 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input159
timestamp 1688980957
transform 1 0 10764 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input160
timestamp 1688980957
transform 1 0 10856 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input161
timestamp 1688980957
transform 1 0 11132 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input162
timestamp 1688980957
transform 1 0 12144 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input163
timestamp 1688980957
transform 1 0 11500 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input164
timestamp 1688980957
transform 1 0 11132 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input165
timestamp 1688980957
transform 1 0 11868 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input166
timestamp 1688980957
transform 1 0 11684 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input167
timestamp 1688980957
transform 1 0 12236 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input168
timestamp 1688980957
transform 1 0 11960 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input169
timestamp 1688980957
transform 1 0 12604 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input170
timestamp 1688980957
transform 1 0 12788 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__buf_1  input171
timestamp 1688980957
transform 1 0 13708 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input172
timestamp 1688980957
transform 1 0 13156 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  input173
timestamp 1688980957
transform 1 0 14076 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input174
timestamp 1688980957
transform 1 0 15456 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input175
timestamp 1688980957
transform 1 0 13432 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input176
timestamp 1688980957
transform 1 0 17848 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input177
timestamp 1688980957
transform 1 0 18676 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input178
timestamp 1688980957
transform 1 0 15916 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input179
timestamp 1688980957
transform 1 0 16928 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  input180
timestamp 1688980957
transform 1 0 13524 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  input181
timestamp 1688980957
transform 1 0 14444 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  input182
timestamp 1688980957
transform 1 0 14076 0 1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  input183
timestamp 1688980957
transform 1 0 15640 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input184
timestamp 1688980957
transform 1 0 16192 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input185
timestamp 1688980957
transform 1 0 14168 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input186
timestamp 1688980957
transform 1 0 14628 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input187
timestamp 1688980957
transform 1 0 14904 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input188
timestamp 1688980957
transform 1 0 15180 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  inst_clk_buf
timestamp 1688980957
transform 1 0 15088 0 1 42432
box -38 -48 1878 592
use sky130_fd_sc_hd__clkbuf_1  Inst_Config_accessConfig_access._0_
timestamp 1688980957
transform 1 0 21160 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_Config_accessConfig_access._1_
timestamp 1688980957
transform 1 0 21344 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_Config_accessConfig_access._2_
timestamp 1688980957
transform 1 0 19228 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_Config_accessConfig_access._3_
timestamp 1688980957
transform 1 0 19688 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_A0_OutPass4_frame_config_mux._0_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 19228 0 -1 17408
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_A0_OutPass4_frame_config_mux._1_
timestamp 1688980957
transform 1 0 14260 0 1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_A0_OutPass4_frame_config_mux._2_
timestamp 1688980957
transform 1 0 18676 0 -1 18496
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_A0_OutPass4_frame_config_mux._3_
timestamp 1688980957
transform 1 0 14812 0 1 34816
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst0._2_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 20976 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst0._3_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 20792 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst0._4_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 20700 0 1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 19688 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 18952 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst1._2_
timestamp 1688980957
transform 1 0 15732 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst1._3_
timestamp 1688980957
transform 1 0 16008 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst1._4_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 15456 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 14812 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 16284 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst2._2_
timestamp 1688980957
transform 1 0 19964 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst2._3_
timestamp 1688980957
transform 1 0 20976 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst2._4_
timestamp 1688980957
transform 1 0 20332 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 19228 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 20700 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst3._2_
timestamp 1688980957
transform 1 0 15916 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst3._3_
timestamp 1688980957
transform 1 0 17664 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst3._4_
timestamp 1688980957
transform 1 0 16652 0 -1 35904
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 15272 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 16284 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_A1_OutPass4_frame_config_mux._0_
timestamp 1688980957
transform 1 0 19228 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_A1_OutPass4_frame_config_mux._1_
timestamp 1688980957
transform 1 0 17296 0 1 15232
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_A1_OutPass4_frame_config_mux._2_
timestamp 1688980957
transform 1 0 18676 0 -1 35904
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_A1_OutPass4_frame_config_mux._3_
timestamp 1688980957
transform 1 0 16652 0 -1 36992
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst0._2_
timestamp 1688980957
transform 1 0 20240 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst0._3_
timestamp 1688980957
transform 1 0 20884 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst0._4_
timestamp 1688980957
transform 1 0 20884 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 19596 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 20608 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst1._2_
timestamp 1688980957
transform 1 0 18308 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst1._3_
timestamp 1688980957
transform 1 0 19044 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst1._4_
timestamp 1688980957
transform 1 0 18768 0 1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 17020 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 18768 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst2._2_
timestamp 1688980957
transform 1 0 18860 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst2._3_
timestamp 1688980957
transform 1 0 20332 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst2._4_
timestamp 1688980957
transform 1 0 20608 0 1 34816
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 19228 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 20608 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst3._2_
timestamp 1688980957
transform 1 0 17204 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst3._3_
timestamp 1688980957
transform 1 0 17940 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst3._4_
timestamp 1688980957
transform 1 0 18124 0 -1 36992
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 16560 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 17664 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_C_OutPass4_frame_config_mux._0_
timestamp 1688980957
transform 1 0 17664 0 1 13056
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_C_OutPass4_frame_config_mux._1_
timestamp 1688980957
transform 1 0 19228 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_C_OutPass4_frame_config_mux._2_
timestamp 1688980957
transform 1 0 19412 0 -1 14144
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_C_OutPass4_frame_config_mux._3_
timestamp 1688980957
transform 1 0 19228 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst0._2_
timestamp 1688980957
transform 1 0 18952 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst0._3_
timestamp 1688980957
transform 1 0 19412 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst0._4_
timestamp 1688980957
transform 1 0 19688 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 19228 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 20056 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst1._2_
timestamp 1688980957
transform 1 0 20608 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst1._3_
timestamp 1688980957
transform 1 0 18952 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst1._4_
timestamp 1688980957
transform 1 0 20884 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 19596 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 21068 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst2._2_
timestamp 1688980957
transform 1 0 20424 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst2._3_
timestamp 1688980957
transform 1 0 20240 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst2._4_
timestamp 1688980957
transform 1 0 21252 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 21344 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 21344 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst3._2_
timestamp 1688980957
transform 1 0 20332 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst3._3_
timestamp 1688980957
transform 1 0 20608 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst3._4_
timestamp 1688980957
transform 1 0 20700 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 19688 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 20516 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_D0_OutPass4_frame_config_mux._0_
timestamp 1688980957
transform 1 0 17296 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_D0_OutPass4_frame_config_mux._1_
timestamp 1688980957
transform 1 0 16468 0 1 32640
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_D0_OutPass4_frame_config_mux._2_
timestamp 1688980957
transform 1 0 17756 0 -1 26112
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_D0_OutPass4_frame_config_mux._3_
timestamp 1688980957
transform 1 0 15824 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst0._2_
timestamp 1688980957
transform 1 0 19136 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst0._3_
timestamp 1688980957
transform 1 0 18400 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst0._4_
timestamp 1688980957
transform 1 0 18768 0 -1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 17848 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 18676 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst1._2_
timestamp 1688980957
transform 1 0 17296 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst1._3_
timestamp 1688980957
transform 1 0 18584 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst1._4_
timestamp 1688980957
transform 1 0 17940 0 1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 16652 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 18308 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst2._2_
timestamp 1688980957
transform 1 0 19228 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst2._3_
timestamp 1688980957
transform 1 0 19780 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst2._4_
timestamp 1688980957
transform 1 0 19412 0 1 25024
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 18308 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 19504 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst3._2_
timestamp 1688980957
transform 1 0 17388 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst3._3_
timestamp 1688980957
transform 1 0 18032 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst3._4_
timestamp 1688980957
transform 1 0 17296 0 1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 16192 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 17664 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_D1_OutPass4_frame_config_mux._0_
timestamp 1688980957
transform 1 0 17848 0 -1 22848
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_D1_OutPass4_frame_config_mux._1_
timestamp 1688980957
transform 1 0 17664 0 1 28288
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_D1_OutPass4_frame_config_mux._2_
timestamp 1688980957
transform 1 0 19596 0 -1 25024
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_D1_OutPass4_frame_config_mux._3_
timestamp 1688980957
transform 1 0 16652 0 -1 29376
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst0._2_
timestamp 1688980957
transform 1 0 18860 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst0._3_
timestamp 1688980957
transform 1 0 18860 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst0._4_
timestamp 1688980957
transform 1 0 21252 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 18308 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 19228 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst1._2_
timestamp 1688980957
transform 1 0 19136 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst1._3_
timestamp 1688980957
transform 1 0 19872 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst1._4_
timestamp 1688980957
transform 1 0 19228 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 19596 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 20148 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst2._2_
timestamp 1688980957
transform 1 0 20976 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst2._3_
timestamp 1688980957
transform 1 0 20424 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst2._4_
timestamp 1688980957
transform 1 0 20700 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 20056 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 20700 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst3._2_
timestamp 1688980957
transform 1 0 17388 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst3._3_
timestamp 1688980957
transform 1 0 18860 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst3._4_
timestamp 1688980957
transform 1 0 18492 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 17204 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 17940 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_D2_OutPass4_frame_config_mux._0_
timestamp 1688980957
transform 1 0 19412 0 1 21760
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_D2_OutPass4_frame_config_mux._1_
timestamp 1688980957
transform 1 0 16652 0 -1 31552
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_D2_OutPass4_frame_config_mux._2_
timestamp 1688980957
transform 1 0 19228 0 1 23936
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_D2_OutPass4_frame_config_mux._3_
timestamp 1688980957
transform 1 0 15640 0 1 30464
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst0._2_
timestamp 1688980957
transform 1 0 20056 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst0._3_
timestamp 1688980957
transform 1 0 20884 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst0._4_
timestamp 1688980957
transform 1 0 20976 0 -1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 21344 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 20976 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst1._2_
timestamp 1688980957
transform 1 0 17756 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst1._3_
timestamp 1688980957
transform 1 0 18400 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst1._4_
timestamp 1688980957
transform 1 0 18124 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 17388 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 18124 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst2._2_
timestamp 1688980957
transform 1 0 21344 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst2._3_
timestamp 1688980957
transform 1 0 19044 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst2._4_
timestamp 1688980957
transform 1 0 20976 0 -1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 19320 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 20700 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst3._2_
timestamp 1688980957
transform 1 0 16560 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst3._3_
timestamp 1688980957
transform 1 0 16284 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst3._4_
timestamp 1688980957
transform 1 0 16836 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 16008 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 17112 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_D3_OutPass4_frame_config_mux._0_
timestamp 1688980957
transform 1 0 19228 0 1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_D3_OutPass4_frame_config_mux._1_
timestamp 1688980957
transform 1 0 19228 0 1 27200
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_D3_OutPass4_frame_config_mux._2_
timestamp 1688980957
transform 1 0 19044 0 -1 19584
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_FAB2RAM_D3_OutPass4_frame_config_mux._3_
timestamp 1688980957
transform 1 0 16284 0 1 33728
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst0._2_
timestamp 1688980957
transform 1 0 18768 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst0._3_
timestamp 1688980957
transform 1 0 20884 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst0._4_
timestamp 1688980957
transform 1 0 20516 0 -1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 18860 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 19228 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst1._2_
timestamp 1688980957
transform 1 0 20332 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst1._3_
timestamp 1688980957
transform 1 0 20792 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst1._4_
timestamp 1688980957
transform 1 0 20976 0 -1 27200
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 19688 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 20608 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst2._2_
timestamp 1688980957
transform 1 0 20608 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst2._3_
timestamp 1688980957
transform 1 0 20332 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst2._4_
timestamp 1688980957
transform 1 0 20884 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 18584 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 20608 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst3._2_
timestamp 1688980957
transform 1 0 18216 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst3._3_
timestamp 1688980957
transform 1 0 18768 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst3._4_
timestamp 1688980957
transform 1 0 17848 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 16744 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 18492 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  Inst_RAM2FAB_D0_InPass4_frame_config_mux._0_
timestamp 1688980957
transform 1 0 19964 0 1 10880
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_RAM2FAB_D0_InPass4_frame_config_mux._1_
timestamp 1688980957
transform 1 0 17204 0 -1 11968
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_RAM2FAB_D0_InPass4_frame_config_mux._2_
timestamp 1688980957
transform 1 0 19964 0 -1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_RAM2FAB_D0_InPass4_frame_config_mux._3_
timestamp 1688980957
transform 1 0 16928 0 -1 8704
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst0._2_
timestamp 1688980957
transform 1 0 19688 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst0._3_
timestamp 1688980957
transform 1 0 19964 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_4  Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst0._4_ dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 20148 0 -1 11968
box -38 -48 1234 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 19412 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 20976 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst1._2_
timestamp 1688980957
transform 1 0 16928 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst1._3_
timestamp 1688980957
transform 1 0 18216 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_4  Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst1._4_
timestamp 1688980957
transform 1 0 17480 0 1 10880
box -38 -48 1234 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 18492 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 18676 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst2._2_
timestamp 1688980957
transform 1 0 19412 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst2._3_
timestamp 1688980957
transform 1 0 20884 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_4  Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst2._4_
timestamp 1688980957
transform 1 0 19688 0 1 6528
box -38 -48 1234 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 18860 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 21344 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst3._2_
timestamp 1688980957
transform 1 0 17664 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst3._3_
timestamp 1688980957
transform 1 0 18492 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_4  Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst3._4_
timestamp 1688980957
transform 1 0 16652 0 -1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 16652 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 18768 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  Inst_RAM2FAB_D1_InPass4_frame_config_mux._0_
timestamp 1688980957
transform 1 0 16652 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_RAM2FAB_D1_InPass4_frame_config_mux._1_
timestamp 1688980957
transform 1 0 17112 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_RAM2FAB_D1_InPass4_frame_config_mux._2_
timestamp 1688980957
transform 1 0 19872 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_RAM2FAB_D1_InPass4_frame_config_mux._3_
timestamp 1688980957
transform 1 0 16560 0 1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst0._2_
timestamp 1688980957
transform 1 0 15824 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst0._3_
timestamp 1688980957
transform 1 0 16836 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_4  Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst0._4_
timestamp 1688980957
transform 1 0 16652 0 -1 6528
box -38 -48 1234 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 16560 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 17112 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst1._2_
timestamp 1688980957
transform 1 0 17572 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst1._3_
timestamp 1688980957
transform 1 0 18676 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_4  Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst1._4_
timestamp 1688980957
transform 1 0 17480 0 -1 4352
box -38 -48 1234 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 17848 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 18584 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst2._2_
timestamp 1688980957
transform 1 0 18584 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst2._3_
timestamp 1688980957
transform 1 0 20608 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_4  Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst2._4_
timestamp 1688980957
transform 1 0 17940 0 1 7616
box -38 -48 1234 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 20884 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 18032 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst3._2_
timestamp 1688980957
transform 1 0 17848 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst3._3_
timestamp 1688980957
transform 1 0 16008 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst3._4_
timestamp 1688980957
transform 1 0 15640 0 1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 16284 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 18124 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  Inst_RAM2FAB_D2_InPass4_frame_config_mux._0_
timestamp 1688980957
transform 1 0 14260 0 -1 5440
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_RAM2FAB_D2_InPass4_frame_config_mux._1_
timestamp 1688980957
transform 1 0 19964 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_RAM2FAB_D2_InPass4_frame_config_mux._2_
timestamp 1688980957
transform 1 0 19596 0 -1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_RAM2FAB_D2_InPass4_frame_config_mux._3_
timestamp 1688980957
transform 1 0 14168 0 1 4352
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst0._2_
timestamp 1688980957
transform 1 0 13708 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst0._3_
timestamp 1688980957
transform 1 0 15732 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst0._4_
timestamp 1688980957
transform 1 0 14260 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 15732 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 15548 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst1._2_
timestamp 1688980957
transform 1 0 15180 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst1._3_
timestamp 1688980957
transform 1 0 16284 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_4  Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst1._4_
timestamp 1688980957
transform 1 0 17480 0 1 5440
box -38 -48 1234 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 14628 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 14352 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst2._2_
timestamp 1688980957
transform 1 0 15456 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst2._3_
timestamp 1688980957
transform 1 0 17940 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst2._4_
timestamp 1688980957
transform 1 0 20884 0 -1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 14628 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 14076 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst3._2_
timestamp 1688980957
transform 1 0 16008 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst3._3_
timestamp 1688980957
transform 1 0 16284 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst3._4_
timestamp 1688980957
transform 1 0 14904 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 14444 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 15640 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__dfxtp_1  Inst_RAM2FAB_D3_InPass4_frame_config_mux._0_
timestamp 1688980957
transform 1 0 14260 0 -1 6528
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_RAM2FAB_D3_InPass4_frame_config_mux._1_
timestamp 1688980957
transform 1 0 19228 0 1 3264
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_RAM2FAB_D3_InPass4_frame_config_mux._2_
timestamp 1688980957
transform 1 0 19412 0 1 7616
box -38 -48 1510 592
use sky130_fd_sc_hd__dfxtp_1  Inst_RAM2FAB_D3_InPass4_frame_config_mux._3_
timestamp 1688980957
transform 1 0 17756 0 -1 9792
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst0._2_
timestamp 1688980957
transform 1 0 13708 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst0._3_
timestamp 1688980957
transform 1 0 14996 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst0._4_
timestamp 1688980957
transform 1 0 14352 0 -1 7616
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 13984 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst0.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 15456 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst1._2_
timestamp 1688980957
transform 1 0 19504 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst1._3_
timestamp 1688980957
transform 1 0 18860 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_4  Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst1._4_
timestamp 1688980957
transform 1 0 18676 0 -1 3264
box -38 -48 1234 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 14168 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst1.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 21068 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst2._2_
timestamp 1688980957
transform 1 0 21344 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst2._3_
timestamp 1688980957
transform 1 0 19320 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst2._4_
timestamp 1688980957
transform 1 0 20884 0 -1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 20884 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst2.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 21344 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst3._2_
timestamp 1688980957
transform 1 0 18216 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst3._3_
timestamp 1688980957
transform 1 0 18584 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst3._4_
timestamp 1688980957
transform 1 0 17940 0 1 9792
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 17480 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst3.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 19228 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit0 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 14260 0 -1 8704
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit1
timestamp 1688980957
transform 1 0 15456 0 1 8704
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit2
timestamp 1688980957
transform 1 0 4876 0 -1 30464
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit3
timestamp 1688980957
transform 1 0 4876 0 -1 29376
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit4
timestamp 1688980957
transform 1 0 4692 0 -1 11968
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit5
timestamp 1688980957
transform 1 0 6072 0 1 11968
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit6
timestamp 1688980957
transform 1 0 9752 0 1 26112
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit7
timestamp 1688980957
transform 1 0 12880 0 -1 26112
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit8
timestamp 1688980957
transform 1 0 7452 0 1 32640
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit9
timestamp 1688980957
transform 1 0 9016 0 -1 33728
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit10
timestamp 1688980957
transform 1 0 4876 0 -1 35904
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit11
timestamp 1688980957
transform 1 0 6256 0 1 34816
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit12
timestamp 1688980957
transform 1 0 4876 0 -1 5440
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit13
timestamp 1688980957
transform 1 0 6532 0 1 5440
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit14
timestamp 1688980957
transform 1 0 7636 0 -1 34816
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit15
timestamp 1688980957
transform 1 0 9292 0 1 33728
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit16
timestamp 1688980957
transform 1 0 6992 0 -1 35904
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit17
timestamp 1688980957
transform 1 0 8924 0 1 35904
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit18
timestamp 1688980957
transform 1 0 4048 0 1 20672
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit19
timestamp 1688980957
transform 1 0 4876 0 -1 19584
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit20
timestamp 1688980957
transform 1 0 6716 0 1 38080
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit21
timestamp 1688980957
transform 1 0 7268 0 -1 36992
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit22
timestamp 1688980957
transform 1 0 9660 0 -1 38080
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit23
timestamp 1688980957
transform 1 0 10028 0 -1 36992
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit24
timestamp 1688980957
transform 1 0 14628 0 -1 16320
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit25
timestamp 1688980957
transform 1 0 16836 0 1 16320
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit26
timestamp 1688980957
transform 1 0 5336 0 1 38080
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit27
timestamp 1688980957
transform 1 0 6348 0 -1 39168
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit28
timestamp 1688980957
transform 1 0 4876 0 -1 16320
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit29
timestamp 1688980957
transform 1 0 6808 0 -1 18496
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit30
timestamp 1688980957
transform 1 0 9016 0 1 32640
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame0_bit31
timestamp 1688980957
transform 1 0 9752 0 -1 31552
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit0
timestamp 1688980957
transform 1 0 16652 0 -1 16320
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit1
timestamp 1688980957
transform 1 0 17664 0 1 17408
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit2
timestamp 1688980957
transform 1 0 7268 0 -1 32640
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit3
timestamp 1688980957
transform 1 0 7452 0 1 31552
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit4
timestamp 1688980957
transform 1 0 7452 0 1 18496
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit5
timestamp 1688980957
transform 1 0 8924 0 1 17408
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit6
timestamp 1688980957
transform 1 0 14628 0 -1 33728
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit7
timestamp 1688980957
transform 1 0 14904 0 1 33728
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit8
timestamp 1688980957
transform 1 0 16652 0 -1 14144
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit9
timestamp 1688980957
transform 1 0 16100 0 1 13056
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit10
timestamp 1688980957
transform 1 0 4048 0 -1 36992
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit11
timestamp 1688980957
transform 1 0 4876 0 1 34816
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit12
timestamp 1688980957
transform 1 0 4692 0 1 11968
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit13
timestamp 1688980957
transform 1 0 6072 0 1 13056
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit14
timestamp 1688980957
transform 1 0 9936 0 1 27200
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit15
timestamp 1688980957
transform 1 0 11592 0 -1 28288
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit16
timestamp 1688980957
transform 1 0 14076 0 1 8704
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit17
timestamp 1688980957
transform 1 0 16008 0 1 9792
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit18
timestamp 1688980957
transform 1 0 3220 0 -1 34816
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit19
timestamp 1688980957
transform 1 0 4600 0 -1 38080
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit20
timestamp 1688980957
transform 1 0 4876 0 -1 15232
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit21
timestamp 1688980957
transform 1 0 7452 0 1 16320
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit22
timestamp 1688980957
transform 1 0 10028 0 -1 27200
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit23
timestamp 1688980957
transform 1 0 11408 0 1 28288
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit24
timestamp 1688980957
transform 1 0 14996 0 1 11968
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit25
timestamp 1688980957
transform 1 0 15548 0 1 10880
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit26
timestamp 1688980957
transform 1 0 4600 0 -1 33728
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit27
timestamp 1688980957
transform 1 0 6348 0 1 33728
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit28
timestamp 1688980957
transform 1 0 8096 0 -1 16320
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit29
timestamp 1688980957
transform 1 0 6992 0 1 14144
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit30
timestamp 1688980957
transform 1 0 11500 0 -1 26112
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame1_bit31
timestamp 1688980957
transform 1 0 11500 0 -1 25024
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit0
timestamp 1688980957
transform 1 0 14996 0 -1 25024
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit1
timestamp 1688980957
transform 1 0 16652 0 -1 23936
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit2
timestamp 1688980957
transform 1 0 2852 0 -1 31552
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit3
timestamp 1688980957
transform 1 0 3312 0 -1 30464
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit4
timestamp 1688980957
transform 1 0 1564 0 1 27200
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit5
timestamp 1688980957
transform 1 0 3772 0 1 26112
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit6
timestamp 1688980957
transform 1 0 13432 0 -1 30464
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit7
timestamp 1688980957
transform 1 0 14076 0 1 30464
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit8
timestamp 1688980957
transform 1 0 16652 0 1 20672
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit9
timestamp 1688980957
transform 1 0 16744 0 -1 20672
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit10
timestamp 1688980957
transform 1 0 1564 0 -1 29376
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit11
timestamp 1688980957
transform 1 0 2208 0 1 28288
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit12
timestamp 1688980957
transform 1 0 6624 0 -1 26112
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit13
timestamp 1688980957
transform 1 0 9660 0 -1 26112
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit14
timestamp 1688980957
transform 1 0 13984 0 -1 32640
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit15
timestamp 1688980957
transform 1 0 16008 0 1 31552
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit16
timestamp 1688980957
transform 1 0 12052 0 -1 18496
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit17
timestamp 1688980957
transform 1 0 14352 0 -1 19584
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit18
timestamp 1688980957
transform 1 0 3772 0 -1 39168
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit19
timestamp 1688980957
transform 1 0 3864 0 1 38080
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit20
timestamp 1688980957
transform 1 0 4508 0 1 19584
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit21
timestamp 1688980957
transform 1 0 4692 0 1 18496
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit22
timestamp 1688980957
transform 1 0 11224 0 1 35904
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit23
timestamp 1688980957
transform 1 0 11776 0 -1 35904
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit24
timestamp 1688980957
transform 1 0 7544 0 -1 21760
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit25
timestamp 1688980957
transform 1 0 8924 0 1 20672
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit26
timestamp 1688980957
transform 1 0 1472 0 -1 21760
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit27
timestamp 1688980957
transform 1 0 2300 0 1 19584
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit28
timestamp 1688980957
transform 1 0 1656 0 1 38080
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit29
timestamp 1688980957
transform 1 0 2208 0 1 35904
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit30
timestamp 1688980957
transform 1 0 12328 0 1 36992
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame2_bit31
timestamp 1688980957
transform 1 0 12972 0 -1 38080
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit0
timestamp 1688980957
transform 1 0 11868 0 -1 16320
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit1
timestamp 1688980957
transform 1 0 12420 0 1 16320
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit2
timestamp 1688980957
transform 1 0 4876 0 -1 14144
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit3
timestamp 1688980957
transform 1 0 5704 0 1 17408
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit4
timestamp 1688980957
transform 1 0 2116 0 1 8704
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit5
timestamp 1688980957
transform 1 0 5060 0 1 9792
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit6
timestamp 1688980957
transform 1 0 12052 0 -1 15232
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit7
timestamp 1688980957
transform 1 0 13248 0 -1 16320
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit8
timestamp 1688980957
transform 1 0 8924 0 1 16320
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit9
timestamp 1688980957
transform 1 0 10028 0 -1 18496
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit10
timestamp 1688980957
transform 1 0 2392 0 -1 17408
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit11
timestamp 1688980957
transform 1 0 3496 0 -1 19584
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit12
timestamp 1688980957
transform 1 0 2300 0 1 14144
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit13
timestamp 1688980957
transform 1 0 4232 0 1 14144
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit14
timestamp 1688980957
transform 1 0 12604 0 1 17408
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit15
timestamp 1688980957
transform 1 0 13892 0 -1 18496
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit16
timestamp 1688980957
transform 1 0 15088 0 1 25024
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit17
timestamp 1688980957
transform 1 0 16468 0 1 25024
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit18
timestamp 1688980957
transform 1 0 1840 0 -1 34816
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit19
timestamp 1688980957
transform 1 0 2300 0 1 32640
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit20
timestamp 1688980957
transform 1 0 1656 0 -1 26112
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit21
timestamp 1688980957
transform 1 0 2300 0 1 25024
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit22
timestamp 1688980957
transform 1 0 15180 0 -1 29376
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit23
timestamp 1688980957
transform 1 0 16008 0 1 28288
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit24
timestamp 1688980957
transform 1 0 14904 0 -1 22848
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit25
timestamp 1688980957
transform 1 0 17296 0 1 21760
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit26
timestamp 1688980957
transform 1 0 3220 0 -1 29376
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit27
timestamp 1688980957
transform 1 0 3864 0 1 28288
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit28
timestamp 1688980957
transform 1 0 7452 0 1 26112
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit29
timestamp 1688980957
transform 1 0 9568 0 -1 25024
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit30
timestamp 1688980957
transform 1 0 14812 0 -1 30464
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame3_bit31
timestamp 1688980957
transform 1 0 14444 0 -1 31552
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit0
timestamp 1688980957
transform 1 0 9384 0 1 9792
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit1
timestamp 1688980957
transform 1 0 7452 0 1 11968
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit2
timestamp 1688980957
transform 1 0 1656 0 -1 11968
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit3
timestamp 1688980957
transform 1 0 2208 0 1 13056
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit4
timestamp 1688980957
transform 1 0 4140 0 1 7616
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit5
timestamp 1688980957
transform 1 0 3772 0 1 8704
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit6
timestamp 1688980957
transform 1 0 12052 0 -1 13056
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit7
timestamp 1688980957
transform 1 0 12604 0 1 11968
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit8
timestamp 1688980957
transform 1 0 9200 0 1 15232
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit9
timestamp 1688980957
transform 1 0 10028 0 -1 15232
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit10
timestamp 1688980957
transform 1 0 2300 0 1 18496
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit11
timestamp 1688980957
transform 1 0 2392 0 -1 18496
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit12
timestamp 1688980957
transform 1 0 4324 0 -1 6528
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit13
timestamp 1688980957
transform 1 0 4784 0 -1 8704
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit14
timestamp 1688980957
transform 1 0 11500 0 -1 8704
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit15
timestamp 1688980957
transform 1 0 11960 0 1 8704
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit16
timestamp 1688980957
transform 1 0 7452 0 1 13056
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit17
timestamp 1688980957
transform 1 0 8648 0 -1 15232
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit18
timestamp 1688980957
transform 1 0 2300 0 1 7616
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit19
timestamp 1688980957
transform 1 0 2300 0 1 9792
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit20
timestamp 1688980957
transform 1 0 1564 0 -1 15232
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit21
timestamp 1688980957
transform 1 0 3220 0 -1 14144
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit22
timestamp 1688980957
transform 1 0 14076 0 1 14144
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit23
timestamp 1688980957
transform 1 0 14536 0 1 15232
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit24
timestamp 1688980957
transform 1 0 13432 0 -1 13056
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit25
timestamp 1688980957
transform 1 0 14812 0 -1 13056
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit26
timestamp 1688980957
transform 1 0 4232 0 1 27200
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit27
timestamp 1688980957
transform 1 0 5612 0 1 27200
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit28
timestamp 1688980957
transform 1 0 4692 0 -1 13056
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit29
timestamp 1688980957
transform 1 0 5612 0 1 14144
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit30
timestamp 1688980957
transform 1 0 11040 0 1 22848
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame4_bit31
timestamp 1688980957
transform 1 0 12420 0 1 22848
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit0
timestamp 1688980957
transform 1 0 9292 0 -1 6528
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit1
timestamp 1688980957
transform 1 0 9568 0 1 6528
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit2
timestamp 1688980957
transform 1 0 3772 0 1 3264
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit3
timestamp 1688980957
transform 1 0 3036 0 -1 3264
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit4
timestamp 1688980957
transform 1 0 1564 0 1 3264
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit5
timestamp 1688980957
transform 1 0 1564 0 -1 4352
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit6
timestamp 1688980957
transform 1 0 14076 0 1 10880
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit7
timestamp 1688980957
transform 1 0 14536 0 -1 10880
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit8
timestamp 1688980957
transform 1 0 8648 0 -1 13056
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit9
timestamp 1688980957
transform 1 0 10028 0 -1 13056
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit10
timestamp 1688980957
transform 1 0 1380 0 1 15232
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit11
timestamp 1688980957
transform 1 0 1840 0 1 16320
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit12
timestamp 1688980957
transform 1 0 3864 0 1 4352
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit13
timestamp 1688980957
transform 1 0 3496 0 -1 5440
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit14
timestamp 1688980957
transform 1 0 7360 0 -1 9792
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit15
timestamp 1688980957
transform 1 0 9016 0 1 8704
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit16
timestamp 1688980957
transform 1 0 8004 0 -1 8704
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit17
timestamp 1688980957
transform 1 0 9568 0 1 7616
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit18
timestamp 1688980957
transform 1 0 1656 0 -1 3264
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit19
timestamp 1688980957
transform 1 0 2944 0 -1 4352
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit20
timestamp 1688980957
transform 1 0 1472 0 -1 6528
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit21
timestamp 1688980957
transform 1 0 2300 0 1 6528
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit22
timestamp 1688980957
transform 1 0 11684 0 1 13056
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit23
timestamp 1688980957
transform 1 0 11868 0 -1 14144
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit24
timestamp 1688980957
transform 1 0 10028 0 -1 10880
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit25
timestamp 1688980957
transform 1 0 10028 0 -1 11968
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit26
timestamp 1688980957
transform 1 0 6440 0 -1 8704
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit27
timestamp 1688980957
transform 1 0 6992 0 1 8704
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit28
timestamp 1688980957
transform 1 0 2300 0 1 11968
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit29
timestamp 1688980957
transform 1 0 2300 0 1 10880
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit30
timestamp 1688980957
transform 1 0 10580 0 1 8704
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame5_bit31
timestamp 1688980957
transform 1 0 12880 0 -1 8704
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit0
timestamp 1688980957
transform 1 0 2852 0 -1 21760
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit1
timestamp 1688980957
transform 1 0 3772 0 1 22848
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit2
timestamp 1688980957
transform 1 0 11500 0 -1 20672
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit3
timestamp 1688980957
transform 1 0 10028 0 -1 19584
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit4
timestamp 1688980957
transform 1 0 12604 0 1 19584
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit5
timestamp 1688980957
transform 1 0 14076 0 1 20672
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit6
timestamp 1688980957
transform 1 0 14996 0 -1 20672
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit7
timestamp 1688980957
transform 1 0 4416 0 -1 25024
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit8
timestamp 1688980957
transform 1 0 4876 0 -1 23936
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit9
timestamp 1688980957
transform 1 0 6808 0 -1 22848
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit10
timestamp 1688980957
transform 1 0 7176 0 1 23936
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit11
timestamp 1688980957
transform 1 0 7452 0 1 22848
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit12
timestamp 1688980957
transform 1 0 10120 0 1 23936
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit13
timestamp 1688980957
transform 1 0 14076 0 1 27200
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit14
timestamp 1688980957
transform 1 0 13984 0 -1 28288
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit15
timestamp 1688980957
transform 1 0 16008 0 1 26112
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit16
timestamp 1688980957
transform 1 0 10948 0 1 6528
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit17
timestamp 1688980957
transform 1 0 11500 0 -1 7616
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit18
timestamp 1688980957
transform 1 0 5612 0 1 8704
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit19
timestamp 1688980957
transform 1 0 4784 0 -1 7616
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit20
timestamp 1688980957
transform 1 0 3312 0 -1 11968
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit21
timestamp 1688980957
transform 1 0 7268 0 -1 10880
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit22
timestamp 1688980957
transform 1 0 9936 0 -1 17408
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit23
timestamp 1688980957
transform 1 0 10672 0 1 17408
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit24
timestamp 1688980957
transform 1 0 7452 0 1 10880
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit25
timestamp 1688980957
transform 1 0 8648 0 -1 10880
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit26
timestamp 1688980957
transform 1 0 2116 0 -1 5440
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit27
timestamp 1688980957
transform 1 0 2300 0 1 4352
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit28
timestamp 1688980957
transform 1 0 5244 0 1 4352
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit29
timestamp 1688980957
transform 1 0 4324 0 -1 4352
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit30
timestamp 1688980957
transform 1 0 6072 0 1 6528
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame6_bit31
timestamp 1688980957
transform 1 0 7452 0 1 6528
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit0
timestamp 1688980957
transform 1 0 12420 0 1 23936
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit1
timestamp 1688980957
transform 1 0 14812 0 -1 23936
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit2
timestamp 1688980957
transform 1 0 13156 0 -1 25024
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit3
timestamp 1688980957
transform 1 0 1564 0 1 33728
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit4
timestamp 1688980957
transform 1 0 3772 0 1 32640
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit5
timestamp 1688980957
transform 1 0 7176 0 -1 33728
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit6
timestamp 1688980957
transform 1 0 4876 0 -1 27200
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit7
timestamp 1688980957
transform 1 0 4324 0 1 25024
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit8
timestamp 1688980957
transform 1 0 8280 0 -1 27200
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit9
timestamp 1688980957
transform 1 0 9752 0 1 29376
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit10
timestamp 1688980957
transform 1 0 11500 0 -1 29376
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit11
timestamp 1688980957
transform 1 0 11500 0 -1 31552
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit12
timestamp 1688980957
transform 1 0 15180 0 -1 17408
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit13
timestamp 1688980957
transform 1 0 16652 0 -1 18496
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit14
timestamp 1688980957
transform 1 0 4876 0 -1 31552
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit15
timestamp 1688980957
transform 1 0 6348 0 -1 30464
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit16
timestamp 1688980957
transform 1 0 6072 0 1 18496
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit17
timestamp 1688980957
transform 1 0 7452 0 -1 19584
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit18
timestamp 1688980957
transform 1 0 12604 0 1 32640
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit19
timestamp 1688980957
transform 1 0 12604 0 -1 32640
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit20
timestamp 1688980957
transform 1 0 9108 0 1 21760
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit21
timestamp 1688980957
transform 1 0 9660 0 1 22848
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit22
timestamp 1688980957
transform 1 0 1380 0 1 30464
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit23
timestamp 1688980957
transform 1 0 1656 0 -1 30464
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit24
timestamp 1688980957
transform 1 0 1472 0 -1 19584
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit25
timestamp 1688980957
transform 1 0 2300 0 1 20672
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit26
timestamp 1688980957
transform 1 0 9016 0 -1 28288
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit27
timestamp 1688980957
transform 1 0 9660 0 1 28288
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit28
timestamp 1688980957
transform 1 0 10580 0 1 21760
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit29
timestamp 1688980957
transform 1 0 11224 0 1 20672
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit30
timestamp 1688980957
transform 1 0 4232 0 -1 21760
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame7_bit31
timestamp 1688980957
transform 1 0 6532 0 1 21760
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit0
timestamp 1688980957
transform 1 0 18308 0 -1 13056
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit1
timestamp 1688980957
transform 1 0 19504 0 -1 30464
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit2
timestamp 1688980957
transform 1 0 19596 0 1 13056
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit3
timestamp 1688980957
transform 1 0 19596 0 -1 32640
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit4
timestamp 1688980957
transform 1 0 19964 0 -1 8704
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit5
timestamp 1688980957
transform 1 0 19596 0 1 8704
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit6
timestamp 1688980957
transform 1 0 19504 0 -1 9792
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit7
timestamp 1688980957
transform 1 0 19504 0 -1 10880
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit8
timestamp 1688980957
transform 1 0 15732 0 1 18496
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit9
timestamp 1688980957
transform 1 0 16652 0 -1 19584
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit10
timestamp 1688980957
transform 1 0 1380 0 -1 31552
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit11
timestamp 1688980957
transform 1 0 1564 0 -1 32640
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit12
timestamp 1688980957
transform 1 0 7084 0 1 28288
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit13
timestamp 1688980957
transform 1 0 7636 0 -1 28288
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit14
timestamp 1688980957
transform 1 0 10672 0 1 33728
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit15
timestamp 1688980957
transform 1 0 11500 0 -1 33728
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit16
timestamp 1688980957
transform 1 0 12972 0 -1 34816
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit17
timestamp 1688980957
transform 1 0 14352 0 -1 34816
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit18
timestamp 1688980957
transform 1 0 2668 0 -1 36992
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit19
timestamp 1688980957
transform 1 0 1472 0 1 36992
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit20
timestamp 1688980957
transform 1 0 1380 0 1 26112
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit21
timestamp 1688980957
transform 1 0 1656 0 1 23936
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit22
timestamp 1688980957
transform 1 0 7452 0 1 29376
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit23
timestamp 1688980957
transform 1 0 8556 0 -1 30464
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit24
timestamp 1688980957
transform 1 0 7452 0 1 35904
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit25
timestamp 1688980957
transform 1 0 8648 0 -1 36992
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit26
timestamp 1688980957
transform 1 0 1380 0 -1 23936
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit27
timestamp 1688980957
transform 1 0 1656 0 1 22848
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit28
timestamp 1688980957
transform 1 0 1472 0 1 39168
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit29
timestamp 1688980957
transform 1 0 1932 0 -1 39168
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit30
timestamp 1688980957
transform 1 0 9384 0 1 18496
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame8_bit31
timestamp 1688980957
transform 1 0 10028 0 -1 20672
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit0
timestamp 1688980957
transform 1 0 14076 0 1 6528
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit1
timestamp 1688980957
transform 1 0 19228 0 1 5440
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit2
timestamp 1688980957
transform 1 0 18492 0 -1 6528
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit3
timestamp 1688980957
transform 1 0 12880 0 -1 5440
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit4
timestamp 1688980957
transform 1 0 14076 0 1 7616
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit5
timestamp 1688980957
transform 1 0 19504 0 -1 5440
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit6
timestamp 1688980957
transform 1 0 19228 0 1 9792
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit7
timestamp 1688980957
transform 1 0 17296 0 -1 10880
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit8
timestamp 1688980957
transform 1 0 17572 0 1 23936
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit9
timestamp 1688980957
transform 1 0 16836 0 -1 32640
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit10
timestamp 1688980957
transform 1 0 19228 0 -1 26112
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit11
timestamp 1688980957
transform 1 0 16652 0 -1 27200
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit12
timestamp 1688980957
transform 1 0 19320 0 -1 22848
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit13
timestamp 1688980957
transform 1 0 18308 0 -1 29376
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit14
timestamp 1688980957
transform 1 0 19596 0 -1 23936
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit15
timestamp 1688980957
transform 1 0 17112 0 -1 28288
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit16
timestamp 1688980957
transform 1 0 19596 0 -1 21760
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit17
timestamp 1688980957
transform 1 0 18124 0 -1 31552
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit18
timestamp 1688980957
transform 1 0 19504 0 1 22848
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit19
timestamp 1688980957
transform 1 0 16652 0 -1 30464
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit20
timestamp 1688980957
transform 1 0 19228 0 1 18496
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit21
timestamp 1688980957
transform 1 0 19596 0 -1 27200
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit22
timestamp 1688980957
transform 1 0 19504 0 -1 20672
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit23
timestamp 1688980957
transform 1 0 17204 0 -1 34816
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit24
timestamp 1688980957
transform 1 0 19596 0 -1 16320
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit25
timestamp 1688980957
transform 1 0 14536 0 -1 38080
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit26
timestamp 1688980957
transform 1 0 19320 0 1 16320
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit27
timestamp 1688980957
transform 1 0 16284 0 1 34816
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit28
timestamp 1688980957
transform 1 0 19504 0 1 14144
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit29
timestamp 1688980957
transform 1 0 17756 0 -1 15232
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit30
timestamp 1688980957
transform 1 0 19228 0 1 34816
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame9_bit31
timestamp 1688980957
transform 1 0 16836 0 1 35904
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame10_bit24
timestamp 1688980957
transform 1 0 18768 0 -1 11968
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame10_bit25
timestamp 1688980957
transform 1 0 16836 0 1 11968
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame10_bit26
timestamp 1688980957
transform 1 0 18584 0 -1 8704
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame10_bit27
timestamp 1688980957
transform 1 0 16836 0 1 8704
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame10_bit28
timestamp 1688980957
transform 1 0 16100 0 1 5440
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame10_bit29
timestamp 1688980957
transform 1 0 18124 0 -1 5440
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame10_bit30
timestamp 1688980957
transform 1 0 18584 0 -1 7616
box -38 -48 1418 592
use sky130_fd_sc_hd__dlxbp_1  Inst_RAM_IO_ConfigMem.Inst_frame10_bit31
timestamp 1688980957
transform 1 0 16284 0 1 7616
box -38 -48 1418 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM_IO_switch_matrix._32_
timestamp 1688980957
transform 1 0 4508 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM_IO_switch_matrix._33_
timestamp 1688980957
transform 1 0 3956 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  Inst_RAM_IO_switch_matrix._34_
timestamp 1688980957
transform 1 0 3772 0 1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM_IO_switch_matrix._35_
timestamp 1688980957
transform 1 0 6348 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM_IO_switch_matrix._36_
timestamp 1688980957
transform 1 0 5980 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  Inst_RAM_IO_switch_matrix._37_
timestamp 1688980957
transform 1 0 5428 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM_IO_switch_matrix._38_
timestamp 1688980957
transform 1 0 5980 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM_IO_switch_matrix._39_
timestamp 1688980957
transform 1 0 5704 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  Inst_RAM_IO_switch_matrix._40_
timestamp 1688980957
transform 1 0 10580 0 -1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  Inst_RAM_IO_switch_matrix._41_
timestamp 1688980957
transform 1 0 10396 0 1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM_IO_switch_matrix._42_
timestamp 1688980957
transform 1 0 10396 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  Inst_RAM_IO_switch_matrix._43_
timestamp 1688980957
transform 1 0 10672 0 -1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  Inst_RAM_IO_switch_matrix._44_
timestamp 1688980957
transform 1 0 10948 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  Inst_RAM_IO_switch_matrix._45_
timestamp 1688980957
transform 1 0 11408 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  Inst_RAM_IO_switch_matrix._46_
timestamp 1688980957
transform 1 0 11684 0 1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  Inst_RAM_IO_switch_matrix._47_
timestamp 1688980957
transform 1 0 11500 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_A0_I0 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 12420 0 -1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_A0_I0_395 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 13340 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_A0_I1_396
timestamp 1688980957
transform 1 0 4324 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_A0_I1
timestamp 1688980957
transform 1 0 3772 0 1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_A0_I2_397
timestamp 1688980957
transform 1 0 6440 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_A0_I2 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 5888 0 1 19584
box -38 -48 1694 592
use sky130_fd_sc_hd__conb_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_A0_I3_398
timestamp 1688980957
transform 1 0 13156 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_A0_I3
timestamp 1688980957
transform 1 0 11592 0 1 34816
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_A1_I0_399
timestamp 1688980957
transform 1 0 10580 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_A1_I0
timestamp 1688980957
transform 1 0 8924 0 -1 21760
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_A1_I1
timestamp 1688980957
transform 1 0 3772 0 -1 20672
box -38 -48 1694 592
use sky130_fd_sc_hd__conb_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_A1_I1_400
timestamp 1688980957
transform 1 0 1840 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_A1_I2_401
timestamp 1688980957
transform 1 0 1472 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_A1_I2
timestamp 1688980957
transform 1 0 2024 0 1 34816
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_A1_I3
timestamp 1688980957
transform 1 0 12880 0 -1 36992
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_A1_I3_402
timestamp 1688980957
transform 1 0 14076 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_C_I0_403
timestamp 1688980957
transform 1 0 18584 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_C_I0
timestamp 1688980957
transform 1 0 16652 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_C_I1
timestamp 1688980957
transform 1 0 7268 0 -1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_C_I1_404
timestamp 1688980957
transform 1 0 8280 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_C_I2_405
timestamp 1688980957
transform 1 0 8924 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_C_I2
timestamp 1688980957
transform 1 0 8188 0 -1 18496
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_C_I3
timestamp 1688980957
transform 1 0 14536 0 1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_C_I3_409
timestamp 1688980957
transform 1 0 15456 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_D0_I0
timestamp 1688980957
transform 1 0 15364 0 1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_D0_I1
timestamp 1688980957
transform 1 0 2668 0 -1 33728
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_D0_I2
timestamp 1688980957
transform 1 0 3036 0 -1 26112
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_D0_I3
timestamp 1688980957
transform 1 0 14076 0 1 28288
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_D1_I0
timestamp 1688980957
transform 1 0 15364 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_D1_I1
timestamp 1688980957
transform 1 0 3772 0 -1 28288
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_D1_I2
timestamp 1688980957
transform 1 0 8924 0 1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_D1_I3
timestamp 1688980957
transform 1 0 14076 0 1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_D2_I0
timestamp 1688980957
transform 1 0 15364 0 1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_D2_I1
timestamp 1688980957
transform 1 0 3772 0 1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_D2_I2
timestamp 1688980957
transform 1 0 2576 0 -1 27200
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_D2_I3
timestamp 1688980957
transform 1 0 13248 0 -1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_D3_I0
timestamp 1688980957
transform 1 0 16652 0 -1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_D3_I1
timestamp 1688980957
transform 1 0 2116 0 -1 28288
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_D3_I2
timestamp 1688980957
transform 1 0 8004 0 -1 26112
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_FAB2RAM_D3_I3
timestamp 1688980957
transform 1 0 14076 0 1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS1_BEG0
timestamp 1688980957
transform 1 0 14904 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__conb_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS1_BEG0_406
timestamp 1688980957
transform 1 0 16008 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__conb_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS1_BEG1_407
timestamp 1688980957
transform 1 0 6440 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS1_BEG1
timestamp 1688980957
transform 1 0 5980 0 1 36992
box -38 -48 1694 592
use sky130_fd_sc_hd__conb_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS1_BEG2_408
timestamp 1688980957
transform 1 0 7176 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS1_BEG2
timestamp 1688980957
transform 1 0 7176 0 1 17408
box -38 -48 1694 592
use sky130_fd_sc_hd__conb_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS1_BEG3_394
timestamp 1688980957
transform 1 0 10764 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS1_BEG3
timestamp 1688980957
transform 1 0 9752 0 1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS2_BEG0
timestamp 1688980957
transform 1 0 8924 0 -1 32640
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS2_BEG1
timestamp 1688980957
transform 1 0 5612 0 1 35904
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS2_BEG2
timestamp 1688980957
transform 1 0 6348 0 -1 6528
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS2_BEG3
timestamp 1688980957
transform 1 0 9016 0 -1 34816
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS2_BEG4
timestamp 1688980957
transform 1 0 8924 0 1 34816
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS2_BEG5
timestamp 1688980957
transform 1 0 5980 0 1 20672
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS2_BEG6
timestamp 1688980957
transform 1 0 6900 0 -1 38080
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS2_BEG7
timestamp 1688980957
transform 1 0 10028 0 1 36992
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS4_BEG0
timestamp 1688980957
transform 1 0 14904 0 -1 14144
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS4_BEG1
timestamp 1688980957
transform 1 0 4600 0 -1 34816
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS4_BEG2
timestamp 1688980957
transform 1 0 6532 0 -1 14144
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS4_BEG3
timestamp 1688980957
transform 1 0 11316 0 1 27200
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS4_BEG4
timestamp 1688980957
transform 1 0 14352 0 1 9792
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS4_BEG5
timestamp 1688980957
transform 1 0 4692 0 1 33728
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS4_BEG6
timestamp 1688980957
transform 1 0 6992 0 -1 17408
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS4_BEG7
timestamp 1688980957
transform 1 0 11500 0 -1 27200
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS4_BEG8
timestamp 1688980957
transform 1 0 14812 0 -1 11968
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS4_BEG9
timestamp 1688980957
transform 1 0 5244 0 1 32640
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS4_BEG10
timestamp 1688980957
transform 1 0 6440 0 1 15232
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS4_BEG11
timestamp 1688980957
transform 1 0 11316 0 1 25024
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS4_BEG12
timestamp 1688980957
transform 1 0 14628 0 -1 9792
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS4_BEG13
timestamp 1688980957
transform 1 0 5152 0 1 29376
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS4_BEG14
timestamp 1688980957
transform 1 0 6440 0 -1 13056
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_J_NS4_BEG15
timestamp 1688980957
transform 1 0 11132 0 1 26112
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_N1BEG0
timestamp 1688980957
transform 1 0 16008 0 1 19584
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_N1BEG1
timestamp 1688980957
transform 1 0 1748 0 1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_N1BEG2
timestamp 1688980957
transform 1 0 7176 0 1 27200
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_N1BEG3
timestamp 1688980957
transform 1 0 10396 0 1 32640
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_N2BEG0
timestamp 1688980957
transform 1 0 12972 0 -1 33728
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_N2BEG1
timestamp 1688980957
transform 1 0 1748 0 -1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_N2BEG2
timestamp 1688980957
transform 1 0 1656 0 -1 25024
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_N2BEG3
timestamp 1688980957
transform 1 0 7360 0 -1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_N2BEG4
timestamp 1688980957
transform 1 0 8372 0 -1 35904
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_N2BEG5
timestamp 1688980957
transform 1 0 1472 0 -1 22848
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_N2BEG6
timestamp 1688980957
transform 1 0 1932 0 -1 38080
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_N2BEG7
timestamp 1688980957
transform 1 0 9752 0 1 19584
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_S1BEG0
timestamp 1688980957
transform 1 0 16008 0 1 17408
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_S1BEG1
timestamp 1688980957
transform 1 0 5888 0 1 30464
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_S1BEG2
timestamp 1688980957
transform 1 0 7360 0 -1 20672
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_S1BEG3
timestamp 1688980957
transform 1 0 12328 0 1 31552
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_S2BEG0
timestamp 1688980957
transform 1 0 9660 0 -1 22848
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_S2BEG1
timestamp 1688980957
transform 1 0 1840 0 1 29376
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_S2BEG2
timestamp 1688980957
transform 1 0 2116 0 -1 20672
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_S2BEG3
timestamp 1688980957
transform 1 0 9292 0 -1 29376
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_S2BEG4
timestamp 1688980957
transform 1 0 11500 0 -1 21760
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_S2BEG5
timestamp 1688980957
transform 1 0 4876 0 1 21760
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_2  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_S2BEG6
timestamp 1688980957
transform 1 0 3128 0 -1 22848
box -38 -48 1694 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_S2BEG7
timestamp 1688980957
transform 1 0 11040 0 1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W1BEG0
timestamp 1688980957
transform 1 0 11132 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W1BEG1
timestamp 1688980957
transform 1 0 6164 0 1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W1BEG2
timestamp 1688980957
transform 1 0 7360 0 -1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W1BEG3
timestamp 1688980957
transform 1 0 10304 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W2BEG0
timestamp 1688980957
transform 1 0 9200 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W2BEG1
timestamp 1688980957
transform 1 0 2392 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W2BEG2
timestamp 1688980957
transform 1 0 4048 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W2BEG3
timestamp 1688980957
transform 1 0 7544 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W2BEG4
timestamp 1688980957
transform 1 0 9476 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W2BEG5
timestamp 1688980957
transform 1 0 1748 0 1 5440
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W2BEG6
timestamp 1688980957
transform 1 0 2300 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W2BEG7
timestamp 1688980957
transform 1 0 12604 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W2BEGb0
timestamp 1688980957
transform 1 0 9752 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W2BEGb1
timestamp 1688980957
transform 1 0 1748 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W2BEGb2
timestamp 1688980957
transform 1 0 4140 0 1 6528
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W2BEGb3
timestamp 1688980957
transform 1 0 8740 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W2BEGb4
timestamp 1688980957
transform 1 0 9384 0 -1 8704
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W2BEGb5
timestamp 1688980957
transform 1 0 2024 0 -1 7616
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W2BEGb6
timestamp 1688980957
transform 1 0 2300 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W2BEGb7
timestamp 1688980957
transform 1 0 11776 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W6BEG0
timestamp 1688980957
transform 1 0 14076 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W6BEG1
timestamp 1688980957
transform 1 0 6348 0 -1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W6BEG2
timestamp 1688980957
transform 1 0 6348 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W6BEG3
timestamp 1688980957
transform 1 0 12052 0 1 21760
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W6BEG4
timestamp 1688980957
transform 1 0 12144 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W6BEG5
timestamp 1688980957
transform 1 0 4968 0 1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W6BEG6
timestamp 1688980957
transform 1 0 4876 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W6BEG7
timestamp 1688980957
transform 1 0 12052 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W6BEG8
timestamp 1688980957
transform 1 0 9476 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W6BEG9
timestamp 1688980957
transform 1 0 3772 0 -1 18496
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W6BEG10
timestamp 1688980957
transform 1 0 4048 0 1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_W6BEG11
timestamp 1688980957
transform 1 0 14076 0 1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_WW4BEG0
timestamp 1688980957
transform 1 0 11132 0 1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_WW4BEG1
timestamp 1688980957
transform 1 0 6624 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_WW4BEG2
timestamp 1688980957
transform 1 0 3772 0 1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_WW4BEG3
timestamp 1688980957
transform 1 0 12052 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_WW4BEG4
timestamp 1688980957
transform 1 0 9844 0 1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_WW4BEG5
timestamp 1688980957
transform 1 0 2208 0 -1 16320
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_WW4BEG6
timestamp 1688980957
transform 1 0 4324 0 -1 10880
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_WW4BEG7
timestamp 1688980957
transform 1 0 12420 0 -1 11968
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_WW4BEG8
timestamp 1688980957
transform 1 0 9844 0 1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_WW4BEG9
timestamp 1688980957
transform 1 0 3772 0 -1 17408
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_WW4BEG10
timestamp 1688980957
transform 1 0 4324 0 -1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_WW4BEG11
timestamp 1688980957
transform 1 0 11684 0 1 9792
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_WW4BEG12
timestamp 1688980957
transform 1 0 8832 0 -1 14144
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_WW4BEG13
timestamp 1688980957
transform 1 0 2300 0 -1 13056
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_WW4BEG14
timestamp 1688980957
transform 1 0 2944 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux41_buf_WW4BEG15
timestamp 1688980957
transform 1 0 13708 0 -1 15232
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_2  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG0.cus_mux21_inst._2_
timestamp 1688980957
transform 1 0 14076 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG0.cus_mux21_inst._3_
timestamp 1688980957
transform 1 0 14536 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG0.cus_mux21_inst._4_
timestamp 1688980957
transform 1 0 14076 0 1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG0.cus_mux21_inst.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 14720 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG0.cus_mux21_inst.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 14628 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG0.cus_mux41_buf_inst0
timestamp 1688980957
transform 1 0 12880 0 -1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG0.cus_mux41_buf_inst1
timestamp 1688980957
transform 1 0 12880 0 -1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_2  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG1.cus_mux21_inst._2_
timestamp 1688980957
transform 1 0 6900 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG1.cus_mux21_inst._3_
timestamp 1688980957
transform 1 0 7176 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG1.cus_mux21_inst._4_
timestamp 1688980957
transform 1 0 7728 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG1.cus_mux21_inst.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 6348 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG1.cus_mux21_inst.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 6992 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG1.cus_mux41_buf_inst0
timestamp 1688980957
transform 1 0 3680 0 -1 32640
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG1.cus_mux41_buf_inst1
timestamp 1688980957
transform 1 0 4968 0 1 31552
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_2  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG2.cus_mux21_inst._2_
timestamp 1688980957
transform 1 0 8004 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG2.cus_mux21_inst._3_
timestamp 1688980957
transform 1 0 9660 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG2.cus_mux21_inst._4_
timestamp 1688980957
transform 1 0 8924 0 1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG2.cus_mux21_inst.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 6348 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG2.cus_mux21_inst.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 7728 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG2.cus_mux41_buf_inst0
timestamp 1688980957
transform 1 0 5336 0 1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG2.cus_mux41_buf_inst1
timestamp 1688980957
transform 1 0 5704 0 1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_2  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG3.cus_mux21_inst._2_
timestamp 1688980957
transform 1 0 12144 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG3.cus_mux21_inst._3_
timestamp 1688980957
transform 1 0 12880 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG3.cus_mux21_inst._4_
timestamp 1688980957
transform 1 0 11684 0 1 30464
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG3.cus_mux21_inst.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 12420 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG3.cus_mux21_inst.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 12696 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG3.cus_mux41_buf_inst0
timestamp 1688980957
transform 1 0 11500 0 -1 30464
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG3.cus_mux41_buf_inst1
timestamp 1688980957
transform 1 0 11132 0 1 29376
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_2  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG0.cus_mux21_inst._2_
timestamp 1688980957
transform 1 0 15272 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG0.cus_mux21_inst._3_
timestamp 1688980957
transform 1 0 16100 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG0.cus_mux21_inst._4_
timestamp 1688980957
transform 1 0 15732 0 -1 19584
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG0.cus_mux21_inst.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 15824 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG0.cus_mux21_inst.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 16100 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG0.cus_mux41_buf_inst0
timestamp 1688980957
transform 1 0 14076 0 1 19584
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG0.cus_mux41_buf_inst1
timestamp 1688980957
transform 1 0 13064 0 -1 20672
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_2  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG1.cus_mux21_inst._2_
timestamp 1688980957
transform 1 0 7360 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG1.cus_mux21_inst._3_
timestamp 1688980957
transform 1 0 7912 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_4  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG1.cus_mux21_inst._4_
timestamp 1688980957
transform 1 0 8188 0 -1 22848
box -38 -48 1234 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG1.cus_mux21_inst.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 6808 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG1.cus_mux21_inst.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 7176 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG1.cus_mux41_buf_inst0
timestamp 1688980957
transform 1 0 4692 0 1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG1.cus_mux41_buf_inst1
timestamp 1688980957
transform 1 0 5244 0 1 22848
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_2  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG2.cus_mux21_inst._2_
timestamp 1688980957
transform 1 0 10488 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG2.cus_mux21_inst._3_
timestamp 1688980957
transform 1 0 11500 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG2.cus_mux21_inst._4_
timestamp 1688980957
transform 1 0 10764 0 -1 23936
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG2.cus_mux21_inst.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 9844 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG2.cus_mux21_inst.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 10212 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG2.cus_mux41_buf_inst0
timestamp 1688980957
transform 1 0 7636 0 -1 25024
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG2.cus_mux41_buf_inst1
timestamp 1688980957
transform 1 0 7728 0 -1 23936
box -38 -48 1970 592
use sky130_fd_sc_hd__inv_2  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG3.cus_mux21_inst._2_
timestamp 1688980957
transform 1 0 16192 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG3.cus_mux21_inst._3_
timestamp 1688980957
transform 1 0 16192 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__o21ai_2  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG3.cus_mux21_inst._4_
timestamp 1688980957
transform 1 0 15456 0 -1 26112
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG3.cus_mux21_inst.break_comb_loop_inst0._0_
timestamp 1688980957
transform 1 0 15916 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG3.cus_mux21_inst.break_comb_loop_inst1._0_
timestamp 1688980957
transform 1 0 15640 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG3.cus_mux41_buf_inst0
timestamp 1688980957
transform 1 0 14076 0 1 26112
box -38 -48 1970 592
use sky130_fd_sc_hd__mux4_1  Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG3.cus_mux41_buf_inst1
timestamp 1688980957
transform 1 0 13708 0 -1 27200
box -38 -48 1970 592
use sky130_fd_sc_hd__clkbuf_1  N4BEG_outbuf_0._0_
timestamp 1688980957
transform 1 0 6348 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  N4BEG_outbuf_1._0_
timestamp 1688980957
transform 1 0 6808 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  N4BEG_outbuf_2._0_
timestamp 1688980957
transform 1 0 5152 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  N4BEG_outbuf_3._0_
timestamp 1688980957
transform 1 0 8096 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  N4BEG_outbuf_4._0_
timestamp 1688980957
transform 1 0 6992 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  N4BEG_outbuf_5._0_
timestamp 1688980957
transform 1 0 5980 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  N4BEG_outbuf_6._0_
timestamp 1688980957
transform 1 0 7084 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  N4BEG_outbuf_7._0_
timestamp 1688980957
transform 1 0 7176 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  N4BEG_outbuf_8._0_
timestamp 1688980957
transform 1 0 9476 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  N4BEG_outbuf_9._0_
timestamp 1688980957
transform 1 0 8924 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  N4BEG_outbuf_10._0_
timestamp 1688980957
transform 1 0 9200 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  N4BEG_outbuf_11._0_
timestamp 1688980957
transform 1 0 8924 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  N4END_inbuf_0._0_
timestamp 1688980957
transform 1 0 6808 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  N4END_inbuf_1._0_
timestamp 1688980957
transform 1 0 6624 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  N4END_inbuf_2._0_
timestamp 1688980957
transform 1 0 7360 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  N4END_inbuf_3._0_
timestamp 1688980957
transform 1 0 6992 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  N4END_inbuf_4._0_
timestamp 1688980957
transform 1 0 7728 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  N4END_inbuf_5._0_
timestamp 1688980957
transform 1 0 7360 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  N4END_inbuf_6._0_
timestamp 1688980957
transform 1 0 8096 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  N4END_inbuf_7._0_
timestamp 1688980957
transform 1 0 7728 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  N4END_inbuf_8._0_
timestamp 1688980957
transform 1 0 8464 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  N4END_inbuf_9._0_
timestamp 1688980957
transform 1 0 8096 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  N4END_inbuf_10._0_
timestamp 1688980957
transform 1 0 8464 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  N4END_inbuf_11._0_
timestamp 1688980957
transform 1 0 8832 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output189
timestamp 1688980957
transform 1 0 21252 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output190
timestamp 1688980957
transform 1 0 21068 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output191
timestamp 1688980957
transform 1 0 20700 0 1 9792
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output192
timestamp 1688980957
transform 1 0 21068 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output193
timestamp 1688980957
transform 1 0 21252 0 -1 16320
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output194
timestamp 1688980957
transform 1 0 21068 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output195
timestamp 1688980957
transform 1 0 21252 0 -1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output196
timestamp 1688980957
transform 1 0 21252 0 1 17408
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output197
timestamp 1688980957
transform 1 0 21068 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output198
timestamp 1688980957
transform 1 0 21252 0 1 14144
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output199
timestamp 1688980957
transform 1 0 21252 0 -1 15232
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output200
timestamp 1688980957
transform 1 0 21068 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output201
timestamp 1688980957
transform 1 0 20884 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output202
timestamp 1688980957
transform 1 0 20516 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output203
timestamp 1688980957
transform 1 0 20700 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output204
timestamp 1688980957
transform 1 0 21252 0 1 11968
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output205
timestamp 1688980957
transform 1 0 21068 0 -1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output206
timestamp 1688980957
transform 1 0 21068 0 1 25024
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output207
timestamp 1688980957
transform 1 0 21252 0 -1 26112
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output208
timestamp 1688980957
transform 1 0 21068 0 1 26112
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output209
timestamp 1688980957
transform 1 0 21252 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output210
timestamp 1688980957
transform 1 0 20884 0 -1 22848
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output211
timestamp 1688980957
transform 1 0 21068 0 1 22848
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output212
timestamp 1688980957
transform 1 0 21252 0 1 23936
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output213
timestamp 1688980957
transform 1 0 21252 0 -1 20672
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output214
timestamp 1688980957
transform 1 0 20884 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output215
timestamp 1688980957
transform 1 0 20332 0 1 20672
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output216
timestamp 1688980957
transform 1 0 20884 0 1 21760
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output217
timestamp 1688980957
transform 1 0 21068 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output218
timestamp 1688980957
transform 1 0 21252 0 1 18496
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output219
timestamp 1688980957
transform 1 0 21068 0 -1 19584
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output220
timestamp 1688980957
transform 1 0 21252 0 1 19584
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output221
timestamp 1688980957
transform 1 0 21252 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output222
timestamp 1688980957
transform 1 0 21252 0 -1 32640
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output223
timestamp 1688980957
transform 1 0 20332 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output224
timestamp 1688980957
transform 1 0 20884 0 -1 33728
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output225
timestamp 1688980957
transform 1 0 21252 0 1 33728
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output226
timestamp 1688980957
transform 1 0 21068 0 -1 34816
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output227
timestamp 1688980957
transform 1 0 21252 0 1 34816
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output228
timestamp 1688980957
transform 1 0 21252 0 -1 35904
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output229
timestamp 1688980957
transform 1 0 21068 0 1 35904
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output230
timestamp 1688980957
transform 1 0 21252 0 -1 36992
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output231
timestamp 1688980957
transform 1 0 21068 0 1 36992
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output232
timestamp 1688980957
transform 1 0 20884 0 1 27200
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output233
timestamp 1688980957
transform 1 0 21252 0 -1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output234
timestamp 1688980957
transform 1 0 21252 0 1 38080
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output235
timestamp 1688980957
transform 1 0 21068 0 -1 39168
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output236
timestamp 1688980957
transform 1 0 21252 0 1 39168
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output237
timestamp 1688980957
transform 1 0 21068 0 -1 40256
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output238
timestamp 1688980957
transform 1 0 21252 0 1 40256
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output239
timestamp 1688980957
transform 1 0 21252 0 -1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output240
timestamp 1688980957
transform 1 0 21068 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output241
timestamp 1688980957
transform 1 0 20700 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output242
timestamp 1688980957
transform 1 0 19964 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output243
timestamp 1688980957
transform 1 0 20884 0 -1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output244
timestamp 1688980957
transform 1 0 20332 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output245
timestamp 1688980957
transform 1 0 20884 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output246
timestamp 1688980957
transform 1 0 21252 0 1 28288
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output247
timestamp 1688980957
transform 1 0 21068 0 -1 29376
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output248
timestamp 1688980957
transform 1 0 21252 0 1 29376
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output249
timestamp 1688980957
transform 1 0 21068 0 -1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output250
timestamp 1688980957
transform 1 0 21068 0 1 30464
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output251
timestamp 1688980957
transform 1 0 21252 0 -1 31552
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output252
timestamp 1688980957
transform 1 0 21068 0 1 31552
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output253
timestamp 1688980957
transform 1 0 16652 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output254
timestamp 1688980957
transform 1 0 19228 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output255
timestamp 1688980957
transform 1 0 19228 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output256
timestamp 1688980957
transform 1 0 19780 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output257
timestamp 1688980957
transform 1 0 19780 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output258
timestamp 1688980957
transform 1 0 20332 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output259
timestamp 1688980957
transform 1 0 19412 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output260
timestamp 1688980957
transform 1 0 20884 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output261
timestamp 1688980957
transform 1 0 20332 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output262
timestamp 1688980957
transform 1 0 20332 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output263
timestamp 1688980957
transform 1 0 20884 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output264
timestamp 1688980957
transform 1 0 17204 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output265
timestamp 1688980957
transform 1 0 17572 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output266
timestamp 1688980957
transform 1 0 17756 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output267
timestamp 1688980957
transform 1 0 17020 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output268
timestamp 1688980957
transform 1 0 17940 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output269
timestamp 1688980957
transform 1 0 17572 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output270
timestamp 1688980957
transform 1 0 18492 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output271
timestamp 1688980957
transform 1 0 18124 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output272
timestamp 1688980957
transform 1 0 18124 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output273
timestamp 1688980957
transform 1 0 2024 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output274
timestamp 1688980957
transform 1 0 2944 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output275
timestamp 1688980957
transform 1 0 2576 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output276
timestamp 1688980957
transform 1 0 2392 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output277
timestamp 1688980957
transform 1 0 3128 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output278
timestamp 1688980957
transform 1 0 2024 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output279
timestamp 1688980957
transform 1 0 3312 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output280
timestamp 1688980957
transform 1 0 3772 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output281
timestamp 1688980957
transform 1 0 4324 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output282
timestamp 1688980957
transform 1 0 3864 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output283
timestamp 1688980957
transform 1 0 4876 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output284
timestamp 1688980957
transform 1 0 4416 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output285
timestamp 1688980957
transform 1 0 3772 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output286
timestamp 1688980957
transform 1 0 5060 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output287
timestamp 1688980957
transform 1 0 4508 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output288
timestamp 1688980957
transform 1 0 5428 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output289
timestamp 1688980957
transform 1 0 5612 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output290
timestamp 1688980957
transform 1 0 4968 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output291
timestamp 1688980957
transform 1 0 4140 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output292
timestamp 1688980957
transform 1 0 5520 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output293
timestamp 1688980957
transform 1 0 6348 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output294
timestamp 1688980957
transform 1 0 7360 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output295
timestamp 1688980957
transform 1 0 7912 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output296
timestamp 1688980957
transform 1 0 8280 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output297
timestamp 1688980957
transform 1 0 8464 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output298
timestamp 1688980957
transform 1 0 9292 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output299
timestamp 1688980957
transform 1 0 8924 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output300
timestamp 1688980957
transform 1 0 6072 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output301
timestamp 1688980957
transform 1 0 6624 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output302
timestamp 1688980957
transform 1 0 7268 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output303
timestamp 1688980957
transform 1 0 6440 0 -1 43520
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output304
timestamp 1688980957
transform 1 0 7176 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output305
timestamp 1688980957
transform 1 0 6900 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output306
timestamp 1688980957
transform 1 0 8004 0 1 41344
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output307
timestamp 1688980957
transform 1 0 6992 0 -1 43520
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output308
timestamp 1688980957
transform 1 0 7728 0 1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output309
timestamp 1688980957
transform 1 0 9200 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output310
timestamp 1688980957
transform 1 0 9844 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output311
timestamp 1688980957
transform 1 0 8280 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output312
timestamp 1688980957
transform 1 0 9752 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output313
timestamp 1688980957
transform 1 0 11500 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output314
timestamp 1688980957
transform 1 0 12052 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output315
timestamp 1688980957
transform 1 0 11868 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output316
timestamp 1688980957
transform 1 0 12236 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output317
timestamp 1688980957
transform 1 0 12788 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output318
timestamp 1688980957
transform 1 0 13156 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output319
timestamp 1688980957
transform 1 0 13524 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output320
timestamp 1688980957
transform 1 0 13156 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output321
timestamp 1688980957
transform 1 0 9568 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output322
timestamp 1688980957
transform 1 0 10304 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output323
timestamp 1688980957
transform 1 0 8924 0 1 1088
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output324
timestamp 1688980957
transform 1 0 10856 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output325
timestamp 1688980957
transform 1 0 9292 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output326
timestamp 1688980957
transform 1 0 10672 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output327
timestamp 1688980957
transform 1 0 11040 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output328
timestamp 1688980957
transform 1 0 11500 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output329
timestamp 1688980957
transform 1 0 14076 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output330
timestamp 1688980957
transform 1 0 15548 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output331
timestamp 1688980957
transform 1 0 15916 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output332
timestamp 1688980957
transform 1 0 15364 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output333
timestamp 1688980957
transform 1 0 16468 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output334
timestamp 1688980957
transform 1 0 16652 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output335
timestamp 1688980957
transform 1 0 17204 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output336
timestamp 1688980957
transform 1 0 13708 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output337
timestamp 1688980957
transform 1 0 14628 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output338
timestamp 1688980957
transform 1 0 14260 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_2  output339
timestamp 1688980957
transform 1 0 14812 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output340
timestamp 1688980957
transform 1 0 14812 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output341
timestamp 1688980957
transform 1 0 16652 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output342
timestamp 1688980957
transform 1 0 15364 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output343
timestamp 1688980957
transform 1 0 15916 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output344
timestamp 1688980957
transform 1 0 15916 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__buf_1  output345
timestamp 1688980957
transform 1 0 18860 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_4  output346
timestamp 1688980957
transform 1 0 3128 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output347
timestamp 1688980957
transform 1 0 3772 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output348
timestamp 1688980957
transform 1 0 4416 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output349
timestamp 1688980957
transform 1 0 5152 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output350
timestamp 1688980957
transform 1 0 2484 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output351
timestamp 1688980957
transform 1 0 2484 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output352
timestamp 1688980957
transform 1 0 3128 0 1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output353
timestamp 1688980957
transform 1 0 5704 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output354
timestamp 1688980957
transform 1 0 1380 0 1 1088
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output355
timestamp 1688980957
transform 1 0 3772 0 -1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output356
timestamp 1688980957
transform 1 0 5980 0 1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output357
timestamp 1688980957
transform 1 0 1932 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output358
timestamp 1688980957
transform 1 0 1932 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output359
timestamp 1688980957
transform 1 0 6348 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output360
timestamp 1688980957
transform 1 0 6900 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output361
timestamp 1688980957
transform 1 0 5612 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output362
timestamp 1688980957
transform 1 0 1380 0 -1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output363
timestamp 1688980957
transform 1 0 4232 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output364
timestamp 1688980957
transform 1 0 1380 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output365
timestamp 1688980957
transform 1 0 1748 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output366
timestamp 1688980957
transform 1 0 1656 0 -1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output367
timestamp 1688980957
transform 1 0 1380 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output368
timestamp 1688980957
transform 1 0 1380 0 -1 18496
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output369
timestamp 1688980957
transform 1 0 1564 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output370
timestamp 1688980957
transform 1 0 6348 0 -1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output371
timestamp 1688980957
transform 1 0 1564 0 -1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output372
timestamp 1688980957
transform 1 0 1380 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output373
timestamp 1688980957
transform 1 0 1564 0 1 13056
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output374
timestamp 1688980957
transform 1 0 3772 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output375
timestamp 1688980957
transform 1 0 4324 0 1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output376
timestamp 1688980957
transform 1 0 1564 0 1 14144
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output377
timestamp 1688980957
transform 1 0 4140 0 -1 16320
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output378
timestamp 1688980957
transform 1 0 6348 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output379
timestamp 1688980957
transform 1 0 1380 0 -1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output380
timestamp 1688980957
transform 1 0 4140 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output381
timestamp 1688980957
transform 1 0 1380 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output382
timestamp 1688980957
transform 1 0 3128 0 1 15232
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output383
timestamp 1688980957
transform 1 0 1564 0 -1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output384
timestamp 1688980957
transform 1 0 1380 0 -1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output385
timestamp 1688980957
transform 1 0 3772 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output386
timestamp 1688980957
transform 1 0 4232 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output387
timestamp 1688980957
transform 1 0 1380 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output388
timestamp 1688980957
transform 1 0 4324 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output389
timestamp 1688980957
transform 1 0 1472 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output390
timestamp 1688980957
transform 1 0 6808 0 1 10880
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output391
timestamp 1688980957
transform 1 0 4140 0 1 11968
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output392
timestamp 1688980957
transform 1 0 1380 0 1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_4  output393
timestamp 1688980957
transform 1 0 1748 0 1 9792
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1688980957
transform 1 0 1104 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1688980957
transform -1 0 21896 0 1 1088
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1688980957
transform 1 0 1104 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1688980957
transform -1 0 21896 0 -1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1688980957
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1688980957
transform -1 0 21896 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1688980957
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1688980957
transform -1 0 21896 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1688980957
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1688980957
transform -1 0 21896 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1688980957
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1688980957
transform -1 0 21896 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1688980957
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1688980957
transform -1 0 21896 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1688980957
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1688980957
transform -1 0 21896 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1688980957
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1688980957
transform -1 0 21896 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1688980957
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1688980957
transform -1 0 21896 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1688980957
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1688980957
transform -1 0 21896 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1688980957
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1688980957
transform -1 0 21896 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1688980957
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1688980957
transform -1 0 21896 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1688980957
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1688980957
transform -1 0 21896 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1688980957
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1688980957
transform -1 0 21896 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1688980957
transform 1 0 1104 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1688980957
transform -1 0 21896 0 -1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1688980957
transform 1 0 1104 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1688980957
transform -1 0 21896 0 1 9792
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1688980957
transform 1 0 1104 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1688980957
transform -1 0 21896 0 -1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1688980957
transform 1 0 1104 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1688980957
transform -1 0 21896 0 1 10880
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1688980957
transform 1 0 1104 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1688980957
transform -1 0 21896 0 -1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1688980957
transform 1 0 1104 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1688980957
transform -1 0 21896 0 1 11968
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1688980957
transform 1 0 1104 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1688980957
transform -1 0 21896 0 -1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1688980957
transform 1 0 1104 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1688980957
transform -1 0 21896 0 1 13056
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1688980957
transform 1 0 1104 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1688980957
transform -1 0 21896 0 -1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1688980957
transform 1 0 1104 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1688980957
transform -1 0 21896 0 1 14144
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1688980957
transform 1 0 1104 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1688980957
transform -1 0 21896 0 -1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1688980957
transform 1 0 1104 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1688980957
transform -1 0 21896 0 1 15232
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1688980957
transform 1 0 1104 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1688980957
transform -1 0 21896 0 -1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1688980957
transform 1 0 1104 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1688980957
transform -1 0 21896 0 1 16320
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1688980957
transform 1 0 1104 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1688980957
transform -1 0 21896 0 -1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1688980957
transform 1 0 1104 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1688980957
transform -1 0 21896 0 1 17408
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1688980957
transform 1 0 1104 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1688980957
transform -1 0 21896 0 -1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1688980957
transform 1 0 1104 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1688980957
transform -1 0 21896 0 1 18496
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1688980957
transform 1 0 1104 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1688980957
transform -1 0 21896 0 -1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1688980957
transform 1 0 1104 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1688980957
transform -1 0 21896 0 1 19584
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_70
timestamp 1688980957
transform 1 0 1104 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_71
timestamp 1688980957
transform -1 0 21896 0 -1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_72
timestamp 1688980957
transform 1 0 1104 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_73
timestamp 1688980957
transform -1 0 21896 0 1 20672
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_74
timestamp 1688980957
transform 1 0 1104 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_75
timestamp 1688980957
transform -1 0 21896 0 -1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_76
timestamp 1688980957
transform 1 0 1104 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_77
timestamp 1688980957
transform -1 0 21896 0 1 21760
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_78
timestamp 1688980957
transform 1 0 1104 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_79
timestamp 1688980957
transform -1 0 21896 0 -1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_80
timestamp 1688980957
transform 1 0 1104 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_81
timestamp 1688980957
transform -1 0 21896 0 1 22848
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_82
timestamp 1688980957
transform 1 0 1104 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_83
timestamp 1688980957
transform -1 0 21896 0 -1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_84
timestamp 1688980957
transform 1 0 1104 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_85
timestamp 1688980957
transform -1 0 21896 0 1 23936
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_86
timestamp 1688980957
transform 1 0 1104 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_87
timestamp 1688980957
transform -1 0 21896 0 -1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_88
timestamp 1688980957
transform 1 0 1104 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_89
timestamp 1688980957
transform -1 0 21896 0 1 25024
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_90
timestamp 1688980957
transform 1 0 1104 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_91
timestamp 1688980957
transform -1 0 21896 0 -1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_92
timestamp 1688980957
transform 1 0 1104 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_93
timestamp 1688980957
transform -1 0 21896 0 1 26112
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_94
timestamp 1688980957
transform 1 0 1104 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_95
timestamp 1688980957
transform -1 0 21896 0 -1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_96
timestamp 1688980957
transform 1 0 1104 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_97
timestamp 1688980957
transform -1 0 21896 0 1 27200
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_98
timestamp 1688980957
transform 1 0 1104 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_99
timestamp 1688980957
transform -1 0 21896 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_100
timestamp 1688980957
transform 1 0 1104 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_101
timestamp 1688980957
transform -1 0 21896 0 1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_102
timestamp 1688980957
transform 1 0 1104 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_103
timestamp 1688980957
transform -1 0 21896 0 -1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_104
timestamp 1688980957
transform 1 0 1104 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_105
timestamp 1688980957
transform -1 0 21896 0 1 29376
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_106
timestamp 1688980957
transform 1 0 1104 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_107
timestamp 1688980957
transform -1 0 21896 0 -1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_108
timestamp 1688980957
transform 1 0 1104 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_109
timestamp 1688980957
transform -1 0 21896 0 1 30464
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_110
timestamp 1688980957
transform 1 0 1104 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_111
timestamp 1688980957
transform -1 0 21896 0 -1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_112
timestamp 1688980957
transform 1 0 1104 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_113
timestamp 1688980957
transform -1 0 21896 0 1 31552
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_114
timestamp 1688980957
transform 1 0 1104 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_115
timestamp 1688980957
transform -1 0 21896 0 -1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_116
timestamp 1688980957
transform 1 0 1104 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_117
timestamp 1688980957
transform -1 0 21896 0 1 32640
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_118
timestamp 1688980957
transform 1 0 1104 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_119
timestamp 1688980957
transform -1 0 21896 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_120
timestamp 1688980957
transform 1 0 1104 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_121
timestamp 1688980957
transform -1 0 21896 0 1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_122
timestamp 1688980957
transform 1 0 1104 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_123
timestamp 1688980957
transform -1 0 21896 0 -1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_124
timestamp 1688980957
transform 1 0 1104 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_125
timestamp 1688980957
transform -1 0 21896 0 1 34816
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_126
timestamp 1688980957
transform 1 0 1104 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_127
timestamp 1688980957
transform -1 0 21896 0 -1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_128
timestamp 1688980957
transform 1 0 1104 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_129
timestamp 1688980957
transform -1 0 21896 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_130
timestamp 1688980957
transform 1 0 1104 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_131
timestamp 1688980957
transform -1 0 21896 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_132
timestamp 1688980957
transform 1 0 1104 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_133
timestamp 1688980957
transform -1 0 21896 0 1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_134
timestamp 1688980957
transform 1 0 1104 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_135
timestamp 1688980957
transform -1 0 21896 0 -1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_136
timestamp 1688980957
transform 1 0 1104 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_137
timestamp 1688980957
transform -1 0 21896 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_138
timestamp 1688980957
transform 1 0 1104 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_139
timestamp 1688980957
transform -1 0 21896 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_140
timestamp 1688980957
transform 1 0 1104 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_141
timestamp 1688980957
transform -1 0 21896 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_142
timestamp 1688980957
transform 1 0 1104 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_143
timestamp 1688980957
transform -1 0 21896 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_144
timestamp 1688980957
transform 1 0 1104 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_145
timestamp 1688980957
transform -1 0 21896 0 1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_146
timestamp 1688980957
transform 1 0 1104 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_147
timestamp 1688980957
transform -1 0 21896 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_148
timestamp 1688980957
transform 1 0 1104 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_149
timestamp 1688980957
transform -1 0 21896 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_150
timestamp 1688980957
transform 1 0 1104 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_151
timestamp 1688980957
transform -1 0 21896 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_152
timestamp 1688980957
transform 1 0 1104 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_153
timestamp 1688980957
transform -1 0 21896 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_154
timestamp 1688980957
transform 1 0 1104 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_155
timestamp 1688980957
transform -1 0 21896 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  S4BEG_outbuf_0._0_
timestamp 1688980957
transform 1 0 13524 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  S4BEG_outbuf_1._0_
timestamp 1688980957
transform 1 0 14628 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  S4BEG_outbuf_2._0_
timestamp 1688980957
transform 1 0 14076 0 -1 42432
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_2  S4BEG_outbuf_3._0_
timestamp 1688980957
transform 1 0 14996 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  S4BEG_outbuf_4._0_
timestamp 1688980957
transform 1 0 15364 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  S4BEG_outbuf_5._0_
timestamp 1688980957
transform 1 0 14444 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  S4BEG_outbuf_6._0_
timestamp 1688980957
transform 1 0 15732 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  S4BEG_outbuf_7._0_
timestamp 1688980957
transform 1 0 14812 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  S4BEG_outbuf_8._0_
timestamp 1688980957
transform 1 0 16100 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  S4BEG_outbuf_9._0_
timestamp 1688980957
transform 1 0 15180 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  S4BEG_outbuf_10._0_
timestamp 1688980957
transform 1 0 16652 0 -1 42432
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  S4BEG_outbuf_11._0_
timestamp 1688980957
transform 1 0 15548 0 1 41344
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  S4END_inbuf_0._0_
timestamp 1688980957
transform 1 0 14444 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  S4END_inbuf_1._0_
timestamp 1688980957
transform 1 0 12880 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  S4END_inbuf_2._0_
timestamp 1688980957
transform 1 0 14720 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  S4END_inbuf_3._0_
timestamp 1688980957
transform 1 0 14812 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  S4END_inbuf_4._0_
timestamp 1688980957
transform 1 0 15088 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  S4END_inbuf_5._0_
timestamp 1688980957
transform 1 0 15364 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  S4END_inbuf_6._0_
timestamp 1688980957
transform 1 0 15916 0 -1 43520
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  S4END_inbuf_7._0_
timestamp 1688980957
transform 1 0 18676 0 1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  S4END_inbuf_8._0_
timestamp 1688980957
transform 1 0 15916 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  S4END_inbuf_9._0_
timestamp 1688980957
transform 1 0 17020 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  S4END_inbuf_10._0_
timestamp 1688980957
transform 1 0 16192 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  S4END_inbuf_11._0_
timestamp 1688980957
transform 1 0 17296 0 -1 42432
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_0._0_
timestamp 1688980957
transform 1 0 15640 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_1._0_
timestamp 1688980957
transform 1 0 15916 0 1 35904
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_2._0_
timestamp 1688980957
transform 1 0 16100 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_3._0_
timestamp 1688980957
transform 1 0 16284 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_4._0_
timestamp 1688980957
transform 1 0 16652 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__dlymetal6s2s_1  strobe_inbuf_5._0_
timestamp 1688980957
transform 1 0 17112 0 1 18496
box -38 -48 958 592
use sky130_fd_sc_hd__buf_1  strobe_inbuf_6._0_
timestamp 1688980957
transform 1 0 16836 0 -1 28288
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_7._0_
timestamp 1688980957
transform 1 0 17020 0 -1 33728
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_8._0_
timestamp 1688980957
transform 1 0 17388 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_inbuf_9._0_
timestamp 1688980957
transform 1 0 17296 0 1 38080
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  strobe_inbuf_10._0_
timestamp 1688980957
transform 1 0 17664 0 -1 13056
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  strobe_inbuf_11._0_
timestamp 1688980957
transform 1 0 21068 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  strobe_inbuf_12._0_
timestamp 1688980957
transform 1 0 18768 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  strobe_inbuf_13._0_
timestamp 1688980957
transform 1 0 20976 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  strobe_inbuf_14._0_
timestamp 1688980957
transform 1 0 20240 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  strobe_inbuf_15._0_
timestamp 1688980957
transform 1 0 20700 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  strobe_inbuf_16._0_
timestamp 1688980957
transform 1 0 20608 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  strobe_inbuf_17._0_
timestamp 1688980957
transform 1 0 21068 0 1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  strobe_inbuf_18._0_
timestamp 1688980957
transform 1 0 20700 0 -1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  strobe_inbuf_19._0_
timestamp 1688980957
transform 1 0 19872 0 -1 3264
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_0._0_
timestamp 1688980957
transform 1 0 15916 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_1._0_
timestamp 1688980957
transform 1 0 16192 0 -1 36992
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_2._0_
timestamp 1688980957
transform 1 0 16468 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_3._0_
timestamp 1688980957
transform 1 0 16744 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_4._0_
timestamp 1688980957
transform 1 0 17020 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_5._0_
timestamp 1688980957
transform 1 0 17296 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_6._0_
timestamp 1688980957
transform 1 0 17572 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_7._0_
timestamp 1688980957
transform 1 0 18124 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_8._0_
timestamp 1688980957
transform 1 0 17480 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_9._0_
timestamp 1688980957
transform 1 0 17664 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_10._0_
timestamp 1688980957
transform 1 0 18400 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_11._0_
timestamp 1688980957
transform 1 0 19228 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_12._0_
timestamp 1688980957
transform 1 0 20056 0 1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_13._0_
timestamp 1688980957
transform 1 0 20516 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_14._0_
timestamp 1688980957
transform 1 0 18860 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_15._0_
timestamp 1688980957
transform 1 0 19780 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_16._0_
timestamp 1688980957
transform 1 0 20056 0 -1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_17._0_
timestamp 1688980957
transform 1 0 19688 0 -1 41344
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_18._0_
timestamp 1688980957
transform 1 0 18584 0 -1 40256
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  strobe_outbuf_19._0_
timestamp 1688980957
transform 1 0 18860 0 1 39168
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_156 dependencies/pdks/sky130A/libs.ref/sky130_fd_sc_hd/mag
timestamp 1688980957
transform 1 0 3680 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_157
timestamp 1688980957
transform 1 0 6256 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_158
timestamp 1688980957
transform 1 0 8832 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_159
timestamp 1688980957
transform 1 0 11408 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_160
timestamp 1688980957
transform 1 0 13984 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_161
timestamp 1688980957
transform 1 0 16560 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_162
timestamp 1688980957
transform 1 0 19136 0 1 1088
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_163
timestamp 1688980957
transform 1 0 6256 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_164
timestamp 1688980957
transform 1 0 11408 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_165
timestamp 1688980957
transform 1 0 16560 0 -1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_166
timestamp 1688980957
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_167
timestamp 1688980957
transform 1 0 8832 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_168
timestamp 1688980957
transform 1 0 13984 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_169
timestamp 1688980957
transform 1 0 19136 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_170
timestamp 1688980957
transform 1 0 6256 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_171
timestamp 1688980957
transform 1 0 11408 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_172
timestamp 1688980957
transform 1 0 16560 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_173
timestamp 1688980957
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_174
timestamp 1688980957
transform 1 0 8832 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_175
timestamp 1688980957
transform 1 0 13984 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_176
timestamp 1688980957
transform 1 0 19136 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_177
timestamp 1688980957
transform 1 0 6256 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_178
timestamp 1688980957
transform 1 0 11408 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_179
timestamp 1688980957
transform 1 0 16560 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_180
timestamp 1688980957
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_181
timestamp 1688980957
transform 1 0 8832 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_182
timestamp 1688980957
transform 1 0 13984 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_183
timestamp 1688980957
transform 1 0 19136 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_184
timestamp 1688980957
transform 1 0 6256 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_185
timestamp 1688980957
transform 1 0 11408 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_186
timestamp 1688980957
transform 1 0 16560 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_187
timestamp 1688980957
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_188
timestamp 1688980957
transform 1 0 8832 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_189
timestamp 1688980957
transform 1 0 13984 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_190
timestamp 1688980957
transform 1 0 19136 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_191
timestamp 1688980957
transform 1 0 6256 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_192
timestamp 1688980957
transform 1 0 11408 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_193
timestamp 1688980957
transform 1 0 16560 0 -1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_194
timestamp 1688980957
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_195
timestamp 1688980957
transform 1 0 8832 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_196
timestamp 1688980957
transform 1 0 13984 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_197
timestamp 1688980957
transform 1 0 19136 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_198
timestamp 1688980957
transform 1 0 6256 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_199
timestamp 1688980957
transform 1 0 11408 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_200
timestamp 1688980957
transform 1 0 16560 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_201
timestamp 1688980957
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_202
timestamp 1688980957
transform 1 0 8832 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_203
timestamp 1688980957
transform 1 0 13984 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_204
timestamp 1688980957
transform 1 0 19136 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_205
timestamp 1688980957
transform 1 0 6256 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_206
timestamp 1688980957
transform 1 0 11408 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_207
timestamp 1688980957
transform 1 0 16560 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_208
timestamp 1688980957
transform 1 0 3680 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_209
timestamp 1688980957
transform 1 0 8832 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_210
timestamp 1688980957
transform 1 0 13984 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_211
timestamp 1688980957
transform 1 0 19136 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_212
timestamp 1688980957
transform 1 0 6256 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_213
timestamp 1688980957
transform 1 0 11408 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_214
timestamp 1688980957
transform 1 0 16560 0 -1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_215
timestamp 1688980957
transform 1 0 3680 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_216
timestamp 1688980957
transform 1 0 8832 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_217
timestamp 1688980957
transform 1 0 13984 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_218
timestamp 1688980957
transform 1 0 19136 0 1 9792
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_219
timestamp 1688980957
transform 1 0 6256 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_220
timestamp 1688980957
transform 1 0 11408 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_221
timestamp 1688980957
transform 1 0 16560 0 -1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_222
timestamp 1688980957
transform 1 0 3680 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_223
timestamp 1688980957
transform 1 0 8832 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_224
timestamp 1688980957
transform 1 0 13984 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_225
timestamp 1688980957
transform 1 0 19136 0 1 10880
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_226
timestamp 1688980957
transform 1 0 6256 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_227
timestamp 1688980957
transform 1 0 11408 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_228
timestamp 1688980957
transform 1 0 16560 0 -1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_229
timestamp 1688980957
transform 1 0 3680 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_230
timestamp 1688980957
transform 1 0 8832 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_231
timestamp 1688980957
transform 1 0 13984 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_232
timestamp 1688980957
transform 1 0 19136 0 1 11968
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_233
timestamp 1688980957
transform 1 0 6256 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_234
timestamp 1688980957
transform 1 0 11408 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_235
timestamp 1688980957
transform 1 0 16560 0 -1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_236
timestamp 1688980957
transform 1 0 3680 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_237
timestamp 1688980957
transform 1 0 8832 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_238
timestamp 1688980957
transform 1 0 13984 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_239
timestamp 1688980957
transform 1 0 19136 0 1 13056
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_240
timestamp 1688980957
transform 1 0 6256 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_241
timestamp 1688980957
transform 1 0 11408 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_242
timestamp 1688980957
transform 1 0 16560 0 -1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_243
timestamp 1688980957
transform 1 0 3680 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_244
timestamp 1688980957
transform 1 0 8832 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_245
timestamp 1688980957
transform 1 0 13984 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_246
timestamp 1688980957
transform 1 0 19136 0 1 14144
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_247
timestamp 1688980957
transform 1 0 6256 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_248
timestamp 1688980957
transform 1 0 11408 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_249
timestamp 1688980957
transform 1 0 16560 0 -1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_250
timestamp 1688980957
transform 1 0 3680 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_251
timestamp 1688980957
transform 1 0 8832 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_252
timestamp 1688980957
transform 1 0 13984 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_253
timestamp 1688980957
transform 1 0 19136 0 1 15232
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_254
timestamp 1688980957
transform 1 0 6256 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_255
timestamp 1688980957
transform 1 0 11408 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_256
timestamp 1688980957
transform 1 0 16560 0 -1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_257
timestamp 1688980957
transform 1 0 3680 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_258
timestamp 1688980957
transform 1 0 8832 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_259
timestamp 1688980957
transform 1 0 13984 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_260
timestamp 1688980957
transform 1 0 19136 0 1 16320
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_261
timestamp 1688980957
transform 1 0 6256 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_262
timestamp 1688980957
transform 1 0 11408 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_263
timestamp 1688980957
transform 1 0 16560 0 -1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_264
timestamp 1688980957
transform 1 0 3680 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_265
timestamp 1688980957
transform 1 0 8832 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_266
timestamp 1688980957
transform 1 0 13984 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_267
timestamp 1688980957
transform 1 0 19136 0 1 17408
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_268
timestamp 1688980957
transform 1 0 6256 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_269
timestamp 1688980957
transform 1 0 11408 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_270
timestamp 1688980957
transform 1 0 16560 0 -1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_271
timestamp 1688980957
transform 1 0 3680 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_272
timestamp 1688980957
transform 1 0 8832 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_273
timestamp 1688980957
transform 1 0 13984 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_274
timestamp 1688980957
transform 1 0 19136 0 1 18496
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_275
timestamp 1688980957
transform 1 0 6256 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_276
timestamp 1688980957
transform 1 0 11408 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_277
timestamp 1688980957
transform 1 0 16560 0 -1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_278
timestamp 1688980957
transform 1 0 3680 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_279
timestamp 1688980957
transform 1 0 8832 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_280
timestamp 1688980957
transform 1 0 13984 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_281
timestamp 1688980957
transform 1 0 19136 0 1 19584
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_282
timestamp 1688980957
transform 1 0 6256 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_283
timestamp 1688980957
transform 1 0 11408 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_284
timestamp 1688980957
transform 1 0 16560 0 -1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_285
timestamp 1688980957
transform 1 0 3680 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_286
timestamp 1688980957
transform 1 0 8832 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_287
timestamp 1688980957
transform 1 0 13984 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_288
timestamp 1688980957
transform 1 0 19136 0 1 20672
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_289
timestamp 1688980957
transform 1 0 6256 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_290
timestamp 1688980957
transform 1 0 11408 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_291
timestamp 1688980957
transform 1 0 16560 0 -1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_292
timestamp 1688980957
transform 1 0 3680 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_293
timestamp 1688980957
transform 1 0 8832 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_294
timestamp 1688980957
transform 1 0 13984 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_295
timestamp 1688980957
transform 1 0 19136 0 1 21760
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_296
timestamp 1688980957
transform 1 0 6256 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_297
timestamp 1688980957
transform 1 0 11408 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_298
timestamp 1688980957
transform 1 0 16560 0 -1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_299
timestamp 1688980957
transform 1 0 3680 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_300
timestamp 1688980957
transform 1 0 8832 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_301
timestamp 1688980957
transform 1 0 13984 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_302
timestamp 1688980957
transform 1 0 19136 0 1 22848
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_303
timestamp 1688980957
transform 1 0 6256 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_304
timestamp 1688980957
transform 1 0 11408 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_305
timestamp 1688980957
transform 1 0 16560 0 -1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_306
timestamp 1688980957
transform 1 0 3680 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_307
timestamp 1688980957
transform 1 0 8832 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_308
timestamp 1688980957
transform 1 0 13984 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_309
timestamp 1688980957
transform 1 0 19136 0 1 23936
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_310
timestamp 1688980957
transform 1 0 6256 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_311
timestamp 1688980957
transform 1 0 11408 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_312
timestamp 1688980957
transform 1 0 16560 0 -1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_313
timestamp 1688980957
transform 1 0 3680 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_314
timestamp 1688980957
transform 1 0 8832 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_315
timestamp 1688980957
transform 1 0 13984 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_316
timestamp 1688980957
transform 1 0 19136 0 1 25024
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_317
timestamp 1688980957
transform 1 0 6256 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_318
timestamp 1688980957
transform 1 0 11408 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_319
timestamp 1688980957
transform 1 0 16560 0 -1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_320
timestamp 1688980957
transform 1 0 3680 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_321
timestamp 1688980957
transform 1 0 8832 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_322
timestamp 1688980957
transform 1 0 13984 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_323
timestamp 1688980957
transform 1 0 19136 0 1 26112
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_324
timestamp 1688980957
transform 1 0 6256 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_325
timestamp 1688980957
transform 1 0 11408 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_326
timestamp 1688980957
transform 1 0 16560 0 -1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_327
timestamp 1688980957
transform 1 0 3680 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_328
timestamp 1688980957
transform 1 0 8832 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_329
timestamp 1688980957
transform 1 0 13984 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_330
timestamp 1688980957
transform 1 0 19136 0 1 27200
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_331
timestamp 1688980957
transform 1 0 6256 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_332
timestamp 1688980957
transform 1 0 11408 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_333
timestamp 1688980957
transform 1 0 16560 0 -1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_334
timestamp 1688980957
transform 1 0 3680 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_335
timestamp 1688980957
transform 1 0 8832 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_336
timestamp 1688980957
transform 1 0 13984 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_337
timestamp 1688980957
transform 1 0 19136 0 1 28288
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_338
timestamp 1688980957
transform 1 0 6256 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_339
timestamp 1688980957
transform 1 0 11408 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_340
timestamp 1688980957
transform 1 0 16560 0 -1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_341
timestamp 1688980957
transform 1 0 3680 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_342
timestamp 1688980957
transform 1 0 8832 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_343
timestamp 1688980957
transform 1 0 13984 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_344
timestamp 1688980957
transform 1 0 19136 0 1 29376
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_345
timestamp 1688980957
transform 1 0 6256 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_346
timestamp 1688980957
transform 1 0 11408 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_347
timestamp 1688980957
transform 1 0 16560 0 -1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_348
timestamp 1688980957
transform 1 0 3680 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_349
timestamp 1688980957
transform 1 0 8832 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_350
timestamp 1688980957
transform 1 0 13984 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_351
timestamp 1688980957
transform 1 0 19136 0 1 30464
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_352
timestamp 1688980957
transform 1 0 6256 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_353
timestamp 1688980957
transform 1 0 11408 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_354
timestamp 1688980957
transform 1 0 16560 0 -1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_355
timestamp 1688980957
transform 1 0 3680 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_356
timestamp 1688980957
transform 1 0 8832 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_357
timestamp 1688980957
transform 1 0 13984 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_358
timestamp 1688980957
transform 1 0 19136 0 1 31552
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_359
timestamp 1688980957
transform 1 0 6256 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_360
timestamp 1688980957
transform 1 0 11408 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_361
timestamp 1688980957
transform 1 0 16560 0 -1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_362
timestamp 1688980957
transform 1 0 3680 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_363
timestamp 1688980957
transform 1 0 8832 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_364
timestamp 1688980957
transform 1 0 13984 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_365
timestamp 1688980957
transform 1 0 19136 0 1 32640
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_366
timestamp 1688980957
transform 1 0 6256 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_367
timestamp 1688980957
transform 1 0 11408 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_368
timestamp 1688980957
transform 1 0 16560 0 -1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_369
timestamp 1688980957
transform 1 0 3680 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_370
timestamp 1688980957
transform 1 0 8832 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_371
timestamp 1688980957
transform 1 0 13984 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_372
timestamp 1688980957
transform 1 0 19136 0 1 33728
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_373
timestamp 1688980957
transform 1 0 6256 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_374
timestamp 1688980957
transform 1 0 11408 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_375
timestamp 1688980957
transform 1 0 16560 0 -1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_376
timestamp 1688980957
transform 1 0 3680 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_377
timestamp 1688980957
transform 1 0 8832 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_378
timestamp 1688980957
transform 1 0 13984 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_379
timestamp 1688980957
transform 1 0 19136 0 1 34816
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_380
timestamp 1688980957
transform 1 0 6256 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_381
timestamp 1688980957
transform 1 0 11408 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_382
timestamp 1688980957
transform 1 0 16560 0 -1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_383
timestamp 1688980957
transform 1 0 3680 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_384
timestamp 1688980957
transform 1 0 8832 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_385
timestamp 1688980957
transform 1 0 13984 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_386
timestamp 1688980957
transform 1 0 19136 0 1 35904
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_387
timestamp 1688980957
transform 1 0 6256 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_388
timestamp 1688980957
transform 1 0 11408 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_389
timestamp 1688980957
transform 1 0 16560 0 -1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_390
timestamp 1688980957
transform 1 0 3680 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_391
timestamp 1688980957
transform 1 0 8832 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_392
timestamp 1688980957
transform 1 0 13984 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_393
timestamp 1688980957
transform 1 0 19136 0 1 36992
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_394
timestamp 1688980957
transform 1 0 6256 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_395
timestamp 1688980957
transform 1 0 11408 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_396
timestamp 1688980957
transform 1 0 16560 0 -1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_397
timestamp 1688980957
transform 1 0 3680 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_398
timestamp 1688980957
transform 1 0 8832 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_399
timestamp 1688980957
transform 1 0 13984 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_400
timestamp 1688980957
transform 1 0 19136 0 1 38080
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_401
timestamp 1688980957
transform 1 0 6256 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_402
timestamp 1688980957
transform 1 0 11408 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_403
timestamp 1688980957
transform 1 0 16560 0 -1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_404
timestamp 1688980957
transform 1 0 3680 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_405
timestamp 1688980957
transform 1 0 8832 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_406
timestamp 1688980957
transform 1 0 13984 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_407
timestamp 1688980957
transform 1 0 19136 0 1 39168
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_408
timestamp 1688980957
transform 1 0 6256 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_409
timestamp 1688980957
transform 1 0 11408 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_410
timestamp 1688980957
transform 1 0 16560 0 -1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_411
timestamp 1688980957
transform 1 0 3680 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_412
timestamp 1688980957
transform 1 0 8832 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_413
timestamp 1688980957
transform 1 0 13984 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_414
timestamp 1688980957
transform 1 0 19136 0 1 40256
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_415
timestamp 1688980957
transform 1 0 6256 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_416
timestamp 1688980957
transform 1 0 11408 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_417
timestamp 1688980957
transform 1 0 16560 0 -1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_418
timestamp 1688980957
transform 1 0 3680 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_419
timestamp 1688980957
transform 1 0 8832 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_420
timestamp 1688980957
transform 1 0 13984 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_421
timestamp 1688980957
transform 1 0 19136 0 1 41344
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_422
timestamp 1688980957
transform 1 0 6256 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_423
timestamp 1688980957
transform 1 0 11408 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_424
timestamp 1688980957
transform 1 0 16560 0 -1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_425
timestamp 1688980957
transform 1 0 3680 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_426
timestamp 1688980957
transform 1 0 8832 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_427
timestamp 1688980957
transform 1 0 13984 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_428
timestamp 1688980957
transform 1 0 19136 0 1 42432
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_429
timestamp 1688980957
transform 1 0 3680 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_430
timestamp 1688980957
transform 1 0 6256 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_431
timestamp 1688980957
transform 1 0 8832 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_432
timestamp 1688980957
transform 1 0 11408 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_433
timestamp 1688980957
transform 1 0 13984 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_434
timestamp 1688980957
transform 1 0 16560 0 -1 43520
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_435
timestamp 1688980957
transform 1 0 19136 0 -1 43520
box -38 -48 130 592
<< labels >>
flabel metal3 s 22840 9256 23300 9376 0 FreeSans 480 0 0 0 Config_accessC_bit0
port 0 nsew signal tristate
flabel metal3 s 22840 9800 23300 9920 0 FreeSans 480 0 0 0 Config_accessC_bit1
port 1 nsew signal tristate
flabel metal3 s 22840 10344 23300 10464 0 FreeSans 480 0 0 0 Config_accessC_bit2
port 2 nsew signal tristate
flabel metal3 s 22840 10888 23300 11008 0 FreeSans 480 0 0 0 Config_accessC_bit3
port 3 nsew signal tristate
flabel metal3 s -300 17960 160 18080 0 FreeSans 480 0 0 0 E1END[0]
port 4 nsew signal input
flabel metal3 s -300 18232 160 18352 0 FreeSans 480 0 0 0 E1END[1]
port 5 nsew signal input
flabel metal3 s -300 18504 160 18624 0 FreeSans 480 0 0 0 E1END[2]
port 6 nsew signal input
flabel metal3 s -300 18776 160 18896 0 FreeSans 480 0 0 0 E1END[3]
port 7 nsew signal input
flabel metal3 s -300 21224 160 21344 0 FreeSans 480 0 0 0 E2END[0]
port 8 nsew signal input
flabel metal3 s -300 21496 160 21616 0 FreeSans 480 0 0 0 E2END[1]
port 9 nsew signal input
flabel metal3 s -300 21768 160 21888 0 FreeSans 480 0 0 0 E2END[2]
port 10 nsew signal input
flabel metal3 s -300 22040 160 22160 0 FreeSans 480 0 0 0 E2END[3]
port 11 nsew signal input
flabel metal3 s -300 22312 160 22432 0 FreeSans 480 0 0 0 E2END[4]
port 12 nsew signal input
flabel metal3 s -300 22584 160 22704 0 FreeSans 480 0 0 0 E2END[5]
port 13 nsew signal input
flabel metal3 s -300 22856 160 22976 0 FreeSans 480 0 0 0 E2END[6]
port 14 nsew signal input
flabel metal3 s -300 23128 160 23248 0 FreeSans 480 0 0 0 E2END[7]
port 15 nsew signal input
flabel metal3 s -300 19048 160 19168 0 FreeSans 480 0 0 0 E2MID[0]
port 16 nsew signal input
flabel metal3 s -300 19320 160 19440 0 FreeSans 480 0 0 0 E2MID[1]
port 17 nsew signal input
flabel metal3 s -300 19592 160 19712 0 FreeSans 480 0 0 0 E2MID[2]
port 18 nsew signal input
flabel metal3 s -300 19864 160 19984 0 FreeSans 480 0 0 0 E2MID[3]
port 19 nsew signal input
flabel metal3 s -300 20136 160 20256 0 FreeSans 480 0 0 0 E2MID[4]
port 20 nsew signal input
flabel metal3 s -300 20408 160 20528 0 FreeSans 480 0 0 0 E2MID[5]
port 21 nsew signal input
flabel metal3 s -300 20680 160 20800 0 FreeSans 480 0 0 0 E2MID[6]
port 22 nsew signal input
flabel metal3 s -300 20952 160 21072 0 FreeSans 480 0 0 0 E2MID[7]
port 23 nsew signal input
flabel metal3 s -300 27752 160 27872 0 FreeSans 480 0 0 0 E6END[0]
port 24 nsew signal input
flabel metal3 s -300 30472 160 30592 0 FreeSans 480 0 0 0 E6END[10]
port 25 nsew signal input
flabel metal3 s -300 30744 160 30864 0 FreeSans 480 0 0 0 E6END[11]
port 26 nsew signal input
flabel metal3 s -300 28024 160 28144 0 FreeSans 480 0 0 0 E6END[1]
port 27 nsew signal input
flabel metal3 s -300 28296 160 28416 0 FreeSans 480 0 0 0 E6END[2]
port 28 nsew signal input
flabel metal3 s -300 28568 160 28688 0 FreeSans 480 0 0 0 E6END[3]
port 29 nsew signal input
flabel metal3 s -300 28840 160 28960 0 FreeSans 480 0 0 0 E6END[4]
port 30 nsew signal input
flabel metal3 s -300 29112 160 29232 0 FreeSans 480 0 0 0 E6END[5]
port 31 nsew signal input
flabel metal3 s -300 29384 160 29504 0 FreeSans 480 0 0 0 E6END[6]
port 32 nsew signal input
flabel metal3 s -300 29656 160 29776 0 FreeSans 480 0 0 0 E6END[7]
port 33 nsew signal input
flabel metal3 s -300 29928 160 30048 0 FreeSans 480 0 0 0 E6END[8]
port 34 nsew signal input
flabel metal3 s -300 30200 160 30320 0 FreeSans 480 0 0 0 E6END[9]
port 35 nsew signal input
flabel metal3 s -300 23400 160 23520 0 FreeSans 480 0 0 0 EE4END[0]
port 36 nsew signal input
flabel metal3 s -300 26120 160 26240 0 FreeSans 480 0 0 0 EE4END[10]
port 37 nsew signal input
flabel metal3 s -300 26392 160 26512 0 FreeSans 480 0 0 0 EE4END[11]
port 38 nsew signal input
flabel metal3 s -300 26664 160 26784 0 FreeSans 480 0 0 0 EE4END[12]
port 39 nsew signal input
flabel metal3 s -300 26936 160 27056 0 FreeSans 480 0 0 0 EE4END[13]
port 40 nsew signal input
flabel metal3 s -300 27208 160 27328 0 FreeSans 480 0 0 0 EE4END[14]
port 41 nsew signal input
flabel metal3 s -300 27480 160 27600 0 FreeSans 480 0 0 0 EE4END[15]
port 42 nsew signal input
flabel metal3 s -300 23672 160 23792 0 FreeSans 480 0 0 0 EE4END[1]
port 43 nsew signal input
flabel metal3 s -300 23944 160 24064 0 FreeSans 480 0 0 0 EE4END[2]
port 44 nsew signal input
flabel metal3 s -300 24216 160 24336 0 FreeSans 480 0 0 0 EE4END[3]
port 45 nsew signal input
flabel metal3 s -300 24488 160 24608 0 FreeSans 480 0 0 0 EE4END[4]
port 46 nsew signal input
flabel metal3 s -300 24760 160 24880 0 FreeSans 480 0 0 0 EE4END[5]
port 47 nsew signal input
flabel metal3 s -300 25032 160 25152 0 FreeSans 480 0 0 0 EE4END[6]
port 48 nsew signal input
flabel metal3 s -300 25304 160 25424 0 FreeSans 480 0 0 0 EE4END[7]
port 49 nsew signal input
flabel metal3 s -300 25576 160 25696 0 FreeSans 480 0 0 0 EE4END[8]
port 50 nsew signal input
flabel metal3 s -300 25848 160 25968 0 FreeSans 480 0 0 0 EE4END[9]
port 51 nsew signal input
flabel metal3 s 22840 15784 23300 15904 0 FreeSans 480 0 0 0 FAB2RAM_A0_O0
port 52 nsew signal tristate
flabel metal3 s 22840 16328 23300 16448 0 FreeSans 480 0 0 0 FAB2RAM_A0_O1
port 53 nsew signal tristate
flabel metal3 s 22840 16872 23300 16992 0 FreeSans 480 0 0 0 FAB2RAM_A0_O2
port 54 nsew signal tristate
flabel metal3 s 22840 17416 23300 17536 0 FreeSans 480 0 0 0 FAB2RAM_A0_O3
port 55 nsew signal tristate
flabel metal3 s 22840 13608 23300 13728 0 FreeSans 480 0 0 0 FAB2RAM_A1_O0
port 56 nsew signal tristate
flabel metal3 s 22840 14152 23300 14272 0 FreeSans 480 0 0 0 FAB2RAM_A1_O1
port 57 nsew signal tristate
flabel metal3 s 22840 14696 23300 14816 0 FreeSans 480 0 0 0 FAB2RAM_A1_O2
port 58 nsew signal tristate
flabel metal3 s 22840 15240 23300 15360 0 FreeSans 480 0 0 0 FAB2RAM_A1_O3
port 59 nsew signal tristate
flabel metal3 s 22840 11432 23300 11552 0 FreeSans 480 0 0 0 FAB2RAM_C_O0
port 60 nsew signal tristate
flabel metal3 s 22840 11976 23300 12096 0 FreeSans 480 0 0 0 FAB2RAM_C_O1
port 61 nsew signal tristate
flabel metal3 s 22840 12520 23300 12640 0 FreeSans 480 0 0 0 FAB2RAM_C_O2
port 62 nsew signal tristate
flabel metal3 s 22840 13064 23300 13184 0 FreeSans 480 0 0 0 FAB2RAM_C_O3
port 63 nsew signal tristate
flabel metal3 s 22840 24488 23300 24608 0 FreeSans 480 0 0 0 FAB2RAM_D0_O0
port 64 nsew signal tristate
flabel metal3 s 22840 25032 23300 25152 0 FreeSans 480 0 0 0 FAB2RAM_D0_O1
port 65 nsew signal tristate
flabel metal3 s 22840 25576 23300 25696 0 FreeSans 480 0 0 0 FAB2RAM_D0_O2
port 66 nsew signal tristate
flabel metal3 s 22840 26120 23300 26240 0 FreeSans 480 0 0 0 FAB2RAM_D0_O3
port 67 nsew signal tristate
flabel metal3 s 22840 22312 23300 22432 0 FreeSans 480 0 0 0 FAB2RAM_D1_O0
port 68 nsew signal tristate
flabel metal3 s 22840 22856 23300 22976 0 FreeSans 480 0 0 0 FAB2RAM_D1_O1
port 69 nsew signal tristate
flabel metal3 s 22840 23400 23300 23520 0 FreeSans 480 0 0 0 FAB2RAM_D1_O2
port 70 nsew signal tristate
flabel metal3 s 22840 23944 23300 24064 0 FreeSans 480 0 0 0 FAB2RAM_D1_O3
port 71 nsew signal tristate
flabel metal3 s 22840 20136 23300 20256 0 FreeSans 480 0 0 0 FAB2RAM_D2_O0
port 72 nsew signal tristate
flabel metal3 s 22840 20680 23300 20800 0 FreeSans 480 0 0 0 FAB2RAM_D2_O1
port 73 nsew signal tristate
flabel metal3 s 22840 21224 23300 21344 0 FreeSans 480 0 0 0 FAB2RAM_D2_O2
port 74 nsew signal tristate
flabel metal3 s 22840 21768 23300 21888 0 FreeSans 480 0 0 0 FAB2RAM_D2_O3
port 75 nsew signal tristate
flabel metal3 s 22840 17960 23300 18080 0 FreeSans 480 0 0 0 FAB2RAM_D3_O0
port 76 nsew signal tristate
flabel metal3 s 22840 18504 23300 18624 0 FreeSans 480 0 0 0 FAB2RAM_D3_O1
port 77 nsew signal tristate
flabel metal3 s 22840 19048 23300 19168 0 FreeSans 480 0 0 0 FAB2RAM_D3_O2
port 78 nsew signal tristate
flabel metal3 s 22840 19592 23300 19712 0 FreeSans 480 0 0 0 FAB2RAM_D3_O3
port 79 nsew signal tristate
flabel metal3 s -300 31016 160 31136 0 FreeSans 480 0 0 0 FrameData[0]
port 80 nsew signal input
flabel metal3 s -300 33736 160 33856 0 FreeSans 480 0 0 0 FrameData[10]
port 81 nsew signal input
flabel metal3 s -300 34008 160 34128 0 FreeSans 480 0 0 0 FrameData[11]
port 82 nsew signal input
flabel metal3 s -300 34280 160 34400 0 FreeSans 480 0 0 0 FrameData[12]
port 83 nsew signal input
flabel metal3 s -300 34552 160 34672 0 FreeSans 480 0 0 0 FrameData[13]
port 84 nsew signal input
flabel metal3 s -300 34824 160 34944 0 FreeSans 480 0 0 0 FrameData[14]
port 85 nsew signal input
flabel metal3 s -300 35096 160 35216 0 FreeSans 480 0 0 0 FrameData[15]
port 86 nsew signal input
flabel metal3 s -300 35368 160 35488 0 FreeSans 480 0 0 0 FrameData[16]
port 87 nsew signal input
flabel metal3 s -300 35640 160 35760 0 FreeSans 480 0 0 0 FrameData[17]
port 88 nsew signal input
flabel metal3 s -300 35912 160 36032 0 FreeSans 480 0 0 0 FrameData[18]
port 89 nsew signal input
flabel metal3 s -300 36184 160 36304 0 FreeSans 480 0 0 0 FrameData[19]
port 90 nsew signal input
flabel metal3 s -300 31288 160 31408 0 FreeSans 480 0 0 0 FrameData[1]
port 91 nsew signal input
flabel metal3 s -300 36456 160 36576 0 FreeSans 480 0 0 0 FrameData[20]
port 92 nsew signal input
flabel metal3 s -300 36728 160 36848 0 FreeSans 480 0 0 0 FrameData[21]
port 93 nsew signal input
flabel metal3 s -300 37000 160 37120 0 FreeSans 480 0 0 0 FrameData[22]
port 94 nsew signal input
flabel metal3 s -300 37272 160 37392 0 FreeSans 480 0 0 0 FrameData[23]
port 95 nsew signal input
flabel metal3 s -300 37544 160 37664 0 FreeSans 480 0 0 0 FrameData[24]
port 96 nsew signal input
flabel metal3 s -300 37816 160 37936 0 FreeSans 480 0 0 0 FrameData[25]
port 97 nsew signal input
flabel metal3 s -300 38088 160 38208 0 FreeSans 480 0 0 0 FrameData[26]
port 98 nsew signal input
flabel metal3 s -300 38360 160 38480 0 FreeSans 480 0 0 0 FrameData[27]
port 99 nsew signal input
flabel metal3 s -300 38632 160 38752 0 FreeSans 480 0 0 0 FrameData[28]
port 100 nsew signal input
flabel metal3 s -300 38904 160 39024 0 FreeSans 480 0 0 0 FrameData[29]
port 101 nsew signal input
flabel metal3 s -300 31560 160 31680 0 FreeSans 480 0 0 0 FrameData[2]
port 102 nsew signal input
flabel metal3 s -300 39176 160 39296 0 FreeSans 480 0 0 0 FrameData[30]
port 103 nsew signal input
flabel metal3 s -300 39448 160 39568 0 FreeSans 480 0 0 0 FrameData[31]
port 104 nsew signal input
flabel metal3 s -300 31832 160 31952 0 FreeSans 480 0 0 0 FrameData[3]
port 105 nsew signal input
flabel metal3 s -300 32104 160 32224 0 FreeSans 480 0 0 0 FrameData[4]
port 106 nsew signal input
flabel metal3 s -300 32376 160 32496 0 FreeSans 480 0 0 0 FrameData[5]
port 107 nsew signal input
flabel metal3 s -300 32648 160 32768 0 FreeSans 480 0 0 0 FrameData[6]
port 108 nsew signal input
flabel metal3 s -300 32920 160 33040 0 FreeSans 480 0 0 0 FrameData[7]
port 109 nsew signal input
flabel metal3 s -300 33192 160 33312 0 FreeSans 480 0 0 0 FrameData[8]
port 110 nsew signal input
flabel metal3 s -300 33464 160 33584 0 FreeSans 480 0 0 0 FrameData[9]
port 111 nsew signal input
flabel metal3 s 22840 26664 23300 26784 0 FreeSans 480 0 0 0 FrameData_O[0]
port 112 nsew signal tristate
flabel metal3 s 22840 32104 23300 32224 0 FreeSans 480 0 0 0 FrameData_O[10]
port 113 nsew signal tristate
flabel metal3 s 22840 32648 23300 32768 0 FreeSans 480 0 0 0 FrameData_O[11]
port 114 nsew signal tristate
flabel metal3 s 22840 33192 23300 33312 0 FreeSans 480 0 0 0 FrameData_O[12]
port 115 nsew signal tristate
flabel metal3 s 22840 33736 23300 33856 0 FreeSans 480 0 0 0 FrameData_O[13]
port 116 nsew signal tristate
flabel metal3 s 22840 34280 23300 34400 0 FreeSans 480 0 0 0 FrameData_O[14]
port 117 nsew signal tristate
flabel metal3 s 22840 34824 23300 34944 0 FreeSans 480 0 0 0 FrameData_O[15]
port 118 nsew signal tristate
flabel metal3 s 22840 35368 23300 35488 0 FreeSans 480 0 0 0 FrameData_O[16]
port 119 nsew signal tristate
flabel metal3 s 22840 35912 23300 36032 0 FreeSans 480 0 0 0 FrameData_O[17]
port 120 nsew signal tristate
flabel metal3 s 22840 36456 23300 36576 0 FreeSans 480 0 0 0 FrameData_O[18]
port 121 nsew signal tristate
flabel metal3 s 22840 37000 23300 37120 0 FreeSans 480 0 0 0 FrameData_O[19]
port 122 nsew signal tristate
flabel metal3 s 22840 27208 23300 27328 0 FreeSans 480 0 0 0 FrameData_O[1]
port 123 nsew signal tristate
flabel metal3 s 22840 37544 23300 37664 0 FreeSans 480 0 0 0 FrameData_O[20]
port 124 nsew signal tristate
flabel metal3 s 22840 38088 23300 38208 0 FreeSans 480 0 0 0 FrameData_O[21]
port 125 nsew signal tristate
flabel metal3 s 22840 38632 23300 38752 0 FreeSans 480 0 0 0 FrameData_O[22]
port 126 nsew signal tristate
flabel metal3 s 22840 39176 23300 39296 0 FreeSans 480 0 0 0 FrameData_O[23]
port 127 nsew signal tristate
flabel metal3 s 22840 39720 23300 39840 0 FreeSans 480 0 0 0 FrameData_O[24]
port 128 nsew signal tristate
flabel metal3 s 22840 40264 23300 40384 0 FreeSans 480 0 0 0 FrameData_O[25]
port 129 nsew signal tristate
flabel metal3 s 22840 40808 23300 40928 0 FreeSans 480 0 0 0 FrameData_O[26]
port 130 nsew signal tristate
flabel metal3 s 22840 41352 23300 41472 0 FreeSans 480 0 0 0 FrameData_O[27]
port 131 nsew signal tristate
flabel metal3 s 22840 41896 23300 42016 0 FreeSans 480 0 0 0 FrameData_O[28]
port 132 nsew signal tristate
flabel metal3 s 22840 42440 23300 42560 0 FreeSans 480 0 0 0 FrameData_O[29]
port 133 nsew signal tristate
flabel metal3 s 22840 27752 23300 27872 0 FreeSans 480 0 0 0 FrameData_O[2]
port 134 nsew signal tristate
flabel metal3 s 22840 42984 23300 43104 0 FreeSans 480 0 0 0 FrameData_O[30]
port 135 nsew signal tristate
flabel metal3 s 22840 43528 23300 43648 0 FreeSans 480 0 0 0 FrameData_O[31]
port 136 nsew signal tristate
flabel metal3 s 22840 28296 23300 28416 0 FreeSans 480 0 0 0 FrameData_O[3]
port 137 nsew signal tristate
flabel metal3 s 22840 28840 23300 28960 0 FreeSans 480 0 0 0 FrameData_O[4]
port 138 nsew signal tristate
flabel metal3 s 22840 29384 23300 29504 0 FreeSans 480 0 0 0 FrameData_O[5]
port 139 nsew signal tristate
flabel metal3 s 22840 29928 23300 30048 0 FreeSans 480 0 0 0 FrameData_O[6]
port 140 nsew signal tristate
flabel metal3 s 22840 30472 23300 30592 0 FreeSans 480 0 0 0 FrameData_O[7]
port 141 nsew signal tristate
flabel metal3 s 22840 31016 23300 31136 0 FreeSans 480 0 0 0 FrameData_O[8]
port 142 nsew signal tristate
flabel metal3 s 22840 31560 23300 31680 0 FreeSans 480 0 0 0 FrameData_O[9]
port 143 nsew signal tristate
flabel metal2 s 16394 -300 16450 160 0 FreeSans 224 90 0 0 FrameStrobe[0]
port 144 nsew signal input
flabel metal2 s 18234 -300 18290 160 0 FreeSans 224 90 0 0 FrameStrobe[10]
port 145 nsew signal input
flabel metal2 s 18418 -300 18474 160 0 FreeSans 224 90 0 0 FrameStrobe[11]
port 146 nsew signal input
flabel metal2 s 18602 -300 18658 160 0 FreeSans 224 90 0 0 FrameStrobe[12]
port 147 nsew signal input
flabel metal2 s 18786 -300 18842 160 0 FreeSans 224 90 0 0 FrameStrobe[13]
port 148 nsew signal input
flabel metal2 s 18970 -300 19026 160 0 FreeSans 224 90 0 0 FrameStrobe[14]
port 149 nsew signal input
flabel metal2 s 19154 -300 19210 160 0 FreeSans 224 90 0 0 FrameStrobe[15]
port 150 nsew signal input
flabel metal2 s 19338 -300 19394 160 0 FreeSans 224 90 0 0 FrameStrobe[16]
port 151 nsew signal input
flabel metal2 s 19522 -300 19578 160 0 FreeSans 224 90 0 0 FrameStrobe[17]
port 152 nsew signal input
flabel metal2 s 19706 -300 19762 160 0 FreeSans 224 90 0 0 FrameStrobe[18]
port 153 nsew signal input
flabel metal2 s 19890 -300 19946 160 0 FreeSans 224 90 0 0 FrameStrobe[19]
port 154 nsew signal input
flabel metal2 s 16578 -300 16634 160 0 FreeSans 224 90 0 0 FrameStrobe[1]
port 155 nsew signal input
flabel metal2 s 16762 -300 16818 160 0 FreeSans 224 90 0 0 FrameStrobe[2]
port 156 nsew signal input
flabel metal2 s 16946 -300 17002 160 0 FreeSans 224 90 0 0 FrameStrobe[3]
port 157 nsew signal input
flabel metal2 s 17130 -300 17186 160 0 FreeSans 224 90 0 0 FrameStrobe[4]
port 158 nsew signal input
flabel metal2 s 17314 -300 17370 160 0 FreeSans 224 90 0 0 FrameStrobe[5]
port 159 nsew signal input
flabel metal2 s 17498 -300 17554 160 0 FreeSans 224 90 0 0 FrameStrobe[6]
port 160 nsew signal input
flabel metal2 s 17682 -300 17738 160 0 FreeSans 224 90 0 0 FrameStrobe[7]
port 161 nsew signal input
flabel metal2 s 17866 -300 17922 160 0 FreeSans 224 90 0 0 FrameStrobe[8]
port 162 nsew signal input
flabel metal2 s 18050 -300 18106 160 0 FreeSans 224 90 0 0 FrameStrobe[9]
port 163 nsew signal input
flabel metal2 s 16394 44540 16450 45000 0 FreeSans 224 90 0 0 FrameStrobe_O[0]
port 164 nsew signal tristate
flabel metal2 s 18234 44540 18290 45000 0 FreeSans 224 90 0 0 FrameStrobe_O[10]
port 165 nsew signal tristate
flabel metal2 s 18418 44540 18474 45000 0 FreeSans 224 90 0 0 FrameStrobe_O[11]
port 166 nsew signal tristate
flabel metal2 s 18602 44540 18658 45000 0 FreeSans 224 90 0 0 FrameStrobe_O[12]
port 167 nsew signal tristate
flabel metal2 s 18786 44540 18842 45000 0 FreeSans 224 90 0 0 FrameStrobe_O[13]
port 168 nsew signal tristate
flabel metal2 s 18970 44540 19026 45000 0 FreeSans 224 90 0 0 FrameStrobe_O[14]
port 169 nsew signal tristate
flabel metal2 s 19154 44540 19210 45000 0 FreeSans 224 90 0 0 FrameStrobe_O[15]
port 170 nsew signal tristate
flabel metal2 s 19338 44540 19394 45000 0 FreeSans 224 90 0 0 FrameStrobe_O[16]
port 171 nsew signal tristate
flabel metal2 s 19522 44540 19578 45000 0 FreeSans 224 90 0 0 FrameStrobe_O[17]
port 172 nsew signal tristate
flabel metal2 s 19706 44540 19762 45000 0 FreeSans 224 90 0 0 FrameStrobe_O[18]
port 173 nsew signal tristate
flabel metal2 s 19890 44540 19946 45000 0 FreeSans 224 90 0 0 FrameStrobe_O[19]
port 174 nsew signal tristate
flabel metal2 s 16578 44540 16634 45000 0 FreeSans 224 90 0 0 FrameStrobe_O[1]
port 175 nsew signal tristate
flabel metal2 s 16762 44540 16818 45000 0 FreeSans 224 90 0 0 FrameStrobe_O[2]
port 176 nsew signal tristate
flabel metal2 s 16946 44540 17002 45000 0 FreeSans 224 90 0 0 FrameStrobe_O[3]
port 177 nsew signal tristate
flabel metal2 s 17130 44540 17186 45000 0 FreeSans 224 90 0 0 FrameStrobe_O[4]
port 178 nsew signal tristate
flabel metal2 s 17314 44540 17370 45000 0 FreeSans 224 90 0 0 FrameStrobe_O[5]
port 179 nsew signal tristate
flabel metal2 s 17498 44540 17554 45000 0 FreeSans 224 90 0 0 FrameStrobe_O[6]
port 180 nsew signal tristate
flabel metal2 s 17682 44540 17738 45000 0 FreeSans 224 90 0 0 FrameStrobe_O[7]
port 181 nsew signal tristate
flabel metal2 s 17866 44540 17922 45000 0 FreeSans 224 90 0 0 FrameStrobe_O[8]
port 182 nsew signal tristate
flabel metal2 s 18050 44540 18106 45000 0 FreeSans 224 90 0 0 FrameStrobe_O[9]
port 183 nsew signal tristate
flabel metal2 s 2962 44540 3018 45000 0 FreeSans 224 90 0 0 N1BEG[0]
port 184 nsew signal tristate
flabel metal2 s 3146 44540 3202 45000 0 FreeSans 224 90 0 0 N1BEG[1]
port 185 nsew signal tristate
flabel metal2 s 3330 44540 3386 45000 0 FreeSans 224 90 0 0 N1BEG[2]
port 186 nsew signal tristate
flabel metal2 s 3514 44540 3570 45000 0 FreeSans 224 90 0 0 N1BEG[3]
port 187 nsew signal tristate
flabel metal2 s 2962 -300 3018 160 0 FreeSans 224 90 0 0 N1END[0]
port 188 nsew signal input
flabel metal2 s 3146 -300 3202 160 0 FreeSans 224 90 0 0 N1END[1]
port 189 nsew signal input
flabel metal2 s 3330 -300 3386 160 0 FreeSans 224 90 0 0 N1END[2]
port 190 nsew signal input
flabel metal2 s 3514 -300 3570 160 0 FreeSans 224 90 0 0 N1END[3]
port 191 nsew signal input
flabel metal2 s 3698 44540 3754 45000 0 FreeSans 224 90 0 0 N2BEG[0]
port 192 nsew signal tristate
flabel metal2 s 3882 44540 3938 45000 0 FreeSans 224 90 0 0 N2BEG[1]
port 193 nsew signal tristate
flabel metal2 s 4066 44540 4122 45000 0 FreeSans 224 90 0 0 N2BEG[2]
port 194 nsew signal tristate
flabel metal2 s 4250 44540 4306 45000 0 FreeSans 224 90 0 0 N2BEG[3]
port 195 nsew signal tristate
flabel metal2 s 4434 44540 4490 45000 0 FreeSans 224 90 0 0 N2BEG[4]
port 196 nsew signal tristate
flabel metal2 s 4618 44540 4674 45000 0 FreeSans 224 90 0 0 N2BEG[5]
port 197 nsew signal tristate
flabel metal2 s 4802 44540 4858 45000 0 FreeSans 224 90 0 0 N2BEG[6]
port 198 nsew signal tristate
flabel metal2 s 4986 44540 5042 45000 0 FreeSans 224 90 0 0 N2BEG[7]
port 199 nsew signal tristate
flabel metal2 s 5170 44540 5226 45000 0 FreeSans 224 90 0 0 N2BEGb[0]
port 200 nsew signal tristate
flabel metal2 s 5354 44540 5410 45000 0 FreeSans 224 90 0 0 N2BEGb[1]
port 201 nsew signal tristate
flabel metal2 s 5538 44540 5594 45000 0 FreeSans 224 90 0 0 N2BEGb[2]
port 202 nsew signal tristate
flabel metal2 s 5722 44540 5778 45000 0 FreeSans 224 90 0 0 N2BEGb[3]
port 203 nsew signal tristate
flabel metal2 s 5906 44540 5962 45000 0 FreeSans 224 90 0 0 N2BEGb[4]
port 204 nsew signal tristate
flabel metal2 s 6090 44540 6146 45000 0 FreeSans 224 90 0 0 N2BEGb[5]
port 205 nsew signal tristate
flabel metal2 s 6274 44540 6330 45000 0 FreeSans 224 90 0 0 N2BEGb[6]
port 206 nsew signal tristate
flabel metal2 s 6458 44540 6514 45000 0 FreeSans 224 90 0 0 N2BEGb[7]
port 207 nsew signal tristate
flabel metal2 s 5170 -300 5226 160 0 FreeSans 224 90 0 0 N2END[0]
port 208 nsew signal input
flabel metal2 s 5354 -300 5410 160 0 FreeSans 224 90 0 0 N2END[1]
port 209 nsew signal input
flabel metal2 s 5538 -300 5594 160 0 FreeSans 224 90 0 0 N2END[2]
port 210 nsew signal input
flabel metal2 s 5722 -300 5778 160 0 FreeSans 224 90 0 0 N2END[3]
port 211 nsew signal input
flabel metal2 s 5906 -300 5962 160 0 FreeSans 224 90 0 0 N2END[4]
port 212 nsew signal input
flabel metal2 s 6090 -300 6146 160 0 FreeSans 224 90 0 0 N2END[5]
port 213 nsew signal input
flabel metal2 s 6274 -300 6330 160 0 FreeSans 224 90 0 0 N2END[6]
port 214 nsew signal input
flabel metal2 s 6458 -300 6514 160 0 FreeSans 224 90 0 0 N2END[7]
port 215 nsew signal input
flabel metal2 s 3698 -300 3754 160 0 FreeSans 224 90 0 0 N2MID[0]
port 216 nsew signal input
flabel metal2 s 3882 -300 3938 160 0 FreeSans 224 90 0 0 N2MID[1]
port 217 nsew signal input
flabel metal2 s 4066 -300 4122 160 0 FreeSans 224 90 0 0 N2MID[2]
port 218 nsew signal input
flabel metal2 s 4250 -300 4306 160 0 FreeSans 224 90 0 0 N2MID[3]
port 219 nsew signal input
flabel metal2 s 4434 -300 4490 160 0 FreeSans 224 90 0 0 N2MID[4]
port 220 nsew signal input
flabel metal2 s 4618 -300 4674 160 0 FreeSans 224 90 0 0 N2MID[5]
port 221 nsew signal input
flabel metal2 s 4802 -300 4858 160 0 FreeSans 224 90 0 0 N2MID[6]
port 222 nsew signal input
flabel metal2 s 4986 -300 5042 160 0 FreeSans 224 90 0 0 N2MID[7]
port 223 nsew signal input
flabel metal2 s 6642 44540 6698 45000 0 FreeSans 224 90 0 0 N4BEG[0]
port 224 nsew signal tristate
flabel metal2 s 8482 44540 8538 45000 0 FreeSans 224 90 0 0 N4BEG[10]
port 225 nsew signal tristate
flabel metal2 s 8666 44540 8722 45000 0 FreeSans 224 90 0 0 N4BEG[11]
port 226 nsew signal tristate
flabel metal2 s 8850 44540 8906 45000 0 FreeSans 224 90 0 0 N4BEG[12]
port 227 nsew signal tristate
flabel metal2 s 9034 44540 9090 45000 0 FreeSans 224 90 0 0 N4BEG[13]
port 228 nsew signal tristate
flabel metal2 s 9218 44540 9274 45000 0 FreeSans 224 90 0 0 N4BEG[14]
port 229 nsew signal tristate
flabel metal2 s 9402 44540 9458 45000 0 FreeSans 224 90 0 0 N4BEG[15]
port 230 nsew signal tristate
flabel metal2 s 6826 44540 6882 45000 0 FreeSans 224 90 0 0 N4BEG[1]
port 231 nsew signal tristate
flabel metal2 s 7010 44540 7066 45000 0 FreeSans 224 90 0 0 N4BEG[2]
port 232 nsew signal tristate
flabel metal2 s 7194 44540 7250 45000 0 FreeSans 224 90 0 0 N4BEG[3]
port 233 nsew signal tristate
flabel metal2 s 7378 44540 7434 45000 0 FreeSans 224 90 0 0 N4BEG[4]
port 234 nsew signal tristate
flabel metal2 s 7562 44540 7618 45000 0 FreeSans 224 90 0 0 N4BEG[5]
port 235 nsew signal tristate
flabel metal2 s 7746 44540 7802 45000 0 FreeSans 224 90 0 0 N4BEG[6]
port 236 nsew signal tristate
flabel metal2 s 7930 44540 7986 45000 0 FreeSans 224 90 0 0 N4BEG[7]
port 237 nsew signal tristate
flabel metal2 s 8114 44540 8170 45000 0 FreeSans 224 90 0 0 N4BEG[8]
port 238 nsew signal tristate
flabel metal2 s 8298 44540 8354 45000 0 FreeSans 224 90 0 0 N4BEG[9]
port 239 nsew signal tristate
flabel metal2 s 6642 -300 6698 160 0 FreeSans 224 90 0 0 N4END[0]
port 240 nsew signal input
flabel metal2 s 8482 -300 8538 160 0 FreeSans 224 90 0 0 N4END[10]
port 241 nsew signal input
flabel metal2 s 8666 -300 8722 160 0 FreeSans 224 90 0 0 N4END[11]
port 242 nsew signal input
flabel metal2 s 8850 -300 8906 160 0 FreeSans 224 90 0 0 N4END[12]
port 243 nsew signal input
flabel metal2 s 9034 -300 9090 160 0 FreeSans 224 90 0 0 N4END[13]
port 244 nsew signal input
flabel metal2 s 9218 -300 9274 160 0 FreeSans 224 90 0 0 N4END[14]
port 245 nsew signal input
flabel metal2 s 9402 -300 9458 160 0 FreeSans 224 90 0 0 N4END[15]
port 246 nsew signal input
flabel metal2 s 6826 -300 6882 160 0 FreeSans 224 90 0 0 N4END[1]
port 247 nsew signal input
flabel metal2 s 7010 -300 7066 160 0 FreeSans 224 90 0 0 N4END[2]
port 248 nsew signal input
flabel metal2 s 7194 -300 7250 160 0 FreeSans 224 90 0 0 N4END[3]
port 249 nsew signal input
flabel metal2 s 7378 -300 7434 160 0 FreeSans 224 90 0 0 N4END[4]
port 250 nsew signal input
flabel metal2 s 7562 -300 7618 160 0 FreeSans 224 90 0 0 N4END[5]
port 251 nsew signal input
flabel metal2 s 7746 -300 7802 160 0 FreeSans 224 90 0 0 N4END[6]
port 252 nsew signal input
flabel metal2 s 7930 -300 7986 160 0 FreeSans 224 90 0 0 N4END[7]
port 253 nsew signal input
flabel metal2 s 8114 -300 8170 160 0 FreeSans 224 90 0 0 N4END[8]
port 254 nsew signal input
flabel metal2 s 8298 -300 8354 160 0 FreeSans 224 90 0 0 N4END[9]
port 255 nsew signal input
flabel metal3 s 22840 7080 23300 7200 0 FreeSans 480 0 0 0 RAM2FAB_D0_I0
port 256 nsew signal input
flabel metal3 s 22840 7624 23300 7744 0 FreeSans 480 0 0 0 RAM2FAB_D0_I1
port 257 nsew signal input
flabel metal3 s 22840 8168 23300 8288 0 FreeSans 480 0 0 0 RAM2FAB_D0_I2
port 258 nsew signal input
flabel metal3 s 22840 8712 23300 8832 0 FreeSans 480 0 0 0 RAM2FAB_D0_I3
port 259 nsew signal input
flabel metal3 s 22840 4904 23300 5024 0 FreeSans 480 0 0 0 RAM2FAB_D1_I0
port 260 nsew signal input
flabel metal3 s 22840 5448 23300 5568 0 FreeSans 480 0 0 0 RAM2FAB_D1_I1
port 261 nsew signal input
flabel metal3 s 22840 5992 23300 6112 0 FreeSans 480 0 0 0 RAM2FAB_D1_I2
port 262 nsew signal input
flabel metal3 s 22840 6536 23300 6656 0 FreeSans 480 0 0 0 RAM2FAB_D1_I3
port 263 nsew signal input
flabel metal3 s 22840 2728 23300 2848 0 FreeSans 480 0 0 0 RAM2FAB_D2_I0
port 264 nsew signal input
flabel metal3 s 22840 3272 23300 3392 0 FreeSans 480 0 0 0 RAM2FAB_D2_I1
port 265 nsew signal input
flabel metal3 s 22840 3816 23300 3936 0 FreeSans 480 0 0 0 RAM2FAB_D2_I2
port 266 nsew signal input
flabel metal3 s 22840 4360 23300 4480 0 FreeSans 480 0 0 0 RAM2FAB_D2_I3
port 267 nsew signal input
flabel metal3 s 22840 552 23300 672 0 FreeSans 480 0 0 0 RAM2FAB_D3_I0
port 268 nsew signal input
flabel metal3 s 22840 1096 23300 1216 0 FreeSans 480 0 0 0 RAM2FAB_D3_I1
port 269 nsew signal input
flabel metal3 s 22840 1640 23300 1760 0 FreeSans 480 0 0 0 RAM2FAB_D3_I2
port 270 nsew signal input
flabel metal3 s 22840 2184 23300 2304 0 FreeSans 480 0 0 0 RAM2FAB_D3_I3
port 271 nsew signal input
flabel metal2 s 9586 -300 9642 160 0 FreeSans 224 90 0 0 S1BEG[0]
port 272 nsew signal tristate
flabel metal2 s 9770 -300 9826 160 0 FreeSans 224 90 0 0 S1BEG[1]
port 273 nsew signal tristate
flabel metal2 s 9954 -300 10010 160 0 FreeSans 224 90 0 0 S1BEG[2]
port 274 nsew signal tristate
flabel metal2 s 10138 -300 10194 160 0 FreeSans 224 90 0 0 S1BEG[3]
port 275 nsew signal tristate
flabel metal2 s 9586 44540 9642 45000 0 FreeSans 224 90 0 0 S1END[0]
port 276 nsew signal input
flabel metal2 s 9770 44540 9826 45000 0 FreeSans 224 90 0 0 S1END[1]
port 277 nsew signal input
flabel metal2 s 9954 44540 10010 45000 0 FreeSans 224 90 0 0 S1END[2]
port 278 nsew signal input
flabel metal2 s 10138 44540 10194 45000 0 FreeSans 224 90 0 0 S1END[3]
port 279 nsew signal input
flabel metal2 s 11794 -300 11850 160 0 FreeSans 224 90 0 0 S2BEG[0]
port 280 nsew signal tristate
flabel metal2 s 11978 -300 12034 160 0 FreeSans 224 90 0 0 S2BEG[1]
port 281 nsew signal tristate
flabel metal2 s 12162 -300 12218 160 0 FreeSans 224 90 0 0 S2BEG[2]
port 282 nsew signal tristate
flabel metal2 s 12346 -300 12402 160 0 FreeSans 224 90 0 0 S2BEG[3]
port 283 nsew signal tristate
flabel metal2 s 12530 -300 12586 160 0 FreeSans 224 90 0 0 S2BEG[4]
port 284 nsew signal tristate
flabel metal2 s 12714 -300 12770 160 0 FreeSans 224 90 0 0 S2BEG[5]
port 285 nsew signal tristate
flabel metal2 s 12898 -300 12954 160 0 FreeSans 224 90 0 0 S2BEG[6]
port 286 nsew signal tristate
flabel metal2 s 13082 -300 13138 160 0 FreeSans 224 90 0 0 S2BEG[7]
port 287 nsew signal tristate
flabel metal2 s 10322 -300 10378 160 0 FreeSans 224 90 0 0 S2BEGb[0]
port 288 nsew signal tristate
flabel metal2 s 10506 -300 10562 160 0 FreeSans 224 90 0 0 S2BEGb[1]
port 289 nsew signal tristate
flabel metal2 s 10690 -300 10746 160 0 FreeSans 224 90 0 0 S2BEGb[2]
port 290 nsew signal tristate
flabel metal2 s 10874 -300 10930 160 0 FreeSans 224 90 0 0 S2BEGb[3]
port 291 nsew signal tristate
flabel metal2 s 11058 -300 11114 160 0 FreeSans 224 90 0 0 S2BEGb[4]
port 292 nsew signal tristate
flabel metal2 s 11242 -300 11298 160 0 FreeSans 224 90 0 0 S2BEGb[5]
port 293 nsew signal tristate
flabel metal2 s 11426 -300 11482 160 0 FreeSans 224 90 0 0 S2BEGb[6]
port 294 nsew signal tristate
flabel metal2 s 11610 -300 11666 160 0 FreeSans 224 90 0 0 S2BEGb[7]
port 295 nsew signal tristate
flabel metal2 s 10322 44540 10378 45000 0 FreeSans 224 90 0 0 S2END[0]
port 296 nsew signal input
flabel metal2 s 10506 44540 10562 45000 0 FreeSans 224 90 0 0 S2END[1]
port 297 nsew signal input
flabel metal2 s 10690 44540 10746 45000 0 FreeSans 224 90 0 0 S2END[2]
port 298 nsew signal input
flabel metal2 s 10874 44540 10930 45000 0 FreeSans 224 90 0 0 S2END[3]
port 299 nsew signal input
flabel metal2 s 11058 44540 11114 45000 0 FreeSans 224 90 0 0 S2END[4]
port 300 nsew signal input
flabel metal2 s 11242 44540 11298 45000 0 FreeSans 224 90 0 0 S2END[5]
port 301 nsew signal input
flabel metal2 s 11426 44540 11482 45000 0 FreeSans 224 90 0 0 S2END[6]
port 302 nsew signal input
flabel metal2 s 11610 44540 11666 45000 0 FreeSans 224 90 0 0 S2END[7]
port 303 nsew signal input
flabel metal2 s 11794 44540 11850 45000 0 FreeSans 224 90 0 0 S2MID[0]
port 304 nsew signal input
flabel metal2 s 11978 44540 12034 45000 0 FreeSans 224 90 0 0 S2MID[1]
port 305 nsew signal input
flabel metal2 s 12162 44540 12218 45000 0 FreeSans 224 90 0 0 S2MID[2]
port 306 nsew signal input
flabel metal2 s 12346 44540 12402 45000 0 FreeSans 224 90 0 0 S2MID[3]
port 307 nsew signal input
flabel metal2 s 12530 44540 12586 45000 0 FreeSans 224 90 0 0 S2MID[4]
port 308 nsew signal input
flabel metal2 s 12714 44540 12770 45000 0 FreeSans 224 90 0 0 S2MID[5]
port 309 nsew signal input
flabel metal2 s 12898 44540 12954 45000 0 FreeSans 224 90 0 0 S2MID[6]
port 310 nsew signal input
flabel metal2 s 13082 44540 13138 45000 0 FreeSans 224 90 0 0 S2MID[7]
port 311 nsew signal input
flabel metal2 s 13266 -300 13322 160 0 FreeSans 224 90 0 0 S4BEG[0]
port 312 nsew signal tristate
flabel metal2 s 15106 -300 15162 160 0 FreeSans 224 90 0 0 S4BEG[10]
port 313 nsew signal tristate
flabel metal2 s 15290 -300 15346 160 0 FreeSans 224 90 0 0 S4BEG[11]
port 314 nsew signal tristate
flabel metal2 s 15474 -300 15530 160 0 FreeSans 224 90 0 0 S4BEG[12]
port 315 nsew signal tristate
flabel metal2 s 15658 -300 15714 160 0 FreeSans 224 90 0 0 S4BEG[13]
port 316 nsew signal tristate
flabel metal2 s 15842 -300 15898 160 0 FreeSans 224 90 0 0 S4BEG[14]
port 317 nsew signal tristate
flabel metal2 s 16026 -300 16082 160 0 FreeSans 224 90 0 0 S4BEG[15]
port 318 nsew signal tristate
flabel metal2 s 13450 -300 13506 160 0 FreeSans 224 90 0 0 S4BEG[1]
port 319 nsew signal tristate
flabel metal2 s 13634 -300 13690 160 0 FreeSans 224 90 0 0 S4BEG[2]
port 320 nsew signal tristate
flabel metal2 s 13818 -300 13874 160 0 FreeSans 224 90 0 0 S4BEG[3]
port 321 nsew signal tristate
flabel metal2 s 14002 -300 14058 160 0 FreeSans 224 90 0 0 S4BEG[4]
port 322 nsew signal tristate
flabel metal2 s 14186 -300 14242 160 0 FreeSans 224 90 0 0 S4BEG[5]
port 323 nsew signal tristate
flabel metal2 s 14370 -300 14426 160 0 FreeSans 224 90 0 0 S4BEG[6]
port 324 nsew signal tristate
flabel metal2 s 14554 -300 14610 160 0 FreeSans 224 90 0 0 S4BEG[7]
port 325 nsew signal tristate
flabel metal2 s 14738 -300 14794 160 0 FreeSans 224 90 0 0 S4BEG[8]
port 326 nsew signal tristate
flabel metal2 s 14922 -300 14978 160 0 FreeSans 224 90 0 0 S4BEG[9]
port 327 nsew signal tristate
flabel metal2 s 13266 44540 13322 45000 0 FreeSans 224 90 0 0 S4END[0]
port 328 nsew signal input
flabel metal2 s 15106 44540 15162 45000 0 FreeSans 224 90 0 0 S4END[10]
port 329 nsew signal input
flabel metal2 s 15290 44540 15346 45000 0 FreeSans 224 90 0 0 S4END[11]
port 330 nsew signal input
flabel metal2 s 15474 44540 15530 45000 0 FreeSans 224 90 0 0 S4END[12]
port 331 nsew signal input
flabel metal2 s 15658 44540 15714 45000 0 FreeSans 224 90 0 0 S4END[13]
port 332 nsew signal input
flabel metal2 s 15842 44540 15898 45000 0 FreeSans 224 90 0 0 S4END[14]
port 333 nsew signal input
flabel metal2 s 16026 44540 16082 45000 0 FreeSans 224 90 0 0 S4END[15]
port 334 nsew signal input
flabel metal2 s 13450 44540 13506 45000 0 FreeSans 224 90 0 0 S4END[1]
port 335 nsew signal input
flabel metal2 s 13634 44540 13690 45000 0 FreeSans 224 90 0 0 S4END[2]
port 336 nsew signal input
flabel metal2 s 13818 44540 13874 45000 0 FreeSans 224 90 0 0 S4END[3]
port 337 nsew signal input
flabel metal2 s 14002 44540 14058 45000 0 FreeSans 224 90 0 0 S4END[4]
port 338 nsew signal input
flabel metal2 s 14186 44540 14242 45000 0 FreeSans 224 90 0 0 S4END[5]
port 339 nsew signal input
flabel metal2 s 14370 44540 14426 45000 0 FreeSans 224 90 0 0 S4END[6]
port 340 nsew signal input
flabel metal2 s 14554 44540 14610 45000 0 FreeSans 224 90 0 0 S4END[7]
port 341 nsew signal input
flabel metal2 s 14738 44540 14794 45000 0 FreeSans 224 90 0 0 S4END[8]
port 342 nsew signal input
flabel metal2 s 14922 44540 14978 45000 0 FreeSans 224 90 0 0 S4END[9]
port 343 nsew signal input
flabel metal2 s 16210 -300 16266 160 0 FreeSans 224 90 0 0 UserCLK
port 344 nsew signal input
flabel metal2 s 16210 44540 16266 45000 0 FreeSans 224 90 0 0 UserCLKo
port 345 nsew signal tristate
flabel metal4 s 6142 1040 6462 43568 0 FreeSans 1920 90 0 0 VGND
port 346 nsew ground bidirectional
flabel metal4 s 11340 1040 11660 43568 0 FreeSans 1920 90 0 0 VGND
port 346 nsew ground bidirectional
flabel metal4 s 16538 1040 16858 43568 0 FreeSans 1920 90 0 0 VGND
port 346 nsew ground bidirectional
flabel metal4 s 21736 1040 22056 43568 0 FreeSans 1920 90 0 0 VGND
port 346 nsew ground bidirectional
flabel metal4 s 3543 1040 3863 43568 0 FreeSans 1920 90 0 0 VPWR
port 347 nsew power bidirectional
flabel metal4 s 8741 1040 9061 43568 0 FreeSans 1920 90 0 0 VPWR
port 347 nsew power bidirectional
flabel metal4 s 13939 1040 14259 43568 0 FreeSans 1920 90 0 0 VPWR
port 347 nsew power bidirectional
flabel metal4 s 19137 1040 19457 43568 0 FreeSans 1920 90 0 0 VPWR
port 347 nsew power bidirectional
flabel metal3 s -300 4904 160 5024 0 FreeSans 480 0 0 0 W1BEG[0]
port 348 nsew signal tristate
flabel metal3 s -300 5176 160 5296 0 FreeSans 480 0 0 0 W1BEG[1]
port 349 nsew signal tristate
flabel metal3 s -300 5448 160 5568 0 FreeSans 480 0 0 0 W1BEG[2]
port 350 nsew signal tristate
flabel metal3 s -300 5720 160 5840 0 FreeSans 480 0 0 0 W1BEG[3]
port 351 nsew signal tristate
flabel metal3 s -300 5992 160 6112 0 FreeSans 480 0 0 0 W2BEG[0]
port 352 nsew signal tristate
flabel metal3 s -300 6264 160 6384 0 FreeSans 480 0 0 0 W2BEG[1]
port 353 nsew signal tristate
flabel metal3 s -300 6536 160 6656 0 FreeSans 480 0 0 0 W2BEG[2]
port 354 nsew signal tristate
flabel metal3 s -300 6808 160 6928 0 FreeSans 480 0 0 0 W2BEG[3]
port 355 nsew signal tristate
flabel metal3 s -300 7080 160 7200 0 FreeSans 480 0 0 0 W2BEG[4]
port 356 nsew signal tristate
flabel metal3 s -300 7352 160 7472 0 FreeSans 480 0 0 0 W2BEG[5]
port 357 nsew signal tristate
flabel metal3 s -300 7624 160 7744 0 FreeSans 480 0 0 0 W2BEG[6]
port 358 nsew signal tristate
flabel metal3 s -300 7896 160 8016 0 FreeSans 480 0 0 0 W2BEG[7]
port 359 nsew signal tristate
flabel metal3 s -300 8168 160 8288 0 FreeSans 480 0 0 0 W2BEGb[0]
port 360 nsew signal tristate
flabel metal3 s -300 8440 160 8560 0 FreeSans 480 0 0 0 W2BEGb[1]
port 361 nsew signal tristate
flabel metal3 s -300 8712 160 8832 0 FreeSans 480 0 0 0 W2BEGb[2]
port 362 nsew signal tristate
flabel metal3 s -300 8984 160 9104 0 FreeSans 480 0 0 0 W2BEGb[3]
port 363 nsew signal tristate
flabel metal3 s -300 9256 160 9376 0 FreeSans 480 0 0 0 W2BEGb[4]
port 364 nsew signal tristate
flabel metal3 s -300 9528 160 9648 0 FreeSans 480 0 0 0 W2BEGb[5]
port 365 nsew signal tristate
flabel metal3 s -300 9800 160 9920 0 FreeSans 480 0 0 0 W2BEGb[6]
port 366 nsew signal tristate
flabel metal3 s -300 10072 160 10192 0 FreeSans 480 0 0 0 W2BEGb[7]
port 367 nsew signal tristate
flabel metal3 s -300 14696 160 14816 0 FreeSans 480 0 0 0 W6BEG[0]
port 368 nsew signal tristate
flabel metal3 s -300 17416 160 17536 0 FreeSans 480 0 0 0 W6BEG[10]
port 369 nsew signal tristate
flabel metal3 s -300 17688 160 17808 0 FreeSans 480 0 0 0 W6BEG[11]
port 370 nsew signal tristate
flabel metal3 s -300 14968 160 15088 0 FreeSans 480 0 0 0 W6BEG[1]
port 371 nsew signal tristate
flabel metal3 s -300 15240 160 15360 0 FreeSans 480 0 0 0 W6BEG[2]
port 372 nsew signal tristate
flabel metal3 s -300 15512 160 15632 0 FreeSans 480 0 0 0 W6BEG[3]
port 373 nsew signal tristate
flabel metal3 s -300 15784 160 15904 0 FreeSans 480 0 0 0 W6BEG[4]
port 374 nsew signal tristate
flabel metal3 s -300 16056 160 16176 0 FreeSans 480 0 0 0 W6BEG[5]
port 375 nsew signal tristate
flabel metal3 s -300 16328 160 16448 0 FreeSans 480 0 0 0 W6BEG[6]
port 376 nsew signal tristate
flabel metal3 s -300 16600 160 16720 0 FreeSans 480 0 0 0 W6BEG[7]
port 377 nsew signal tristate
flabel metal3 s -300 16872 160 16992 0 FreeSans 480 0 0 0 W6BEG[8]
port 378 nsew signal tristate
flabel metal3 s -300 17144 160 17264 0 FreeSans 480 0 0 0 W6BEG[9]
port 379 nsew signal tristate
flabel metal3 s -300 10344 160 10464 0 FreeSans 480 0 0 0 WW4BEG[0]
port 380 nsew signal tristate
flabel metal3 s -300 13064 160 13184 0 FreeSans 480 0 0 0 WW4BEG[10]
port 381 nsew signal tristate
flabel metal3 s -300 13336 160 13456 0 FreeSans 480 0 0 0 WW4BEG[11]
port 382 nsew signal tristate
flabel metal3 s -300 13608 160 13728 0 FreeSans 480 0 0 0 WW4BEG[12]
port 383 nsew signal tristate
flabel metal3 s -300 13880 160 14000 0 FreeSans 480 0 0 0 WW4BEG[13]
port 384 nsew signal tristate
flabel metal3 s -300 14152 160 14272 0 FreeSans 480 0 0 0 WW4BEG[14]
port 385 nsew signal tristate
flabel metal3 s -300 14424 160 14544 0 FreeSans 480 0 0 0 WW4BEG[15]
port 386 nsew signal tristate
flabel metal3 s -300 10616 160 10736 0 FreeSans 480 0 0 0 WW4BEG[1]
port 387 nsew signal tristate
flabel metal3 s -300 10888 160 11008 0 FreeSans 480 0 0 0 WW4BEG[2]
port 388 nsew signal tristate
flabel metal3 s -300 11160 160 11280 0 FreeSans 480 0 0 0 WW4BEG[3]
port 389 nsew signal tristate
flabel metal3 s -300 11432 160 11552 0 FreeSans 480 0 0 0 WW4BEG[4]
port 390 nsew signal tristate
flabel metal3 s -300 11704 160 11824 0 FreeSans 480 0 0 0 WW4BEG[5]
port 391 nsew signal tristate
flabel metal3 s -300 11976 160 12096 0 FreeSans 480 0 0 0 WW4BEG[6]
port 392 nsew signal tristate
flabel metal3 s -300 12248 160 12368 0 FreeSans 480 0 0 0 WW4BEG[7]
port 393 nsew signal tristate
flabel metal3 s -300 12520 160 12640 0 FreeSans 480 0 0 0 WW4BEG[8]
port 394 nsew signal tristate
flabel metal3 s -300 12792 160 12912 0 FreeSans 480 0 0 0 WW4BEG[9]
port 395 nsew signal tristate
rlabel via1 11580 43520 11580 43520 0 VGND
rlabel metal1 11500 42976 11500 42976 0 VPWR
rlabel metal2 21482 9231 21482 9231 0 Config_accessC_bit0
rlabel metal3 22594 9860 22594 9860 0 Config_accessC_bit1
rlabel metal2 20930 10319 20930 10319 0 Config_accessC_bit2
rlabel metal1 21850 10778 21850 10778 0 Config_accessC_bit3
rlabel metal3 820 18020 820 18020 0 E1END[0]
rlabel metal3 1004 18292 1004 18292 0 E1END[1]
rlabel metal3 544 18564 544 18564 0 E1END[2]
rlabel metal3 636 18836 636 18836 0 E1END[3]
rlabel metal3 820 21284 820 21284 0 E2END[0]
rlabel metal3 452 21556 452 21556 0 E2END[1]
rlabel metal3 682 21828 682 21828 0 E2END[2]
rlabel metal3 774 22100 774 22100 0 E2END[3]
rlabel metal3 1234 22372 1234 22372 0 E2END[4]
rlabel metal3 636 22644 636 22644 0 E2END[5]
rlabel metal3 728 22916 728 22916 0 E2END[6]
rlabel metal2 2806 23409 2806 23409 0 E2END[7]
rlabel metal2 2898 19227 2898 19227 0 E2MID[0]
rlabel metal2 3266 19091 3266 19091 0 E2MID[1]
rlabel metal3 958 19652 958 19652 0 E2MID[2]
rlabel metal3 452 19924 452 19924 0 E2MID[3]
rlabel metal3 820 20196 820 20196 0 E2MID[4]
rlabel metal2 3266 21165 3266 21165 0 E2MID[5]
rlabel metal3 728 20740 728 20740 0 E2MID[6]
rlabel metal3 452 21012 452 21012 0 E2MID[7]
rlabel metal3 452 27812 452 27812 0 E6END[0]
rlabel metal2 1610 32708 1610 32708 0 E6END[10]
rlabel metal2 4094 30957 4094 30957 0 E6END[11]
rlabel metal2 2990 28611 2990 28611 0 E6END[1]
rlabel metal3 774 28356 774 28356 0 E6END[2]
rlabel metal2 3818 28679 3818 28679 0 E6END[3]
rlabel metal3 452 28900 452 28900 0 E6END[4]
rlabel metal3 820 29172 820 29172 0 E6END[5]
rlabel metal2 3542 29529 3542 29529 0 E6END[6]
rlabel metal2 2806 30209 2806 30209 0 E6END[7]
rlabel metal3 452 29988 452 29988 0 E6END[8]
rlabel metal3 751 30260 751 30260 0 E6END[9]
rlabel metal3 774 23460 774 23460 0 EE4END[0]
rlabel metal3 406 26180 406 26180 0 EE4END[10]
rlabel metal3 958 26452 958 26452 0 EE4END[11]
rlabel metal3 682 26724 682 26724 0 EE4END[12]
rlabel metal3 728 26996 728 26996 0 EE4END[13]
rlabel metal3 728 27268 728 27268 0 EE4END[14]
rlabel metal3 820 27540 820 27540 0 EE4END[15]
rlabel metal3 452 23732 452 23732 0 EE4END[1]
rlabel metal3 866 24004 866 24004 0 EE4END[2]
rlabel metal3 452 24276 452 24276 0 EE4END[3]
rlabel metal2 3266 24905 3266 24905 0 EE4END[4]
rlabel metal3 498 24820 498 24820 0 EE4END[5]
rlabel metal3 820 25092 820 25092 0 EE4END[6]
rlabel metal2 2806 25789 2806 25789 0 EE4END[7]
rlabel metal2 3082 25993 3082 25993 0 EE4END[8]
rlabel metal3 1441 25908 1441 25908 0 EE4END[9]
rlabel metal3 22180 15844 22180 15844 0 FAB2RAM_A0_O0
rlabel metal3 22525 16388 22525 16388 0 FAB2RAM_A0_O1
rlabel metal3 22180 16932 22180 16932 0 FAB2RAM_A0_O2
rlabel metal3 22548 17476 22548 17476 0 FAB2RAM_A0_O3
rlabel metal3 22180 13668 22180 13668 0 FAB2RAM_A1_O0
rlabel metal3 22548 14212 22548 14212 0 FAB2RAM_A1_O1
rlabel metal3 22180 14756 22180 14756 0 FAB2RAM_A1_O2
rlabel metal3 22732 15300 22732 15300 0 FAB2RAM_A1_O3
rlabel metal3 21996 11492 21996 11492 0 FAB2RAM_C_O0
rlabel metal3 22548 12036 22548 12036 0 FAB2RAM_C_O1
rlabel metal3 21996 12580 21996 12580 0 FAB2RAM_C_O2
rlabel metal3 22548 13124 22548 13124 0 FAB2RAM_C_O3
rlabel metal3 22180 24548 22180 24548 0 FAB2RAM_D0_O0
rlabel metal3 22594 25092 22594 25092 0 FAB2RAM_D0_O1
rlabel metal3 22180 25636 22180 25636 0 FAB2RAM_D0_O2
rlabel metal3 22594 26180 22594 26180 0 FAB2RAM_D0_O3
rlabel metal2 21482 22287 21482 22287 0 FAB2RAM_D1_O0
rlabel metal1 21666 22746 21666 22746 0 FAB2RAM_D1_O1
rlabel metal1 21528 23290 21528 23290 0 FAB2RAM_D1_O2
rlabel metal3 22548 24004 22548 24004 0 FAB2RAM_D1_O3
rlabel metal3 22180 20196 22180 20196 0 FAB2RAM_D2_O0
rlabel metal3 22548 20740 22548 20740 0 FAB2RAM_D2_O1
rlabel metal1 20792 21114 20792 21114 0 FAB2RAM_D2_O2
rlabel metal1 21666 21862 21666 21862 0 FAB2RAM_D2_O3
rlabel metal3 22180 18020 22180 18020 0 FAB2RAM_D3_O0
rlabel metal3 22548 18564 22548 18564 0 FAB2RAM_D3_O1
rlabel metal3 22180 19108 22180 19108 0 FAB2RAM_D3_O2
rlabel metal3 22548 19652 22548 19652 0 FAB2RAM_D3_O3
rlabel metal3 1418 31076 1418 31076 0 FrameData[0]
rlabel metal2 3174 34697 3174 34697 0 FrameData[10]
rlabel metal2 4094 34527 4094 34527 0 FrameData[11]
rlabel metal3 1441 34340 1441 34340 0 FrameData[12]
rlabel metal3 820 34612 820 34612 0 FrameData[13]
rlabel metal3 475 34884 475 34884 0 FrameData[14]
rlabel metal2 3082 36193 3082 36193 0 FrameData[15]
rlabel metal3 1671 35428 1671 35428 0 FrameData[16]
rlabel metal3 222 35700 222 35700 0 FrameData[17]
rlabel metal3 567 35972 567 35972 0 FrameData[18]
rlabel metal2 2898 36720 2898 36720 0 FrameData[19]
rlabel metal3 1970 31348 1970 31348 0 FrameData[1]
rlabel metal3 1671 36516 1671 36516 0 FrameData[20]
rlabel metal3 475 36788 475 36788 0 FrameData[21]
rlabel metal3 751 37060 751 37060 0 FrameData[22]
rlabel metal2 2714 39695 2714 39695 0 FrameData[23]
rlabel metal3 728 37604 728 37604 0 FrameData[24]
rlabel metal3 452 37876 452 37876 0 FrameData[25]
rlabel metal1 1978 41038 1978 41038 0 FrameData[26]
rlabel metal3 1096 38420 1096 38420 0 FrameData[27]
rlabel metal3 636 38692 636 38692 0 FrameData[28]
rlabel metal3 728 38964 728 38964 0 FrameData[29]
rlabel metal2 1472 32572 1472 32572 0 FrameData[2]
rlabel metal3 1556 39236 1556 39236 0 FrameData[30]
rlabel metal2 2806 40307 2806 40307 0 FrameData[31]
rlabel metal3 452 31892 452 31892 0 FrameData[3]
rlabel metal3 1004 32164 1004 32164 0 FrameData[4]
rlabel metal3 1004 32436 1004 32436 0 FrameData[5]
rlabel metal2 2990 33337 2990 33337 0 FrameData[6]
rlabel metal2 3358 33473 3358 33473 0 FrameData[7]
rlabel metal3 820 33252 820 33252 0 FrameData[8]
rlabel metal3 3404 33592 3404 33592 0 FrameData[9]
rlabel metal3 22180 26724 22180 26724 0 FrameData_O[0]
rlabel metal3 22180 32164 22180 32164 0 FrameData_O[10]
rlabel metal3 22525 32708 22525 32708 0 FrameData_O[11]
rlabel metal3 22088 33252 22088 33252 0 FrameData_O[12]
rlabel metal3 22548 33796 22548 33796 0 FrameData_O[13]
rlabel metal3 22180 34340 22180 34340 0 FrameData_O[14]
rlabel metal3 22548 34884 22548 34884 0 FrameData_O[15]
rlabel metal3 22180 35428 22180 35428 0 FrameData_O[16]
rlabel metal3 22594 35972 22594 35972 0 FrameData_O[17]
rlabel metal3 22180 36516 22180 36516 0 FrameData_O[18]
rlabel metal3 22594 37060 22594 37060 0 FrameData_O[19]
rlabel metal3 22548 27268 22548 27268 0 FrameData_O[1]
rlabel metal3 22180 37604 22180 37604 0 FrameData_O[20]
rlabel metal3 22548 38148 22548 38148 0 FrameData_O[21]
rlabel metal3 22180 38692 22180 38692 0 FrameData_O[22]
rlabel metal3 22548 39236 22548 39236 0 FrameData_O[23]
rlabel metal3 22180 39780 22180 39780 0 FrameData_O[24]
rlabel metal3 22548 40324 22548 40324 0 FrameData_O[25]
rlabel metal3 22548 40868 22548 40868 0 FrameData_O[26]
rlabel metal3 22594 41412 22594 41412 0 FrameData_O[27]
rlabel metal1 21436 41786 21436 41786 0 FrameData_O[28]
rlabel metal1 21206 42330 21206 42330 0 FrameData_O[29]
rlabel metal3 21996 27812 21996 27812 0 FrameData_O[2]
rlabel metal2 20562 42415 20562 42415 0 FrameData_O[30]
rlabel metal1 21896 42262 21896 42262 0 FrameData_O[31]
rlabel metal3 22548 28356 22548 28356 0 FrameData_O[3]
rlabel metal3 22180 28900 22180 28900 0 FrameData_O[4]
rlabel metal3 22548 29444 22548 29444 0 FrameData_O[5]
rlabel metal3 22180 29988 22180 29988 0 FrameData_O[6]
rlabel metal3 22594 30532 22594 30532 0 FrameData_O[7]
rlabel metal3 22180 31076 22180 31076 0 FrameData_O[8]
rlabel metal1 21850 31654 21850 31654 0 FrameData_O[9]
rlabel metal2 18676 1326 18676 1326 0 FrameStrobe[0]
rlabel metal2 18315 68 18315 68 0 FrameStrobe[10]
rlabel metal2 18499 68 18499 68 0 FrameStrobe[11]
rlabel metal2 18630 636 18630 636 0 FrameStrobe[12]
rlabel metal2 18814 1044 18814 1044 0 FrameStrobe[13]
rlabel metal2 18998 976 18998 976 0 FrameStrobe[14]
rlabel metal2 19129 68 19129 68 0 FrameStrobe[15]
rlabel metal2 19419 68 19419 68 0 FrameStrobe[16]
rlabel metal2 19603 68 19603 68 0 FrameStrobe[17]
rlabel metal2 19787 68 19787 68 0 FrameStrobe[18]
rlabel metal2 20109 68 20109 68 0 FrameStrobe[19]
rlabel metal2 16659 68 16659 68 0 FrameStrobe[1]
rlabel metal2 16843 68 16843 68 0 FrameStrobe[2]
rlabel metal2 16974 143 16974 143 0 FrameStrobe[3]
rlabel metal2 17211 68 17211 68 0 FrameStrobe[4]
rlabel metal1 15686 1258 15686 1258 0 FrameStrobe[5]
rlabel metal2 17579 68 17579 68 0 FrameStrobe[6]
rlabel metal2 17710 670 17710 670 0 FrameStrobe[7]
rlabel metal2 17894 1010 17894 1010 0 FrameStrobe[8]
rlabel metal2 18078 1316 18078 1316 0 FrameStrobe[9]
rlabel metal2 16422 43921 16422 43921 0 FrameStrobe_O[0]
rlabel metal1 19481 42738 19481 42738 0 FrameStrobe_O[10]
rlabel metal2 18446 43972 18446 43972 0 FrameStrobe_O[11]
rlabel metal2 18630 44193 18630 44193 0 FrameStrobe_O[12]
rlabel metal2 18814 44261 18814 44261 0 FrameStrobe_O[13]
rlabel metal2 18998 44074 18998 44074 0 FrameStrobe_O[14]
rlabel metal2 19182 43904 19182 43904 0 FrameStrobe_O[15]
rlabel metal2 19366 44193 19366 44193 0 FrameStrobe_O[16]
rlabel metal2 19550 43700 19550 43700 0 FrameStrobe_O[17]
rlabel metal2 19734 43904 19734 43904 0 FrameStrobe_O[18]
rlabel metal2 19918 44057 19918 44057 0 FrameStrobe_O[19]
rlabel metal1 17204 43418 17204 43418 0 FrameStrobe_O[1]
rlabel metal2 17802 43622 17802 43622 0 FrameStrobe_O[2]
rlabel metal1 17710 42330 17710 42330 0 FrameStrobe_O[3]
rlabel metal2 17158 43700 17158 43700 0 FrameStrobe_O[4]
rlabel metal2 17342 43938 17342 43938 0 FrameStrobe_O[5]
rlabel metal2 17526 43700 17526 43700 0 FrameStrobe_O[6]
rlabel metal2 17710 43836 17710 43836 0 FrameStrobe_O[7]
rlabel metal2 17894 43649 17894 43649 0 FrameStrobe_O[8]
rlabel metal2 18078 43904 18078 43904 0 FrameStrobe_O[9]
rlabel metal1 21390 6800 21390 6800 0 Inst_Config_accessConfig_access.ConfigBits\[0\]
rlabel metal1 21114 8466 21114 8466 0 Inst_Config_accessConfig_access.ConfigBits\[1\]
rlabel metal1 20056 9690 20056 9690 0 Inst_Config_accessConfig_access.ConfigBits\[2\]
rlabel metal1 20240 10778 20240 10778 0 Inst_Config_accessConfig_access.ConfigBits\[3\]
rlabel metal1 20700 16218 20700 16218 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.ConfigBits\[0\]
rlabel metal1 16054 37264 16054 37264 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.ConfigBits\[1\]
rlabel metal1 20378 17578 20378 17578 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.ConfigBits\[2\]
rlabel metal1 17204 35258 17204 35258 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.ConfigBits\[3\]
rlabel metal1 19734 17646 19734 17646 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.I\[0\]
rlabel metal1 7498 37230 7498 37230 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.I\[1\]
rlabel metal1 18476 18326 18476 18326 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.I\[2\]
rlabel metal1 14290 34986 14290 34986 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.I\[3\]
rlabel metal1 19182 17204 19182 17204 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.Q\[0\]
rlabel metal1 16468 37230 16468 37230 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.Q\[1\]
rlabel metal1 20838 17170 20838 17170 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.Q\[2\]
rlabel metal1 16376 34578 16376 34578 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.Q\[3\]
rlabel metal1 20930 16082 20930 16082 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst0.AIN\[0\]
rlabel metal1 21022 15504 21022 15504 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst0.AIN\[1\]
rlabel metal2 21114 16388 21114 16388 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst0._0_
rlabel metal2 20930 16150 20930 16150 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst0._1_
rlabel metal1 15318 36890 15318 36890 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst1.AIN\[0\]
rlabel metal1 16284 37230 16284 37230 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst1.AIN\[1\]
rlabel metal1 15778 36754 15778 36754 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst1._0_
rlabel metal1 16100 36822 16100 36822 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst1._1_
rlabel metal1 20010 17612 20010 17612 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst2.AIN\[0\]
rlabel metal1 21206 17204 21206 17204 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst2.AIN\[1\]
rlabel metal1 20286 17714 20286 17714 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst2._0_
rlabel metal1 20884 16966 20884 16966 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst2._1_
rlabel metal1 15640 34578 15640 34578 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst3.AIN\[0\]
rlabel metal1 16376 34714 16376 34714 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst3.AIN\[1\]
rlabel metal2 16054 35190 16054 35190 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst3._0_
rlabel metal1 17526 35666 17526 35666 0 Inst_FAB2RAM_A0_OutPass4_frame_config_mux.cus_mux21_inst3._1_
rlabel metal1 20930 14484 20930 14484 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.ConfigBits\[0\]
rlabel metal1 18860 15470 18860 15470 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.ConfigBits\[1\]
rlabel metal1 20332 35258 20332 35258 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.ConfigBits\[2\]
rlabel metal1 18170 36618 18170 36618 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.ConfigBits\[3\]
rlabel metal1 19683 15470 19683 15470 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.I\[0\]
rlabel metal1 17204 15470 17204 15470 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.I\[1\]
rlabel metal1 18614 35734 18614 35734 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.I\[2\]
rlabel metal1 16734 36754 16734 36754 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.I\[3\]
rlabel metal1 20792 14994 20792 14994 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.Q\[0\]
rlabel metal2 18722 15844 18722 15844 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.Q\[1\]
rlabel metal1 20424 35530 20424 35530 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.Q\[2\]
rlabel metal1 17986 36890 17986 36890 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.Q\[3\]
rlabel metal1 20286 14960 20286 14960 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst0.AIN\[0\]
rlabel metal1 21114 14960 21114 14960 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst0.AIN\[1\]
rlabel metal1 21022 14348 21022 14348 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst0._0_
rlabel metal1 21114 14450 21114 14450 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst0._1_
rlabel metal1 17710 15674 17710 15674 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst1.AIN\[0\]
rlabel metal1 19274 16116 19274 16116 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst1.AIN\[1\]
rlabel metal1 18676 15674 18676 15674 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst1._0_
rlabel metal1 19090 15606 19090 15606 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst1._1_
rlabel metal1 18998 35054 18998 35054 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst2.AIN\[0\]
rlabel viali 20562 36756 20562 36756 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst2.AIN\[1\]
rlabel metal1 19734 34952 19734 34952 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst2._0_
rlabel metal1 21068 35054 21068 35054 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst2._1_
rlabel metal2 16606 36618 16606 36618 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst3.AIN\[0\]
rlabel metal1 18170 37196 18170 37196 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst3.AIN\[1\]
rlabel metal1 17848 36754 17848 36754 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst3._0_
rlabel metal1 18446 36822 18446 36822 0 Inst_FAB2RAM_A1_OutPass4_frame_config_mux.cus_mux21_inst3._1_
rlabel via1 19550 12818 19550 12818 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.ConfigBits\[0\]
rlabel metal1 20102 30022 20102 30022 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.ConfigBits\[1\]
rlabel metal1 20976 12818 20976 12818 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.ConfigBits\[2\]
rlabel metal1 20700 32878 20700 32878 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.ConfigBits\[3\]
rlabel metal1 18257 13294 18257 13294 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.I\[0\]
rlabel metal1 19637 30634 19637 30634 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.I\[1\]
rlabel metal1 19913 13906 19913 13906 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.I\[2\]
rlabel metal1 19637 32810 19637 32810 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.I\[3\]
rlabel metal1 20286 12852 20286 12852 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.Q\[0\]
rlabel metal1 21022 32538 21022 32538 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.Q\[1\]
rlabel metal2 21160 13124 21160 13124 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.Q\[2\]
rlabel metal1 20792 32742 20792 32742 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.Q\[3\]
rlabel metal1 19136 13498 19136 13498 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst0.AIN\[0\]
rlabel metal1 19642 12240 19642 12240 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst0.AIN\[1\]
rlabel metal2 19826 13396 19826 13396 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst0._0_
rlabel metal1 19780 12410 19780 12410 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst0._1_
rlabel metal1 19688 31450 19688 31450 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst1.AIN\[0\]
rlabel metal1 21390 33014 21390 33014 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst1.AIN\[1\]
rlabel metal1 20884 29818 20884 29818 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst1._0_
rlabel metal1 20148 29682 20148 29682 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst1._1_
rlabel metal1 20470 12886 20470 12886 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst2.AIN\[0\]
rlabel metal1 20930 11866 20930 11866 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst2.AIN\[1\]
rlabel metal1 20976 12682 20976 12682 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst2._0_
rlabel metal1 21252 12750 21252 12750 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst2._1_
rlabel metal1 20056 33354 20056 33354 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst3.AIN\[0\]
rlabel metal1 20792 33966 20792 33966 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst3.AIN\[1\]
rlabel metal2 20792 32878 20792 32878 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst3._0_
rlabel metal1 20930 32946 20930 32946 0 Inst_FAB2RAM_C_OutPass4_frame_config_mux.cus_mux21_inst3._1_
rlabel metal1 18768 24786 18768 24786 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.ConfigBits\[0\]
rlabel metal1 17986 32844 17986 32844 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.ConfigBits\[1\]
rlabel metal1 19734 25262 19734 25262 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.ConfigBits\[2\]
rlabel metal1 17526 26826 17526 26826 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.ConfigBits\[3\]
rlabel metal1 17516 24786 17516 24786 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.I\[0\]
rlabel metal1 16882 33456 16882 33456 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.I\[1\]
rlabel via2 4554 25755 4554 25755 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.I\[2\]
rlabel metal1 16192 28050 16192 28050 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.I\[3\]
rlabel metal1 18814 24922 18814 24922 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.Q\[0\]
rlabel metal1 18446 32878 18446 32878 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.Q\[1\]
rlabel metal2 19182 26146 19182 26146 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.Q\[2\]
rlabel metal1 17894 27404 17894 27404 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.Q\[3\]
rlabel metal1 19090 24786 19090 24786 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst0.AIN\[0\]
rlabel metal1 18676 25262 18676 25262 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst0.AIN\[1\]
rlabel metal1 19090 24650 19090 24650 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst0._0_
rlabel metal1 18860 24718 18860 24718 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst0._1_
rlabel metal1 17342 33524 17342 33524 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst1.AIN\[0\]
rlabel metal1 18768 32878 18768 32878 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst1.AIN\[1\]
rlabel metal2 18078 33184 18078 33184 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst1._0_
rlabel metal1 18354 32946 18354 32946 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst1._1_
rlabel metal1 19274 26384 19274 26384 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst2.AIN\[0\]
rlabel metal1 20010 25330 20010 25330 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst2.AIN\[1\]
rlabel metal2 19550 25908 19550 25908 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst2._0_
rlabel metal1 19826 25330 19826 25330 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst2._1_
rlabel metal1 16928 26350 16928 26350 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst3.AIN\[0\]
rlabel metal1 18262 26996 18262 26996 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst3.AIN\[1\]
rlabel metal1 17480 26554 17480 26554 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst3._0_
rlabel metal2 18170 27302 18170 27302 0 Inst_FAB2RAM_D0_OutPass4_frame_config_mux.cus_mux21_inst3._1_
rlabel metal1 18906 23052 18906 23052 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.ConfigBits\[0\]
rlabel metal1 19274 28492 19274 28492 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.ConfigBits\[1\]
rlabel metal1 20700 24174 20700 24174 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.ConfigBits\[2\]
rlabel metal1 18354 28050 18354 28050 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.ConfigBits\[3\]
rlabel via1 18165 22610 18165 22610 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.I\[0\]
rlabel metal1 17326 28458 17326 28458 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.I\[1\]
rlabel metal1 20286 25228 20286 25228 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.I\[2\]
rlabel metal1 17250 29614 17250 29614 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.I\[3\]
rlabel metal2 19458 22848 19458 22848 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.Q\[0\]
rlabel metal1 20378 28628 20378 28628 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.Q\[1\]
rlabel metal1 20976 24922 20976 24922 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.Q\[2\]
rlabel metal1 18124 29274 18124 29274 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.Q\[3\]
rlabel metal1 18630 21998 18630 21998 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst0.AIN\[0\]
rlabel metal1 19182 23086 19182 23086 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst0.AIN\[1\]
rlabel metal1 19596 21862 19596 21862 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst0._0_
rlabel metal1 19090 22712 19090 22712 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst0._1_
rlabel metal1 19182 28084 19182 28084 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst1.AIN\[0\]
rlabel metal1 20148 28526 20148 28526 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst1.AIN\[1\]
rlabel metal1 19320 28186 19320 28186 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst1._0_
rlabel metal1 19780 28594 19780 28594 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst1._1_
rlabel metal2 20102 25636 20102 25636 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst2.AIN\[0\]
rlabel metal1 20700 25262 20700 25262 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst2.AIN\[1\]
rlabel metal1 20976 24378 20976 24378 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst2._0_
rlabel metal1 20838 24242 20838 24242 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst2._1_
rlabel metal1 17342 28526 17342 28526 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst3.AIN\[0\]
rlabel metal1 19090 28118 19090 28118 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst3.AIN\[1\]
rlabel metal1 18630 28084 18630 28084 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst3._0_
rlabel metal1 18906 27982 18906 27982 0 Inst_FAB2RAM_D1_OutPass4_frame_config_mux.cus_mux21_inst3._1_
rlabel metal1 20976 21522 20976 21522 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.ConfigBits\[0\]
rlabel metal1 18446 31756 18446 31756 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.ConfigBits\[1\]
rlabel metal1 19090 23630 19090 23630 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.ConfigBits\[2\]
rlabel metal1 16836 29614 16836 29614 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.ConfigBits\[3\]
rlabel metal1 17250 23256 17250 23256 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.I\[0\]
rlabel metal1 7130 30600 7130 30600 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.I\[1\]
rlabel metal1 19458 23698 19458 23698 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.I\[2\]
rlabel metal2 16238 29444 16238 29444 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.I\[3\]
rlabel metal1 20930 21862 20930 21862 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.Q\[0\]
rlabel metal1 18216 31450 18216 31450 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.Q\[1\]
rlabel metal1 20608 24038 20608 24038 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.Q\[2\]
rlabel metal1 17204 30702 17204 30702 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.Q\[3\]
rlabel metal1 20700 20910 20700 20910 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst0.AIN\[0\]
rlabel metal1 21160 19822 21160 19822 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst0.AIN\[1\]
rlabel metal1 20378 21114 20378 21114 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst0._0_
rlabel metal1 21206 19754 21206 19754 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst0._1_
rlabel metal1 17802 30736 17802 30736 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst1.AIN\[0\]
rlabel metal1 18630 31858 18630 31858 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst1.AIN\[1\]
rlabel metal1 18078 30770 18078 30770 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst1._0_
rlabel metal1 18492 30770 18492 30770 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst1._1_
rlabel metal1 21390 23732 21390 23732 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst2.AIN\[0\]
rlabel metal2 19274 23987 19274 23987 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst2.AIN\[1\]
rlabel metal1 21298 23562 21298 23562 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst2._0_
rlabel metal1 20792 23630 20792 23630 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst2._1_
rlabel metal1 16468 29614 16468 29614 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst3.AIN\[0\]
rlabel metal1 16514 30260 16514 30260 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst3.AIN\[1\]
rlabel metal1 16836 29750 16836 29750 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst3._0_
rlabel metal1 16790 29682 16790 29682 0 Inst_FAB2RAM_D2_OutPass4_frame_config_mux.cus_mux21_inst3._1_
rlabel metal1 20470 18598 20470 18598 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.ConfigBits\[0\]
rlabel metal1 20838 26962 20838 26962 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.ConfigBits\[1\]
rlabel metal1 21022 18734 21022 18734 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.ConfigBits\[2\]
rlabel metal1 17940 33966 17940 33966 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.ConfigBits\[3\]
rlabel metal2 19090 20570 19090 20570 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.I\[0\]
rlabel metal1 19918 28016 19918 28016 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.I\[1\]
rlabel metal1 18630 19822 18630 19822 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.I\[2\]
rlabel metal1 16785 33898 16785 33898 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.I\[3\]
rlabel metal1 20332 20026 20332 20026 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.Q\[0\]
rlabel metal1 20746 27574 20746 27574 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.Q\[1\]
rlabel metal1 20838 18292 20838 18292 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.Q\[2\]
rlabel metal1 18583 33966 18583 33966 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.Q\[3\]
rlabel metal1 18860 19346 18860 19346 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst0.AIN\[0\]
rlabel metal1 21114 17680 21114 17680 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst0.AIN\[1\]
rlabel metal1 20332 19210 20332 19210 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst0._0_
rlabel metal1 20930 19278 20930 19278 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst0._1_
rlabel metal1 20378 26316 20378 26316 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst1.AIN\[0\]
rlabel metal1 20976 26350 20976 26350 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst1.AIN\[1\]
rlabel metal2 20470 26656 20470 26656 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst1._0_
rlabel metal1 21114 26554 21114 26554 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst1._1_
rlabel metal1 20148 18734 20148 18734 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst2.AIN\[0\]
rlabel metal1 20608 18258 20608 18258 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst2.AIN\[1\]
rlabel metal1 20884 18802 20884 18802 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst2._0_
rlabel metal2 20562 18530 20562 18530 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst2._1_
rlabel metal1 18170 33966 18170 33966 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst3.AIN\[0\]
rlabel metal1 18998 33932 18998 33932 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst3.AIN\[1\]
rlabel metal1 18078 33898 18078 33898 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst3._0_
rlabel metal1 18170 34068 18170 34068 0 Inst_FAB2RAM_D3_OutPass4_frame_config_mux.cus_mux21_inst3._1_
rlabel metal1 20286 11628 20286 11628 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.ConfigBits\[0\]
rlabel metal1 17802 12070 17802 12070 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.ConfigBits\[1\]
rlabel metal1 19688 6766 19688 6766 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.ConfigBits\[2\]
rlabel metal1 17526 8806 17526 8806 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.ConfigBits\[3\]
rlabel metal2 21022 11407 21022 11407 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.O\[0\]
rlabel metal1 2576 9554 2576 9554 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.O\[1\]
rlabel metal1 20562 6936 20562 6936 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.O\[2\]
rlabel metal1 14122 14926 14122 14926 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.O\[3\]
rlabel metal1 21206 8976 21206 8976 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.Q\[0\]
rlabel metal1 18860 11118 18860 11118 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.Q\[1\]
rlabel metal1 21482 5678 21482 5678 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.Q\[2\]
rlabel metal1 18676 8602 18676 8602 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.Q\[3\]
rlabel metal2 19734 11186 19734 11186 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst0.AIN\[0\]
rlabel metal2 21022 9809 21022 9809 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst0.AIN\[1\]
rlabel metal2 19826 11526 19826 11526 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst0._0_
rlabel metal1 21022 11764 21022 11764 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst0._1_
rlabel metal1 16974 11764 16974 11764 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst1.AIN\[0\]
rlabel metal1 18584 11322 18584 11322 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst1.AIN\[1\]
rlabel metal2 17894 11322 17894 11322 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst1._0_
rlabel metal2 18354 11594 18354 11594 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst1._1_
rlabel metal1 19458 6732 19458 6732 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst2.AIN\[0\]
rlabel metal1 21252 5882 21252 5882 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst2.AIN\[1\]
rlabel metal1 20102 6800 20102 6800 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst2._0_
rlabel metal1 20654 6800 20654 6800 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst2._1_
rlabel metal1 17204 7854 17204 7854 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst3.AIN\[0\]
rlabel metal1 18768 8942 18768 8942 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst3.AIN\[1\]
rlabel metal1 17388 7378 17388 7378 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst3._0_
rlabel metal1 17618 7412 17618 7412 0 Inst_RAM2FAB_D0_InPass4_frame_config_mux.cus_mux21_inst3._1_
rlabel metal2 17158 6052 17158 6052 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.ConfigBits\[0\]
rlabel metal2 18722 4726 18722 4726 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.ConfigBits\[1\]
rlabel metal1 19826 7174 19826 7174 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.ConfigBits\[2\]
rlabel metal1 17250 7480 17250 7480 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.ConfigBits\[3\]
rlabel metal1 9890 7310 9890 7310 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.O\[0\]
rlabel metal1 2392 16082 2392 16082 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.O\[1\]
rlabel metal1 2484 10574 2484 10574 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.O\[2\]
rlabel metal1 12972 10574 12972 10574 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.O\[3\]
rlabel metal1 17526 4114 17526 4114 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.Q\[0\]
rlabel metal1 18676 4590 18676 4590 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.Q\[1\]
rlabel metal1 21114 6426 21114 6426 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.Q\[2\]
rlabel metal1 18032 6970 18032 6970 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.Q\[3\]
rlabel metal1 16836 4726 16836 4726 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst0.AIN\[0\]
rlabel metal1 17066 3978 17066 3978 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst0.AIN\[1\]
rlabel metal1 16514 5882 16514 5882 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst0._0_
rlabel metal1 17250 4794 17250 4794 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst0._1_
rlabel metal1 17756 3502 17756 3502 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst1.AIN\[0\]
rlabel metal1 18906 4148 18906 4148 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst1.AIN\[1\]
rlabel metal1 17802 3706 17802 3706 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst1._0_
rlabel metal1 18446 4080 18446 4080 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst1._1_
rlabel metal1 20930 5576 20930 5576 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst2.AIN\[0\]
rlabel metal2 18078 6256 18078 6256 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst2.AIN\[1\]
rlabel metal1 18630 6970 18630 6970 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst2._0_
rlabel metal1 19826 7854 19826 7854 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst2._1_
rlabel metal1 17894 7344 17894 7344 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst3.AIN\[0\]
rlabel metal1 16238 7276 16238 7276 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst3.AIN\[1\]
rlabel metal2 17986 7786 17986 7786 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst3._0_
rlabel metal2 16146 7599 16146 7599 0 Inst_RAM2FAB_D1_InPass4_frame_config_mux.cus_mux21_inst3._1_
rlabel metal1 14904 6630 14904 6630 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.ConfigBits\[0\]
rlabel metal2 17618 5542 17618 5542 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.ConfigBits\[1\]
rlabel metal1 20240 6086 20240 6086 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.ConfigBits\[2\]
rlabel metal2 14950 5508 14950 5508 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.ConfigBits\[3\]
rlabel metal1 12190 5814 12190 5814 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.O\[0\]
rlabel metal2 18354 5729 18354 5729 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.O\[1\]
rlabel metal2 21206 5967 21206 5967 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.O\[2\]
rlabel metal1 14950 8262 14950 8262 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.O\[3\]
rlabel metal1 15732 5338 15732 5338 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.Q\[0\]
rlabel metal1 14674 3502 14674 3502 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.Q\[1\]
rlabel metal1 14352 3026 14352 3026 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.Q\[2\]
rlabel metal1 15732 4590 15732 4590 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.Q\[3\]
rlabel metal1 15548 4998 15548 4998 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst0.AIN\[0\]
rlabel metal1 15732 5882 15732 5882 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst0.AIN\[1\]
rlabel metal1 14490 5712 14490 5712 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst0._0_
rlabel metal1 14858 5712 14858 5712 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst0._1_
rlabel metal1 14950 3706 14950 3706 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst1.AIN\[0\]
rlabel metal1 14904 3638 14904 3638 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst1.AIN\[1\]
rlabel metal1 15686 4250 15686 4250 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst1._0_
rlabel metal1 16652 4794 16652 4794 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst1._1_
rlabel metal1 14858 3162 14858 3162 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst2.AIN\[0\]
rlabel metal2 14122 3383 14122 3383 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst2.AIN\[1\]
rlabel metal2 15594 4403 15594 4403 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst2._0_
rlabel metal1 21114 5270 21114 5270 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst2._1_
rlabel metal1 14582 4250 14582 4250 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst3.AIN\[0\]
rlabel metal1 16008 4794 16008 4794 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst3.AIN\[1\]
rlabel metal2 16146 5338 16146 5338 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst3._0_
rlabel metal1 16146 5338 16146 5338 0 Inst_RAM2FAB_D2_InPass4_frame_config_mux.cus_mux21_inst3._1_
rlabel metal2 15042 7548 15042 7548 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.ConfigBits\[0\]
rlabel metal1 18906 4658 18906 4658 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.ConfigBits\[1\]
rlabel metal1 20608 9554 20608 9554 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.ConfigBits\[2\]
rlabel metal1 18492 10030 18492 10030 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.ConfigBits\[3\]
rlabel metal1 8878 13940 8878 13940 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.O\[0\]
rlabel metal1 1794 7378 1794 7378 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.O\[1\]
rlabel metal1 2530 8398 2530 8398 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.O\[2\]
rlabel viali 12107 9554 12107 9554 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.O\[3\]
rlabel metal2 15686 6596 15686 6596 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.Q\[0\]
rlabel metal1 20976 3706 20976 3706 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.Q\[1\]
rlabel metal1 21206 6290 21206 6290 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.Q\[2\]
rlabel metal1 19228 9690 19228 9690 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.Q\[3\]
rlabel metal1 13892 6426 13892 6426 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst0.AIN\[0\]
rlabel metal1 15502 6936 15502 6936 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst0.AIN\[1\]
rlabel metal1 14214 6970 14214 6970 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst0._0_
rlabel metal1 15042 7446 15042 7446 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst0._1_
rlabel metal1 15088 3978 15088 3978 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst1.AIN\[0\]
rlabel metal1 20240 4250 20240 4250 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst1.AIN\[1\]
rlabel metal1 19182 3094 19182 3094 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst1._0_
rlabel metal2 19550 3740 19550 3740 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst1._1_
rlabel metal1 21390 7820 21390 7820 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst2.AIN\[0\]
rlabel metal1 21436 6426 21436 6426 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst2.AIN\[1\]
rlabel metal1 21298 8058 21298 8058 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst2._0_
rlabel metal1 20378 9146 20378 9146 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst2._1_
rlabel metal1 18124 8942 18124 8942 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst3.AIN\[0\]
rlabel metal1 19044 9350 19044 9350 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst3.AIN\[1\]
rlabel metal1 18262 9146 18262 9146 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst3._0_
rlabel metal1 18630 9962 18630 9962 0 Inst_RAM2FAB_D3_InPass4_frame_config_mux.cus_mux21_inst3._1_
rlabel metal1 11684 21862 11684 21862 0 Inst_RAM_IO_ConfigMem.ConfigBits\[100\]
rlabel metal1 12190 21114 12190 21114 0 Inst_RAM_IO_ConfigMem.ConfigBits\[101\]
rlabel metal1 5106 21386 5106 21386 0 Inst_RAM_IO_ConfigMem.ConfigBits\[102\]
rlabel metal1 7084 21862 7084 21862 0 Inst_RAM_IO_ConfigMem.ConfigBits\[103\]
rlabel metal2 3910 22100 3910 22100 0 Inst_RAM_IO_ConfigMem.ConfigBits\[104\]
rlabel metal1 3726 22712 3726 22712 0 Inst_RAM_IO_ConfigMem.ConfigBits\[105\]
rlabel metal2 12650 19584 12650 19584 0 Inst_RAM_IO_ConfigMem.ConfigBits\[106\]
rlabel metal2 12466 18972 12466 18972 0 Inst_RAM_IO_ConfigMem.ConfigBits\[107\]
rlabel metal1 14214 19958 14214 19958 0 Inst_RAM_IO_ConfigMem.ConfigBits\[108\]
rlabel metal1 14628 20366 14628 20366 0 Inst_RAM_IO_ConfigMem.ConfigBits\[109\]
rlabel metal1 16100 20230 16100 20230 0 Inst_RAM_IO_ConfigMem.ConfigBits\[110\]
rlabel metal1 5382 24344 5382 24344 0 Inst_RAM_IO_ConfigMem.ConfigBits\[111\]
rlabel metal1 6210 23494 6210 23494 0 Inst_RAM_IO_ConfigMem.ConfigBits\[112\]
rlabel metal1 8096 22474 8096 22474 0 Inst_RAM_IO_ConfigMem.ConfigBits\[113\]
rlabel metal1 8280 24378 8280 24378 0 Inst_RAM_IO_ConfigMem.ConfigBits\[114\]
rlabel metal1 9062 23630 9062 23630 0 Inst_RAM_IO_ConfigMem.ConfigBits\[115\]
rlabel metal2 11178 23868 11178 23868 0 Inst_RAM_IO_ConfigMem.ConfigBits\[116\]
rlabel metal1 14444 26894 14444 26894 0 Inst_RAM_IO_ConfigMem.ConfigBits\[117\]
rlabel metal1 15134 26894 15134 26894 0 Inst_RAM_IO_ConfigMem.ConfigBits\[118\]
rlabel metal2 16238 26044 16238 26044 0 Inst_RAM_IO_ConfigMem.ConfigBits\[119\]
rlabel metal1 11914 6970 11914 6970 0 Inst_RAM_IO_ConfigMem.ConfigBits\[120\]
rlabel metal1 12466 7514 12466 7514 0 Inst_RAM_IO_ConfigMem.ConfigBits\[121\]
rlabel metal1 6762 7990 6762 7990 0 Inst_RAM_IO_ConfigMem.ConfigBits\[122\]
rlabel metal1 6624 7514 6624 7514 0 Inst_RAM_IO_ConfigMem.ConfigBits\[123\]
rlabel metal1 7130 11594 7130 11594 0 Inst_RAM_IO_ConfigMem.ConfigBits\[124\]
rlabel metal1 8464 10778 8464 10778 0 Inst_RAM_IO_ConfigMem.ConfigBits\[125\]
rlabel metal1 10856 16694 10856 16694 0 Inst_RAM_IO_ConfigMem.ConfigBits\[126\]
rlabel metal1 11638 16626 11638 16626 0 Inst_RAM_IO_ConfigMem.ConfigBits\[127\]
rlabel metal1 9200 11254 9200 11254 0 Inst_RAM_IO_ConfigMem.ConfigBits\[128\]
rlabel metal1 10074 10778 10074 10778 0 Inst_RAM_IO_ConfigMem.ConfigBits\[129\]
rlabel metal1 3128 5338 3128 5338 0 Inst_RAM_IO_ConfigMem.ConfigBits\[130\]
rlabel metal1 3496 4794 3496 4794 0 Inst_RAM_IO_ConfigMem.ConfigBits\[131\]
rlabel metal1 5842 4794 5842 4794 0 Inst_RAM_IO_ConfigMem.ConfigBits\[132\]
rlabel metal1 5336 3910 5336 3910 0 Inst_RAM_IO_ConfigMem.ConfigBits\[133\]
rlabel metal1 7682 6970 7682 6970 0 Inst_RAM_IO_ConfigMem.ConfigBits\[134\]
rlabel metal1 8602 6970 8602 6970 0 Inst_RAM_IO_ConfigMem.ConfigBits\[135\]
rlabel metal1 10258 6426 10258 6426 0 Inst_RAM_IO_ConfigMem.ConfigBits\[136\]
rlabel metal1 10672 6970 10672 6970 0 Inst_RAM_IO_ConfigMem.ConfigBits\[137\]
rlabel metal2 2438 4692 2438 4692 0 Inst_RAM_IO_ConfigMem.ConfigBits\[138\]
rlabel metal1 3542 2822 3542 2822 0 Inst_RAM_IO_ConfigMem.ConfigBits\[139\]
rlabel metal1 2760 3706 2760 3706 0 Inst_RAM_IO_ConfigMem.ConfigBits\[140\]
rlabel metal1 2668 4250 2668 4250 0 Inst_RAM_IO_ConfigMem.ConfigBits\[141\]
rlabel metal1 13340 10574 13340 10574 0 Inst_RAM_IO_ConfigMem.ConfigBits\[142\]
rlabel metal1 14168 10574 14168 10574 0 Inst_RAM_IO_ConfigMem.ConfigBits\[143\]
rlabel metal1 9706 12784 9706 12784 0 Inst_RAM_IO_ConfigMem.ConfigBits\[144\]
rlabel metal1 11040 12682 11040 12682 0 Inst_RAM_IO_ConfigMem.ConfigBits\[145\]
rlabel metal2 2438 16694 2438 16694 0 Inst_RAM_IO_ConfigMem.ConfigBits\[146\]
rlabel metal1 2944 16762 2944 16762 0 Inst_RAM_IO_ConfigMem.ConfigBits\[147\]
rlabel metal1 4876 4794 4876 4794 0 Inst_RAM_IO_ConfigMem.ConfigBits\[148\]
rlabel metal1 4968 5338 4968 5338 0 Inst_RAM_IO_ConfigMem.ConfigBits\[149\]
rlabel metal1 8924 9418 8924 9418 0 Inst_RAM_IO_ConfigMem.ConfigBits\[150\]
rlabel metal2 10028 9146 10028 9146 0 Inst_RAM_IO_ConfigMem.ConfigBits\[151\]
rlabel metal1 9568 8330 9568 8330 0 Inst_RAM_IO_ConfigMem.ConfigBits\[152\]
rlabel metal2 10626 8228 10626 8228 0 Inst_RAM_IO_ConfigMem.ConfigBits\[153\]
rlabel metal1 2668 3162 2668 3162 0 Inst_RAM_IO_ConfigMem.ConfigBits\[154\]
rlabel metal1 3634 3910 3634 3910 0 Inst_RAM_IO_ConfigMem.ConfigBits\[155\]
rlabel metal2 3174 8466 3174 8466 0 Inst_RAM_IO_ConfigMem.ConfigBits\[156\]
rlabel metal2 3496 10506 3496 10506 0 Inst_RAM_IO_ConfigMem.ConfigBits\[157\]
rlabel metal1 12604 13498 12604 13498 0 Inst_RAM_IO_ConfigMem.ConfigBits\[158\]
rlabel metal1 12972 14042 12972 14042 0 Inst_RAM_IO_ConfigMem.ConfigBits\[159\]
rlabel metal1 11500 10778 11500 10778 0 Inst_RAM_IO_ConfigMem.ConfigBits\[160\]
rlabel metal2 12374 11322 12374 11322 0 Inst_RAM_IO_ConfigMem.ConfigBits\[161\]
rlabel metal1 7406 8602 7406 8602 0 Inst_RAM_IO_ConfigMem.ConfigBits\[162\]
rlabel metal1 7958 9146 7958 9146 0 Inst_RAM_IO_ConfigMem.ConfigBits\[163\]
rlabel metal1 3634 12410 3634 12410 0 Inst_RAM_IO_ConfigMem.ConfigBits\[164\]
rlabel metal1 3358 11254 3358 11254 0 Inst_RAM_IO_ConfigMem.ConfigBits\[165\]
rlabel metal2 12742 9282 12742 9282 0 Inst_RAM_IO_ConfigMem.ConfigBits\[166\]
rlabel metal1 13616 8602 13616 8602 0 Inst_RAM_IO_ConfigMem.ConfigBits\[167\]
rlabel metal1 10488 10234 10488 10234 0 Inst_RAM_IO_ConfigMem.ConfigBits\[168\]
rlabel metal1 10350 12376 10350 12376 0 Inst_RAM_IO_ConfigMem.ConfigBits\[169\]
rlabel metal2 2622 13940 2622 13940 0 Inst_RAM_IO_ConfigMem.ConfigBits\[170\]
rlabel metal1 3358 13498 3358 13498 0 Inst_RAM_IO_ConfigMem.ConfigBits\[171\]
rlabel metal1 5106 8058 5106 8058 0 Inst_RAM_IO_ConfigMem.ConfigBits\[172\]
rlabel metal1 5244 9146 5244 9146 0 Inst_RAM_IO_ConfigMem.ConfigBits\[173\]
rlabel metal2 13110 12104 13110 12104 0 Inst_RAM_IO_ConfigMem.ConfigBits\[174\]
rlabel metal2 13662 12036 13662 12036 0 Inst_RAM_IO_ConfigMem.ConfigBits\[175\]
rlabel metal1 10396 14518 10396 14518 0 Inst_RAM_IO_ConfigMem.ConfigBits\[176\]
rlabel metal2 11086 14586 11086 14586 0 Inst_RAM_IO_ConfigMem.ConfigBits\[177\]
rlabel metal1 4278 17102 4278 17102 0 Inst_RAM_IO_ConfigMem.ConfigBits\[178\]
rlabel metal2 5014 17238 5014 17238 0 Inst_RAM_IO_ConfigMem.ConfigBits\[179\]
rlabel metal1 5244 6426 5244 6426 0 Inst_RAM_IO_ConfigMem.ConfigBits\[180\]
rlabel metal1 5704 8330 5704 8330 0 Inst_RAM_IO_ConfigMem.ConfigBits\[181\]
rlabel metal1 12512 8602 12512 8602 0 Inst_RAM_IO_ConfigMem.ConfigBits\[182\]
rlabel metal1 12972 9146 12972 9146 0 Inst_RAM_IO_ConfigMem.ConfigBits\[183\]
rlabel metal1 9016 13498 9016 13498 0 Inst_RAM_IO_ConfigMem.ConfigBits\[184\]
rlabel metal2 10074 14348 10074 14348 0 Inst_RAM_IO_ConfigMem.ConfigBits\[185\]
rlabel metal1 3312 8058 3312 8058 0 Inst_RAM_IO_ConfigMem.ConfigBits\[186\]
rlabel metal2 3358 11526 3358 11526 0 Inst_RAM_IO_ConfigMem.ConfigBits\[187\]
rlabel metal1 3118 14858 3118 14858 0 Inst_RAM_IO_ConfigMem.ConfigBits\[188\]
rlabel metal1 4232 14042 4232 14042 0 Inst_RAM_IO_ConfigMem.ConfigBits\[189\]
rlabel metal1 14766 14586 14766 14586 0 Inst_RAM_IO_ConfigMem.ConfigBits\[190\]
rlabel metal1 15272 14926 15272 14926 0 Inst_RAM_IO_ConfigMem.ConfigBits\[191\]
rlabel metal1 14628 12954 14628 12954 0 Inst_RAM_IO_ConfigMem.ConfigBits\[192\]
rlabel metal1 15594 12954 15594 12954 0 Inst_RAM_IO_ConfigMem.ConfigBits\[193\]
rlabel metal1 6854 26894 6854 26894 0 Inst_RAM_IO_ConfigMem.ConfigBits\[194\]
rlabel metal2 7590 27166 7590 27166 0 Inst_RAM_IO_ConfigMem.ConfigBits\[195\]
rlabel metal2 5750 12563 5750 12563 0 Inst_RAM_IO_ConfigMem.ConfigBits\[196\]
rlabel metal1 7084 14586 7084 14586 0 Inst_RAM_IO_ConfigMem.ConfigBits\[197\]
rlabel metal2 12650 22542 12650 22542 0 Inst_RAM_IO_ConfigMem.ConfigBits\[198\]
rlabel metal2 13294 22508 13294 22508 0 Inst_RAM_IO_ConfigMem.ConfigBits\[199\]
rlabel metal1 12880 16218 12880 16218 0 Inst_RAM_IO_ConfigMem.ConfigBits\[200\]
rlabel metal1 13432 16762 13432 16762 0 Inst_RAM_IO_ConfigMem.ConfigBits\[201\]
rlabel metal1 5796 14042 5796 14042 0 Inst_RAM_IO_ConfigMem.ConfigBits\[202\]
rlabel metal1 6486 16626 6486 16626 0 Inst_RAM_IO_ConfigMem.ConfigBits\[203\]
rlabel metal1 4554 8806 4554 8806 0 Inst_RAM_IO_ConfigMem.ConfigBits\[204\]
rlabel metal1 6072 10234 6072 10234 0 Inst_RAM_IO_ConfigMem.ConfigBits\[205\]
rlabel metal1 12926 15130 12926 15130 0 Inst_RAM_IO_ConfigMem.ConfigBits\[206\]
rlabel metal1 13800 15538 13800 15538 0 Inst_RAM_IO_ConfigMem.ConfigBits\[207\]
rlabel metal1 10120 16014 10120 16014 0 Inst_RAM_IO_ConfigMem.ConfigBits\[208\]
rlabel metal1 10810 16014 10810 16014 0 Inst_RAM_IO_ConfigMem.ConfigBits\[209\]
rlabel metal1 3680 17306 3680 17306 0 Inst_RAM_IO_ConfigMem.ConfigBits\[210\]
rlabel metal2 5014 18343 5014 18343 0 Inst_RAM_IO_ConfigMem.ConfigBits\[211\]
rlabel metal1 3864 14586 3864 14586 0 Inst_RAM_IO_ConfigMem.ConfigBits\[212\]
rlabel metal2 5290 15028 5290 15028 0 Inst_RAM_IO_ConfigMem.ConfigBits\[213\]
rlabel metal1 14214 17782 14214 17782 0 Inst_RAM_IO_ConfigMem.ConfigBits\[214\]
rlabel metal2 15318 17884 15318 17884 0 Inst_RAM_IO_ConfigMem.ConfigBits\[215\]
rlabel metal1 16100 24310 16100 24310 0 Inst_RAM_IO_ConfigMem.ConfigBits\[216\]
rlabel metal1 17066 24242 17066 24242 0 Inst_RAM_IO_ConfigMem.ConfigBits\[217\]
rlabel metal2 2898 33898 2898 33898 0 Inst_RAM_IO_ConfigMem.ConfigBits\[218\]
rlabel metal1 3312 33082 3312 33082 0 Inst_RAM_IO_ConfigMem.ConfigBits\[219\]
rlabel metal1 2898 25670 2898 25670 0 Inst_RAM_IO_ConfigMem.ConfigBits\[220\]
rlabel metal2 3358 25704 3358 25704 0 Inst_RAM_IO_ConfigMem.ConfigBits\[221\]
rlabel metal2 16238 28849 16238 28849 0 Inst_RAM_IO_ConfigMem.ConfigBits\[222\]
rlabel metal2 15318 28628 15318 28628 0 Inst_RAM_IO_ConfigMem.ConfigBits\[223\]
rlabel metal1 16008 22134 16008 22134 0 Inst_RAM_IO_ConfigMem.ConfigBits\[224\]
rlabel metal1 16928 22066 16928 22066 0 Inst_RAM_IO_ConfigMem.ConfigBits\[225\]
rlabel metal1 4186 29002 4186 29002 0 Inst_RAM_IO_ConfigMem.ConfigBits\[226\]
rlabel metal1 4646 28118 4646 28118 0 Inst_RAM_IO_ConfigMem.ConfigBits\[227\]
rlabel metal1 9062 25398 9062 25398 0 Inst_RAM_IO_ConfigMem.ConfigBits\[228\]
rlabel metal1 10396 24922 10396 24922 0 Inst_RAM_IO_ConfigMem.ConfigBits\[229\]
rlabel metal1 14766 29784 14766 29784 0 Inst_RAM_IO_ConfigMem.ConfigBits\[230\]
rlabel metal1 15410 29682 15410 29682 0 Inst_RAM_IO_ConfigMem.ConfigBits\[231\]
rlabel metal2 16054 23902 16054 23902 0 Inst_RAM_IO_ConfigMem.ConfigBits\[232\]
rlabel metal1 17158 23154 17158 23154 0 Inst_RAM_IO_ConfigMem.ConfigBits\[233\]
rlabel metal1 4186 30838 4186 30838 0 Inst_RAM_IO_ConfigMem.ConfigBits\[234\]
rlabel metal1 4692 30362 4692 30362 0 Inst_RAM_IO_ConfigMem.ConfigBits\[235\]
rlabel metal1 2622 27003 2622 27003 0 Inst_RAM_IO_ConfigMem.ConfigBits\[236\]
rlabel metal1 4002 26554 4002 26554 0 Inst_RAM_IO_ConfigMem.ConfigBits\[237\]
rlabel metal2 13938 29025 13938 29025 0 Inst_RAM_IO_ConfigMem.ConfigBits\[238\]
rlabel metal2 14490 29852 14490 29852 0 Inst_RAM_IO_ConfigMem.ConfigBits\[239\]
rlabel metal1 17572 21114 17572 21114 0 Inst_RAM_IO_ConfigMem.ConfigBits\[240\]
rlabel metal1 17848 20570 17848 20570 0 Inst_RAM_IO_ConfigMem.ConfigBits\[241\]
rlabel metal2 2714 28458 2714 28458 0 Inst_RAM_IO_ConfigMem.ConfigBits\[242\]
rlabel metal2 2530 28254 2530 28254 0 Inst_RAM_IO_ConfigMem.ConfigBits\[243\]
rlabel metal1 7866 25738 7866 25738 0 Inst_RAM_IO_ConfigMem.ConfigBits\[244\]
rlabel metal1 8602 25976 8602 25976 0 Inst_RAM_IO_ConfigMem.ConfigBits\[245\]
rlabel metal1 14766 31960 14766 31960 0 Inst_RAM_IO_ConfigMem.ConfigBits\[246\]
rlabel metal1 15502 31858 15502 31858 0 Inst_RAM_IO_ConfigMem.ConfigBits\[247\]
rlabel metal2 13110 18802 13110 18802 0 Inst_RAM_IO_ConfigMem.ConfigBits\[248\]
rlabel metal1 13984 19278 13984 19278 0 Inst_RAM_IO_ConfigMem.ConfigBits\[249\]
rlabel metal2 4462 38046 4462 38046 0 Inst_RAM_IO_ConfigMem.ConfigBits\[250\]
rlabel metal2 5014 37740 5014 37740 0 Inst_RAM_IO_ConfigMem.ConfigBits\[251\]
rlabel metal1 5750 19958 5750 19958 0 Inst_RAM_IO_ConfigMem.ConfigBits\[252\]
rlabel metal1 5934 20026 5934 20026 0 Inst_RAM_IO_ConfigMem.ConfigBits\[253\]
rlabel metal2 12282 35734 12282 35734 0 Inst_RAM_IO_ConfigMem.ConfigBits\[254\]
rlabel metal2 12834 35292 12834 35292 0 Inst_RAM_IO_ConfigMem.ConfigBits\[255\]
rlabel metal1 8602 21420 8602 21420 0 Inst_RAM_IO_ConfigMem.ConfigBits\[256\]
rlabel metal1 9890 21114 9890 21114 0 Inst_RAM_IO_ConfigMem.ConfigBits\[257\]
rlabel metal1 3220 21318 3220 21318 0 Inst_RAM_IO_ConfigMem.ConfigBits\[258\]
rlabel metal1 3910 20026 3910 20026 0 Inst_RAM_IO_ConfigMem.ConfigBits\[259\]
rlabel metal2 2714 36652 2714 36652 0 Inst_RAM_IO_ConfigMem.ConfigBits\[260\]
rlabel metal2 2622 35530 2622 35530 0 Inst_RAM_IO_ConfigMem.ConfigBits\[261\]
rlabel metal1 13524 36686 13524 36686 0 Inst_RAM_IO_ConfigMem.ConfigBits\[262\]
rlabel metal1 14214 36686 14214 36686 0 Inst_RAM_IO_ConfigMem.ConfigBits\[263\]
rlabel metal1 17526 16218 17526 16218 0 Inst_RAM_IO_ConfigMem.ConfigBits\[264\]
rlabel via1 17893 17102 17893 17102 0 Inst_RAM_IO_ConfigMem.ConfigBits\[265\]
rlabel metal1 8188 32198 8188 32198 0 Inst_RAM_IO_ConfigMem.ConfigBits\[266\]
rlabel metal2 8510 31484 8510 31484 0 Inst_RAM_IO_ConfigMem.ConfigBits\[267\]
rlabel metal1 8464 18598 8464 18598 0 Inst_RAM_IO_ConfigMem.ConfigBits\[268\]
rlabel metal2 9982 18054 9982 18054 0 Inst_RAM_IO_ConfigMem.ConfigBits\[269\]
rlabel metal1 15226 33048 15226 33048 0 Inst_RAM_IO_ConfigMem.ConfigBits\[270\]
rlabel metal1 15870 32946 15870 32946 0 Inst_RAM_IO_ConfigMem.ConfigBits\[271\]
rlabel metal1 16245 13838 16245 13838 0 Inst_RAM_IO_ConfigMem.ConfigBits\[272\]
rlabel metal1 16882 13498 16882 13498 0 Inst_RAM_IO_ConfigMem.ConfigBits\[273\]
rlabel metal1 5060 36550 5060 36550 0 Inst_RAM_IO_ConfigMem.ConfigBits\[274\]
rlabel metal1 5520 34646 5520 34646 0 Inst_RAM_IO_ConfigMem.ConfigBits\[275\]
rlabel metal2 6532 12886 6532 12886 0 Inst_RAM_IO_ConfigMem.ConfigBits\[276\]
rlabel metal2 7130 13702 7130 13702 0 Inst_RAM_IO_ConfigMem.ConfigBits\[277\]
rlabel metal1 11178 27574 11178 27574 0 Inst_RAM_IO_ConfigMem.ConfigBits\[278\]
rlabel metal2 11914 27608 11914 27608 0 Inst_RAM_IO_ConfigMem.ConfigBits\[279\]
rlabel metal2 15134 9622 15134 9622 0 Inst_RAM_IO_ConfigMem.ConfigBits\[280\]
rlabel metal1 15456 10030 15456 10030 0 Inst_RAM_IO_ConfigMem.ConfigBits\[281\]
rlabel metal2 4278 34272 4278 34272 0 Inst_RAM_IO_ConfigMem.ConfigBits\[282\]
rlabel metal1 5382 33966 5382 33966 0 Inst_RAM_IO_ConfigMem.ConfigBits\[283\]
rlabel metal1 6256 14790 6256 14790 0 Inst_RAM_IO_ConfigMem.ConfigBits\[284\]
rlabel metal2 7590 17000 7590 17000 0 Inst_RAM_IO_ConfigMem.ConfigBits\[285\]
rlabel metal1 11316 26826 11316 26826 0 Inst_RAM_IO_ConfigMem.ConfigBits\[286\]
rlabel metal1 12144 27030 12144 27030 0 Inst_RAM_IO_ConfigMem.ConfigBits\[287\]
rlabel metal1 16054 11686 16054 11686 0 Inst_RAM_IO_ConfigMem.ConfigBits\[288\]
rlabel metal2 16606 11560 16606 11560 0 Inst_RAM_IO_ConfigMem.ConfigBits\[289\]
rlabel metal2 5658 33116 5658 33116 0 Inst_RAM_IO_ConfigMem.ConfigBits\[290\]
rlabel metal2 5842 33082 5842 33082 0 Inst_RAM_IO_ConfigMem.ConfigBits\[291\]
rlabel metal1 8425 15538 8425 15538 0 Inst_RAM_IO_ConfigMem.ConfigBits\[292\]
rlabel metal2 8050 15028 8050 15028 0 Inst_RAM_IO_ConfigMem.ConfigBits\[293\]
rlabel metal2 12558 25500 12558 25500 0 Inst_RAM_IO_ConfigMem.ConfigBits\[294\]
rlabel metal2 11914 25058 11914 25058 0 Inst_RAM_IO_ConfigMem.ConfigBits\[295\]
rlabel metal2 15318 9044 15318 9044 0 Inst_RAM_IO_ConfigMem.ConfigBits\[296\]
rlabel metal1 15870 9146 15870 9146 0 Inst_RAM_IO_ConfigMem.ConfigBits\[297\]
rlabel metal2 5934 29852 5934 29852 0 Inst_RAM_IO_ConfigMem.ConfigBits\[298\]
rlabel metal1 5842 29274 5842 29274 0 Inst_RAM_IO_ConfigMem.ConfigBits\[299\]
rlabel metal1 6164 11866 6164 11866 0 Inst_RAM_IO_ConfigMem.ConfigBits\[300\]
rlabel metal1 7084 12410 7084 12410 0 Inst_RAM_IO_ConfigMem.ConfigBits\[301\]
rlabel metal1 10994 26486 10994 26486 0 Inst_RAM_IO_ConfigMem.ConfigBits\[302\]
rlabel metal2 13938 26180 13938 26180 0 Inst_RAM_IO_ConfigMem.ConfigBits\[303\]
rlabel metal2 8510 32538 8510 32538 0 Inst_RAM_IO_ConfigMem.ConfigBits\[304\]
rlabel metal1 9660 32470 9660 32470 0 Inst_RAM_IO_ConfigMem.ConfigBits\[305\]
rlabel metal1 5888 35802 5888 35802 0 Inst_RAM_IO_ConfigMem.ConfigBits\[306\]
rlabel metal2 7314 35700 7314 35700 0 Inst_RAM_IO_ConfigMem.ConfigBits\[307\]
rlabel metal1 6256 5066 6256 5066 0 Inst_RAM_IO_ConfigMem.ConfigBits\[308\]
rlabel metal1 7268 5882 7268 5882 0 Inst_RAM_IO_ConfigMem.ConfigBits\[309\]
rlabel metal1 8694 34476 8694 34476 0 Inst_RAM_IO_ConfigMem.ConfigBits\[310\]
rlabel metal1 9982 34170 9982 34170 0 Inst_RAM_IO_ConfigMem.ConfigBits\[311\]
rlabel metal2 8050 35292 8050 35292 0 Inst_RAM_IO_ConfigMem.ConfigBits\[312\]
rlabel metal2 9522 35173 9522 35173 0 Inst_RAM_IO_ConfigMem.ConfigBits\[313\]
rlabel metal1 5566 21046 5566 21046 0 Inst_RAM_IO_ConfigMem.ConfigBits\[314\]
rlabel metal2 5934 20196 5934 20196 0 Inst_RAM_IO_ConfigMem.ConfigBits\[315\]
rlabel metal2 7774 37978 7774 37978 0 Inst_RAM_IO_ConfigMem.ConfigBits\[316\]
rlabel metal2 8326 37366 8326 37366 0 Inst_RAM_IO_ConfigMem.ConfigBits\[317\]
rlabel metal2 10718 37468 10718 37468 0 Inst_RAM_IO_ConfigMem.ConfigBits\[318\]
rlabel metal1 10764 36890 10764 36890 0 Inst_RAM_IO_ConfigMem.ConfigBits\[319\]
rlabel metal1 15824 16218 15824 16218 0 Inst_RAM_IO_ConfigMem.ConfigBits\[320\]
rlabel metal1 16514 16626 16514 16626 0 Inst_RAM_IO_ConfigMem.ConfigBits\[321\]
rlabel metal1 6486 38182 6486 38182 0 Inst_RAM_IO_ConfigMem.ConfigBits\[322\]
rlabel metal1 6716 37162 6716 37162 0 Inst_RAM_IO_ConfigMem.ConfigBits\[323\]
rlabel metal1 6578 16218 6578 16218 0 Inst_RAM_IO_ConfigMem.ConfigBits\[324\]
rlabel metal1 7820 17646 7820 17646 0 Inst_RAM_IO_ConfigMem.ConfigBits\[325\]
rlabel metal1 10442 31960 10442 31960 0 Inst_RAM_IO_ConfigMem.ConfigBits\[326\]
rlabel metal1 10902 31450 10902 31450 0 Inst_RAM_IO_ConfigMem.ConfigBits\[327\]
rlabel metal1 16882 18938 16882 18938 0 Inst_RAM_IO_ConfigMem.ConfigBits\[48\]
rlabel metal1 17434 19482 17434 19482 0 Inst_RAM_IO_ConfigMem.ConfigBits\[49\]
rlabel metal2 2438 31654 2438 31654 0 Inst_RAM_IO_ConfigMem.ConfigBits\[50\]
rlabel metal2 2990 31994 2990 31994 0 Inst_RAM_IO_ConfigMem.ConfigBits\[51\]
rlabel metal2 8142 28084 8142 28084 0 Inst_RAM_IO_ConfigMem.ConfigBits\[52\]
rlabel metal2 7774 27608 7774 27608 0 Inst_RAM_IO_ConfigMem.ConfigBits\[53\]
rlabel metal2 10994 33388 10994 33388 0 Inst_RAM_IO_ConfigMem.ConfigBits\[54\]
rlabel metal2 11270 33082 11270 33082 0 Inst_RAM_IO_ConfigMem.ConfigBits\[55\]
rlabel metal2 13846 33898 13846 33898 0 Inst_RAM_IO_ConfigMem.ConfigBits\[56\]
rlabel metal1 13570 33592 13570 33592 0 Inst_RAM_IO_ConfigMem.ConfigBits\[57\]
rlabel metal2 2438 36074 2438 36074 0 Inst_RAM_IO_ConfigMem.ConfigBits\[58\]
rlabel metal2 2990 36380 2990 36380 0 Inst_RAM_IO_ConfigMem.ConfigBits\[59\]
rlabel metal2 2438 25466 2438 25466 0 Inst_RAM_IO_ConfigMem.ConfigBits\[60\]
rlabel metal1 2622 24378 2622 24378 0 Inst_RAM_IO_ConfigMem.ConfigBits\[61\]
rlabel metal1 8096 29070 8096 29070 0 Inst_RAM_IO_ConfigMem.ConfigBits\[62\]
rlabel metal2 8602 29580 8602 29580 0 Inst_RAM_IO_ConfigMem.ConfigBits\[63\]
rlabel metal1 8924 35598 8924 35598 0 Inst_RAM_IO_ConfigMem.ConfigBits\[64\]
rlabel metal2 9660 35598 9660 35598 0 Inst_RAM_IO_ConfigMem.ConfigBits\[65\]
rlabel metal2 2346 23018 2346 23018 0 Inst_RAM_IO_ConfigMem.ConfigBits\[66\]
rlabel metal1 2300 22678 2300 22678 0 Inst_RAM_IO_ConfigMem.ConfigBits\[67\]
rlabel metal1 2576 37774 2576 37774 0 Inst_RAM_IO_ConfigMem.ConfigBits\[68\]
rlabel metal2 3174 38284 3174 38284 0 Inst_RAM_IO_ConfigMem.ConfigBits\[69\]
rlabel metal2 10442 19414 10442 19414 0 Inst_RAM_IO_ConfigMem.ConfigBits\[70\]
rlabel metal1 10718 19822 10718 19822 0 Inst_RAM_IO_ConfigMem.ConfigBits\[71\]
rlabel metal1 13524 23630 13524 23630 0 Inst_RAM_IO_ConfigMem.ConfigBits\[72\]
rlabel metal1 14214 23630 14214 23630 0 Inst_RAM_IO_ConfigMem.ConfigBits\[73\]
rlabel metal1 14214 24718 14214 24718 0 Inst_RAM_IO_ConfigMem.ConfigBits\[74\]
rlabel metal1 3496 32266 3496 32266 0 Inst_RAM_IO_ConfigMem.ConfigBits\[75\]
rlabel metal1 5566 32334 5566 32334 0 Inst_RAM_IO_ConfigMem.ConfigBits\[76\]
rlabel metal1 7682 33286 7682 33286 0 Inst_RAM_IO_ConfigMem.ConfigBits\[77\]
rlabel metal2 6026 25908 6026 25908 0 Inst_RAM_IO_ConfigMem.ConfigBits\[78\]
rlabel metal2 6946 25194 6946 25194 0 Inst_RAM_IO_ConfigMem.ConfigBits\[79\]
rlabel metal2 9338 26588 9338 26588 0 Inst_RAM_IO_ConfigMem.ConfigBits\[80\]
rlabel metal1 11306 29750 11306 29750 0 Inst_RAM_IO_ConfigMem.ConfigBits\[81\]
rlabel metal1 12650 29274 12650 29274 0 Inst_RAM_IO_ConfigMem.ConfigBits\[82\]
rlabel metal1 12236 31110 12236 31110 0 Inst_RAM_IO_ConfigMem.ConfigBits\[83\]
rlabel metal2 16238 17510 16238 17510 0 Inst_RAM_IO_ConfigMem.ConfigBits\[84\]
rlabel metal2 16606 17816 16606 17816 0 Inst_RAM_IO_ConfigMem.ConfigBits\[85\]
rlabel metal2 5934 30940 5934 30940 0 Inst_RAM_IO_ConfigMem.ConfigBits\[86\]
rlabel metal2 7406 30532 7406 30532 0 Inst_RAM_IO_ConfigMem.ConfigBits\[87\]
rlabel metal2 7130 19652 7130 19652 0 Inst_RAM_IO_ConfigMem.ConfigBits\[88\]
rlabel metal1 8234 19482 8234 19482 0 Inst_RAM_IO_ConfigMem.ConfigBits\[89\]
rlabel metal2 13386 32300 13386 32300 0 Inst_RAM_IO_ConfigMem.ConfigBits\[90\]
rlabel metal1 13294 31790 13294 31790 0 Inst_RAM_IO_ConfigMem.ConfigBits\[91\]
rlabel metal1 10120 22202 10120 22202 0 Inst_RAM_IO_ConfigMem.ConfigBits\[92\]
rlabel metal1 10488 22678 10488 22678 0 Inst_RAM_IO_ConfigMem.ConfigBits\[93\]
rlabel metal2 2346 30124 2346 30124 0 Inst_RAM_IO_ConfigMem.ConfigBits\[94\]
rlabel metal1 2576 29614 2576 29614 0 Inst_RAM_IO_ConfigMem.ConfigBits\[95\]
rlabel metal2 2530 19924 2530 19924 0 Inst_RAM_IO_ConfigMem.ConfigBits\[96\]
rlabel metal2 2714 20604 2714 20604 0 Inst_RAM_IO_ConfigMem.ConfigBits\[97\]
rlabel metal1 9844 28186 9844 28186 0 Inst_RAM_IO_ConfigMem.ConfigBits\[98\]
rlabel metal1 10580 28730 10580 28730 0 Inst_RAM_IO_ConfigMem.ConfigBits\[99\]
rlabel metal1 16284 19754 16284 19754 0 Inst_RAM_IO_switch_matrix.J_NS1_BEG0
rlabel metal1 8625 31246 8625 31246 0 Inst_RAM_IO_switch_matrix.J_NS1_BEG1
rlabel metal1 8188 18394 8188 18394 0 Inst_RAM_IO_switch_matrix.J_NS1_BEG2
rlabel metal1 12742 31790 12742 31790 0 Inst_RAM_IO_switch_matrix.J_NS1_BEG3
rlabel metal1 9844 22610 9844 22610 0 Inst_RAM_IO_switch_matrix.J_NS2_BEG0
rlabel metal2 3818 9588 3818 9588 0 Inst_RAM_IO_switch_matrix.J_NS2_BEG1
rlabel metal1 5589 6834 5589 6834 0 Inst_RAM_IO_switch_matrix.J_NS2_BEG2
rlabel metal1 11638 24854 11638 24854 0 Inst_RAM_IO_switch_matrix.J_NS2_BEG3
rlabel metal1 13386 20332 13386 20332 0 Inst_RAM_IO_switch_matrix.J_NS2_BEG4
rlabel metal1 5014 6834 5014 6834 0 Inst_RAM_IO_switch_matrix.J_NS2_BEG5
rlabel metal1 4600 19210 4600 19210 0 Inst_RAM_IO_switch_matrix.J_NS2_BEG6
rlabel metal2 14030 37264 14030 37264 0 Inst_RAM_IO_switch_matrix.J_NS2_BEG7
rlabel via1 14835 14926 14835 14926 0 Inst_RAM_IO_switch_matrix.J_NS4_BEG0
rlabel metal1 5658 24208 5658 24208 0 Inst_RAM_IO_switch_matrix.J_NS4_BEG1
rlabel metal1 5796 21318 5796 21318 0 Inst_RAM_IO_switch_matrix.J_NS4_BEG10
rlabel metal1 13110 25126 13110 25126 0 Inst_RAM_IO_switch_matrix.J_NS4_BEG11
rlabel metal1 16192 17510 16192 17510 0 Inst_RAM_IO_switch_matrix.J_NS4_BEG12
rlabel via1 6314 23154 6314 23154 0 Inst_RAM_IO_switch_matrix.J_NS4_BEG13
rlabel metal1 7636 20502 7636 20502 0 Inst_RAM_IO_switch_matrix.J_NS4_BEG14
rlabel metal2 14904 20060 14904 20060 0 Inst_RAM_IO_switch_matrix.J_NS4_BEG15
rlabel metal1 8271 24718 8271 24718 0 Inst_RAM_IO_switch_matrix.J_NS4_BEG2
rlabel metal2 12466 30039 12466 30039 0 Inst_RAM_IO_switch_matrix.J_NS4_BEG3
rlabel via1 15146 17646 15146 17646 0 Inst_RAM_IO_switch_matrix.J_NS4_BEG4
rlabel via1 5451 9554 5451 9554 0 Inst_RAM_IO_switch_matrix.J_NS4_BEG5
rlabel metal2 9890 25092 9890 25092 0 Inst_RAM_IO_switch_matrix.J_NS4_BEG6
rlabel via2 13018 26741 13018 26741 0 Inst_RAM_IO_switch_matrix.J_NS4_BEG7
rlabel metal1 12926 22678 12926 22678 0 Inst_RAM_IO_switch_matrix.J_NS4_BEG8
rlabel metal2 5244 20332 5244 20332 0 Inst_RAM_IO_switch_matrix.J_NS4_BEG9
rlabel metal2 17388 37196 17388 37196 0 Inst_RAM_IO_switch_matrix.N1BEG0
rlabel metal2 1978 41650 1978 41650 0 Inst_RAM_IO_switch_matrix.N1BEG1
rlabel metal1 1334 29274 1334 29274 0 Inst_RAM_IO_switch_matrix.N1BEG2
rlabel metal2 8418 36176 8418 36176 0 Inst_RAM_IO_switch_matrix.N1BEG3
rlabel metal1 14490 33354 14490 33354 0 Inst_RAM_IO_switch_matrix.N2BEG0
rlabel metal2 1702 41276 1702 41276 0 Inst_RAM_IO_switch_matrix.N2BEG1
rlabel metal2 12742 35063 12742 35063 0 Inst_RAM_IO_switch_matrix.N2BEG2
rlabel metal3 5520 40460 5520 40460 0 Inst_RAM_IO_switch_matrix.N2BEG3
rlabel metal2 2116 38420 2116 38420 0 Inst_RAM_IO_switch_matrix.N2BEG4
rlabel metal2 690 34765 690 34765 0 Inst_RAM_IO_switch_matrix.N2BEG5
rlabel metal1 3542 37978 3542 37978 0 Inst_RAM_IO_switch_matrix.N2BEG6
rlabel metal1 11224 20026 11224 20026 0 Inst_RAM_IO_switch_matrix.N2BEG7
rlabel metal3 4623 41548 4623 41548 0 Inst_RAM_IO_switch_matrix.N2BEGb0
rlabel metal1 4416 36346 4416 36346 0 Inst_RAM_IO_switch_matrix.N2BEGb1
rlabel metal3 1380 16796 1380 16796 0 Inst_RAM_IO_switch_matrix.N2BEGb2
rlabel metal1 6210 34714 6210 34714 0 Inst_RAM_IO_switch_matrix.N2BEGb3
rlabel metal1 5842 36890 5842 36890 0 Inst_RAM_IO_switch_matrix.N2BEGb4
rlabel metal4 12604 29580 12604 29580 0 Inst_RAM_IO_switch_matrix.N2BEGb5
rlabel metal2 6026 38454 6026 38454 0 Inst_RAM_IO_switch_matrix.N2BEGb6
rlabel metal2 5750 38420 5750 38420 0 Inst_RAM_IO_switch_matrix.N2BEGb7
rlabel metal2 14674 41004 14674 41004 0 Inst_RAM_IO_switch_matrix.N4BEG0
rlabel metal1 8050 34170 8050 34170 0 Inst_RAM_IO_switch_matrix.N4BEG1
rlabel metal2 1150 27676 1150 27676 0 Inst_RAM_IO_switch_matrix.N4BEG2
rlabel metal1 11500 30906 11500 30906 0 Inst_RAM_IO_switch_matrix.N4BEG3
rlabel metal2 17572 14858 17572 14858 0 Inst_RAM_IO_switch_matrix.S1BEG0
rlabel metal2 9476 17204 9476 17204 0 Inst_RAM_IO_switch_matrix.S1BEG1
rlabel metal2 12650 7803 12650 7803 0 Inst_RAM_IO_switch_matrix.S1BEG2
rlabel metal1 14214 2414 14214 2414 0 Inst_RAM_IO_switch_matrix.S1BEG3
rlabel metal3 14099 9724 14099 9724 0 Inst_RAM_IO_switch_matrix.S2BEG0
rlabel metal2 828 24684 828 24684 0 Inst_RAM_IO_switch_matrix.S2BEG1
rlabel metal1 1702 2346 1702 2346 0 Inst_RAM_IO_switch_matrix.S2BEG2
rlabel metal1 184 25058 184 25058 0 Inst_RAM_IO_switch_matrix.S2BEG3
rlabel metal3 14421 17340 14421 17340 0 Inst_RAM_IO_switch_matrix.S2BEG4
rlabel metal1 690 19788 690 19788 0 Inst_RAM_IO_switch_matrix.S2BEG5
rlabel metal2 966 2519 966 2519 0 Inst_RAM_IO_switch_matrix.S2BEG6
rlabel metal1 16790 15130 16790 15130 0 Inst_RAM_IO_switch_matrix.S2BEG7
rlabel metal4 1564 32564 1564 32564 0 Inst_RAM_IO_switch_matrix.S2BEGb0
rlabel metal1 782 26894 782 26894 0 Inst_RAM_IO_switch_matrix.S2BEGb1
rlabel metal1 8694 3060 8694 3060 0 Inst_RAM_IO_switch_matrix.S2BEGb2
rlabel metal3 1449 34476 1449 34476 0 Inst_RAM_IO_switch_matrix.S2BEGb3
rlabel metal3 18308 34000 18308 34000 0 Inst_RAM_IO_switch_matrix.S2BEGb4
rlabel metal3 17020 19448 17020 19448 0 Inst_RAM_IO_switch_matrix.S2BEGb5
rlabel metal1 22954 952 22954 952 0 Inst_RAM_IO_switch_matrix.S2BEGb6
rlabel metal2 14582 35530 14582 35530 0 Inst_RAM_IO_switch_matrix.S2BEGb7
rlabel metal2 17388 7956 17388 7956 0 Inst_RAM_IO_switch_matrix.S4BEG0
rlabel metal2 8648 7276 8648 7276 0 Inst_RAM_IO_switch_matrix.S4BEG1
rlabel metal2 18630 9962 18630 9962 0 Inst_RAM_IO_switch_matrix.S4BEG2
rlabel via3 18285 4012 18285 4012 0 Inst_RAM_IO_switch_matrix.S4BEG3
rlabel metal2 13018 6528 13018 6528 0 Inst_RAM_IO_switch_matrix.W1BEG0
rlabel metal1 8096 5678 8096 5678 0 Inst_RAM_IO_switch_matrix.W1BEG1
rlabel via2 5474 3043 5474 3043 0 Inst_RAM_IO_switch_matrix.W1BEG2
rlabel metal1 11914 6290 11914 6290 0 Inst_RAM_IO_switch_matrix.W1BEG3
rlabel metal1 10994 6290 10994 6290 0 Inst_RAM_IO_switch_matrix.W2BEG0
rlabel metal1 5842 4114 5842 4114 0 Inst_RAM_IO_switch_matrix.W2BEG1
rlabel metal1 5290 3026 5290 3026 0 Inst_RAM_IO_switch_matrix.W2BEG2
rlabel metal1 8878 7514 8878 7514 0 Inst_RAM_IO_switch_matrix.W2BEG3
rlabel metal1 11224 6290 11224 6290 0 Inst_RAM_IO_switch_matrix.W2BEG4
rlabel metal2 1610 5066 1610 5066 0 Inst_RAM_IO_switch_matrix.W2BEG5
rlabel metal1 9154 7888 9154 7888 0 Inst_RAM_IO_switch_matrix.W2BEG6
rlabel metal2 13754 9146 13754 9146 0 Inst_RAM_IO_switch_matrix.W2BEG7
rlabel metal1 10442 13158 10442 13158 0 Inst_RAM_IO_switch_matrix.W2BEGb0
rlabel metal1 1886 5780 1886 5780 0 Inst_RAM_IO_switch_matrix.W2BEGb1
rlabel metal2 6026 7038 6026 7038 0 Inst_RAM_IO_switch_matrix.W2BEGb2
rlabel metal1 10580 9690 10580 9690 0 Inst_RAM_IO_switch_matrix.W2BEGb3
rlabel metal1 11500 8602 11500 8602 0 Inst_RAM_IO_switch_matrix.W2BEGb4
rlabel metal1 4002 7514 4002 7514 0 Inst_RAM_IO_switch_matrix.W2BEGb5
rlabel metal1 4784 8942 4784 8942 0 Inst_RAM_IO_switch_matrix.W2BEGb6
rlabel metal2 13662 14688 13662 14688 0 Inst_RAM_IO_switch_matrix.W2BEGb7
rlabel metal1 15870 13498 15870 13498 0 Inst_RAM_IO_switch_matrix.W6BEG0
rlabel metal1 4554 26962 4554 26962 0 Inst_RAM_IO_switch_matrix.W6BEG1
rlabel metal1 5152 15674 5152 15674 0 Inst_RAM_IO_switch_matrix.W6BEG10
rlabel metal1 14858 17204 14858 17204 0 Inst_RAM_IO_switch_matrix.W6BEG11
rlabel metal1 1610 13940 1610 13940 0 Inst_RAM_IO_switch_matrix.W6BEG2
rlabel metal1 14260 15470 14260 15470 0 Inst_RAM_IO_switch_matrix.W6BEG3
rlabel metal1 14214 16558 14214 16558 0 Inst_RAM_IO_switch_matrix.W6BEG4
rlabel metal2 6854 17170 6854 17170 0 Inst_RAM_IO_switch_matrix.W6BEG5
rlabel metal1 6946 11322 6946 11322 0 Inst_RAM_IO_switch_matrix.W6BEG6
rlabel metal2 9246 15912 9246 15912 0 Inst_RAM_IO_switch_matrix.W6BEG7
rlabel metal1 11316 16218 11316 16218 0 Inst_RAM_IO_switch_matrix.W6BEG8
rlabel metal1 3128 15470 3128 15470 0 Inst_RAM_IO_switch_matrix.W6BEG9
rlabel metal1 3726 6290 3726 6290 0 Inst_RAM_IO_switch_matrix.WW4BEG0
rlabel metal1 7130 9588 7130 9588 0 Inst_RAM_IO_switch_matrix.WW4BEG1
rlabel viali 8602 7849 8602 7849 0 Inst_RAM_IO_switch_matrix.WW4BEG10
rlabel metal2 2254 9639 2254 9639 0 Inst_RAM_IO_switch_matrix.WW4BEG11
rlabel metal1 10764 13906 10764 13906 0 Inst_RAM_IO_switch_matrix.WW4BEG12
rlabel metal1 5014 12886 5014 12886 0 Inst_RAM_IO_switch_matrix.WW4BEG13
rlabel metal1 5382 15130 5382 15130 0 Inst_RAM_IO_switch_matrix.WW4BEG14
rlabel metal1 15548 14382 15548 14382 0 Inst_RAM_IO_switch_matrix.WW4BEG15
rlabel metal1 6854 11084 6854 11084 0 Inst_RAM_IO_switch_matrix.WW4BEG2
rlabel metal1 2254 12172 2254 12172 0 Inst_RAM_IO_switch_matrix.WW4BEG3
rlabel metal1 6762 10642 6762 10642 0 Inst_RAM_IO_switch_matrix.WW4BEG4
rlabel metal1 8740 13294 8740 13294 0 Inst_RAM_IO_switch_matrix.WW4BEG5
rlabel metal1 5014 10778 5014 10778 0 Inst_RAM_IO_switch_matrix.WW4BEG6
rlabel metal2 8234 12002 8234 12002 0 Inst_RAM_IO_switch_matrix.WW4BEG7
rlabel metal1 11408 13906 11408 13906 0 Inst_RAM_IO_switch_matrix.WW4BEG8
rlabel metal1 4002 15538 4002 15538 0 Inst_RAM_IO_switch_matrix.WW4BEG9
rlabel metal1 14858 23834 14858 23834 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG0.cus_mux21_inst.A0
rlabel metal1 14812 22746 14812 22746 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG0.cus_mux21_inst.A1
rlabel metal1 14812 24378 14812 24378 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG0.cus_mux21_inst.AIN\[0\]
rlabel metal1 14720 23290 14720 23290 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG0.cus_mux21_inst.AIN\[1\]
rlabel metal2 14306 24650 14306 24650 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG0.cus_mux21_inst._0_
rlabel metal1 14674 24276 14674 24276 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG0.cus_mux21_inst._1_
rlabel metal1 6072 32402 6072 32402 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG1.cus_mux21_inst.A0
rlabel metal1 7038 31994 7038 31994 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG1.cus_mux21_inst.A1
rlabel metal1 6670 32538 6670 32538 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG1.cus_mux21_inst.AIN\[0\]
rlabel metal1 7222 32538 7222 32538 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG1.cus_mux21_inst.AIN\[1\]
rlabel metal1 6854 33082 6854 33082 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG1.cus_mux21_inst._0_
rlabel metal1 7360 33082 7360 33082 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG1.cus_mux21_inst._1_
rlabel metal1 6578 25908 6578 25908 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG2.cus_mux21_inst.A0
rlabel metal1 7774 25262 7774 25262 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG2.cus_mux21_inst.A1
rlabel metal1 8050 25364 8050 25364 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG2.cus_mux21_inst.AIN\[0\]
rlabel metal1 8602 25126 8602 25126 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG2.cus_mux21_inst.AIN\[1\]
rlabel metal2 8142 25908 8142 25908 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG2.cus_mux21_inst._0_
rlabel metal1 9522 26384 9522 26384 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG2.cus_mux21_inst._1_
rlabel metal1 13018 30362 13018 30362 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG3.cus_mux21_inst.A0
rlabel metal1 12972 29818 12972 29818 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG3.cus_mux21_inst.A1
rlabel metal1 12466 30770 12466 30770 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG3.cus_mux21_inst.AIN\[0\]
rlabel metal1 12926 30838 12926 30838 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG3.cus_mux21_inst.AIN\[1\]
rlabel metal1 12052 30634 12052 30634 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG3.cus_mux21_inst._0_
rlabel metal1 12190 30770 12190 30770 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_N4BEG3.cus_mux21_inst._1_
rlabel metal1 16008 20026 16008 20026 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG0.cus_mux21_inst.A0
rlabel metal1 16008 18258 16008 18258 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG0.cus_mux21_inst.A1
rlabel metal1 15502 19210 15502 19210 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG0.cus_mux21_inst.AIN\[0\]
rlabel metal1 16192 18394 16192 18394 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG0.cus_mux21_inst.AIN\[1\]
rlabel metal2 15410 19142 15410 19142 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG0.cus_mux21_inst._0_
rlabel metal2 16330 20094 16330 20094 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG0.cus_mux21_inst._1_
rlabel metal1 6808 23698 6808 23698 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG1.cus_mux21_inst.A0
rlabel metal1 7268 23086 7268 23086 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG1.cus_mux21_inst.A1
rlabel metal1 7406 23664 7406 23664 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG1.cus_mux21_inst.AIN\[0\]
rlabel metal1 8096 21998 8096 21998 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG1.cus_mux21_inst.AIN\[1\]
rlabel metal1 8050 22610 8050 22610 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG1.cus_mux21_inst._0_
rlabel metal1 8372 22066 8372 22066 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG1.cus_mux21_inst._1_
rlabel metal2 9522 24480 9522 24480 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG2.cus_mux21_inst.A0
rlabel metal1 10028 23698 10028 23698 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG2.cus_mux21_inst.A1
rlabel metal1 10534 23732 10534 23732 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG2.cus_mux21_inst.AIN\[0\]
rlabel metal1 10718 23494 10718 23494 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG2.cus_mux21_inst.AIN\[1\]
rlabel metal1 10810 23698 10810 23698 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG2.cus_mux21_inst._0_
rlabel metal1 11546 23766 11546 23766 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG2.cus_mux21_inst._1_
rlabel metal1 16054 26554 16054 26554 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG3.cus_mux21_inst.A0
rlabel metal1 15732 26962 15732 26962 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG3.cus_mux21_inst.A1
rlabel metal1 16238 26928 16238 26928 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG3.cus_mux21_inst.AIN\[0\]
rlabel metal1 16422 25942 16422 25942 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG3.cus_mux21_inst.AIN\[1\]
rlabel metal1 15732 25874 15732 25874 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG3.cus_mux21_inst._0_
rlabel metal1 16192 25942 16192 25942 0 Inst_RAM_IO_switch_matrix.inst_cus_mux81_buf_S4BEG3.cus_mux21_inst._1_
rlabel metal1 2530 42704 2530 42704 0 N1BEG[0]
rlabel metal2 3174 43972 3174 43972 0 N1BEG[1]
rlabel metal1 2990 42772 2990 42772 0 N1BEG[2]
rlabel metal1 3128 43350 3128 43350 0 N1BEG[3]
rlabel metal2 2622 663 2622 663 0 N1END[0]
rlabel metal2 3227 68 3227 68 0 N1END[1]
rlabel metal1 2714 1292 2714 1292 0 N1END[2]
rlabel metal2 3489 68 3489 68 0 N1END[3]
rlabel metal1 3496 42738 3496 42738 0 N2BEG[0]
rlabel metal2 2254 43639 2254 43639 0 N2BEG[1]
rlabel metal1 3818 42330 3818 42330 0 N2BEG[2]
rlabel metal1 4232 42330 4232 42330 0 N2BEG[3]
rlabel metal2 4462 43904 4462 43904 0 N2BEG[4]
rlabel metal1 4462 42738 4462 42738 0 N2BEG[5]
rlabel metal1 4968 42330 4968 42330 0 N2BEG[6]
rlabel metal1 4922 42738 4922 42738 0 N2BEG[7]
rlabel metal1 4600 43418 4600 43418 0 N2BEGb[0]
rlabel metal2 5382 43972 5382 43972 0 N2BEGb[1]
rlabel metal1 5244 43350 5244 43350 0 N2BEGb[2]
rlabel metal2 5750 43904 5750 43904 0 N2BEGb[3]
rlabel metal2 5934 43972 5934 43972 0 N2BEGb[4]
rlabel metal1 5704 42874 5704 42874 0 N2BEGb[5]
rlabel metal1 4738 43078 4738 43078 0 N2BEGb[6]
rlabel metal1 6302 42670 6302 42670 0 N2BEGb[7]
rlabel metal2 5198 534 5198 534 0 N2END[0]
rlabel metal2 5382 704 5382 704 0 N2END[1]
rlabel metal2 5619 68 5619 68 0 N2END[2]
rlabel metal2 5750 398 5750 398 0 N2END[3]
rlabel metal2 5934 1214 5934 1214 0 N2END[4]
rlabel metal2 6118 534 6118 534 0 N2END[5]
rlabel metal2 6249 68 6249 68 0 N2END[6]
rlabel metal2 6486 534 6486 534 0 N2END[7]
rlabel metal2 3726 704 3726 704 0 N2MID[0]
rlabel metal2 3910 1010 3910 1010 0 N2MID[1]
rlabel metal2 4094 636 4094 636 0 N2MID[2]
rlabel metal2 4278 636 4278 636 0 N2MID[3]
rlabel metal2 4462 1010 4462 1010 0 N2MID[4]
rlabel metal2 4646 738 4646 738 0 N2MID[5]
rlabel metal2 4883 68 4883 68 0 N2MID[6]
rlabel metal2 5014 704 5014 704 0 N2MID[7]
rlabel metal1 6624 42330 6624 42330 0 N4BEG[0]
rlabel metal1 8142 43350 8142 43350 0 N4BEG[10]
rlabel metal1 8464 43418 8464 43418 0 N4BEG[11]
rlabel metal2 8694 43163 8694 43163 0 N4BEG[12]
rlabel metal1 8878 43418 8878 43418 0 N4BEG[13]
rlabel metal2 9246 43632 9246 43632 0 N4BEG[14]
rlabel metal1 9292 43418 9292 43418 0 N4BEG[15]
rlabel metal1 6670 42738 6670 42738 0 N4BEG[1]
rlabel metal2 7038 43632 7038 43632 0 N4BEG[2]
rlabel metal2 7222 43428 7222 43428 0 N4BEG[3]
rlabel metal1 7130 43418 7130 43418 0 N4BEG[4]
rlabel metal2 7590 43632 7590 43632 0 N4BEG[5]
rlabel metal1 7452 42058 7452 42058 0 N4BEG[6]
rlabel metal2 7958 42986 7958 42986 0 N4BEG[7]
rlabel metal1 7682 43078 7682 43078 0 N4BEG[8]
rlabel metal1 8188 42738 8188 42738 0 N4BEG[9]
rlabel metal4 644 21216 644 21216 0 N4BEG_outbuf_0.A
rlabel metal1 6164 40970 6164 40970 0 N4BEG_outbuf_0.X
rlabel metal3 828 2176 828 2176 0 N4BEG_outbuf_1.A
rlabel metal1 5658 41616 5658 41616 0 N4BEG_outbuf_1.X
rlabel metal3 17963 19380 17963 19380 0 N4BEG_outbuf_10.A
rlabel metal1 9982 41650 9982 41650 0 N4BEG_outbuf_10.X
rlabel metal3 15801 21148 15801 21148 0 N4BEG_outbuf_11.A
rlabel via1 9434 41582 9434 41582 0 N4BEG_outbuf_11.X
rlabel metal4 1288 18700 1288 18700 0 N4BEG_outbuf_2.A
rlabel metal2 5658 41140 5658 41140 0 N4BEG_outbuf_2.X
rlabel metal2 7222 1581 7222 1581 0 N4BEG_outbuf_3.A
rlabel metal1 6210 41140 6210 41140 0 N4BEG_outbuf_3.X
rlabel metal2 12558 15980 12558 15980 0 N4BEG_outbuf_4.A
rlabel metal1 7498 41072 7498 41072 0 N4BEG_outbuf_4.X
rlabel metal2 14306 6919 14306 6919 0 N4BEG_outbuf_5.A
rlabel metal1 6118 41786 6118 41786 0 N4BEG_outbuf_5.X
rlabel metal2 14490 1428 14490 1428 0 N4BEG_outbuf_6.A
rlabel metal1 7866 40698 7866 40698 0 N4BEG_outbuf_6.X
rlabel metal3 7567 1836 7567 1836 0 N4BEG_outbuf_7.A
rlabel metal1 7682 41616 7682 41616 0 N4BEG_outbuf_7.X
rlabel metal3 21137 19380 21137 19380 0 N4BEG_outbuf_8.A
rlabel metal1 8280 41582 8280 41582 0 N4BEG_outbuf_8.X
rlabel metal1 8556 1734 8556 1734 0 N4BEG_outbuf_9.A
rlabel metal1 8740 41582 8740 41582 0 N4BEG_outbuf_9.X
rlabel metal2 6670 670 6670 670 0 N4END[0]
rlabel metal2 8510 755 8510 755 0 N4END[10]
rlabel metal2 8694 670 8694 670 0 N4END[11]
rlabel metal2 8878 806 8878 806 0 N4END[12]
rlabel metal2 9062 143 9062 143 0 N4END[13]
rlabel metal2 9246 1554 9246 1554 0 N4END[14]
rlabel metal2 9430 415 9430 415 0 N4END[15]
rlabel metal2 6854 704 6854 704 0 N4END[1]
rlabel metal2 7091 68 7091 68 0 N4END[2]
rlabel metal2 7222 636 7222 636 0 N4END[3]
rlabel metal2 7459 68 7459 68 0 N4END[4]
rlabel metal2 7590 806 7590 806 0 N4END[5]
rlabel metal2 7774 942 7774 942 0 N4END[6]
rlabel metal2 7905 68 7905 68 0 N4END[7]
rlabel metal2 8004 3026 8004 3026 0 N4END[8]
rlabel metal1 8234 3026 8234 3026 0 N4END[9]
rlabel metal3 21237 7140 21237 7140 0 RAM2FAB_D0_I0
rlabel metal3 22525 7684 22525 7684 0 RAM2FAB_D0_I1
rlabel metal3 21789 8228 21789 8228 0 RAM2FAB_D0_I2
rlabel metal3 22525 8772 22525 8772 0 RAM2FAB_D0_I3
rlabel metal1 13570 3060 13570 3060 0 RAM2FAB_D1_I0
rlabel metal3 22525 5508 22525 5508 0 RAM2FAB_D1_I1
rlabel metal3 21237 6052 21237 6052 0 RAM2FAB_D1_I2
rlabel metal3 22525 6596 22525 6596 0 RAM2FAB_D1_I3
rlabel metal3 21996 2788 21996 2788 0 RAM2FAB_D2_I0
rlabel metal3 22525 3332 22525 3332 0 RAM2FAB_D2_I1
rlabel metal3 21536 3876 21536 3876 0 RAM2FAB_D2_I2
rlabel metal3 16008 1836 16008 1836 0 RAM2FAB_D2_I3
rlabel metal3 20869 612 20869 612 0 RAM2FAB_D3_I0
rlabel metal3 22525 1156 22525 1156 0 RAM2FAB_D3_I1
rlabel metal3 21904 1700 21904 1700 0 RAM2FAB_D3_I2
rlabel metal3 22617 2244 22617 2244 0 RAM2FAB_D3_I3
rlabel metal2 9614 908 9614 908 0 S1BEG[0]
rlabel metal2 9851 68 9851 68 0 S1BEG[1]
rlabel metal2 10035 68 10035 68 0 S1BEG[2]
rlabel metal2 10166 908 10166 908 0 S1BEG[3]
rlabel metal2 9614 43598 9614 43598 0 S1END[0]
rlabel metal2 9798 44193 9798 44193 0 S1END[1]
rlabel metal2 9982 43938 9982 43938 0 S1END[2]
rlabel metal2 10166 43938 10166 43938 0 S1END[3]
rlabel metal2 11769 68 11769 68 0 S2BEG[0]
rlabel metal2 12006 908 12006 908 0 S2BEG[1]
rlabel metal2 12190 636 12190 636 0 S2BEG[2]
rlabel metal2 12374 806 12374 806 0 S2BEG[3]
rlabel metal2 12558 636 12558 636 0 S2BEG[4]
rlabel metal2 12742 670 12742 670 0 S2BEG[5]
rlabel metal2 12926 364 12926 364 0 S2BEG[6]
rlabel metal2 13110 908 13110 908 0 S2BEG[7]
rlabel metal2 10350 1486 10350 1486 0 S2BEGb[0]
rlabel metal2 10534 908 10534 908 0 S2BEGb[1]
rlabel metal2 10718 670 10718 670 0 S2BEGb[2]
rlabel metal2 10955 68 10955 68 0 S2BEGb[3]
rlabel metal2 11086 670 11086 670 0 S2BEGb[4]
rlabel metal2 11217 68 11217 68 0 S2BEGb[5]
rlabel metal2 11507 68 11507 68 0 S2BEGb[6]
rlabel metal2 11638 483 11638 483 0 S2BEGb[7]
rlabel metal2 10350 44074 10350 44074 0 S2END[0]
rlabel metal2 10534 43921 10534 43921 0 S2END[1]
rlabel metal2 10718 44193 10718 44193 0 S2END[2]
rlabel metal2 10902 44074 10902 44074 0 S2END[3]
rlabel metal2 11086 43717 11086 43717 0 S2END[4]
rlabel metal2 11270 44125 11270 44125 0 S2END[5]
rlabel metal2 11454 44074 11454 44074 0 S2END[6]
rlabel metal2 11638 44193 11638 44193 0 S2END[7]
rlabel metal2 11822 43598 11822 43598 0 S2MID[0]
rlabel metal2 12006 43904 12006 43904 0 S2MID[1]
rlabel metal2 12190 44142 12190 44142 0 S2MID[2]
rlabel metal2 12374 44193 12374 44193 0 S2MID[3]
rlabel metal2 12558 44057 12558 44057 0 S2MID[4]
rlabel metal2 12742 43938 12742 43938 0 S2MID[5]
rlabel metal2 12926 44193 12926 44193 0 S2MID[6]
rlabel metal2 13110 44057 13110 44057 0 S2MID[7]
rlabel metal2 13294 806 13294 806 0 S4BEG[0]
rlabel metal2 15081 68 15081 68 0 S4BEG[10]
rlabel metal2 15318 1758 15318 1758 0 S4BEG[11]
rlabel metal2 15555 68 15555 68 0 S4BEG[12]
rlabel metal2 15686 1350 15686 1350 0 S4BEG[13]
rlabel metal1 16422 2890 16422 2890 0 S4BEG[14]
rlabel metal1 16744 2822 16744 2822 0 S4BEG[15]
rlabel metal2 13478 908 13478 908 0 S4BEG[1]
rlabel metal2 13662 772 13662 772 0 S4BEG[2]
rlabel metal2 13846 483 13846 483 0 S4BEG[3]
rlabel metal2 14030 738 14030 738 0 S4BEG[4]
rlabel metal2 14267 68 14267 68 0 S4BEG[5]
rlabel metal2 14398 755 14398 755 0 S4BEG[6]
rlabel metal2 14582 687 14582 687 0 S4BEG[7]
rlabel metal2 14819 68 14819 68 0 S4BEG[8]
rlabel metal2 14950 772 14950 772 0 S4BEG[9]
rlabel metal1 13570 42262 13570 42262 0 S4BEG_outbuf_0.A
rlabel metal1 14766 39882 14766 39882 0 S4BEG_outbuf_0.X
rlabel metal1 14674 42160 14674 42160 0 S4BEG_outbuf_1.A
rlabel metal3 18239 2652 18239 2652 0 S4BEG_outbuf_1.X
rlabel metal1 16514 41786 16514 41786 0 S4BEG_outbuf_10.A
rlabel metal2 20424 33388 20424 33388 0 S4BEG_outbuf_10.X
rlabel metal1 15548 41582 15548 41582 0 S4BEG_outbuf_11.A
rlabel metal2 14306 21692 14306 21692 0 S4BEG_outbuf_11.X
rlabel metal1 14490 42262 14490 42262 0 S4BEG_outbuf_2.A
rlabel metal4 17480 17340 17480 17340 0 S4BEG_outbuf_2.X
rlabel metal1 14996 42262 14996 42262 0 S4BEG_outbuf_3.A
rlabel metal3 17687 884 17687 884 0 S4BEG_outbuf_3.X
rlabel metal1 15364 42194 15364 42194 0 S4BEG_outbuf_4.A
rlabel metal1 19274 12614 19274 12614 0 S4BEG_outbuf_4.X
rlabel metal1 14904 41582 14904 41582 0 S4BEG_outbuf_5.A
rlabel metal3 19780 9452 19780 9452 0 S4BEG_outbuf_5.X
rlabel metal1 15870 42194 15870 42194 0 S4BEG_outbuf_6.A
rlabel metal3 16652 29036 16652 29036 0 S4BEG_outbuf_6.X
rlabel metal1 15364 41514 15364 41514 0 S4BEG_outbuf_7.A
rlabel metal3 14306 34476 14306 34476 0 S4BEG_outbuf_7.X
rlabel metal1 16008 41786 16008 41786 0 S4BEG_outbuf_8.A
rlabel metal3 15341 32844 15341 32844 0 S4BEG_outbuf_8.X
rlabel metal1 15318 41650 15318 41650 0 S4BEG_outbuf_9.A
rlabel metal1 18170 7514 18170 7514 0 S4BEG_outbuf_9.X
rlabel metal2 13294 43870 13294 43870 0 S4END[0]
rlabel metal1 15226 41038 15226 41038 0 S4END[10]
rlabel metal2 15318 44261 15318 44261 0 S4END[11]
rlabel metal2 15502 43632 15502 43632 0 S4END[12]
rlabel metal2 15686 44261 15686 44261 0 S4END[13]
rlabel metal1 16008 41106 16008 41106 0 S4END[14]
rlabel metal2 16054 43700 16054 43700 0 S4END[15]
rlabel metal2 13478 44057 13478 44057 0 S4END[1]
rlabel metal2 13662 44193 13662 44193 0 S4END[2]
rlabel metal2 13846 43598 13846 43598 0 S4END[3]
rlabel metal2 14030 44193 14030 44193 0 S4END[4]
rlabel metal2 14214 44193 14214 44193 0 S4END[5]
rlabel metal2 14398 43054 14398 43054 0 S4END[6]
rlabel metal1 14720 41106 14720 41106 0 S4END[7]
rlabel metal1 14720 41174 14720 41174 0 S4END[8]
rlabel metal1 15318 41106 15318 41106 0 S4END[9]
rlabel metal1 19504 13906 19504 13906 0 UserCLK
rlabel metal1 17664 40698 17664 40698 0 UserCLKo
rlabel metal3 383 4964 383 4964 0 W1BEG[0]
rlabel metal2 4094 4352 4094 4352 0 W1BEG[1]
rlabel metal2 4186 5508 4186 5508 0 W1BEG[2]
rlabel metal2 4094 5831 4094 5831 0 W1BEG[3]
rlabel metal2 2898 2295 2898 2295 0 W2BEG[0]
rlabel metal3 682 6324 682 6324 0 W2BEG[1]
rlabel metal3 1303 6596 1303 6596 0 W2BEG[2]
rlabel metal2 4094 6477 4094 6477 0 W2BEG[3]
rlabel metal2 1610 2145 1610 2145 0 W2BEG[4]
rlabel metal3 2154 7412 2154 7412 0 W2BEG[5]
rlabel metal3 1441 7684 1441 7684 0 W2BEG[6]
rlabel metal2 2346 2689 2346 2689 0 W2BEG[7]
rlabel metal2 2668 2278 2668 2278 0 W2BEGb[0]
rlabel metal3 2476 8500 2476 8500 0 W2BEGb[1]
rlabel metal3 774 8772 774 8772 0 W2BEGb[2]
rlabel metal3 2430 9044 2430 9044 0 W2BEGb[3]
rlabel metal1 1518 2074 1518 2074 0 W2BEGb[4]
rlabel metal3 1740 9588 1740 9588 0 W2BEGb[5]
rlabel metal3 912 9860 912 9860 0 W2BEGb[6]
rlabel metal2 3174 5440 3174 5440 0 W2BEGb[7]
rlabel metal3 544 14756 544 14756 0 W6BEG[0]
rlabel metal3 475 17476 475 17476 0 W6BEG[10]
rlabel metal3 475 17748 475 17748 0 W6BEG[11]
rlabel metal3 291 15028 291 15028 0 W6BEG[1]
rlabel metal3 866 15300 866 15300 0 W6BEG[2]
rlabel metal3 567 15572 567 15572 0 W6BEG[3]
rlabel metal3 866 15844 866 15844 0 W6BEG[4]
rlabel metal3 199 16116 199 16116 0 W6BEG[5]
rlabel via2 4002 16405 4002 16405 0 W6BEG[6]
rlabel metal2 3634 16711 3634 16711 0 W6BEG[7]
rlabel metal3 958 16932 958 16932 0 W6BEG[8]
rlabel metal3 774 17204 774 17204 0 W6BEG[9]
rlabel metal3 3404 10268 3404 10268 0 WW4BEG[0]
rlabel metal1 2392 8602 2392 8602 0 WW4BEG[10]
rlabel metal3 2292 13396 2292 13396 0 WW4BEG[11]
rlabel metal3 567 13668 567 13668 0 WW4BEG[12]
rlabel metal3 774 13940 774 13940 0 WW4BEG[13]
rlabel metal3 912 14212 912 14212 0 WW4BEG[14]
rlabel metal3 1004 14484 1004 14484 0 WW4BEG[15]
rlabel metal2 4002 10455 4002 10455 0 WW4BEG[1]
rlabel metal3 3588 10880 3588 10880 0 WW4BEG[2]
rlabel metal3 1487 11220 1487 11220 0 WW4BEG[3]
rlabel metal3 590 11492 590 11492 0 WW4BEG[4]
rlabel metal3 475 11764 475 11764 0 WW4BEG[5]
rlabel metal2 4094 11679 4094 11679 0 WW4BEG[6]
rlabel metal2 4002 12359 4002 12359 0 WW4BEG[7]
rlabel metal1 3450 5134 3450 5134 0 WW4BEG[8]
rlabel metal3 1464 12852 1464 12852 0 WW4BEG[9]
rlabel metal2 20286 26724 20286 26724 0 data_inbuf_0.X
rlabel metal1 20562 28084 20562 28084 0 data_inbuf_1.X
rlabel metal1 20194 31824 20194 31824 0 data_inbuf_10.X
rlabel metal2 18906 33252 18906 33252 0 data_inbuf_11.X
rlabel metal2 19182 33762 19182 33762 0 data_inbuf_12.X
rlabel metal1 19872 34170 19872 34170 0 data_inbuf_13.X
rlabel metal1 19642 34612 19642 34612 0 data_inbuf_14.X
rlabel metal1 19228 34714 19228 34714 0 data_inbuf_15.X
rlabel metal1 20010 34578 20010 34578 0 data_inbuf_16.X
rlabel metal2 18446 35802 18446 35802 0 data_inbuf_17.X
rlabel metal1 21114 36720 21114 36720 0 data_inbuf_18.X
rlabel metal1 19918 37196 19918 37196 0 data_inbuf_19.X
rlabel metal1 20056 27914 20056 27914 0 data_inbuf_2.X
rlabel metal1 20102 37434 20102 37434 0 data_inbuf_20.X
rlabel metal1 20654 37434 20654 37434 0 data_inbuf_21.X
rlabel metal1 20378 37434 20378 37434 0 data_inbuf_22.X
rlabel metal2 18630 38148 18630 38148 0 data_inbuf_23.X
rlabel metal1 20056 37978 20056 37978 0 data_inbuf_24.X
rlabel metal1 18446 38522 18446 38522 0 data_inbuf_25.X
rlabel metal1 19734 39032 19734 39032 0 data_inbuf_26.X
rlabel metal2 18078 39780 18078 39780 0 data_inbuf_27.X
rlabel metal1 20286 39610 20286 39610 0 data_inbuf_28.X
rlabel metal2 19872 39882 19872 39882 0 data_inbuf_29.X
rlabel metal1 20654 29172 20654 29172 0 data_inbuf_3.X
rlabel metal1 17434 40460 17434 40460 0 data_inbuf_30.X
rlabel metal1 18906 40630 18906 40630 0 data_inbuf_31.X
rlabel metal1 20654 29274 20654 29274 0 data_inbuf_4.X
rlabel metal1 20286 29580 20286 29580 0 data_inbuf_5.X
rlabel metal1 19136 30362 19136 30362 0 data_inbuf_6.X
rlabel metal1 20194 31450 20194 31450 0 data_inbuf_7.X
rlabel metal1 19182 30566 19182 30566 0 data_inbuf_8.X
rlabel metal1 19458 31824 19458 31824 0 data_inbuf_9.X
rlabel metal2 20102 26792 20102 26792 0 data_outbuf_0.X
rlabel metal1 20470 28186 20470 28186 0 data_outbuf_1.X
rlabel metal2 20010 32232 20010 32232 0 data_outbuf_10.X
rlabel metal1 19964 33626 19964 33626 0 data_outbuf_11.X
rlabel metal1 20608 34102 20608 34102 0 data_outbuf_12.X
rlabel metal1 20378 34714 20378 34714 0 data_outbuf_13.X
rlabel metal1 19458 34476 19458 34476 0 data_outbuf_14.X
rlabel metal1 19964 35802 19964 35802 0 data_outbuf_15.X
rlabel metal1 19826 34714 19826 34714 0 data_outbuf_16.X
rlabel viali 20282 36142 20282 36142 0 data_outbuf_17.X
rlabel metal1 20976 36890 20976 36890 0 data_outbuf_18.X
rlabel metal2 19734 37604 19734 37604 0 data_outbuf_19.X
rlabel metal1 20930 28492 20930 28492 0 data_outbuf_2.X
rlabel metal1 20608 37706 20608 37706 0 data_outbuf_20.X
rlabel metal1 20654 37978 20654 37978 0 data_outbuf_21.X
rlabel metal1 20654 38454 20654 38454 0 data_outbuf_22.X
rlabel metal1 20240 38522 20240 38522 0 data_outbuf_23.X
rlabel metal1 21068 40018 21068 40018 0 data_outbuf_24.X
rlabel metal2 18814 39202 18814 39202 0 data_outbuf_25.X
rlabel metal1 20516 39270 20516 39270 0 data_outbuf_26.X
rlabel metal2 19182 40290 19182 40290 0 data_outbuf_27.X
rlabel metal2 19734 39321 19734 39321 0 data_outbuf_28.X
rlabel metal1 20470 40052 20470 40052 0 data_outbuf_29.X
rlabel metal2 20470 29410 20470 29410 0 data_outbuf_3.X
rlabel metal1 20746 40052 20746 40052 0 data_outbuf_30.X
rlabel metal1 18814 41140 18814 41140 0 data_outbuf_31.X
rlabel metal1 20654 29750 20654 29750 0 data_outbuf_4.X
rlabel metal1 20378 29818 20378 29818 0 data_outbuf_5.X
rlabel metal1 20792 31178 20792 31178 0 data_outbuf_6.X
rlabel metal1 20930 31994 20930 31994 0 data_outbuf_7.X
rlabel metal1 20286 31926 20286 31926 0 data_outbuf_8.X
rlabel metal1 19596 31994 19596 31994 0 data_outbuf_9.X
rlabel metal1 12788 21658 12788 21658 0 net1
rlabel metal1 3496 23290 3496 23290 0 net10
rlabel metal1 17756 14926 17756 14926 0 net100
rlabel metal1 2484 1190 2484 1190 0 net101
rlabel metal1 3450 2040 3450 2040 0 net102
rlabel metal1 2944 1326 2944 1326 0 net103
rlabel metal2 12972 30804 12972 30804 0 net104
rlabel metal3 14812 17476 14812 17476 0 net105
rlabel metal1 2622 1428 2622 1428 0 net106
rlabel metal1 5428 2618 5428 2618 0 net107
rlabel metal3 20700 816 20700 816 0 net108
rlabel metal3 6716 17884 6716 17884 0 net109
rlabel metal2 3266 23800 3266 23800 0 net11
rlabel metal1 8142 2346 8142 2346 0 net110
rlabel metal3 7935 37332 7935 37332 0 net111
rlabel metal2 9798 14144 9798 14144 0 net112
rlabel metal3 14444 13736 14444 13736 0 net113
rlabel metal1 4186 2074 4186 2074 0 net114
rlabel metal1 3910 6664 3910 6664 0 net115
rlabel metal3 1748 12988 1748 12988 0 net116
rlabel metal1 4784 2074 4784 2074 0 net117
rlabel metal1 7222 20774 7222 20774 0 net118
rlabel metal1 598 13668 598 13668 0 net119
rlabel via2 4002 23613 4002 23613 0 net12
rlabel metal4 5520 15980 5520 15980 0 net120
rlabel metal1 14306 13430 14306 13430 0 net121
rlabel metal2 8234 2618 8234 2618 0 net122
rlabel metal2 7820 2414 7820 2414 0 net123
rlabel metal1 8556 2414 8556 2414 0 net124
rlabel metal3 8303 2244 8303 2244 0 net125
rlabel metal1 8832 2006 8832 2006 0 net126
rlabel metal2 8050 1700 8050 1700 0 net127
rlabel metal1 5704 1326 5704 1326 0 net128
rlabel metal3 7337 1292 7337 1292 0 net129
rlabel metal1 5842 19448 5842 19448 0 net13
rlabel metal4 10396 9180 10396 9180 0 net130
rlabel metal1 7222 3366 7222 3366 0 net131
rlabel metal1 6762 1938 6762 1938 0 net132
rlabel metal1 7544 2414 7544 2414 0 net133
rlabel metal1 7268 2006 7268 2006 0 net134
rlabel metal1 7728 2414 7728 2414 0 net135
rlabel metal1 7774 2074 7774 2074 0 net136
rlabel metal2 19734 7395 19734 7395 0 net137
rlabel metal1 18630 6630 18630 6630 0 net138
rlabel metal1 19228 6766 19228 6766 0 net139
rlabel metal2 4048 18802 4048 18802 0 net14
rlabel metal1 18308 9894 18308 9894 0 net140
rlabel metal1 16790 4522 16790 4522 0 net141
rlabel metal1 18078 3536 18078 3536 0 net142
rlabel metal2 15134 5015 15134 5015 0 net143
rlabel metal1 16590 6698 16590 6698 0 net144
rlabel metal2 15962 5083 15962 5083 0 net145
rlabel metal2 17250 4335 17250 4335 0 net146
rlabel metal2 20010 3774 20010 3774 0 net147
rlabel metal1 14674 4080 14674 4080 0 net148
rlabel via1 14577 6290 14577 6290 0 net149
rlabel metal1 3634 19958 3634 19958 0 net15
rlabel via2 18446 3723 18446 3723 0 net150
rlabel metal1 19534 7786 19534 7786 0 net151
rlabel via1 18073 9554 18073 9554 0 net152
rlabel metal1 15652 16626 15652 16626 0 net153
rlabel metal2 7360 38828 7360 38828 0 net154
rlabel metal1 10442 17544 10442 17544 0 net155
rlabel metal1 10994 33422 10994 33422 0 net156
rlabel metal1 9936 42602 9936 42602 0 net157
rlabel metal3 6417 36788 6417 36788 0 net158
rlabel metal3 10741 35836 10741 35836 0 net159
rlabel metal1 1702 20026 1702 20026 0 net16
rlabel metal3 10097 42364 10097 42364 0 net160
rlabel metal1 9062 35054 9062 35054 0 net161
rlabel metal2 11914 26248 11914 26248 0 net162
rlabel metal2 7912 40188 7912 40188 0 net163
rlabel metal1 10718 37230 10718 37230 0 net164
rlabel metal1 11638 37638 11638 37638 0 net165
rlabel metal1 5796 36006 5796 36006 0 net166
rlabel metal1 920 42602 920 42602 0 net167
rlabel metal1 10810 34680 10810 34680 0 net168
rlabel metal1 12834 42568 12834 42568 0 net169
rlabel via2 1702 18819 1702 18819 0 net17
rlabel metal4 12972 27056 12972 27056 0 net170
rlabel metal2 13938 43367 13938 43367 0 net171
rlabel metal1 13202 42534 13202 42534 0 net172
rlabel metal3 19228 19652 19228 19652 0 net173
rlabel metal1 15824 40970 15824 40970 0 net174
rlabel metal1 18630 42670 18630 42670 0 net175
rlabel metal1 16242 41578 16242 41578 0 net176
rlabel metal1 17250 42126 17250 42126 0 net177
rlabel metal1 16652 41242 16652 41242 0 net178
rlabel metal1 17158 40902 17158 40902 0 net179
rlabel metal1 3404 22134 3404 22134 0 net18
rlabel metal1 13754 42636 13754 42636 0 net180
rlabel metal4 14444 28492 14444 28492 0 net181
rlabel metal2 13846 42296 13846 42296 0 net182
rlabel metal1 14674 42704 14674 42704 0 net183
rlabel metal1 13110 42636 13110 42636 0 net184
rlabel metal1 13984 41786 13984 41786 0 net185
rlabel metal2 14720 42636 14720 42636 0 net186
rlabel metal1 14996 41242 14996 41242 0 net187
rlabel metal1 15410 41242 15410 41242 0 net188
rlabel metal1 21252 6630 21252 6630 0 net189
rlabel metal1 3588 21114 3588 21114 0 net19
rlabel metal1 21298 8602 21298 8602 0 net190
rlabel metal1 20562 10030 20562 10030 0 net191
rlabel metal1 20976 10710 20976 10710 0 net192
rlabel metal1 21298 16116 21298 16116 0 net193
rlabel metal1 20608 16490 20608 16490 0 net194
rlabel metal1 21298 17238 21298 17238 0 net195
rlabel metal3 20010 20740 20010 20740 0 net196
rlabel metal1 21206 13974 21206 13974 0 net197
rlabel metal1 21206 14382 21206 14382 0 net198
rlabel metal2 22678 18564 22678 18564 0 net199
rlabel metal1 5934 21862 5934 21862 0 net2
rlabel metal2 2254 21845 2254 21845 0 net20
rlabel metal2 21160 18836 21160 18836 0 net200
rlabel metal1 20608 12614 20608 12614 0 net201
rlabel metal1 20378 16966 20378 16966 0 net202
rlabel metal1 21206 12886 21206 12886 0 net203
rlabel metal1 22862 32164 22862 32164 0 net204
rlabel metal1 20102 24582 20102 24582 0 net205
rlabel metal1 21252 25262 21252 25262 0 net206
rlabel metal2 19642 25704 19642 25704 0 net207
rlabel metal1 21206 26384 21206 26384 0 net208
rlabel metal1 21390 22474 21390 22474 0 net209
rlabel metal2 7222 24956 7222 24956 0 net21
rlabel metal1 20884 22610 20884 22610 0 net210
rlabel metal1 21114 23086 21114 23086 0 net211
rlabel metal1 21114 24174 21114 24174 0 net212
rlabel metal1 21298 20468 21298 20468 0 net213
rlabel metal1 20976 30838 20976 30838 0 net214
rlabel metal2 20700 20740 20700 20740 0 net215
rlabel metal1 21206 22066 21206 22066 0 net216
rlabel metal1 21206 18360 21206 18360 0 net217
rlabel metal1 22034 18734 22034 18734 0 net218
rlabel metal1 21160 18938 21160 18938 0 net219
rlabel metal3 2346 20672 2346 20672 0 net22
rlabel metal2 20378 20434 20378 20434 0 net220
rlabel metal1 21344 27098 21344 27098 0 net221
rlabel metal1 21298 32436 21298 32436 0 net222
rlabel metal1 20102 33558 20102 33558 0 net223
rlabel metal2 21022 34510 21022 34510 0 net224
rlabel metal2 21298 34884 21298 34884 0 net225
rlabel metal1 21022 34646 21022 34646 0 net226
rlabel metal1 21298 35088 21298 35088 0 net227
rlabel metal1 21206 35666 21206 35666 0 net228
rlabel metal1 20792 36074 20792 36074 0 net229
rlabel metal2 9430 30430 9430 30430 0 net23
rlabel metal1 21298 36788 21298 36788 0 net230
rlabel metal1 21160 37230 21160 37230 0 net231
rlabel metal2 21022 27914 21022 27914 0 net232
rlabel metal1 21252 37842 21252 37842 0 net233
rlabel metal1 21298 38284 21298 38284 0 net234
rlabel metal1 21206 39032 21206 39032 0 net235
rlabel metal1 20654 39066 20654 39066 0 net236
rlabel metal1 21206 40120 21206 40120 0 net237
rlabel metal1 20700 39542 20700 39542 0 net238
rlabel metal1 21068 40698 21068 40698 0 net239
rlabel metal1 2852 33558 2852 33558 0 net24
rlabel metal1 20608 40630 20608 40630 0 net240
rlabel metal1 19458 39542 19458 39542 0 net241
rlabel metal1 20654 39882 20654 39882 0 net242
rlabel metal1 20930 28084 20930 28084 0 net243
rlabel metal1 20470 40154 20470 40154 0 net244
rlabel metal1 18722 40902 18722 40902 0 net245
rlabel metal1 21298 28492 21298 28492 0 net246
rlabel metal1 21022 29206 21022 29206 0 net247
rlabel metal1 21206 29614 21206 29614 0 net248
rlabel metal1 21114 30294 21114 30294 0 net249
rlabel metal2 8142 17986 8142 17986 0 net25
rlabel metal2 21298 31212 21298 31212 0 net250
rlabel metal2 21344 32844 21344 32844 0 net251
rlabel metal1 21160 31790 21160 31790 0 net252
rlabel metal1 15916 40154 15916 40154 0 net253
rlabel metal1 18308 40358 18308 40358 0 net254
rlabel metal1 20194 39304 20194 39304 0 net255
rlabel metal1 17848 40630 17848 40630 0 net256
rlabel metal2 19412 40970 19412 40970 0 net257
rlabel metal2 18078 40239 18078 40239 0 net258
rlabel metal2 17526 40749 17526 40749 0 net259
rlabel metal1 7590 31960 7590 31960 0 net26
rlabel metal1 20516 40902 20516 40902 0 net260
rlabel metal1 18400 40154 18400 40154 0 net261
rlabel metal2 18630 40477 18630 40477 0 net262
rlabel metal2 19458 40154 19458 40154 0 net263
rlabel metal1 18998 42296 18998 42296 0 net264
rlabel metal1 18124 41242 18124 41242 0 net265
rlabel metal1 20010 41242 20010 41242 0 net266
rlabel metal1 21206 41242 21206 41242 0 net267
rlabel metal1 18584 41786 18584 41786 0 net268
rlabel metal1 17848 40902 17848 40902 0 net269
rlabel metal2 3358 28832 3358 28832 0 net27
rlabel metal2 17802 40375 17802 40375 0 net270
rlabel metal1 17802 41242 17802 41242 0 net271
rlabel metal1 19458 40120 19458 40120 0 net272
rlabel via2 16606 41021 16606 41021 0 net273
rlabel metal1 2346 42602 2346 42602 0 net274
rlabel metal2 2714 42194 2714 42194 0 net275
rlabel metal2 2530 42262 2530 42262 0 net276
rlabel metal1 3128 42670 3128 42670 0 net277
rlabel metal1 2300 42330 2300 42330 0 net278
rlabel metal1 3266 41786 3266 41786 0 net279
rlabel metal2 1794 31076 1794 31076 0 net28
rlabel metal1 3864 41786 3864 41786 0 net280
rlabel metal1 9246 42296 9246 42296 0 net281
rlabel metal2 2806 42466 2806 42466 0 net282
rlabel metal1 4922 42228 4922 42228 0 net283
rlabel metal1 5060 41242 5060 41242 0 net284
rlabel metal1 4186 41786 4186 41786 0 net285
rlabel metal1 4692 41786 4692 41786 0 net286
rlabel metal2 4094 41973 4094 41973 0 net287
rlabel metal1 5106 41786 5106 41786 0 net288
rlabel metal2 5520 41820 5520 41820 0 net289
rlabel metal1 8004 27370 8004 27370 0 net29
rlabel metal1 5474 41208 5474 41208 0 net290
rlabel metal2 6026 39491 6026 39491 0 net291
rlabel metal1 6026 39610 6026 39610 0 net292
rlabel metal2 5750 41956 5750 41956 0 net293
rlabel metal1 9798 41548 9798 41548 0 net294
rlabel metal1 8878 41446 8878 41446 0 net295
rlabel metal1 9568 41990 9568 41990 0 net296
rlabel metal2 10626 42772 10626 42772 0 net297
rlabel metal1 8970 41684 8970 41684 0 net298
rlabel metal1 11546 32538 11546 32538 0 net299
rlabel metal1 9384 18394 9384 18394 0 net3
rlabel metal2 15180 26588 15180 26588 0 net30
rlabel metal1 5566 41786 5566 41786 0 net300
rlabel metal1 5750 41208 5750 41208 0 net301
rlabel metal1 6256 42058 6256 42058 0 net302
rlabel metal1 7360 40970 7360 40970 0 net303
rlabel metal2 6026 42432 6026 42432 0 net304
rlabel via2 8418 41259 8418 41259 0 net305
rlabel metal1 7820 41514 7820 41514 0 net306
rlabel metal1 7590 41786 7590 41786 0 net307
rlabel metal1 8234 41786 8234 41786 0 net308
rlabel metal2 9706 2414 9706 2414 0 net309
rlabel metal1 17388 17578 17388 17578 0 net31
rlabel metal1 9936 1326 9936 1326 0 net310
rlabel metal2 9430 1054 9430 1054 0 net311
rlabel metal1 10810 1938 10810 1938 0 net312
rlabel metal1 12052 1326 12052 1326 0 net313
rlabel metal1 12190 1904 12190 1904 0 net314
rlabel metal1 11822 1326 11822 1326 0 net315
rlabel metal1 12374 1360 12374 1360 0 net316
rlabel metal2 12742 2822 12742 2822 0 net317
rlabel metal2 13202 2482 13202 2482 0 net318
rlabel metal2 12466 1836 12466 1836 0 net319
rlabel metal1 1978 29546 1978 29546 0 net32
rlabel metal1 13110 1938 13110 1938 0 net320
rlabel metal1 9614 2992 9614 2992 0 net321
rlabel metal2 10488 2822 10488 2822 0 net322
rlabel metal2 8556 2278 8556 2278 0 net323
rlabel metal1 10994 2040 10994 2040 0 net324
rlabel metal2 9476 1326 9476 1326 0 net325
rlabel metal1 10718 1326 10718 1326 0 net326
rlabel metal1 10902 2618 10902 2618 0 net327
rlabel metal1 11454 2006 11454 2006 0 net328
rlabel metal1 14030 1326 14030 1326 0 net329
rlabel metal2 1610 23001 1610 23001 0 net33
rlabel metal1 15824 3094 15824 3094 0 net330
rlabel metal1 16698 3434 16698 3434 0 net331
rlabel metal1 15502 2414 15502 2414 0 net332
rlabel metal1 16606 2448 16606 2448 0 net333
rlabel metal1 16790 2992 16790 2992 0 net334
rlabel metal1 17710 3094 17710 3094 0 net335
rlabel metal1 13846 2040 13846 2040 0 net336
rlabel metal1 14858 2822 14858 2822 0 net337
rlabel metal2 15226 1768 15226 1768 0 net338
rlabel metal1 15134 2414 15134 2414 0 net339
rlabel via1 2714 26979 2714 26979 0 net34
rlabel metal2 14950 2652 14950 2652 0 net340
rlabel metal1 16606 1326 16606 1326 0 net341
rlabel metal1 15364 2822 15364 2822 0 net342
rlabel metal1 15916 2006 15916 2006 0 net343
rlabel viali 16045 2414 16045 2414 0 net344
rlabel metal1 18906 40528 18906 40528 0 net345
rlabel metal1 3726 2346 3726 2346 0 net346
rlabel metal2 3910 2587 3910 2587 0 net347
rlabel metal1 4922 3094 4922 3094 0 net348
rlabel metal1 11822 3672 11822 3672 0 net349
rlabel metal1 1978 28424 1978 28424 0 net35
rlabel metal1 2576 1938 2576 1938 0 net350
rlabel metal2 2622 2686 2622 2686 0 net351
rlabel metal1 4140 3162 4140 3162 0 net352
rlabel metal1 5842 6392 5842 6392 0 net353
rlabel metal2 1518 1003 1518 1003 0 net354
rlabel metal2 3450 5338 3450 5338 0 net355
rlabel metal1 6210 5610 6210 5610 0 net356
rlabel metal1 1886 2414 1886 2414 0 net357
rlabel metal1 2024 2006 2024 2006 0 net358
rlabel metal2 1518 5984 1518 5984 0 net359
rlabel metal3 7452 23256 7452 23256 0 net36
rlabel metal1 6302 7446 6302 7446 0 net360
rlabel metal1 6072 7786 6072 7786 0 net361
rlabel metal2 1518 2669 1518 2669 0 net362
rlabel metal1 4048 8058 4048 8058 0 net363
rlabel metal2 1518 5321 1518 5321 0 net364
rlabel metal2 1886 4845 1886 4845 0 net365
rlabel via2 1794 13923 1794 13923 0 net366
rlabel metal2 1518 16286 1518 16286 0 net367
rlabel metal2 1978 17731 1978 17731 0 net368
rlabel metal1 598 22066 598 22066 0 net369
rlabel metal1 4784 28050 4784 28050 0 net37
rlabel viali 6477 11730 6477 11730 0 net370
rlabel metal2 13754 14127 13754 14127 0 net371
rlabel metal2 15272 13396 15272 13396 0 net372
rlabel metal2 2162 14297 2162 14297 0 net373
rlabel metal3 5014 14348 5014 14348 0 net374
rlabel metal1 4462 16490 4462 16490 0 net375
rlabel metal2 1242 15674 1242 15674 0 net376
rlabel metal1 3588 15674 3588 15674 0 net377
rlabel metal1 3496 6426 3496 6426 0 net378
rlabel metal2 1518 8211 1518 8211 0 net379
rlabel metal1 7774 26010 7774 26010 0 net38
rlabel metal1 3174 9350 3174 9350 0 net380
rlabel metal3 3565 9588 3565 9588 0 net381
rlabel metal1 5704 13498 5704 13498 0 net382
rlabel metal1 1472 10710 1472 10710 0 net383
rlabel metal2 15686 13889 15686 13889 0 net384
rlabel metal1 6946 9452 6946 9452 0 net385
rlabel metal2 8188 9860 8188 9860 0 net386
rlabel metal1 1518 6732 1518 6732 0 net387
rlabel metal1 5474 9962 5474 9962 0 net388
rlabel metal1 1472 7446 1472 7446 0 net389
rlabel metal2 15088 31756 15088 31756 0 net39
rlabel metal1 6946 11152 6946 11152 0 net390
rlabel metal1 4278 12104 4278 12104 0 net391
rlabel metal1 1840 7786 1840 7786 0 net392
rlabel metal1 2162 12376 2162 12376 0 net393
rlabel metal2 10718 32028 10718 32028 0 net394
rlabel metal1 13478 18938 13478 18938 0 net395
rlabel metal1 4646 37298 4646 37298 0 net396
rlabel metal1 6532 19822 6532 19822 0 net397
rlabel metal2 12558 35326 12558 35326 0 net398
rlabel metal1 10580 21318 10580 21318 0 net399
rlabel metal1 2070 17782 2070 17782 0 net4
rlabel metal1 1702 24378 1702 24378 0 net40
rlabel metal1 2254 20434 2254 20434 0 net400
rlabel metal1 2346 35054 2346 35054 0 net401
rlabel metal1 14076 36346 14076 36346 0 net402
rlabel metal1 18814 17204 18814 17204 0 net403
rlabel metal1 8372 30906 8372 30906 0 net404
rlabel metal1 8786 18326 8786 18326 0 net405
rlabel metal1 16054 16082 16054 16082 0 net406
rlabel metal1 6578 37230 6578 37230 0 net407
rlabel metal1 7636 17646 7636 17646 0 net408
rlabel metal1 15594 32402 15594 32402 0 net409
rlabel metal2 5382 26180 5382 26180 0 net41
rlabel metal2 5566 28237 5566 28237 0 net42
rlabel metal1 7222 21930 7222 21930 0 net43
rlabel metal1 2990 28050 2990 28050 0 net44
rlabel via2 2530 26843 2530 26843 0 net45
rlabel metal2 14168 31756 14168 31756 0 net46
rlabel metal1 15364 24174 15364 24174 0 net47
rlabel metal1 4002 33456 4002 33456 0 net48
rlabel metal1 19550 26928 19550 26928 0 net49
rlabel via2 1610 20315 1610 20315 0 net5
rlabel metal2 19688 28900 19688 28900 0 net50
rlabel metal1 2467 18258 2467 18258 0 net51
rlabel metal3 15916 33592 15916 33592 0 net52
rlabel metal1 19550 32368 19550 32368 0 net53
rlabel metal1 1702 39032 1702 39032 0 net54
rlabel metal1 16283 31790 16283 31790 0 net55
rlabel via1 15409 25262 15409 25262 0 net56
rlabel metal2 1702 40239 1702 40239 0 net57
rlabel metal1 19872 36754 19872 36754 0 net58
rlabel metal1 17756 33082 17756 33082 0 net59
rlabel metal1 2990 21862 2990 21862 0 net6
rlabel via1 19825 30226 19825 30226 0 net60
rlabel metal1 17940 18734 17940 18734 0 net61
rlabel metal2 1610 40052 1610 40052 0 net62
rlabel metal1 20010 20434 20010 20434 0 net63
rlabel metal2 2622 39525 2622 39525 0 net64
rlabel metal1 19625 16082 19625 16082 0 net65
rlabel metal3 1932 39780 1932 39780 0 net66
rlabel metal3 2300 17884 2300 17884 0 net67
rlabel metal1 18262 39372 18262 39372 0 net68
rlabel metal1 1931 38318 1931 38318 0 net69
rlabel metal1 5060 21862 5060 21862 0 net7
rlabel via1 18077 14994 18077 14994 0 net70
rlabel metal1 21022 13498 21022 13498 0 net71
rlabel via2 2254 41531 2254 41531 0 net72
rlabel metal3 14260 15164 14260 15164 0 net73
rlabel metal2 1886 33779 1886 33779 0 net74
rlabel metal3 2277 21148 2277 21148 0 net75
rlabel metal2 1702 34459 1702 34459 0 net76
rlabel viali 19541 10000 19541 10000 0 net77
rlabel metal1 19550 10676 19550 10676 0 net78
rlabel metal1 16513 18734 16513 18734 0 net79
rlabel metal1 11684 35054 11684 35054 0 net8
rlabel metal1 13018 12750 13018 12750 0 net80
rlabel metal1 21160 1258 21160 1258 0 net81
rlabel metal1 17342 12818 17342 12818 0 net82
rlabel metal3 15709 2380 15709 2380 0 net83
rlabel metal3 15824 2516 15824 2516 0 net84
rlabel metal1 20976 3026 20976 3026 0 net85
rlabel metal1 20010 3026 20010 3026 0 net86
rlabel metal1 20792 3502 20792 3502 0 net87
rlabel metal1 20608 3026 20608 3026 0 net88
rlabel metal3 15249 1972 15249 1972 0 net89
rlabel metal3 2714 21080 2714 21080 0 net9
rlabel metal2 21436 2380 21436 2380 0 net90
rlabel metal1 20700 3094 20700 3094 0 net91
rlabel metal2 17066 1785 17066 1785 0 net92
rlabel metal1 1702 36210 1702 36210 0 net93
rlabel metal1 21206 1870 21206 1870 0 net94
rlabel via2 17618 2499 17618 2499 0 net95
rlabel metal1 6348 8398 6348 8398 0 net96
rlabel metal2 20102 2621 20102 2621 0 net97
rlabel metal1 21988 1326 21988 1326 0 net98
rlabel metal1 1978 38794 1978 38794 0 net99
rlabel metal1 15916 39066 15916 39066 0 strobe_inbuf_0.X
rlabel metal1 16192 36346 16192 36346 0 strobe_inbuf_1.X
rlabel metal2 17986 13209 17986 13209 0 strobe_inbuf_10.X
rlabel metal1 21344 2074 21344 2074 0 strobe_inbuf_11.X
rlabel metal1 20332 2618 20332 2618 0 strobe_inbuf_12.X
rlabel metal2 21896 33252 21896 33252 0 strobe_inbuf_13.X
rlabel metal3 19412 20876 19412 20876 0 strobe_inbuf_14.X
rlabel metal1 21758 3570 21758 3570 0 strobe_inbuf_15.X
rlabel metal3 20861 19788 20861 19788 0 strobe_inbuf_16.X
rlabel metal3 22402 20876 22402 20876 0 strobe_inbuf_17.X
rlabel metal1 20976 2074 20976 2074 0 strobe_inbuf_18.X
rlabel metal3 19665 32844 19665 32844 0 strobe_inbuf_19.X
rlabel metal1 16100 38522 16100 38522 0 strobe_inbuf_2.X
rlabel metal1 16560 40902 16560 40902 0 strobe_inbuf_3.X
rlabel metal1 16974 40970 16974 40970 0 strobe_inbuf_4.X
rlabel metal2 17526 40052 17526 40052 0 strobe_inbuf_5.X
rlabel metal2 17066 28543 17066 28543 0 strobe_inbuf_6.X
rlabel metal1 17112 33626 17112 33626 0 strobe_inbuf_7.X
rlabel metal1 17572 39610 17572 39610 0 strobe_inbuf_8.X
rlabel metal1 17526 38522 17526 38522 0 strobe_inbuf_9.X
rlabel metal1 16146 39610 16146 39610 0 strobe_outbuf_0.X
rlabel metal1 16330 36890 16330 36890 0 strobe_outbuf_1.X
rlabel metal2 18354 41004 18354 41004 0 strobe_outbuf_10.X
rlabel metal1 19366 41480 19366 41480 0 strobe_outbuf_11.X
rlabel metal3 18630 41004 18630 41004 0 strobe_outbuf_12.X
rlabel metal1 19412 41090 19412 41090 0 strobe_outbuf_13.X
rlabel metal1 18262 40052 18262 40052 0 strobe_outbuf_14.X
rlabel metal1 19136 39814 19136 39814 0 strobe_outbuf_15.X
rlabel metal1 20148 39066 20148 39066 0 strobe_outbuf_16.X
rlabel metal1 18630 40018 18630 40018 0 strobe_outbuf_17.X
rlabel metal1 18722 40154 18722 40154 0 strobe_outbuf_18.X
rlabel metal1 19274 39610 19274 39610 0 strobe_outbuf_19.X
rlabel metal1 18354 41106 18354 41106 0 strobe_outbuf_2.X
rlabel metal3 19941 41276 19941 41276 0 strobe_outbuf_3.X
rlabel metal1 20930 41106 20930 41106 0 strobe_outbuf_4.X
rlabel metal1 18906 41548 18906 41548 0 strobe_outbuf_5.X
rlabel metal1 18078 41130 18078 41130 0 strobe_outbuf_6.X
rlabel metal1 18078 40086 18078 40086 0 strobe_outbuf_7.X
rlabel metal1 17572 40154 17572 40154 0 strobe_outbuf_8.X
rlabel metal1 18170 39270 18170 39270 0 strobe_outbuf_9.X
<< properties >>
string FIXED_BBOX 0 0 23000 44700
<< end >>
